VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sram_ifc
  CLASS BLOCK ;
  FOREIGN sram_ifc ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 400.000 ;
  PIN addr_r[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 57.840 150.000 58.440 ;
    END
  END addr_r[0]
  PIN addr_r[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 360.440 150.000 361.040 ;
    END
  END addr_r[10]
  PIN addr_r[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 200.640 150.000 201.240 ;
    END
  END addr_r[11]
  PIN addr_r[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 55.290 396.000 55.570 400.000 ;
    END
  END addr_r[12]
  PIN addr_r[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 316.240 150.000 316.840 ;
    END
  END addr_r[13]
  PIN addr_r[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END addr_r[1]
  PIN addr_r[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.390 396.000 48.670 400.000 ;
    END
  END addr_r[2]
  PIN addr_r[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 140.390 0.000 140.670 4.000 ;
    END
  END addr_r[3]
  PIN addr_r[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END addr_r[4]
  PIN addr_r[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END addr_r[5]
  PIN addr_r[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END addr_r[6]
  PIN addr_r[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END addr_r[7]
  PIN addr_r[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 46.090 0.000 46.370 4.000 ;
    END
  END addr_r[8]
  PIN addr_r[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 299.240 4.000 299.840 ;
    END
  END addr_r[9]
  PIN addr_w[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END addr_w[0]
  PIN addr_w[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END addr_w[10]
  PIN addr_w[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 251.640 4.000 252.240 ;
    END
  END addr_w[11]
  PIN addr_w[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 44.240 150.000 44.840 ;
    END
  END addr_w[12]
  PIN addr_w[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END addr_w[13]
  PIN addr_w[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END addr_w[1]
  PIN addr_w[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 173.440 150.000 174.040 ;
    END
  END addr_w[2]
  PIN addr_w[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 0.040 150.000 0.640 ;
    END
  END addr_w[3]
  PIN addr_w[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 78.240 150.000 78.840 ;
    END
  END addr_w[4]
  PIN addr_w[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END addr_w[5]
  PIN addr_w[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END addr_w[6]
  PIN addr_w[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.490 0.000 18.770 4.000 ;
    END
  END addr_w[7]
  PIN addr_w[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 268.640 4.000 269.240 ;
    END
  END addr_w[8]
  PIN addr_w[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 258.440 4.000 259.040 ;
    END
  END addr_w[9]
  PIN baseaddr_r_sync[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 248.240 150.000 248.840 ;
    END
  END baseaddr_r_sync[0]
  PIN baseaddr_r_sync[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.690 396.000 73.970 400.000 ;
    END
  END baseaddr_r_sync[1]
  PIN baseaddr_r_sync[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 108.840 150.000 109.440 ;
    END
  END baseaddr_r_sync[2]
  PIN baseaddr_r_sync[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END baseaddr_r_sync[3]
  PIN baseaddr_r_sync[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 153.040 150.000 153.640 ;
    END
  END baseaddr_r_sync[4]
  PIN baseaddr_r_sync[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 101.290 0.000 101.570 4.000 ;
    END
  END baseaddr_r_sync[5]
  PIN baseaddr_r_sync[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 132.640 150.000 133.240 ;
    END
  END baseaddr_r_sync[6]
  PIN baseaddr_r_sync[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END baseaddr_r_sync[7]
  PIN baseaddr_r_sync[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 82.890 396.000 83.170 400.000 ;
    END
  END baseaddr_r_sync[8]
  PIN baseaddr_w_sync[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END baseaddr_w_sync[0]
  PIN baseaddr_w_sync[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 367.240 150.000 367.840 ;
    END
  END baseaddr_w_sync[1]
  PIN baseaddr_w_sync[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.990 0.000 30.270 4.000 ;
    END
  END baseaddr_w_sync[2]
  PIN baseaddr_w_sync[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END baseaddr_w_sync[3]
  PIN baseaddr_w_sync[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 4.690 396.000 4.970 400.000 ;
    END
  END baseaddr_w_sync[4]
  PIN baseaddr_w_sync[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 117.390 396.000 117.670 400.000 ;
    END
  END baseaddr_w_sync[5]
  PIN baseaddr_w_sync[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.290 0.000 124.570 4.000 ;
    END
  END baseaddr_w_sync[6]
  PIN baseaddr_w_sync[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END baseaddr_w_sync[7]
  PIN baseaddr_w_sync[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 61.240 150.000 61.840 ;
    END
  END baseaddr_w_sync[8]
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END clk
  PIN conf[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.390 396.000 71.670 400.000 ;
    END
  END conf[0]
  PIN conf[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 92.090 0.000 92.370 4.000 ;
    END
  END conf[1]
  PIN conf[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 227.840 150.000 228.440 ;
    END
  END conf[2]
  PIN csb
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 95.240 150.000 95.840 ;
    END
  END csb
  PIN csb0_sync
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 138.090 396.000 138.370 400.000 ;
    END
  END csb0_sync
  PIN csb1_sync
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 292.440 4.000 293.040 ;
    END
  END csb1_sync
  PIN d_fabric_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 68.040 150.000 68.640 ;
    END
  END d_fabric_in[0]
  PIN d_fabric_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 10.240 150.000 10.840 ;
    END
  END d_fabric_in[10]
  PIN d_fabric_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.690 396.000 50.970 400.000 ;
    END
  END d_fabric_in[11]
  PIN d_fabric_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 391.040 150.000 391.640 ;
    END
  END d_fabric_in[12]
  PIN d_fabric_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END d_fabric_in[13]
  PIN d_fabric_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END d_fabric_in[14]
  PIN d_fabric_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END d_fabric_in[15]
  PIN d_fabric_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 87.490 396.000 87.770 400.000 ;
    END
  END d_fabric_in[16]
  PIN d_fabric_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 384.240 150.000 384.840 ;
    END
  END d_fabric_in[17]
  PIN d_fabric_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 333.240 150.000 333.840 ;
    END
  END d_fabric_in[18]
  PIN d_fabric_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 140.390 396.000 140.670 400.000 ;
    END
  END d_fabric_in[19]
  PIN d_fabric_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END d_fabric_in[1]
  PIN d_fabric_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 103.590 0.000 103.870 4.000 ;
    END
  END d_fabric_in[20]
  PIN d_fabric_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 323.040 150.000 323.640 ;
    END
  END d_fabric_in[21]
  PIN d_fabric_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 74.840 150.000 75.440 ;
    END
  END d_fabric_in[22]
  PIN d_fabric_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 282.240 150.000 282.840 ;
    END
  END d_fabric_in[23]
  PIN d_fabric_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 187.040 4.000 187.640 ;
    END
  END d_fabric_in[24]
  PIN d_fabric_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 101.290 396.000 101.570 400.000 ;
    END
  END d_fabric_in[25]
  PIN d_fabric_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 360.440 4.000 361.040 ;
    END
  END d_fabric_in[26]
  PIN d_fabric_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END d_fabric_in[27]
  PIN d_fabric_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 265.240 150.000 265.840 ;
    END
  END d_fabric_in[28]
  PIN d_fabric_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 299.240 150.000 299.840 ;
    END
  END d_fabric_in[29]
  PIN d_fabric_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END d_fabric_in[2]
  PIN d_fabric_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 102.040 150.000 102.640 ;
    END
  END d_fabric_in[30]
  PIN d_fabric_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END d_fabric_in[31]
  PIN d_fabric_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 27.240 150.000 27.840 ;
    END
  END d_fabric_in[3]
  PIN d_fabric_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 89.790 396.000 90.070 400.000 ;
    END
  END d_fabric_in[4]
  PIN d_fabric_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.790 396.000 67.070 400.000 ;
    END
  END d_fabric_in[5]
  PIN d_fabric_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END d_fabric_in[6]
  PIN d_fabric_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 397.840 150.000 398.440 ;
    END
  END d_fabric_in[7]
  PIN d_fabric_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END d_fabric_in[8]
  PIN d_fabric_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END d_fabric_in[9]
  PIN d_fabric_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END d_fabric_out[0]
  PIN d_fabric_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END d_fabric_out[10]
  PIN d_fabric_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 3.440 150.000 4.040 ;
    END
  END d_fabric_out[11]
  PIN d_fabric_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 350.240 150.000 350.840 ;
    END
  END d_fabric_out[12]
  PIN d_fabric_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 75.990 0.000 76.270 4.000 ;
    END
  END d_fabric_out[13]
  PIN d_fabric_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 17.040 150.000 17.640 ;
    END
  END d_fabric_out[14]
  PIN d_fabric_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 9.290 396.000 9.570 400.000 ;
    END
  END d_fabric_out[15]
  PIN d_fabric_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 292.440 150.000 293.040 ;
    END
  END d_fabric_out[16]
  PIN d_fabric_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 62.190 396.000 62.470 400.000 ;
    END
  END d_fabric_out[17]
  PIN d_fabric_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END d_fabric_out[18]
  PIN d_fabric_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 159.840 150.000 160.440 ;
    END
  END d_fabric_out[19]
  PIN d_fabric_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 147.290 0.000 147.570 4.000 ;
    END
  END d_fabric_out[1]
  PIN d_fabric_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END d_fabric_out[20]
  PIN d_fabric_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END d_fabric_out[21]
  PIN d_fabric_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END d_fabric_out[22]
  PIN d_fabric_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END d_fabric_out[23]
  PIN d_fabric_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 234.640 150.000 235.240 ;
    END
  END d_fabric_out[24]
  PIN d_fabric_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END d_fabric_out[25]
  PIN d_fabric_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END d_fabric_out[26]
  PIN d_fabric_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END d_fabric_out[27]
  PIN d_fabric_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 11.590 396.000 11.870 400.000 ;
    END
  END d_fabric_out[28]
  PIN d_fabric_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END d_fabric_out[29]
  PIN d_fabric_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END d_fabric_out[2]
  PIN d_fabric_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 27.690 396.000 27.970 400.000 ;
    END
  END d_fabric_out[30]
  PIN d_fabric_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 149.590 396.000 149.870 400.000 ;
    END
  END d_fabric_out[31]
  PIN d_fabric_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 105.890 396.000 106.170 400.000 ;
    END
  END d_fabric_out[3]
  PIN d_fabric_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 34.040 150.000 34.640 ;
    END
  END d_fabric_out[4]
  PIN d_fabric_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 343.440 150.000 344.040 ;
    END
  END d_fabric_out[5]
  PIN d_fabric_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 326.440 150.000 327.040 ;
    END
  END d_fabric_out[6]
  PIN d_fabric_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 268.640 150.000 269.240 ;
    END
  END d_fabric_out[7]
  PIN d_fabric_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END d_fabric_out[8]
  PIN d_fabric_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END d_fabric_out[9]
  PIN d_sram_in[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END d_sram_in[0]
  PIN d_sram_in[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 217.640 150.000 218.240 ;
    END
  END d_sram_in[10]
  PIN d_sram_in[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 210.840 150.000 211.440 ;
    END
  END d_sram_in[11]
  PIN d_sram_in[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 32.290 396.000 32.570 400.000 ;
    END
  END d_sram_in[12]
  PIN d_sram_in[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END d_sram_in[13]
  PIN d_sram_in[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END d_sram_in[14]
  PIN d_sram_in[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END d_sram_in[15]
  PIN d_sram_in[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 190.440 150.000 191.040 ;
    END
  END d_sram_in[16]
  PIN d_sram_in[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 142.840 150.000 143.440 ;
    END
  END d_sram_in[17]
  PIN d_sram_in[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END d_sram_in[18]
  PIN d_sram_in[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 374.040 150.000 374.640 ;
    END
  END d_sram_in[19]
  PIN d_sram_in[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END d_sram_in[1]
  PIN d_sram_in[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END d_sram_in[20]
  PIN d_sram_in[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 309.440 150.000 310.040 ;
    END
  END d_sram_in[21]
  PIN d_sram_in[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.190 0.000 85.470 4.000 ;
    END
  END d_sram_in[22]
  PIN d_sram_in[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END d_sram_in[23]
  PIN d_sram_in[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 115.640 150.000 116.240 ;
    END
  END d_sram_in[24]
  PIN d_sram_in[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 128.890 396.000 129.170 400.000 ;
    END
  END d_sram_in[25]
  PIN d_sram_in[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.490 0.000 41.770 4.000 ;
    END
  END d_sram_in[26]
  PIN d_sram_in[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 377.440 4.000 378.040 ;
    END
  END d_sram_in[27]
  PIN d_sram_in[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END d_sram_in[28]
  PIN d_sram_in[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 119.040 150.000 119.640 ;
    END
  END d_sram_in[29]
  PIN d_sram_in[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 34.590 0.000 34.870 4.000 ;
    END
  END d_sram_in[2]
  PIN d_sram_in[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 34.590 396.000 34.870 400.000 ;
    END
  END d_sram_in[30]
  PIN d_sram_in[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 176.840 150.000 177.440 ;
    END
  END d_sram_in[31]
  PIN d_sram_in[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END d_sram_in[3]
  PIN d_sram_in[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 16.190 396.000 16.470 400.000 ;
    END
  END d_sram_in[4]
  PIN d_sram_in[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 207.440 150.000 208.040 ;
    END
  END d_sram_in[5]
  PIN d_sram_in[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END d_sram_in[6]
  PIN d_sram_in[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 40.840 150.000 41.440 ;
    END
  END d_sram_in[7]
  PIN d_sram_in[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 20.440 150.000 21.040 ;
    END
  END d_sram_in[8]
  PIN d_sram_in[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 224.440 150.000 225.040 ;
    END
  END d_sram_in[9]
  PIN d_sram_out[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END d_sram_out[0]
  PIN d_sram_out[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 50.690 0.000 50.970 4.000 ;
    END
  END d_sram_out[10]
  PIN d_sram_out[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END d_sram_out[11]
  PIN d_sram_out[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END d_sram_out[12]
  PIN d_sram_out[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 43.790 396.000 44.070 400.000 ;
    END
  END d_sram_out[13]
  PIN d_sram_out[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END d_sram_out[14]
  PIN d_sram_out[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 121.990 396.000 122.270 400.000 ;
    END
  END d_sram_out[15]
  PIN d_sram_out[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.590 0.000 57.870 4.000 ;
    END
  END d_sram_out[16]
  PIN d_sram_out[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 380.840 150.000 381.440 ;
    END
  END d_sram_out[17]
  PIN d_sram_out[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END d_sram_out[18]
  PIN d_sram_out[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 110.490 396.000 110.770 400.000 ;
    END
  END d_sram_out[19]
  PIN d_sram_out[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 306.040 150.000 306.640 ;
    END
  END d_sram_out[1]
  PIN d_sram_out[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 136.040 150.000 136.640 ;
    END
  END d_sram_out[20]
  PIN d_sram_out[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END d_sram_out[21]
  PIN d_sram_out[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.890 0.000 14.170 4.000 ;
    END
  END d_sram_out[22]
  PIN d_sram_out[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 112.790 396.000 113.070 400.000 ;
    END
  END d_sram_out[23]
  PIN d_sram_out[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 85.040 150.000 85.640 ;
    END
  END d_sram_out[24]
  PIN d_sram_out[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END d_sram_out[25]
  PIN d_sram_out[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 124.290 396.000 124.570 400.000 ;
    END
  END d_sram_out[26]
  PIN d_sram_out[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 125.840 150.000 126.440 ;
    END
  END d_sram_out[27]
  PIN d_sram_out[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 62.190 0.000 62.470 4.000 ;
    END
  END d_sram_out[28]
  PIN d_sram_out[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 142.690 0.000 142.970 4.000 ;
    END
  END d_sram_out[29]
  PIN d_sram_out[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 357.040 150.000 357.640 ;
    END
  END d_sram_out[2]
  PIN d_sram_out[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END d_sram_out[30]
  PIN d_sram_out[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 244.840 4.000 245.440 ;
    END
  END d_sram_out[31]
  PIN d_sram_out[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 193.840 150.000 194.440 ;
    END
  END d_sram_out[3]
  PIN d_sram_out[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.990 0.000 53.270 4.000 ;
    END
  END d_sram_out[4]
  PIN d_sram_out[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 23.090 0.000 23.370 4.000 ;
    END
  END d_sram_out[5]
  PIN d_sram_out[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 146.000 275.440 150.000 276.040 ;
    END
  END d_sram_out[6]
  PIN d_sram_out[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END d_sram_out[7]
  PIN d_sram_out[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END d_sram_out[8]
  PIN d_sram_out[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END d_sram_out[9]
  PIN out_reg
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 94.390 396.000 94.670 400.000 ;
    END
  END out_reg
  PIN reb
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END reb
  PIN w_mask[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 91.840 150.000 92.440 ;
    END
  END w_mask[0]
  PIN w_mask[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 23.090 396.000 23.370 400.000 ;
    END
  END w_mask[10]
  PIN w_mask[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 340.040 150.000 340.640 ;
    END
  END w_mask[11]
  PIN w_mask[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END w_mask[12]
  PIN w_mask[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END w_mask[13]
  PIN w_mask[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END w_mask[14]
  PIN w_mask[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 36.890 0.000 37.170 4.000 ;
    END
  END w_mask[15]
  PIN w_mask[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.990 396.000 99.270 400.000 ;
    END
  END w_mask[16]
  PIN w_mask[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 144.990 396.000 145.270 400.000 ;
    END
  END w_mask[17]
  PIN w_mask[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 285.640 150.000 286.240 ;
    END
  END w_mask[18]
  PIN w_mask[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 115.090 0.000 115.370 4.000 ;
    END
  END w_mask[19]
  PIN w_mask[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 51.040 150.000 51.640 ;
    END
  END w_mask[1]
  PIN w_mask[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END w_mask[20]
  PIN w_mask[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 282.240 4.000 282.840 ;
    END
  END w_mask[21]
  PIN w_mask[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 78.290 396.000 78.570 400.000 ;
    END
  END w_mask[22]
  PIN w_mask[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END w_mask[23]
  PIN w_mask[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 25.390 0.000 25.670 4.000 ;
    END
  END w_mask[24]
  PIN w_mask[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 210.840 4.000 211.440 ;
    END
  END w_mask[25]
  PIN w_mask[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.890 396.000 60.170 400.000 ;
    END
  END w_mask[26]
  PIN w_mask[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END w_mask[27]
  PIN w_mask[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 39.190 396.000 39.470 400.000 ;
    END
  END w_mask[28]
  PIN w_mask[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 133.490 396.000 133.770 400.000 ;
    END
  END w_mask[29]
  PIN w_mask[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 0.090 396.000 0.370 400.000 ;
    END
  END w_mask[2]
  PIN w_mask[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END w_mask[30]
  PIN w_mask[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END w_mask[31]
  PIN w_mask[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 258.440 150.000 259.040 ;
    END
  END w_mask[3]
  PIN w_mask[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 241.440 150.000 242.040 ;
    END
  END w_mask[4]
  PIN w_mask[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 20.790 396.000 21.070 400.000 ;
    END
  END w_mask[5]
  PIN w_mask[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 183.640 150.000 184.240 ;
    END
  END w_mask[6]
  PIN w_mask[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 149.640 150.000 150.240 ;
    END
  END w_mask[7]
  PIN w_mask[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 251.640 150.000 252.240 ;
    END
  END w_mask[8]
  PIN w_mask[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 146.000 166.640 150.000 167.240 ;
    END
  END w_mask[9]
  PIN web
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END web
  PIN web0_sync
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END web0_sync
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 76.505 144.440 78.105 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 143.175 144.440 144.775 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 144.440 389.045 ;
      LAYER met1 ;
        RECT 5.520 10.640 145.290 389.200 ;
      LAYER met2 ;
        RECT 0.650 395.720 4.410 398.325 ;
        RECT 5.250 395.720 9.010 398.325 ;
        RECT 9.850 395.720 11.310 398.325 ;
        RECT 12.150 395.720 15.910 398.325 ;
        RECT 16.750 395.720 20.510 398.325 ;
        RECT 21.350 395.720 22.810 398.325 ;
        RECT 23.650 395.720 27.410 398.325 ;
        RECT 28.250 395.720 32.010 398.325 ;
        RECT 32.850 395.720 34.310 398.325 ;
        RECT 35.150 395.720 38.910 398.325 ;
        RECT 39.750 395.720 43.510 398.325 ;
        RECT 44.350 395.720 48.110 398.325 ;
        RECT 48.950 395.720 50.410 398.325 ;
        RECT 51.250 395.720 55.010 398.325 ;
        RECT 55.850 395.720 59.610 398.325 ;
        RECT 60.450 395.720 61.910 398.325 ;
        RECT 62.750 395.720 66.510 398.325 ;
        RECT 67.350 395.720 71.110 398.325 ;
        RECT 71.950 395.720 73.410 398.325 ;
        RECT 74.250 395.720 78.010 398.325 ;
        RECT 78.850 395.720 82.610 398.325 ;
        RECT 83.450 395.720 87.210 398.325 ;
        RECT 88.050 395.720 89.510 398.325 ;
        RECT 90.350 395.720 94.110 398.325 ;
        RECT 94.950 395.720 98.710 398.325 ;
        RECT 99.550 395.720 101.010 398.325 ;
        RECT 101.850 395.720 105.610 398.325 ;
        RECT 106.450 395.720 110.210 398.325 ;
        RECT 111.050 395.720 112.510 398.325 ;
        RECT 113.350 395.720 117.110 398.325 ;
        RECT 117.950 395.720 121.710 398.325 ;
        RECT 122.550 395.720 124.010 398.325 ;
        RECT 124.850 395.720 128.610 398.325 ;
        RECT 129.450 395.720 133.210 398.325 ;
        RECT 134.050 395.720 137.810 398.325 ;
        RECT 138.650 395.720 140.110 398.325 ;
        RECT 140.950 395.720 144.710 398.325 ;
        RECT 145.550 395.720 149.310 398.325 ;
        RECT 0.090 4.280 149.870 395.720 ;
        RECT 0.650 0.155 2.110 4.280 ;
        RECT 2.950 0.155 6.710 4.280 ;
        RECT 7.550 0.155 11.310 4.280 ;
        RECT 12.150 0.155 13.610 4.280 ;
        RECT 14.450 0.155 18.210 4.280 ;
        RECT 19.050 0.155 22.810 4.280 ;
        RECT 23.650 0.155 25.110 4.280 ;
        RECT 25.950 0.155 29.710 4.280 ;
        RECT 30.550 0.155 34.310 4.280 ;
        RECT 35.150 0.155 36.610 4.280 ;
        RECT 37.450 0.155 41.210 4.280 ;
        RECT 42.050 0.155 45.810 4.280 ;
        RECT 46.650 0.155 50.410 4.280 ;
        RECT 51.250 0.155 52.710 4.280 ;
        RECT 53.550 0.155 57.310 4.280 ;
        RECT 58.150 0.155 61.910 4.280 ;
        RECT 62.750 0.155 64.210 4.280 ;
        RECT 65.050 0.155 68.810 4.280 ;
        RECT 69.650 0.155 73.410 4.280 ;
        RECT 74.250 0.155 75.710 4.280 ;
        RECT 76.550 0.155 80.310 4.280 ;
        RECT 81.150 0.155 84.910 4.280 ;
        RECT 85.750 0.155 89.510 4.280 ;
        RECT 90.350 0.155 91.810 4.280 ;
        RECT 92.650 0.155 96.410 4.280 ;
        RECT 97.250 0.155 101.010 4.280 ;
        RECT 101.850 0.155 103.310 4.280 ;
        RECT 104.150 0.155 107.910 4.280 ;
        RECT 108.750 0.155 112.510 4.280 ;
        RECT 113.350 0.155 114.810 4.280 ;
        RECT 115.650 0.155 119.410 4.280 ;
        RECT 120.250 0.155 124.010 4.280 ;
        RECT 124.850 0.155 126.310 4.280 ;
        RECT 127.150 0.155 130.910 4.280 ;
        RECT 131.750 0.155 135.510 4.280 ;
        RECT 136.350 0.155 140.110 4.280 ;
        RECT 140.950 0.155 142.410 4.280 ;
        RECT 143.250 0.155 147.010 4.280 ;
        RECT 147.850 0.155 149.870 4.280 ;
      LAYER met3 ;
        RECT 4.400 397.440 145.600 398.305 ;
        RECT 0.065 392.040 149.895 397.440 ;
        RECT 4.400 390.640 145.600 392.040 ;
        RECT 0.065 385.240 149.895 390.640 ;
        RECT 4.400 383.840 145.600 385.240 ;
        RECT 0.065 381.840 149.895 383.840 ;
        RECT 0.065 380.440 145.600 381.840 ;
        RECT 0.065 378.440 149.895 380.440 ;
        RECT 4.400 377.040 149.895 378.440 ;
        RECT 0.065 375.040 149.895 377.040 ;
        RECT 4.400 373.640 145.600 375.040 ;
        RECT 0.065 368.240 149.895 373.640 ;
        RECT 4.400 366.840 145.600 368.240 ;
        RECT 0.065 361.440 149.895 366.840 ;
        RECT 4.400 360.040 145.600 361.440 ;
        RECT 0.065 358.040 149.895 360.040 ;
        RECT 4.400 356.640 145.600 358.040 ;
        RECT 0.065 351.240 149.895 356.640 ;
        RECT 4.400 349.840 145.600 351.240 ;
        RECT 0.065 344.440 149.895 349.840 ;
        RECT 4.400 343.040 145.600 344.440 ;
        RECT 0.065 341.040 149.895 343.040 ;
        RECT 4.400 339.640 145.600 341.040 ;
        RECT 0.065 334.240 149.895 339.640 ;
        RECT 4.400 332.840 145.600 334.240 ;
        RECT 0.065 327.440 149.895 332.840 ;
        RECT 4.400 326.040 145.600 327.440 ;
        RECT 0.065 324.040 149.895 326.040 ;
        RECT 0.065 322.640 145.600 324.040 ;
        RECT 0.065 320.640 149.895 322.640 ;
        RECT 4.400 319.240 149.895 320.640 ;
        RECT 0.065 317.240 149.895 319.240 ;
        RECT 4.400 315.840 145.600 317.240 ;
        RECT 0.065 310.440 149.895 315.840 ;
        RECT 4.400 309.040 145.600 310.440 ;
        RECT 0.065 307.040 149.895 309.040 ;
        RECT 0.065 305.640 145.600 307.040 ;
        RECT 0.065 303.640 149.895 305.640 ;
        RECT 4.400 302.240 149.895 303.640 ;
        RECT 0.065 300.240 149.895 302.240 ;
        RECT 4.400 298.840 145.600 300.240 ;
        RECT 0.065 293.440 149.895 298.840 ;
        RECT 4.400 292.040 145.600 293.440 ;
        RECT 0.065 286.640 149.895 292.040 ;
        RECT 4.400 285.240 145.600 286.640 ;
        RECT 0.065 283.240 149.895 285.240 ;
        RECT 4.400 281.840 145.600 283.240 ;
        RECT 0.065 276.440 149.895 281.840 ;
        RECT 4.400 275.040 145.600 276.440 ;
        RECT 0.065 269.640 149.895 275.040 ;
        RECT 4.400 268.240 145.600 269.640 ;
        RECT 0.065 266.240 149.895 268.240 ;
        RECT 4.400 264.840 145.600 266.240 ;
        RECT 0.065 259.440 149.895 264.840 ;
        RECT 4.400 258.040 145.600 259.440 ;
        RECT 0.065 252.640 149.895 258.040 ;
        RECT 4.400 251.240 145.600 252.640 ;
        RECT 0.065 249.240 149.895 251.240 ;
        RECT 0.065 247.840 145.600 249.240 ;
        RECT 0.065 245.840 149.895 247.840 ;
        RECT 4.400 244.440 149.895 245.840 ;
        RECT 0.065 242.440 149.895 244.440 ;
        RECT 4.400 241.040 145.600 242.440 ;
        RECT 0.065 235.640 149.895 241.040 ;
        RECT 4.400 234.240 145.600 235.640 ;
        RECT 0.065 228.840 149.895 234.240 ;
        RECT 4.400 227.440 145.600 228.840 ;
        RECT 0.065 225.440 149.895 227.440 ;
        RECT 4.400 224.040 145.600 225.440 ;
        RECT 0.065 218.640 149.895 224.040 ;
        RECT 4.400 217.240 145.600 218.640 ;
        RECT 0.065 211.840 149.895 217.240 ;
        RECT 4.400 210.440 145.600 211.840 ;
        RECT 0.065 208.440 149.895 210.440 ;
        RECT 4.400 207.040 145.600 208.440 ;
        RECT 0.065 201.640 149.895 207.040 ;
        RECT 4.400 200.240 145.600 201.640 ;
        RECT 0.065 194.840 149.895 200.240 ;
        RECT 4.400 193.440 145.600 194.840 ;
        RECT 0.065 191.440 149.895 193.440 ;
        RECT 0.065 190.040 145.600 191.440 ;
        RECT 0.065 188.040 149.895 190.040 ;
        RECT 4.400 186.640 149.895 188.040 ;
        RECT 0.065 184.640 149.895 186.640 ;
        RECT 4.400 183.240 145.600 184.640 ;
        RECT 0.065 177.840 149.895 183.240 ;
        RECT 4.400 176.440 145.600 177.840 ;
        RECT 0.065 174.440 149.895 176.440 ;
        RECT 0.065 173.040 145.600 174.440 ;
        RECT 0.065 171.040 149.895 173.040 ;
        RECT 4.400 169.640 149.895 171.040 ;
        RECT 0.065 167.640 149.895 169.640 ;
        RECT 4.400 166.240 145.600 167.640 ;
        RECT 0.065 160.840 149.895 166.240 ;
        RECT 4.400 159.440 145.600 160.840 ;
        RECT 0.065 154.040 149.895 159.440 ;
        RECT 4.400 152.640 145.600 154.040 ;
        RECT 0.065 150.640 149.895 152.640 ;
        RECT 4.400 149.240 145.600 150.640 ;
        RECT 0.065 143.840 149.895 149.240 ;
        RECT 4.400 142.440 145.600 143.840 ;
        RECT 0.065 137.040 149.895 142.440 ;
        RECT 4.400 135.640 145.600 137.040 ;
        RECT 0.065 133.640 149.895 135.640 ;
        RECT 4.400 132.240 145.600 133.640 ;
        RECT 0.065 126.840 149.895 132.240 ;
        RECT 4.400 125.440 145.600 126.840 ;
        RECT 0.065 120.040 149.895 125.440 ;
        RECT 4.400 118.640 145.600 120.040 ;
        RECT 0.065 116.640 149.895 118.640 ;
        RECT 0.065 115.240 145.600 116.640 ;
        RECT 0.065 113.240 149.895 115.240 ;
        RECT 4.400 111.840 149.895 113.240 ;
        RECT 0.065 109.840 149.895 111.840 ;
        RECT 4.400 108.440 145.600 109.840 ;
        RECT 0.065 103.040 149.895 108.440 ;
        RECT 4.400 101.640 145.600 103.040 ;
        RECT 0.065 96.240 149.895 101.640 ;
        RECT 4.400 94.840 145.600 96.240 ;
        RECT 0.065 92.840 149.895 94.840 ;
        RECT 4.400 91.440 145.600 92.840 ;
        RECT 0.065 86.040 149.895 91.440 ;
        RECT 4.400 84.640 145.600 86.040 ;
        RECT 0.065 79.240 149.895 84.640 ;
        RECT 4.400 77.840 145.600 79.240 ;
        RECT 0.065 75.840 149.895 77.840 ;
        RECT 4.400 74.440 145.600 75.840 ;
        RECT 0.065 69.040 149.895 74.440 ;
        RECT 4.400 67.640 145.600 69.040 ;
        RECT 0.065 62.240 149.895 67.640 ;
        RECT 4.400 60.840 145.600 62.240 ;
        RECT 0.065 58.840 149.895 60.840 ;
        RECT 0.065 57.440 145.600 58.840 ;
        RECT 0.065 55.440 149.895 57.440 ;
        RECT 4.400 54.040 149.895 55.440 ;
        RECT 0.065 52.040 149.895 54.040 ;
        RECT 4.400 50.640 145.600 52.040 ;
        RECT 0.065 45.240 149.895 50.640 ;
        RECT 4.400 43.840 145.600 45.240 ;
        RECT 0.065 41.840 149.895 43.840 ;
        RECT 0.065 40.440 145.600 41.840 ;
        RECT 0.065 38.440 149.895 40.440 ;
        RECT 4.400 37.040 149.895 38.440 ;
        RECT 0.065 35.040 149.895 37.040 ;
        RECT 4.400 33.640 145.600 35.040 ;
        RECT 0.065 28.240 149.895 33.640 ;
        RECT 4.400 26.840 145.600 28.240 ;
        RECT 0.065 21.440 149.895 26.840 ;
        RECT 4.400 20.040 145.600 21.440 ;
        RECT 0.065 18.040 149.895 20.040 ;
        RECT 4.400 16.640 145.600 18.040 ;
        RECT 0.065 11.240 149.895 16.640 ;
        RECT 4.400 9.840 145.600 11.240 ;
        RECT 0.065 4.440 149.895 9.840 ;
        RECT 4.400 3.040 145.600 4.440 ;
        RECT 0.065 1.040 149.895 3.040 ;
        RECT 0.065 0.175 145.600 1.040 ;
      LAYER met4 ;
        RECT 15.510 10.640 139.545 389.200 ;
      LAYER met5 ;
        RECT 5.520 146.375 144.440 344.770 ;
  END
END sram_ifc
END LIBRARY

