* NGSPICE file created from sram_ifc.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_4 abstract view
.subckt sky130_fd_sc_hd__dfxtp_4 D Q CLK VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_4 abstract view
.subckt sky130_fd_sc_hd__and4_4 A B C D X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_4 abstract view
.subckt sky130_fd_sc_hd__nor4_4 A B C D Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_4 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_4 A1_N A2_N B1 B2 X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C X VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_4 abstract view
.subckt sky130_fd_sc_hd__a32oi_4 A1 A2 A3 B1 B2 Y VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D Y VGND VPWR
.ends

.subckt sram_ifc addr_r[0] addr_r[10] addr_r[11] addr_r[12] addr_r[13] addr_r[1] addr_r[2]
+ addr_r[3] addr_r[4] addr_r[5] addr_r[6] addr_r[7] addr_r[8] addr_r[9] addr_w[0]
+ addr_w[10] addr_w[11] addr_w[12] addr_w[13] addr_w[1] addr_w[2] addr_w[3] addr_w[4]
+ addr_w[5] addr_w[6] addr_w[7] addr_w[8] addr_w[9] baseaddr_r_sync[0] baseaddr_r_sync[1]
+ baseaddr_r_sync[2] baseaddr_r_sync[3] baseaddr_r_sync[4] baseaddr_r_sync[5] baseaddr_r_sync[6]
+ baseaddr_r_sync[7] baseaddr_r_sync[8] baseaddr_w_sync[0] baseaddr_w_sync[1] baseaddr_w_sync[2]
+ baseaddr_w_sync[3] baseaddr_w_sync[4] baseaddr_w_sync[5] baseaddr_w_sync[6] baseaddr_w_sync[7]
+ baseaddr_w_sync[8] clk conf[0] conf[1] conf[2] csb csb0_sync csb1_sync d_fabric_in[0]
+ d_fabric_in[10] d_fabric_in[11] d_fabric_in[12] d_fabric_in[13] d_fabric_in[14]
+ d_fabric_in[15] d_fabric_in[16] d_fabric_in[17] d_fabric_in[18] d_fabric_in[19]
+ d_fabric_in[1] d_fabric_in[20] d_fabric_in[21] d_fabric_in[22] d_fabric_in[23] d_fabric_in[24]
+ d_fabric_in[25] d_fabric_in[26] d_fabric_in[27] d_fabric_in[28] d_fabric_in[29]
+ d_fabric_in[2] d_fabric_in[30] d_fabric_in[31] d_fabric_in[3] d_fabric_in[4] d_fabric_in[5]
+ d_fabric_in[6] d_fabric_in[7] d_fabric_in[8] d_fabric_in[9] d_fabric_out[0] d_fabric_out[10]
+ d_fabric_out[11] d_fabric_out[12] d_fabric_out[13] d_fabric_out[14] d_fabric_out[15]
+ d_fabric_out[16] d_fabric_out[17] d_fabric_out[18] d_fabric_out[19] d_fabric_out[1]
+ d_fabric_out[20] d_fabric_out[21] d_fabric_out[22] d_fabric_out[23] d_fabric_out[24]
+ d_fabric_out[25] d_fabric_out[26] d_fabric_out[27] d_fabric_out[28] d_fabric_out[29]
+ d_fabric_out[2] d_fabric_out[30] d_fabric_out[31] d_fabric_out[3] d_fabric_out[4]
+ d_fabric_out[5] d_fabric_out[6] d_fabric_out[7] d_fabric_out[8] d_fabric_out[9]
+ d_sram_in[0] d_sram_in[10] d_sram_in[11] d_sram_in[12] d_sram_in[13] d_sram_in[14]
+ d_sram_in[15] d_sram_in[16] d_sram_in[17] d_sram_in[18] d_sram_in[19] d_sram_in[1]
+ d_sram_in[20] d_sram_in[21] d_sram_in[22] d_sram_in[23] d_sram_in[24] d_sram_in[25]
+ d_sram_in[26] d_sram_in[27] d_sram_in[28] d_sram_in[29] d_sram_in[2] d_sram_in[30]
+ d_sram_in[31] d_sram_in[3] d_sram_in[4] d_sram_in[5] d_sram_in[6] d_sram_in[7] d_sram_in[8]
+ d_sram_in[9] d_sram_out[0] d_sram_out[10] d_sram_out[11] d_sram_out[12] d_sram_out[13]
+ d_sram_out[14] d_sram_out[15] d_sram_out[16] d_sram_out[17] d_sram_out[18] d_sram_out[19]
+ d_sram_out[1] d_sram_out[20] d_sram_out[21] d_sram_out[22] d_sram_out[23] d_sram_out[24]
+ d_sram_out[25] d_sram_out[26] d_sram_out[27] d_sram_out[28] d_sram_out[29] d_sram_out[2]
+ d_sram_out[30] d_sram_out[31] d_sram_out[3] d_sram_out[4] d_sram_out[5] d_sram_out[6]
+ d_sram_out[7] d_sram_out[8] d_sram_out[9] out_reg reb w_mask[0] w_mask[10] w_mask[11]
+ w_mask[12] w_mask[13] w_mask[14] w_mask[15] w_mask[16] w_mask[17] w_mask[18] w_mask[19]
+ w_mask[1] w_mask[20] w_mask[21] w_mask[22] w_mask[23] w_mask[24] w_mask[25] w_mask[26]
+ w_mask[27] w_mask[28] w_mask[29] w_mask[2] w_mask[30] w_mask[31] w_mask[3] w_mask[4]
+ w_mask[5] w_mask[6] w_mask[7] w_mask[8] w_mask[9] web web0_sync VPWR VGND
XFILLER_100_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_19 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_203 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_111 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_205 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0703__A _0629_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_155 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_133_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_214 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_269 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_280 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_291 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_159 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0613__A _0697_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_354 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1104__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0708__B1 _0707_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_252 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0765__A2_N _0528_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_394 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_36_258 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_239 VGND VPWR sky130_fd_sc_hd__fill_2
X_0985_ _0985_/A _0985_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0523__A _0523_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_24 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_383 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_331 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_364 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_300 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0650__A2 _0623_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_129 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1127__CLK _1127_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_191 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0608__A _0542_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0770_ _0762_/X _1089_/D _0769_/X d_fabric_out[6] VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_5_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_80 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_147 VGND VPWR sky130_fd_sc_hd__decap_4
X_1184_ d_fabric_in[18] _1184_/Q _1187_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_91_150 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0518__A _0587_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0632__A2 _0627_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_300 VGND VPWR sky130_fd_sc_hd__decap_12
X_0968_ _0968_/A _0968_/X VGND VPWR sky130_fd_sc_hd__buf_1
Xclkbuf_4_12_0_clk clkbuf_3_6_0_clk/X _1187_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0899_ _0899_/A _0899_/B _0903_/C _1177_/Q _0899_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0700__B _0700_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_28 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_309 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_277 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_117 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_44 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0871__A2 _0833_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_367 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_135_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0623__A2 _0620_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_198 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1144__D d_sram_out[29] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_139 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0847__C1 _0846_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0862__A2 _0839_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_93 VGND VPWR sky130_fd_sc_hd__decap_8
X_0822_ d_sram_in[0] _0880_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0753_ _0540_/D _0496_/A _0709_/X _0753_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_127_196 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0801__A _0776_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0684_ _0684_/A _0676_/X _0677_/X _0684_/D _0684_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
Xclkbuf_3_1_0_clk clkbuf_3_1_0_clk/A clkbuf_4_3_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_123_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_342 VGND VPWR sky130_fd_sc_hd__decap_12
X_1167_ d_fabric_in[1] _0827_/A _1175_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_161 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_183 VGND VPWR sky130_fd_sc_hd__fill_2
X_1098_ _0798_/X _1098_/Q _1127_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0853__A2 _0946_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_264 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_141 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1030__A2 _1025_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0711__A _0659_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_301 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_367 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_164 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_220 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_174 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1139__D d_sram_out[24] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_166 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0978__D _0991_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0780__A1 _0779_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0780__B2 _1091_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_361 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0994__C _0954_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1021_ _0978_/A _1021_/B _0978_/C _1024_/D _1021_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_93_278 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_131 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0930__B1_N _0873_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0805_ _0799_/X _1102_/Q _0695_/X _0801_/X d_fabric_out[19] VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__1012__A2 _0983_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0531__A _0580_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0736_ _0668_/X _1126_/Q _0501_/X _0735_/X _0736_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_103_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1065__C _1010_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0667_ _0493_/X _0750_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0598_ _0579_/C _0701_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1079__A2 _1040_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1219_ addr_r[7] baseaddr_r_sync[7] _1124_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_25_301 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_194 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0826__A2 _0943_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_312 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0817__A2 _1110_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0616__A _1151_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_94 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_56 VGND VPWR sky130_fd_sc_hd__decap_12
X_0521_ _0512_/X _0740_/B _0677_/C _1127_/Q _0546_/B VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_98_337 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_326 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0753__A1 _0540_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_1004_ _1003_/Y _1024_/D VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0526__A _0525_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_228 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0899__C _0903_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1160__CLK _1201_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_326 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_315 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_208 VGND VPWR sky130_fd_sc_hd__decap_3
X_0719_ _0651_/Y _0719_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_103_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_131 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_123 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_42 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_86 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0602__C _0702_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0735__A1 _0512_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0735__B2 _0771_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_201 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_191 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_289 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1152__D _1160_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_237 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0991__D _0991_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_170 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0671__B1 _0487_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_93 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_192 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1183__CLK _1187_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_145 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_123 VGND VPWR sky130_fd_sc_hd__decap_8
X_0504_ _0504_/A _0505_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_98_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_329 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0703__B _0700_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_229 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_123 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0613__B _0701_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0708__A1 _0705_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1147__D _1155_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_204 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_226 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_373 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0892__B1 _0891_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_270 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_0984_ _0843_/A _0985_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_113_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_170 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_310 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_36 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_192 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_395 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_376 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_398 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0714__A _0713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0938__A1 _1196_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1060__B1 _1057_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_115 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_159 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_118 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_204 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_310 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0874__B1 _0873_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0608__B _0524_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_354 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_240 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_62 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0624__A _0580_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0929__A1 _1188_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1051__B1 _1049_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1221__CLK _1221_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_80 VGND VPWR sky130_fd_sc_hd__decap_12
X_1183_ d_fabric_in[17] _1183_/Q _1187_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_91_162 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0865__B1 _0844_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_398 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0534__A _0580_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_312 VGND VPWR sky130_fd_sc_hd__decap_12
X_0967_ _0945_/Y _0966_/Y _0946_/X _0960_/X w_mask[1] VGND VPWR sky130_fd_sc_hd__a211o_4
X_0898_ _0895_/D _0877_/X _0897_/Y d_sram_in[10] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__0700__C _0656_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_284 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_273 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_159 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_310 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0709__A _0501_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0856__B1 _0855_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_27 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_128_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1033__B1 _1029_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_62 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0619__A _0619_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0847__B1 _0844_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_398 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1160__D _1223_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_184 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_379 VGND VPWR sky130_fd_sc_hd__decap_12
X_0821_ _0663_/A _1114_/Q _1146_/Q _0779_/X d_fabric_out[31] VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_80_93 VGND VPWR sky130_fd_sc_hd__decap_12
X_0752_ _0532_/X _0751_/X _0719_/X _0752_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_0683_ _0509_/B _0683_/B _0681_/X _0683_/D _0684_/D VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_43_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_298 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0529__A _0528_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1117__CLK _1187_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1166_ d_fabric_in[0] d_sram_in[0] _1175_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_302 VGND VPWR sky130_fd_sc_hd__decap_12
X_1097_ _0795_/X _1097_/Q _1142_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_100_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_326 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_121_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_298 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_129 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_184 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_154 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_379 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_232 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_85 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_178 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0780__A2 _1091_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1155__D _1226_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0994__D _0940_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_213 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_202 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_129 VGND VPWR sky130_fd_sc_hd__fill_2
X_1020_ _0998_/X _1018_/X _1019_/X w_mask[10] VGND VPWR sky130_fd_sc_hd__o21ai_4
Xclkbuf_4_11_0_clk clkbuf_3_5_0_clk/X _1161_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_19_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_110 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_198 VGND VPWR sky130_fd_sc_hd__decap_3
X_0804_ _0799_/X _1101_/Q _0594_/A _0801_/X d_fabric_out[18] VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_115_123 VGND VPWR sky130_fd_sc_hd__decap_12
X_0735_ _0512_/X _0677_/B _0739_/D _0695_/X _0771_/B _0735_/X VGND VPWR sky130_fd_sc_hd__a32o_4
X_0666_ _0663_/X _0660_/X _0665_/X d_fabric_out[0] VGND VPWR sky130_fd_sc_hd__a21o_4
X_0597_ _0725_/C _0617_/A _0597_/C _0619_/A VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_84_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_213 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0781__A1_N _0674_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_268 VGND VPWR sky130_fd_sc_hd__decap_4
X_1218_ addr_r[6] baseaddr_r_sync[6] _1124_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_184 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_132 VGND VPWR sky130_fd_sc_hd__fill_2
X_1149_ _1157_/Q _0620_/A _1174_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_25_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_198 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0722__A _0722_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_178 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_86 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_16_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_110 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_0_0_clk clkbuf_3_1_0_clk/A clkbuf_4_0_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_45_85 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_96 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0616__B _0505_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_51 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_68 VGND VPWR sky130_fd_sc_hd__decap_12
X_0520_ _0682_/C _0677_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0753__A2 _0496_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_202 VGND VPWR sky130_fd_sc_hd__fill_2
X_1003_ _0940_/D _1003_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_81_205 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0542__A _0681_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0899__D _1177_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0718_ _0718_/A _0716_/X _0501_/X _0717_/X _0718_/X VGND VPWR sky130_fd_sc_hd__or4_4
X_0649_ _0626_/Y _0632_/X _0636_/Y _0647_/X _0648_/Y _0649_/X VGND VPWR sky130_fd_sc_hd__o41a_4
XFILLER_103_159 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0717__A _0722_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_176 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_143 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_110_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_54 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_98 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0602__D _0602_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_251 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0735__A2 _0677_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_170 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_275 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_205 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0627__A _0562_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_249 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_154 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_112_90 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_198 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0671__A1 _0512_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_146 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_157 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0671__B2 _0771_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_160 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_7 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_240 VGND VPWR sky130_fd_sc_hd__decap_4
X_0503_ _0503_/A _0505_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_86_308 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_129 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_94_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_238 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0703__C _0701_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_135 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_319 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_330 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_208 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_135 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0613__C _0594_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_240 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0910__A _0866_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0708__A2 _0706_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1163__D _1163_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0892__A1 _0827_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_238 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1150__CLK _1127_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0983_ _0982_/X _0983_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_12_190 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0898__B1_N _0897_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_48 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_208 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_219 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_388 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_241 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0714__B _0714_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_285 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0938__A2 _0876_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1060__A1 _0992_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1173__CLK _1187_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_300 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0874__A1 _0872_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_322 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_86 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0905__A _0861_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_252 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_263 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0929__A2 _0926_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1158__D _1221_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1051__A1 _0966_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0640__A _0580_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_93 VGND VPWR sky130_fd_sc_hd__decap_12
X_1182_ d_fabric_in[16] _1182_/Q _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_83_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_333 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0865__A1 _0827_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_293 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0815__A out_reg VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_324 VGND VPWR sky130_fd_sc_hd__decap_12
X_0966_ _0966_/A _0966_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_133_316 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0550__A _0549_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0897_ _0847_/X _0896_/X _0897_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_99_252 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_230 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_403 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0700__D _1130_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1196__CLK _1116_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_300 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_322 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_182 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0856__A1 _0851_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_130 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_241 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0725__A _0725_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_403 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1033__A1 _0945_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_198 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_145 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0619__B _0612_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_171 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_130 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0847__A1 _0880_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0635__A _0526_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_196 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_263 VGND VPWR sky130_fd_sc_hd__decap_12
X_0820_ _0663_/A _1113_/Q _1113_/D _0815_/X d_fabric_out[30] VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_127_110 VGND VPWR sky130_fd_sc_hd__decap_12
X_0751_ _0668_/X _1127_/Q _0635_/C _0751_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_0682_ _0722_/A _0682_/B _0682_/C _1128_/Q _0683_/D VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_36_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_406 VGND VPWR sky130_fd_sc_hd__fill_1
X_1165_ _1165_/D csb1_sync _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1096_ _0793_/X _1096_/Q _1103_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_314 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0545__A _0545_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_154 VGND VPWR sky130_fd_sc_hd__decap_12
X_0949_ _0948_/X _0955_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_106_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0774__B1 _0709_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_277 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_152 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0829__A1 _0880_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_174 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1211__CLK _1174_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_32 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_391 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_110 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0765__B1 _0668_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_236 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1171__D d_fabric_in[5] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_141 VGND VPWR sky130_fd_sc_hd__decap_3
X_0803_ _0799_/X _1100_/Q _0487_/X _0801_/X d_fabric_out[17] VGND VPWR sky130_fd_sc_hd__o22a_4
X_0734_ _0663_/X _1085_/D _0733_/X d_fabric_out[2] VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0756__B1 _0755_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_135 VGND VPWR sky130_fd_sc_hd__decap_12
X_0665_ _0665_/A _0776_/A _0665_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_130_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_330 VGND VPWR sky130_fd_sc_hd__decap_12
X_0596_ _0695_/A _0580_/C _0718_/A _0526_/X _0595_/X _0597_/C VGND VPWR sky130_fd_sc_hd__a2111oi_4
XFILLER_29_119 VGND VPWR sky130_fd_sc_hd__decap_3
X_1217_ addr_r[5] baseaddr_r_sync[5] _1161_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_130 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_280 VGND VPWR sky130_fd_sc_hd__fill_2
X_1148_ _1156_/Q _1148_/Q _1174_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1079_ _0985_/A _1040_/X _1075_/Y _1079_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_33_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0778__A2_N _0496_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0722__B _0492_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_7 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0747__B1 _0695_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_214 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_239 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_306 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0616__C _1146_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1107__CLK _1103_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1166__D d_fabric_in[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_269 VGND VPWR sky130_fd_sc_hd__decap_6
X_1002_ _0998_/X _1001_/X _0996_/X w_mask[7] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_19_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0823__A _1226_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_361 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0542__B _0513_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0717_ _0722_/D _0656_/B _0717_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_131_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_106_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_0648_ _0509_/A _0629_/X _0622_/Y _0648_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XFILLER_97_350 VGND VPWR sky130_fd_sc_hd__fill_2
X_0579_ _0580_/A _0580_/C _0579_/C _1130_/Q _0579_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_57_214 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_100 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0717__B _0656_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_261 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0733__A _0733_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_282 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_10_0_clk clkbuf_3_5_0_clk/X _1221_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_134_263 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0735__A3 _0739_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_258 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0908__A _0903_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_74 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_217 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_280 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_283 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_51 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0671__A2 _0677_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_150 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_194 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0959__B1 _0958_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_172 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_361 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0643__A _0505_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_113_403 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0795__A1_N _0575_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0502_ _0502_/A _0509_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_98_158 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_94_320 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_203 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0553__A _0524_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0703__D _0702_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0728__A _0721_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_239 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0613__D _1141_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0910__B _0910_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_309 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_301 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0638__A _0722_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0892__A2 _0890_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_283 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_294 VGND VPWR sky130_fd_sc_hd__decap_12
X_0982_ _0991_/A _0982_/B _0991_/C _0991_/D _0982_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_66_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_364 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0548__A _0547_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_264 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_297 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1060__A2 _1059_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_266 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_320 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_161 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_334 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0874__A2 _0833_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_272 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0905__B _0904_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_275 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_97 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1051__A2 _1043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1174__D d_fabric_in[8] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_7 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_139 VGND VPWR sky130_fd_sc_hd__fill_2
X_1181_ d_fabric_in[15] _1181_/Q _1226_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_301 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_161 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_356 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0865__A2 _0859_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_197 VGND VPWR sky130_fd_sc_hd__fill_2
X_0965_ _0965_/A _0966_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0896_ _0846_/A _0890_/X _0895_/X _0896_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0831__A _1226_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_306 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1084__D _0712_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_334 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0856__A2 _0833_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0725__B _0544_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_337 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1033__A2 _1032_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0741__A _0544_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1140__CLK _1124_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_109 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_334 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_97 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0619__C _0618_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_291 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_73_153 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0847__A2 _0946_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0916__A _0903_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_304 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0635__B _0635_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_80 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1169__D d_fabric_in[3] VGND VPWR sky130_fd_sc_hd__diode_2
X_0750_ _0750_/A _0750_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0651__A _0500_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_306 VGND VPWR sky130_fd_sc_hd__decap_12
X_0681_ _0681_/A _0492_/C _0722_/C _0487_/X _0681_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_96_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_367 VGND VPWR sky130_fd_sc_hd__decap_12
X_1164_ web web0_sync _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1095_ _0790_/X _1095_/Q _1142_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_326 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_164 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_52_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0545__B _0545_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_223 VGND VPWR sky130_fd_sc_hd__fill_2
X_0948_ _0969_/A _0948_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0561__A _0585_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1163__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_306 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_59 VGND VPWR sky130_fd_sc_hd__fill_2
X_0879_ _1010_/C _1046_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0774__A1 _0580_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_201 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_131 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0829__A2 _0826_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_44 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_133_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_245 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_188 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0765__B2 _0724_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_74 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0646__A _0642_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_123 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_156 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_178 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1186__CLK _1226_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0802_ _0799_/X _1099_/Q _1099_/D _0801_/X d_fabric_out[16] VGND VPWR sky130_fd_sc_hd__o22a_4
X_0733_ _0733_/A _1085_/Q _0733_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0756__A1 _0663_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_147 VGND VPWR sky130_fd_sc_hd__decap_12
X_0664_ out_reg _0776_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_130_117 VGND VPWR sky130_fd_sc_hd__decap_12
X_0595_ _1132_/Q _0583_/C _0595_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_69_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_278 VGND VPWR sky130_fd_sc_hd__decap_12
X_1216_ addr_r[4] baseaddr_r_sync[4] _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0556__A _0581_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_101 VGND VPWR sky130_fd_sc_hd__decap_4
X_1147_ _1155_/Q _1147_/Q _1174_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_111_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_123 VGND VPWR sky130_fd_sc_hd__decap_3
X_1078_ _1032_/X _1070_/X _1076_/X w_mask[29] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_52_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_178 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0722__C _0722_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0747__A1 _0750_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0747__B2 _0496_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_337 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_167 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0616__D _0580_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_86 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_6_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_117 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1182__D d_fabric_in[16] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_226 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_131 VGND VPWR sky130_fd_sc_hd__decap_3
X_1001_ _1000_/X _1001_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_19_175 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_134 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1000__A _0978_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0542__C _0544_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0716_ _0716_/A _0720_/A _0716_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1201__CLK _1201_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_0647_ _0638_/X _0639_/X _0641_/X _0646_/X _0647_/X VGND VPWR sky130_fd_sc_hd__or4_4
X_0578_ _0578_/A _0578_/B _0574_/Y _0578_/D _0578_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XANTENNA__1092__D _1092_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_237 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_259 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_123 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_292 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_19 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_156 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_126 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0733__B _1085_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_294 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_244 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_299 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0908__B _0903_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_70 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0671__A3 _0676_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_140 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_63 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_151 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0959__A1 _0957_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_173 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_300 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0643__B _0643_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_162 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1081__B1 _1079_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1224__CLK _1161_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1177__D d_fabric_in[11] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_7 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_125_220 VGND VPWR sky130_fd_sc_hd__decap_12
X_0501_ _0500_/X _0501_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_94_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_11_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_248 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_207 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_270 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_115 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0834__A _0943_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_137 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1072__B1 _1071_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_209 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1087__D _0754_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_159 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_148 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_218 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0728__B _0728_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_240 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0744__A _0738_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_295 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1063__B1 _1061_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_88 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0810__B1 _0723_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_220 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_275 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_181 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0638__B _0558_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_313 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_262 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0654__A _0690_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0981_ _0981_/A _0991_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1054__B1 _1052_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_129 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_310 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_332 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0868__B1 _0867_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_335 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0564__A _0555_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_245 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0739__A _0722_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_151 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_346 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_357 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_232 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_118_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_215 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_310 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_129 VGND VPWR sky130_fd_sc_hd__decap_8
X_1180_ d_fabric_in[14] _0912_/D _1116_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_313 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1190__D d_fabric_in[24] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_173 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_143 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_368 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_276 VGND VPWR sky130_fd_sc_hd__decap_12
X_0964_ _0981_/A _1021_/B _0940_/C _0940_/D _0965_/A VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_118_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0831__B _0841_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0895_ _0899_/A _0899_/B _0903_/C _0895_/D _0895_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_99_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1092__CLK _1114_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_346 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_165 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_23_221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_210 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0725__C _0725_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_349 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0741__B _0513_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_178 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_125 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_65 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_140 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_302 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_110 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0916__B _0903_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_165 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0635__C _0635_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0932__A _0920_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_123 VGND VPWR sky130_fd_sc_hd__decap_12
X_0680_ _0544_/C _0722_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_115_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1185__D d_fabric_in[19] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_184 VGND VPWR sky130_fd_sc_hd__decap_4
X_1163_ _1163_/D csb0_sync _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1094_ _0788_/X _1094_/Q _1142_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1003__A _0940_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0545__C _0544_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0842__A _0841_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0947_ _0940_/A _0969_/A VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0561__B _0555_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_318 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0774__A2 _0659_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0878_ _0835_/X _1010_/C VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_133_159 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1095__D _0790_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_235 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_68 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_56 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_257 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_126_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_123 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_22 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_109_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_86 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_279 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_121 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0646__B _0643_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_154 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0662__A _0661_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0801_ _0776_/A _0801_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0756__A2 _0754_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0732_ out_reg _0733_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0610__D1 _0609_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0663_ _0663_/A _0663_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_115_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_0594_ _0594_/A _0594_/B _0718_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_130_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_257 VGND VPWR sky130_fd_sc_hd__decap_3
X_1215_ addr_r[3] baseaddr_r_sync[3] _1142_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0837__A _0836_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_260 VGND VPWR sky130_fd_sc_hd__fill_2
X_1146_ d_sram_out[31] _1146_/Q _1221_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0556__B _0490_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_198 VGND VPWR sky130_fd_sc_hd__fill_2
X_1077_ _1025_/X _1070_/X _1076_/X w_mask[28] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_52_157 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1130__CLK _1201_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0572__A _0571_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_218 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0722__D _0722_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0747__A2 _0736_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_404 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_249 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_165 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_187 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_282 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_135 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_66 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_179 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_251 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_231 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_129 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_238 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1153__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1000_ _0978_/A _0991_/B _1024_/C _0991_/D _1000_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_74_260 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_293 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_146 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_0_clk_A clk VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1000__B _0991_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_385 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0542__D _0542_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_251 VGND VPWR sky130_fd_sc_hd__decap_12
X_0715_ _0663_/X _0712_/X _0714_/X d_fabric_out[1] VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_89_319 VGND VPWR sky130_fd_sc_hd__fill_2
X_0646_ _0642_/X _0643_/X _0644_/X _0645_/X _0646_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA_clkbuf_4_9_0_clk_A clkbuf_4_8_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_330 VGND VPWR sky130_fd_sc_hd__fill_1
X_0577_ _0575_/Y _0576_/X _0518_/X _0628_/B _0578_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_111_184 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0567__A _0583_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_227 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_122_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_219 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_271 VGND VPWR sky130_fd_sc_hd__fill_2
X_1129_ d_sram_out[14] _0724_/D _1124_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_25_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_35 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1176__CLK _1185_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0908__C _0908_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_271 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_82 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_190 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_130 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_75 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_152 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0959__A2 _0838_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_174 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_312 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0643__C _0530_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_163 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1081__A1 _1040_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_385 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0940__A _0940_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_232 VGND VPWR sky130_fd_sc_hd__fill_2
X_0500_ _0499_/X _0500_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_98_138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_105 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1193__D d_fabric_in[27] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_363 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_238 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_230 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_105 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_62_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_149 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_127 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1011__A _1009_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1072__A1 _1018_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1199__CLK _1226_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_257 VGND VPWR sky130_fd_sc_hd__decap_12
X_0629_ _0628_/X _0629_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_133_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_193 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_133_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0728__C _0723_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_403 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0744__B _0744_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1063__A1 _1001_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_56 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0810__A1 _0806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0810__B2 _0808_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_287 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_208 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_336 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_241 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_74 VGND VPWR sky130_fd_sc_hd__decap_12
X_0980_ _0968_/X _0979_/X _0975_/Y w_mask[3] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__1054__A1 _0979_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1188__D d_fabric_in[22] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_7 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0670__A _0602_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_182 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1006__A _1005_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0868__A1 _0864_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_344 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_314 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_230 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0845__A _0835_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_35_241 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1098__D _0798_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0580__A _0580_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_224 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_6_0_clk_A clkbuf_3_7_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0739__B _0492_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1214__CLK _1142_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0755__A _0733_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_66 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0490__A _0490_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0795__B1 _1113_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_300 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_322 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_325 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0665__A _0665_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_222 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_288 VGND VPWR sky130_fd_sc_hd__decap_12
X_0963_ _0950_/Y _1021_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0786__B1 _0785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_0894_ _0891_/D _0877_/X _0893_/Y d_sram_in[9] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__0831__C _0835_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_205 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_216 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_174 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0575__A _0724_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_358 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0710__B1 _0709_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_196 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_391 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_188 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_233 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0725__D _0594_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0741__C _0724_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0777__B1 _0776_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_314 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_88 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0916__C _0908_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_177 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_288 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0768__B1 _0766_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_86 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_127_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_62 VGND VPWR sky130_fd_sc_hd__decap_12
X_1162_ _1225_/Q _1162_/Q _1185_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1093_ _0784_/X _1093_/Q _1103_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_45_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_203 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_361 VGND VPWR sky130_fd_sc_hd__decap_12
X_0946_ _0946_/A _0942_/Y _0946_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0561__C _1151_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0759__B1 _0719_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_0877_ _0876_/X _0877_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_126_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_306 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_68 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_56 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_341 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_300 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_2_3_0_clk_A clkbuf_2_3_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_217 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0646__C _0644_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_114 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0943__A _0836_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0989__B1 _0988_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_361 VGND VPWR sky130_fd_sc_hd__decap_12
X_0800_ _0713_/X _0798_/X _0799_/X _1098_/Q d_fabric_out[15] VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__1196__D d_fabric_in[30] VGND VPWR sky130_fd_sc_hd__diode_2
X_0731_ _0750_/A _0718_/X _0730_/X _0594_/A _0711_/X _1085_/D VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_6_251 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0610__C1 _0608_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0662_ _0661_/Y _0663_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_108_190 VGND VPWR sky130_fd_sc_hd__decap_8
X_0593_ _0587_/C _0594_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_123_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_236 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0913__B1 _0912_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_206 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_239 VGND VPWR sky130_fd_sc_hd__fill_2
X_1214_ addr_r[2] baseaddr_r_sync[2] _1142_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_100 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_133 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0837__B _0943_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_155 VGND VPWR sky130_fd_sc_hd__fill_2
X_1145_ d_sram_out[30] _1113_/D _1114_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1014__A _0991_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_272 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0556__C _0504_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1076_ _0985_/A _1035_/X _1075_/Y _1076_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA_clkbuf_4_5_0_clk_A clkbuf_3_2_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_0929_ _1188_/Q _0926_/X _0870_/X d_sram_in[22] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__0747__A3 _0746_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_300 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0904__B1 _0903_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_217 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_261 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_361 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0763__A _0733_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_62 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_219 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_274 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_105_171 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_193 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_155 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_209 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_272 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0673__A _0673_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1000__C _1024_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_263 VGND VPWR sky130_fd_sc_hd__decap_12
X_0714_ _0713_/X _0714_/B _0714_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0645_ _0583_/A _0643_/B _0530_/A _1121_/Q _0645_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__1009__A _1009_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0576_ _0587_/A _0585_/B _0725_/A _0505_/A _0576_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_111_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_217 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0848__A _0847_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0567__B _0580_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_250 VGND VPWR sky130_fd_sc_hd__fill_2
X_1128_ d_sram_out[13] _1128_/Q _1161_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_15_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0583__A _0583_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1059_ _1043_/A _1059_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_15_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_174 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_228 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0908__D _1179_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_209 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_88 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0493__A _0493_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_253 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_120 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_286 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_175 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0643__D _0724_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_87 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_153 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1081__A2 _1043_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_324 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0940__B _0956_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_117 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1120__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_51 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0668__A _0716_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_228 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_1_0_0_clk_A clkbuf_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0577__A1_N _0575_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_0 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1011__B _1028_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1072__A2 _1070_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_172 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_183 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_117_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_406 VGND VPWR sky130_fd_sc_hd__fill_1
X_0628_ _0580_/B _0628_/B _0628_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_131_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_301 VGND VPWR sky130_fd_sc_hd__fill_2
X_0559_ _0554_/Y _0557_/X _1128_/Q _0558_/X _0578_/A VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__0578__A _0578_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_334 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_323 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0728__D _0728_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_250 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_261 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_231 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0744__C _0740_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_2_0_clk_A clkbuf_3_3_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1063__A2 _1059_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_172 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_42_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0810__A2 _1105_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1143__CLK _1103_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_299 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0488__A _1147_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_312 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_323 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_13_0_clk_A clkbuf_3_6_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_348 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_80 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0951__A _0950_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1054__A2 _1043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_280 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0868__A2 _0833_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_356 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_209 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0845__B _0943_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1022__A _1021_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_381 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_245 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0861__A _0861_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1166__CLK _1175_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_289 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0580__B _0580_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_129_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_109 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0739__C _0722_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_24 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_356 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_304 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0755__B _0755_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_264 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_278 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_89 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0771__A _1138_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_306 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0795__B2 _0711_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_228 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_86 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_334 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0946__A _0946_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_123 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0665__B _0776_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_242 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1189__CLK _1187_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_201 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1199__D addr_w[1] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_234 VGND VPWR sky130_fd_sc_hd__decap_12
X_0962_ _0940_/A _0981_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0681__A _0681_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0786__B2 _1093_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0786__A1 _0779_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0893_ _0866_/A _0892_/X _0893_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_64_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_234 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_278 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_109 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1017__A _0978_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_304 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0710__A1 _0685_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_145 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_245 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0591__A _0552_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_306 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0741__D _1130_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0777__A1 _0762_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_158 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_56 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_58_175 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_326 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_134 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0916__D _1181_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0768__A1 _0723_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0768__B2 _0767_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_237 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_7 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_182 VGND VPWR sky130_fd_sc_hd__fill_1
X_1161_ _1224_/Q _1161_/Q _1161_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0676__A _0512_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_145 VGND VPWR sky130_fd_sc_hd__fill_2
X_1092_ _1092_/D _1092_/Q _1114_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_60_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_215 VGND VPWR sky130_fd_sc_hd__decap_8
X_0945_ _0945_/A _0945_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0561__D _0503_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0759__A1 _0757_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_293 VGND VPWR sky130_fd_sc_hd__decap_12
X_0876_ _0920_/B _0876_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1204__CLK _1175_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_1_0_clk_A clkbuf_4_0_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0931__A1 _1190_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0586__A _0585_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_123 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_156 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_318 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_353 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_237 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_50 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0496__A _0496_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_270 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_98 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0646__D _0645_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0989__A1 _0985_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0943__B _0943_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_80 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1227__CLK _1142_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0730_ _1117_/Q _0548_/X _0719_/X _0729_/X _0730_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__0610__B1 _0688_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_263 VGND VPWR sky130_fd_sc_hd__decap_12
X_0661_ out_reg _0661_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0592_ _0579_/C _0617_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0913__A1 _1172_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_367 VGND VPWR sky130_fd_sc_hd__decap_12
X_1213_ addr_r[1] baseaddr_r_sync[1] _1161_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_27_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_112 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_77_281 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0837__C _0835_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_51 VGND VPWR sky130_fd_sc_hd__decap_8
X_1144_ d_sram_out[29] _0678_/A _1175_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1014__B _1021_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1075_ _1066_/B _1074_/X _1048_/C _1075_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_25_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0556__D _0555_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0928_ _1187_/Q _0926_/X _0867_/X d_sram_in[21] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_106_117 VGND VPWR sky130_fd_sc_hd__decap_12
X_0859_ _0955_/D _0946_/A _0859_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_20_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0904__A1 _1170_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_240 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_24 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0763__B _0763_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_373 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_131_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_286 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_123 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0605__A2_N _0562_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_292 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0954__A _0954_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_251 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_398 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1000__D _0991_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0713_ out_reg _0713_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0644_ _0580_/A _0643_/B _0585_/C _0720_/A _0644_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__1009__B _1009_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0575_ _0724_/D _0575_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_111_153 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_354 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0567__C _0530_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1025__A _1024_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0864__A _1171_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_104 VGND VPWR sky130_fd_sc_hd__decap_12
X_1127_ d_sram_out[12] _1127_/Q _1127_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1058_ _0983_/X _1043_/X _1057_/X w_mask[20] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_15_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0583__B _0579_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_265 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_404 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_88_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_284 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_265 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_118 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_110 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_99 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_154 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0940__C _0940_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_245 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0949__A _0948_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_343 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_207 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_240 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0559__A2_N _0557_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0684__A _0684_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1057__B1 _1056_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1011__C _0988_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_181 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0804__B1 _0594_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0859__A _0955_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0627_ _0562_/X _0627_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0578__B _0578_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0558_ _0505_/B _1153_/Q _0725_/A _0505_/A _0558_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_133_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_162 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1095__CLK _1142_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_346 VGND VPWR sky130_fd_sc_hd__decap_12
X_0489_ _0503_/A _0490_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_85_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_210 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0594__A _0594_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_265 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_107 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_287 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0744__D _0743_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_215 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0769__A _0733_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_22 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_379 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_210 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_3_0_clk clkbuf_2_3_0_clk/A clkbuf_3_7_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_83_98 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_91 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_361 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0679__A _0722_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_292 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_154 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_327 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_187 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0845__C _0885_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_393 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_268 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0580__C _0580_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0589__A _0579_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0961__C1 _0960_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_110 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0739__D _0739_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_36 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_368 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_187 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_202 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1110__CLK _1103_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0771__B _0771_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_147 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0894__B1_N _0893_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0499__A _0620_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_270 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_49_346 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_132 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0946__B _0942_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_135 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_146 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_213 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0962__A _0940_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_246 VGND VPWR sky130_fd_sc_hd__decap_12
X_0961_ _0942_/Y _0945_/Y _0946_/X _0960_/X w_mask[0] VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__0681__B _0492_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0786__A2 _0784_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0892_ _0827_/A _0890_/X _0891_/X _0892_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_57_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_213 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1017__B _0982_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_19 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0710__A2 _0708_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1133__CLK _1116_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_308 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_190 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0872__A _1173_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0591__B _0591_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0777__A2 _1090_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_117 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_290 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_58_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0768__A2 _0750_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_71 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_249 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0957__A _0956_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0676__B _0492_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1160_ _1223_/Q _1160_/Q _1201_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1156__CLK _1174_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_124 VGND VPWR sky130_fd_sc_hd__fill_2
X_1091_ _1091_/D _1091_/Q _1127_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_64_157 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_179 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0692__A _0739_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_190 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_385 VGND VPWR sky130_fd_sc_hd__decap_12
X_0944_ _0968_/A _0945_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0759__A2 _0758_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0875_ _0833_/A _0920_/B VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1028__A _1028_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_398 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0931__A2 _0926_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0586__B _0585_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_105 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_124_129 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1179__CLK _1116_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_227 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_146 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0989__A2 _0974_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0943__C _0908_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_98 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_385 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0610__A1 _0675_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0660_ _0487_/X _0496_/X _0659_/X _0660_/X VGND VPWR sky130_fd_sc_hd__a21bo_4
X_0591_ _0552_/Y _0591_/B _0591_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_69_216 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_123_184 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0687__A _0675_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0913__A2 _1046_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_379 VGND VPWR sky130_fd_sc_hd__decap_12
X_1212_ addr_r[0] baseaddr_r_sync[0] _1185_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_77_260 VGND VPWR sky130_fd_sc_hd__fill_2
X_1143_ d_sram_out[28] _0532_/A _1103_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_1_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1014__C _0978_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1074_ _1009_/A _0957_/X _0973_/C _0987_/D _1074_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_37_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_149 VGND VPWR sky130_fd_sc_hd__fill_2
X_0927_ _1186_/Q _0926_/X _0862_/X d_sram_in[20] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_106_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_0858_ _0852_/B _0955_/D VGND VPWR sky130_fd_sc_hd__buf_1
X_0789_ _0779_/X _0788_/X _0785_/X _1094_/Q d_fabric_out[11] VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__0904__A2 _0890_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0597__A _0725_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_208 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_105 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_45_36 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_274 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_296 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_385 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_86 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_298 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_390 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_105 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_285 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_300 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0970__A _0956_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_276 VGND VPWR sky130_fd_sc_hd__decap_12
X_0712_ _0750_/A _0672_/X _0710_/Y _0487_/X _0711_/X _0712_/X VGND VPWR sky130_fd_sc_hd__a32o_4
X_0643_ _0505_/B _0643_/B _0530_/A _0724_/D _0643_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__1009__C _0991_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_110 VGND VPWR sky130_fd_sc_hd__decap_12
X_0574_ _0518_/X _0579_/C _0573_/Y _0574_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__0898__A1 _0895_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_165 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0567__D _1118_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_241 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_403 VGND VPWR sky130_fd_sc_hd__decap_4
X_1126_ d_sram_out[11] _1126_/Q _1127_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_25_116 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_65_296 VGND VPWR sky130_fd_sc_hd__fill_2
X_1057_ _1044_/X _1018_/X _1056_/Y _1057_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_15_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_108 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0583__C _0583_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_119 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_193 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0880__A _0880_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_27 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_38 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0889__A1 _1174_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_187 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1217__CLK _1161_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_68 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_296 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_100 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_300 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_111 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_277 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1101__D _0594_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_144 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0940__D _0940_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0577__B1 _0518_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_355 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0965__A _0965_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_263 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_274 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0684__B _0676_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_222 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_2 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_266 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1057__A1 _1044_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_288 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0804__A1 _0799_/X VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_0_clk clk clkbuf_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_16
XFILLER_87_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_152 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0804__B2 _0801_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_202 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0568__B1 _0567_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0859__B _0946_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0626_ _0682_/C _0686_/C _0626_/C _0626_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_97_141 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_130 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1036__A _0988_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0557_ _0556_/X _0557_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0578__C _0574_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_358 VGND VPWR sky130_fd_sc_hd__decap_8
X_0488_ _1147_/Q _0488_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0875__A _0833_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_274 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0594__B _0594_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1109_ _1141_/Q _1109_/Q _1103_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_13_119 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_53_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0559__B1 _1128_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_257 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_227 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0769__B _1089_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_141 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_34 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0785__A _0663_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0731__B1 _0594_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_266 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_141 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0798__B1 _0797_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0679__B _0682_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_152 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_166 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0695__A _0695_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_255 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_277 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_258 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0789__B1 _0785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0580__D _0580_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0961__B1 _0946_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0589__B _0580_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0609_ _0723_/D _0594_/B _0609_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_37_48 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_159 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0499__B _1147_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_293 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_144 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_361 VGND VPWR sky130_fd_sc_hd__decap_12
X_0960_ _0988_/A _0955_/X _0988_/C _0960_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_32_258 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0681__C _0722_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1085__CLK _1114_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0891_ _0899_/A _0899_/B _0903_/C _0891_/D _0891_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_126_385 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1017__C _0978_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_111 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_133 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_214 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_300 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_2_0_clk clkbuf_2_3_0_clk/A clkbuf_3_5_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_48_69 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_188 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_83 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_171 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_199 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0676__C _0676_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1090_ _1090_/D _0776_/B _1127_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0973__A _0978_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0692__B _0558_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_228 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_0943_ _0836_/Y _0943_/B _0908_/C _1042_/D _0968_/A VGND VPWR sky130_fd_sc_hd__or4_4
X_0874_ _0872_/Y _0833_/A _0873_/X d_sram_in[7] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_114_300 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1028__B _1027_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1100__CLK _1116_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_250 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_272 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1044__A _0843_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0586__C _0587_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0883__A _0883_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_27 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_138 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_209 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_283 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_125 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_169 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1104__D _0675_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_117 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_331 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0943__D _1042_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0610__A2 _0583_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1123__CLK _1127_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0590_ _0682_/C _0628_/B _0509_/A _0578_/Y _0589_/Y _0591_/B VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__0968__A _0968_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_196 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0687__B _0690_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1211_ addr_w[13] _1042_/D _1174_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1142_ d_sram_out[27] _1142_/Q _1142_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1073_ _1022_/X _1070_/X _1071_/X w_mask[27] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__1014__D _1024_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_264 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_128 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_172 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_403 VGND VPWR sky130_fd_sc_hd__decap_4
X_0926_ _0920_/B _0926_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_134_406 VGND VPWR sky130_fd_sc_hd__fill_1
X_0857_ _1170_/Q _0857_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1039__A _0948_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0788_ _0554_/Y _0787_/X _0739_/D _0787_/X _0788_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_141 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0878__A _0835_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0597__B _0617_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_136 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_48 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_98 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1146__CLK _1221_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_264 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_297 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_312 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_183 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0711_ _0659_/A _0711_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_128_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_406 VGND VPWR sky130_fd_sc_hd__fill_1
X_0642_ _0587_/A _0643_/B _0587_/C _0540_/D _0642_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__1009__D _0987_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0573_ _0540_/D _0524_/X _1121_/Q _0587_/C _0573_/Y VGND VPWR sky130_fd_sc_hd__a22oi_4
XANTENNA__0698__A _0697_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0898__A2 _0877_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_188 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_177 VGND VPWR sky130_fd_sc_hd__decap_6
X_1125_ d_sram_out[10] _0720_/A _1103_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_65_275 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_139 VGND VPWR sky130_fd_sc_hd__fill_2
X_1056_ _1048_/B _1056_/B _1048_/C _1056_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__0583__D _0673_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1169__CLK _1187_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0880__B _1046_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_367 VGND VPWR sky130_fd_sc_hd__decap_12
X_0909_ _1171_/Q _0890_/X _0908_/X _0910_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_0_249 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0889__A2 _0877_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_312 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_101 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_236 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0577__B2 _0628_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_301 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_297 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0684__C _0677_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_80 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_234 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1057__A2 _1018_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0981__A _0981_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0804__A2 _1101_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_131 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0568__A1 _0560_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_74 VGND VPWR sky130_fd_sc_hd__decap_12
X_0625_ _0614_/Y _0528_/X _0603_/Y _0571_/X _0626_/C VGND VPWR sky130_fd_sc_hd__o22a_4
X_0556_ _0581_/A _0490_/A _0504_/A _0555_/Y _0556_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_97_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1036__B _1028_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0578__D _0578_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0487_ _1132_/Q _0487_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_264 VGND VPWR sky130_fd_sc_hd__fill_2
X_1108_ _0602_/D _1108_/Q _1124_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1039_ _0948_/X _1021_/B _1024_/C _1003_/Y _1039_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__1202__D addr_w[4] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0891__A _0899_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_153 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_107_236 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0559__B2 _0558_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_46 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_186 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0731__A1 _0750_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0731__B2 _0711_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0788__A2_N _0787_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1112__D _0678_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0798__A1 _1130_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_385 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0679__C _0544_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_164 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_289 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0789__B2 _1094_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0789__A1 _0779_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1207__CLK _1221_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_206 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0961__A1 _0942_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0589__C _0583_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0608_ _0542_/D _0524_/X _0608_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0886__A _0908_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0539_ _0725_/A _0681_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_58_304 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_123 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0499__C _0620_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_304 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1107__D _0543_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_82 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0681__D _0487_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0890_ _1046_/C _0890_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_138_180 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_226 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_248 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_209 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1017__D _1024_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_67_178 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0790__A1_N _0560_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_312 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0934__A1 _1192_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_178 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_126 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_215 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0870__B1 _0848_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_62 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_95 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_301 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0925__A1 _1185_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0676__D _0676_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0973__B _0982_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_398 VGND VPWR sky130_fd_sc_hd__decap_8
X_0942_ _0941_/X _0942_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_13_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_117 VGND VPWR sky130_fd_sc_hd__decap_12
X_0873_ _0872_/Y _0839_/A _0854_/Y _0873_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_62_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_240 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0586__D _1117_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_310 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_170 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1210__D addr_w[12] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_312 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_25 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_262 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_398 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1120__D d_sram_out[5] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_93 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1020__B1 _1019_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1210_ addr_w[12] _0940_/D _1142_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_77_240 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_104 VGND VPWR sky130_fd_sc_hd__fill_2
X_1141_ d_sram_out[26] _1141_/Q _1201_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_92_210 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0984__A _0843_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_126 VGND VPWR sky130_fd_sc_hd__decap_4
X_1072_ _1018_/X _1070_/X _1071_/X w_mask[26] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_92_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_243 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_159 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_354 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_2_1_0_clk clkbuf_1_0_0_clk/X clkbuf_3_3_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_0925_ _1185_/Q _0907_/X _0855_/X d_sram_in[19] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__0906__B1_N _0905_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0856_ _0851_/Y _0833_/X _0855_/X d_sram_in[3] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__1039__B _1021_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0787_ _0496_/A _0787_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1098__CLK _1127_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_304 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1055__A _0955_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0597__C _0597_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_251 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_28_148 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1205__D addr_w[7] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1078__B1 _1076_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_118 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_140 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_245 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1002__B1 _0996_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_178 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1115__D d_sram_out[0] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1069__B1 _1067_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0816__B1 _0722_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_192 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_162 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_335 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0710_ _0685_/X _0708_/Y _0709_/X _0710_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0979__A _0978_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0641_ _0697_/A _0700_/B _0702_/C _1117_/Q _0641_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0572_ _0571_/X _0587_/C VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0698__B _0700_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_346 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_221 VGND VPWR sky130_fd_sc_hd__fill_2
X_1124_ d_sram_out[9] _0673_/A _1124_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_65_254 VGND VPWR sky130_fd_sc_hd__fill_2
X_1055_ _0955_/A _0957_/X _0973_/C _0987_/D _1056_/B VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_80_224 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_246 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_140 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_162 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0807__B1 _0542_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_278 VGND VPWR sky130_fd_sc_hd__fill_2
X_0908_ _0903_/A _0903_/B _0908_/C _1179_/Q _0908_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_134_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_0839_ _0839_/A _0839_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_56_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_243 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_112_32 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_213 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1113__CLK _1114_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_102 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_324 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_135 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_51 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0799__A _0661_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_232 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0684__D _0684_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_4 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_143 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_30_154 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_80 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0568__A2 _0562_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_86 VGND VPWR sky130_fd_sc_hd__decap_12
X_0624_ _0580_/B _0686_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0502__A _0502_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_110 VGND VPWR sky130_fd_sc_hd__decap_8
X_0555_ _1153_/Q _0555_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0486_ reb csb _1165_/D VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_38_210 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1136__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_276 VGND VPWR sky130_fd_sc_hd__decap_12
X_1107_ _0543_/A _1107_/Q _1103_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_53_235 VGND VPWR sky130_fd_sc_hd__decap_3
X_1038_ _0945_/A _1035_/X _1037_/X w_mask[14] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0891__B _0899_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_98 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0731__A2 _0718_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_202 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_279 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0798__A2 _0750_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0679__D _0679_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1159__CLK _1226_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_176 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0992__A _0991_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_330 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_92_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0789__A2 _0788_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0961__A2 _0945_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0589__D _0588_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0607_ _1138_/Q _0530_/A _0688_/A VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_112_240 VGND VPWR sky130_fd_sc_hd__decap_12
X_0538_ _0581_/A _0725_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_85_157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_179 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1213__D addr_r[1] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_310 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_105 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1123__D d_sram_out[8] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_398 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0987__A _0955_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_371 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_105 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_330 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_149 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_363 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_324 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1208__D addr_w[10] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0897__A _0847_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0934__A2 _0932_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_104_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_265 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_287 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_138 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_171 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0870__A1 _0869_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_108_398 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0925__A2 _0907_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_219 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0600__A _0583_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1118__D d_sram_out[3] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_282 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_93 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0973__C _0973_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_300 VGND VPWR sky130_fd_sc_hd__decap_12
X_0941_ _0940_/X _0941_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_13_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_0872_ _1173_/Q _0872_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_70_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_324 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0510__A _1151_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_296 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_285 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_322 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_302 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_117_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_37 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_241 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_115_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_110 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1020__A1 _0998_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1140_ d_sram_out[25] _0602_/D _1124_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_49_92 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_222 VGND VPWR sky130_fd_sc_hd__fill_1
X_1071_ _0985_/A _1032_/X _1066_/Y _1071_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_80_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_160 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_185 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0505__A _0505_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0924_ _1184_/Q _0907_/X _0849_/X d_sram_in[18] VGND VPWR sky130_fd_sc_hd__a21bo_4
X_0855_ _0851_/Y _0839_/X _0854_/Y _0855_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__1039__C _1024_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0786_ _0779_/X _0784_/X _0785_/X _1093_/Q d_fabric_out[10] VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_114_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_316 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1055__B _0957_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0770__B1 _0769_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_285 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1078__A1 _1032_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_300 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1221__D addr_r[9] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_110 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1002__A1 _0998_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0761__B1 _0759_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_230 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_403 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1192__CLK _1114_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_406 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1069__A1 _1015_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0816__A1 _0813_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1131__D d_sram_out[16] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0816__B2 _0815_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_202 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0640_ _0580_/B _0700_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_0571_ _0571_/A _0571_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0698__C _0594_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_135 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0995__A _0995_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0752__B1 _0719_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_1123_ d_sram_out[8] _0502_/A _1127_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1054_ _0979_/X _1043_/X _1052_/X w_mask[19] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_18_182 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0807__A1 _0806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_152 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0807__B2 _0801_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_80_269 VGND VPWR sky130_fd_sc_hd__decap_3
X_0907_ _0920_/B _0907_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_119_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_227 VGND VPWR sky130_fd_sc_hd__decap_12
X_0838_ _0835_/X _0838_/B _0839_/A VGND VPWR sky130_fd_sc_hd__and2_4
X_0769_ _0733_/A _1089_/Q _0769_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1066__A _1066_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_303 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_218 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_403 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1216__D addr_r[4] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_211 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_71_236 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_141 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_103 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_293 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0734__B1 _0733_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_336 VGND VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_2_0_0_clk clkbuf_1_0_0_clk/X clkbuf_3_1_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__1126__D d_sram_out[11] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_62_203 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_93 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_5 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_258 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_15_163 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1088__CLK _1114_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_98 VGND VPWR sky130_fd_sc_hd__decap_12
X_0623_ _1115_/Q _0620_/X _0622_/Y _0623_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_131_208 VGND VPWR sky130_fd_sc_hd__decap_12
X_0554_ _1126_/Q _0554_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_97_199 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_19 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_288 VGND VPWR sky130_fd_sc_hd__decap_12
X_1106_ _1138_/Q _1106_/Q _1127_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_53_214 VGND VPWR sky130_fd_sc_hd__fill_2
X_1037_ _0985_/X _1001_/X _1036_/Y _1037_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_53_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_269 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0891__C _0903_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_188 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_216 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_400 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_115_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_200 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0731__A3 _0730_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_309 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_247 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_280 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_385 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0603__A _0532_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_398 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0707__B1 _0550_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_306 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_353 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_280 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_330 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0513__A _0505_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1103__CLK _1103_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0606_ _0583_/A _0724_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_112_252 VGND VPWR sky130_fd_sc_hd__decap_12
X_0537_ _0526_/X _0532_/X _0676_/C _0546_/C VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_66_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_331 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_300 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_135_322 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_230 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_263 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_117 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_320 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_83 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_300 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1126__CLK _1127_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_239 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0987__B _0957_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_383 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_180 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0508__A _0508_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_23_217 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_171 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0897__B _0896_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_272 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1074__A _1009_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_136 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1224__D addr_r[12] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_239 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0870__A2 _0839_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1149__CLK _1174_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_132 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_110 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_158 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1134__D d_sram_out[19] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_128 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0973__D _0991_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_93 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_194 VGND VPWR sky130_fd_sc_hd__fill_1
X_0940_ _0940_/A _0956_/A _0940_/C _0940_/D _0940_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_9_232 VGND VPWR sky130_fd_sc_hd__decap_12
X_0871_ _0869_/Y _0833_/X _0870_/X d_sram_in[6] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_126_141 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0998__A _0968_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_220 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_180 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0660__B1_N _0659_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_334 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1219__D addr_r[7] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0701__A _0724_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_49 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_220 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_6_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_152 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1129__D d_sram_out[14] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0611__A _0724_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1020__A2 _1018_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_220 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_297 VGND VPWR sky130_fd_sc_hd__fill_2
X_1070_ _1043_/A _1070_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_33_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0505__B _0505_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0923_ _1183_/Q _0876_/X _0844_/X _0922_/Y d_sram_in[17] VGND VPWR sky130_fd_sc_hd__a211o_4
X_0854_ _0854_/A _0854_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1039__D _1003_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0785_ _0663_/A _0785_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0521__A _0512_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_166 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0770__A1 _0762_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_328 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1055__C _0973_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_297 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_223 VGND VPWR sky130_fd_sc_hd__fill_2
X_1199_ addr_w[1] baseaddr_w_sync[1] _1226_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1078__A2 _1070_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_278 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_312 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_197 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_203 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_236 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1002__A2 _1001_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0761__A1 _0675_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_199 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0761__B2 _0760_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_253 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_234 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_256 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1069__A2 _1059_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_289 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0816__A2 _1109_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_62 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0606__A _0583_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0570_ _0523_/A _0503_/A _0571_/A VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__0698__D _0677_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0752__A1 _0532_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_201 VGND VPWR sky130_fd_sc_hd__fill_2
X_1122_ d_sram_out[7] _0580_/D _1127_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_65_245 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_76_80 VGND VPWR sky130_fd_sc_hd__decap_12
X_1053_ _0974_/X _1043_/X _1052_/X w_mask[18] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_80_215 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_131 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0807__A2 _1103_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_197 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0516__A _0504_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0906_ _1178_/Q _0877_/X _0905_/Y d_sram_in[12] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_119_269 VGND VPWR sky130_fd_sc_hd__decap_6
X_0837_ _0836_/Y _0943_/B _0835_/C _0838_/B VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_134_239 VGND VPWR sky130_fd_sc_hd__decap_12
X_0768_ _0723_/D _0750_/X _0766_/X _0767_/X _1089_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__1066__B _1066_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_337 VGND VPWR sky130_fd_sc_hd__decap_12
X_0699_ _0699_/A _0699_/B _0697_/X _0698_/X _0699_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__1082__A csb VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_267 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_104 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_164 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_126 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_337 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_159 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_115_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_315 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0734__A1 _0663_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1142__D d_sram_out[27] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_226 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_6 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_93 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_239 VGND VPWR sky130_fd_sc_hd__decap_12
X_0622_ _0620_/A _0488_/Y _0620_/C _0622_/Y VGND VPWR sky130_fd_sc_hd__nand3_4
X_0553_ _0524_/X _0628_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_1105_ _0723_/D _1105_/Q _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1036_ _0988_/C _1028_/X _1036_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__0891__D _0891_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_178 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_156 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1182__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1227__D conf[1] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_29_212 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_397 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_106_272 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1137__D d_sram_out[22] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0707__A1 _1116_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_137 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_57_71 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_226 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_129_342 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_3 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_171 VGND VPWR sky130_fd_sc_hd__decap_12
X_0605_ _0603_/Y _0562_/X _1142_/Q _0639_/B _0605_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_0536_ _0725_/C _0676_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_112_264 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_343 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_365 VGND VPWR sky130_fd_sc_hd__fill_1
X_1019_ _0985_/X _0992_/X _1011_/Y _1019_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0704__A _0690_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_334 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0937__A1 _1195_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0919__B1_N _0918_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_297 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_126 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0873__B1 _0854_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_74 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_72_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_403 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0625__B1 _0603_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_51 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0614__A _1113_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_312 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0928__A1 _1187_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1050__B1 _1049_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0987__C _0991_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_159 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_395 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_343 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0524__A _0581_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1041__B1 _1037_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0919__A1 _1181_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1220__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1074__B _0957_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0519_ _0518_/X _0682_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_104_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0855__B1 _0854_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_251 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_295 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0609__A _0723_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_151 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1150__D _1158_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_324 VGND VPWR sky130_fd_sc_hd__decap_12
X_0870_ _0869_/Y _0839_/X _0848_/Y _0870_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_70_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1023__B1 _1019_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0519__A _0518_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_170 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_63_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_346 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_379 VGND VPWR sky130_fd_sc_hd__decap_12
X_0999_ _0954_/A _1024_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0701__B _0701_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1116__CLK _1116_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_120 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_123 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0611__B _0617_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_111_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1145__D d_sram_out[30] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_232 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_268 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0819__B1 _0679_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_140 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_379 VGND VPWR sky130_fd_sc_hd__decap_12
X_0922_ _0922_/A _0876_/X _0922_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_0853_ _0827_/A _0946_/A _0844_/X _0852_/X _0854_/A VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_60_3 VGND VPWR sky130_fd_sc_hd__decap_3
X_0784_ _0722_/D _0711_/X _0783_/X _0784_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0521__B _0740_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_178 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1055__D _0987_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_210 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0770__A2 _1089_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1139__CLK _1142_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_202 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_257 VGND VPWR sky130_fd_sc_hd__fill_2
X_1198_ addr_w[0] baseaddr_w_sync[0] _1175_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_91_290 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_184 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_105_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0746__C1 _0745_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0761__A2 _0750_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_351 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_246 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_268 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_290 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_154 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_187 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_51 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_51_62 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0622__A _0620_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0752__A2 _0751_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1121_ d_sram_out[6] _1121_/Q _1201_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1052_ _1044_/X _1015_/X _1048_/Y _1052_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_18_162 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_110 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_290 VGND VPWR sky130_fd_sc_hd__fill_2
X_0905_ _0861_/A _0904_/X _0905_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__0532__A _0532_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_207 VGND VPWR sky130_fd_sc_hd__decap_6
X_0836_ _0835_/A _0836_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_127_281 VGND VPWR sky130_fd_sc_hd__decap_12
X_0767_ _1121_/Q _0659_/A _0709_/X _0767_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__1066__C _1048_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_209 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_349 VGND VPWR sky130_fd_sc_hd__decap_12
X_0698_ _0697_/A _0700_/B _0594_/B _0677_/D _0698_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_102_159 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1082__B web VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_205 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_249 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_105 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_176 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_154 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_127 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0967__C1 _0960_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_98 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0734__A2 _1085_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_308 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_192 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_238 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_7 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0617__A _0617_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_290 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_135 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_30_179 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_375 VGND VPWR sky130_fd_sc_hd__fill_2
X_0621_ _0591_/X _0619_/X _0620_/X _0621_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
X_0552_ _1154_/Q _0552_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_97_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_319 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_235 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_246 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_257 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_268 VGND VPWR sky130_fd_sc_hd__decap_6
X_1104_ _0675_/D _1104_/Q _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_53_227 VGND VPWR sky130_fd_sc_hd__fill_2
X_1035_ _1034_/X _1035_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0527__A _0581_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_290 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_21_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_293 VGND VPWR sky130_fd_sc_hd__fill_1
X_0819_ _0813_/X _1112_/Q _0679_/D _0815_/X d_fabric_out[29] VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_130_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_371 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_308 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_319 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_224 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_312 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0707__A2 _0622_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_121_232 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_105 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1153__D _1161_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_83 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_94 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_238 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_249 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_354 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0604_ _0557_/X _0639_/B VGND VPWR sky130_fd_sc_hd__inv_8
X_0535_ _0700_/A _0725_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_112_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_308 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0615__A2_N _0576_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_385 VGND VPWR sky130_fd_sc_hd__decap_12
X_1018_ _1018_/A _1018_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_34_260 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_219 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0704__B _0704_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0937__A2 _0932_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_346 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_56 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0720__A _0720_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_210 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_330 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_363 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0873__A1 _0872_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_86 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0625__A1 _0614_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0625__B2 _0571_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_74 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_324 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0928__A2 _0926_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1050__A1 _0941_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_142 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1148__D _1156_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0630__A _0594_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0987__D _0987_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1172__CLK _1114_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_141 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_63_355 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_241 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0524__B _0544_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_184 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1041__A1 _0945_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0919__A2 _0907_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0540__A _0681_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1074__C _0973_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0518_ _0587_/A _0518_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_98_285 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_279 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0855__A1 _0851_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_196 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_11 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0791__B1 _0785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_123 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1195__CLK _1185_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_178 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_30 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_127 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_406 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0609__B _0594_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_160 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_245 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1023__A1 _0998_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0782__B1 _0762_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_141 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0535__A _0700_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_117_110 VGND VPWR sky130_fd_sc_hd__decap_12
X_0998_ _0968_/A _0998_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0701__C _0628_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0773__B1 _0719_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_266 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_196 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_132 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_123_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_198 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0611__C _0610_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0764__B1 _0763_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_277 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_247 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_225 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0819__A1 _0813_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1161__D _1224_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0819__B2 _0815_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1210__CLK _1142_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_100 VGND VPWR sky130_fd_sc_hd__fill_2
X_0921_ _0880_/A _0833_/A _0920_/X d_sram_in[16] VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_41_391 VGND VPWR sky130_fd_sc_hd__decap_12
X_0852_ _0851_/A _0852_/B _0852_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0783_ _0720_/A _0750_/A _0783_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_53_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_281 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0521__C _0677_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_141 VGND VPWR sky130_fd_sc_hd__fill_1
X_1197_ d_fabric_in[31] _1197_/Q _1114_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_101_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_144 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_135 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0746__B1 _0651_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_363 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_19_98 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_317 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_86 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_227 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0903__A _0903_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_85 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0622__B _0488_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_306 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1156__D _0841_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_406 VGND VPWR sky130_fd_sc_hd__fill_1
X_1120_ d_sram_out[5] _0677_/D _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_65_225 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_93 VGND VPWR sky130_fd_sc_hd__decap_12
X_1051_ _0966_/A _1043_/X _1049_/X w_mask[17] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_80_206 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_306 VGND VPWR sky130_fd_sc_hd__decap_12
X_0904_ _1170_/Q _0890_/X _0903_/X _0904_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0813__A _0661_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0976__B1 _0975_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0835_ _0835_/A _0883_/A _0835_/C _0835_/X VGND VPWR sky130_fd_sc_hd__or3_4
XANTENNA__1106__CLK _1127_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0532__B _0656_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_293 VGND VPWR sky130_fd_sc_hd__decap_12
X_0766_ _0609_/X _0765_/X _0719_/X _0766_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_0697_ _0697_/A _0700_/B _0580_/C _0580_/D _0697_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_102_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_203 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0900__B1 _0899_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_247 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_58 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_36 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0723__A _0740_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0967__B1 _0946_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_339 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_236 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_8 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0617__B _0616_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_155 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_188 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1129__CLK _1124_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0633__A _0594_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0958__B1 _0833_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_282 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_398 VGND VPWR sky130_fd_sc_hd__decap_8
X_0620_ _0620_/A _1147_/Q _0620_/C _0620_/X VGND VPWR sky130_fd_sc_hd__and3_4
X_0551_ _0509_/X _0546_/Y _0550_/X _0551_/Y VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_97_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_1103_ _0542_/D _1103_/Q _1103_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0808__A _0776_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1034_ _0948_/X _0956_/X _1024_/C _1003_/Y _1034_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0527__B _0490_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_261 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_114 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_147 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0543__A _0543_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_8_0_clk_A clkbuf_4_8_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0818_ _0813_/X _1111_/Q _0532_/A _0815_/X d_fabric_out[28] VGND VPWR sky130_fd_sc_hd__o22a_4
X_0749_ _0663_/X _0747_/X _0748_/X d_fabric_out[3] VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_130_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_320 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_269 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0718__A _0718_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_280 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_138_311 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_32 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_366 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_120_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_191 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_252 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_51 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_323 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_90_312 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0628__A _0580_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_261 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_184 VGND VPWR sky130_fd_sc_hd__decap_12
X_0603_ _0532_/A _0603_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_98_80 VGND VPWR sky130_fd_sc_hd__decap_12
X_0534_ _0580_/A _0700_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_100_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_128 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0538__A _0581_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_301 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_239 VGND VPWR sky130_fd_sc_hd__decap_6
X_1017_ _0978_/A _0982_/B _0978_/C _1024_/D _1018_/A VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_81_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_272 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0704__C _0699_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_118_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0720__B _0506_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0873__A2 _0839_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_209 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0625__A2 _0528_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1050__A2 _1043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_209 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1164__D web VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_172 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_186 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1041__A2 _1040_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_196 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0540__B _0682_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_264 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1074__D _0987_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0517_ _0585_/A _0587_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_100_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_269 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0855__A2 _0839_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_183 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_142 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_175 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_242 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_23 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_5_0_clk_A clkbuf_3_5_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_306 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0791__A1 _0713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_188 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0791__B2 _1095_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_257 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1159__D _1222_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0641__A _0697_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1023__A2 _1022_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_166 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0782__A1 _0779_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0782__B2 _1092_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_245 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_289 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_197 VGND VPWR sky130_fd_sc_hd__fill_2
X_0997_ _0968_/X _0995_/X _0996_/X w_mask[6] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_105_306 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0701__D _1132_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0773__A1 _0771_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0726__A _0544_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1162__CLK _1185_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_144 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0764__A1 _0762_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_361 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_96 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_51 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0819__A2 _1112_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0636__A _0676_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_145 VGND VPWR sky130_fd_sc_hd__fill_2
X_0920_ _1182_/Q _0920_/B _0920_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_60_189 VGND VPWR sky130_fd_sc_hd__fill_2
X_0851_ _0851_/A _0851_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0782_ _0779_/X _1092_/D _0762_/X _1092_/Q d_fabric_out[9] VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__0521__D _1127_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_331 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_109 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_267 VGND VPWR sky130_fd_sc_hd__decap_8
X_1196_ d_fabric_in[30] _1196_/Q _1116_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_51_101 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0546__A _0509_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_123 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1185__CLK _1185_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_219 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0746__A1 _1118_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_223 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_120 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_197 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_145 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_98 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_329 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0903__B _0903_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_97 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_2_2_0_clk_A clkbuf_2_3_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0622__C _0620_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0902__B1_N _0901_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_263 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1172__D d_fabric_in[6] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_237 VGND VPWR sky130_fd_sc_hd__decap_4
X_1050_ _0941_/X _1043_/X _1049_/X w_mask[16] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_80_229 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_123 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_93 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_318 VGND VPWR sky130_fd_sc_hd__decap_12
X_0903_ _0903_/A _0903_/B _0903_/C _1178_/Q _0903_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0976__A1 _0968_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0834_ _0943_/B _0883_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_0765_ _0614_/Y _0528_/X _0668_/X _0724_/D _0765_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_0696_ _0518_/X _0701_/B _0702_/C _0695_/X _0699_/B VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_102_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_4_0_clk_A clkbuf_3_2_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0900__A1 _0851_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_80 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_107 VGND VPWR sky130_fd_sc_hd__decap_3
X_1179_ d_fabric_in[13] _1179_/Q _1116_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_118 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0723__B _0740_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0967__A1 _0945_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1200__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_340 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_172 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_259 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_207 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_123 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_9 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_167 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0914__A _0847_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0633__B _0702_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1080__B1 _1079_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0958__A1 _0883_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1167__D d_fabric_in[1] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_294 VGND VPWR sky130_fd_sc_hd__decap_8
X_0550_ _0549_/Y _0550_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_93_310 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_373 VGND VPWR sky130_fd_sc_hd__decap_12
X_1102_ _0695_/A _1102_/Q _1116_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1033_ _0945_/A _1032_/X _1029_/Y w_mask[13] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_46_270 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_273 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0824__A _0841_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1071__B1 _1066_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0817_ _0813_/X _1110_/Q _0739_/D _0815_/X d_fabric_out[27] VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__1223__CLK _1201_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_220 VGND VPWR sky130_fd_sc_hd__decap_12
X_0748_ _0733_/A _1086_/Q _0748_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_107_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_59 VGND VPWR sky130_fd_sc_hd__fill_2
X_0679_ _0722_/A _0682_/B _0544_/C _0679_/D _0683_/B VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_96_192 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_398 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0718__B _0716_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_292 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_323 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1062__B1 _1061_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_55 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_264 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_286 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_129 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_218 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0628__B _0628_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_357 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_284 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0644__A _0580_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_367 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1053__B1 _1052_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0800__B1 _0799_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_196 VGND VPWR sky130_fd_sc_hd__decap_12
X_0602_ _0697_/A _0701_/B _0702_/C _0602_/D _0612_/B VGND VPWR sky130_fd_sc_hd__and4_4
X_0533_ _0505_/B _0580_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_3_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0867__B1 _0866_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_140 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_184 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_335 VGND VPWR sky130_fd_sc_hd__fill_2
X_1016_ _0998_/X _1015_/X _1012_/X w_mask[9] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_81_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0554__A _1126_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0704__D _0704_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_245 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_134_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0729__A _0550_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1119__CLK _1103_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_1_0_clk_A clkbuf_3_1_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_343 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_218 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_184 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_243 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_265 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_12_0_clk_A clkbuf_3_6_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_80 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0639__A _0723_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_129 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0849__B1 _0848_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_398 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1180__D d_fabric_in[14] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_379 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0540__C _0682_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_243 VGND VPWR sky130_fd_sc_hd__fill_2
X_0516_ _0504_/A _0585_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_100_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_204 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_118 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0549__A _0548_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_237 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_324 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1090__D _1090_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_110 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_120_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_19 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_254 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_35 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0791__A2 _0790_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_107 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1091__CLK _1127_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_143 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0922__A _0922_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_269 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0641__B _0700_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_178 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0782__A2 _1092_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1175__D d_fabric_in[9] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_268 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_184 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0832__A _0831_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0996_ _0985_/X _0979_/X _0988_/Y _0996_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_117_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_329 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1085__D _1085_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0773__A2 _0772_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_26 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_121 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0726__B _0513_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_202 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0742__A _0725_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_77 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_178 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0764__A2 _1088_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_86 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_290 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0636__B _0686_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0652__A _0681_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0850_ _0830_/Y _0833_/X _0849_/X d_sram_in[2] VGND VPWR sky130_fd_sc_hd__o21ai_4
X_0781_ _0674_/A _0496_/X _0676_/D _0496_/X _1092_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_39_3 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_257 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_398 VGND VPWR sky130_fd_sc_hd__decap_8
X_1195_ d_fabric_in[29] _1195_/Q _1185_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0827__A _0827_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0546__B _0546_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_157 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_179 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0562__A _0561_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_0_0_clk_A clkbuf_4_0_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0979_ _0978_/X _0979_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0746__A2 _0548_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_110 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0737__A _1126_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_124 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0903__C _0903_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_190 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_136_251 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_116_80 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0647__A _0638_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_179 VGND VPWR sky130_fd_sc_hd__fill_2
X_0902_ _1177_/Q _0877_/X _0901_/Y d_sram_in[11] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__0976__A2 _0974_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0833_ _0833_/A _0833_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0764_ _0762_/X _1088_/D _0763_/X d_fabric_out[5] VGND VPWR sky130_fd_sc_hd__a21o_4
X_0695_ _0695_/A _0695_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_88_308 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_330 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_385 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0900__A2 _0890_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0557__A _0556_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1152__CLK _1201_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1178_ d_fabric_in[12] _1178_/Q _1187_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XPHY_108 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0723__C _0722_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0967__A2 _0966_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_319 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_352 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_184 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_135 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_102_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_105 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_274 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0914__B _0913_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_149 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1080__A1 _1035_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_15 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0958__A2 _0885_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_7_367 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_124_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1183__D d_fabric_in[17] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1175__CLK _1175_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_322 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_385 VGND VPWR sky130_fd_sc_hd__decap_12
X_1101_ _0594_/A _1101_/Q _1116_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0894__A1 _0891_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_1032_ _1031_/X _1032_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_61_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_285 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_296 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_190 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1001__A _1000_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1071__A1 _0985_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0816_ _0813_/X _1109_/Q _0722_/D _0815_/X d_fabric_out[26] VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__0840__A _0840_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_232 VGND VPWR sky130_fd_sc_hd__decap_12
X_0747_ _0750_/A _0736_/X _0746_/X _0695_/X _0496_/A _0747_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_130_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_149 VGND VPWR sky130_fd_sc_hd__fill_2
X_0678_ _0678_/A _0679_/D VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1093__D _0784_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_238 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0718__C _0501_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_241 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_335 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1062__A1 _0995_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_67 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0750__A _0750_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_232 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_243 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1198__CLK _1175_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_235 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_298 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_276 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0573__B1 _1121_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_268 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_75 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_369 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_403 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0644__B _0643_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1053__A1 _0974_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1178__D d_fabric_in[12] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_379 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0800__B2 _1098_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0800__A1 _0713_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0601_ _0583_/C _0702_/C VGND VPWR sky130_fd_sc_hd__buf_1
X_0532_ _0532_/A _0656_/B _0532_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_112_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0867__A1 _0864_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_347 VGND VPWR sky130_fd_sc_hd__decap_12
X_1015_ _1014_/X _1015_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0835__A _0835_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1088__D _1088_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_80 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0570__A _0523_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_213 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_202 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0729__B _0720_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_355 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_303 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_78 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0745__A _0550_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_380 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_187 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0794__B1 _0785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_300 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_119 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0639__B _0639_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0849__A1 _0830_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_80 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1213__CLK _1161_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_336 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_196 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0655__A _1099_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_110 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0540__D _0540_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_222 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0537__B1 _0676_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_406 VGND VPWR sky130_fd_sc_hd__fill_1
X_0515_ _0682_/B _0740_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_39_300 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0565__A _0585_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_120_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_166 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_266 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_47 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_255 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_299 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0922__B _0876_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0641__C _0702_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0767__B1 _0709_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_190 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_203 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_122_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_236 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1191__D d_fabric_in[25] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_174 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_166 VGND VPWR sky130_fd_sc_hd__fill_2
X_0995_ _0995_/A _0995_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1109__CLK _1103_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_135 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0758__B1 _0687_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_38 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_174 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_131_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0726__C _1113_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_361 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0997__B1 _0996_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0742__B _0544_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0749__B1 _0748_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_89 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_171 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0921__B1 _0920_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_144 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_306 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0636__C _0635_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_74 VGND VPWR sky130_fd_sc_hd__decap_12
X_0780_ _0779_/X _1091_/D _0762_/X _1091_/Q d_fabric_out[8] VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__1186__D d_fabric_in[20] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_206 VGND VPWR sky130_fd_sc_hd__fill_2
X_1194_ d_fabric_in[28] _1194_/Q _1187_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_36_133 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1004__A _1003_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0546__C _0546_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_199 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0843__A _0843_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_361 VGND VPWR sky130_fd_sc_hd__decap_12
X_0978_ _0978_/A _0991_/B _0978_/C _0991_/D _0978_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__1096__D _0793_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_269 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0737__B _0506_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_291 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_155 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_261 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_188 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_294 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_158 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0903__D _1178_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_241 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_217 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0647__B _0639_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_114 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_33_136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_283 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_294 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_158 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0663__A _0663_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_208 VGND VPWR sky130_fd_sc_hd__decap_12
X_0901_ _0854_/A _0901_/B _0901_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_0832_ _0831_/X _0833_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_115_403 VGND VPWR sky130_fd_sc_hd__decap_4
X_0763_ _0733_/A _0763_/B _0763_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0694_ _0700_/A _0700_/B _0583_/C _1126_/Q _0699_/A VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_51_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_141 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0838__A _0835_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_239 VGND VPWR sky130_fd_sc_hd__fill_2
X_1177_ d_fabric_in[11] _1177_/Q _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_71_209 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_109 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0723__D _0723_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_200 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_222 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_364 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0748__A _0733_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_99 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_294 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_147 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_139 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1080__A2 _1070_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_27 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_112_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_51 VGND VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_9_0_clk clkbuf_4_8_0_clk/A _1174_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_87_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_206 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_228 VGND VPWR sky130_fd_sc_hd__fill_2
X_1100_ _1132_/Q _1100_/Q _1116_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_93_334 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_239 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0894__A2 _0877_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_367 VGND VPWR sky130_fd_sc_hd__decap_12
X_1031_ _0981_/A _1021_/B _1024_/C _1003_/Y _1031_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_46_283 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_294 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1071__A2 _1032_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0815_ out_reg _0815_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0746_ _1118_/Q _0548_/X _0651_/Y _0745_/X _0746_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_107_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_117 VGND VPWR sky130_fd_sc_hd__decap_12
X_0677_ _0716_/A _0677_/B _0677_/C _0677_/D _0677_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_69_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_172 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_375 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0718__D _0717_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_264 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1062__A2 _1059_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_79 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0573__B2 _0587_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0573__A1 _0540_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_172 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_150 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_301 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_87 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_323 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_242 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0644__C _0585_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_86 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0941__A _0940_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1053__A2 _1043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_7_110 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0800__A2 _0798_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1142__CLK _1142_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0600_ _0583_/A _0697_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1194__D d_fabric_in[28] VGND VPWR sky130_fd_sc_hd__diode_2
X_0531_ _0580_/C _0656_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_66_312 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0867__A2 _0839_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_3 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_175 VGND VPWR sky130_fd_sc_hd__fill_2
X_1014_ _0991_/A _1021_/B _0978_/C _1024_/D _1014_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0835__B _0883_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_359 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0851__A _0851_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_306 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0570__B _0503_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_118_27 VGND VPWR sky130_fd_sc_hd__decap_4
X_0729_ _0550_/X _0720_/X _0728_/X _0729_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_134_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0729__C _0728_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_220 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0745__B _0745_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_253 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_201 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_56 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_392 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1165__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_199 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0794__B2 _1096_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0794__A1 _0713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_20 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_385 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0849__A2 _0839_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_153 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0655__B _0771_/B VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_270 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1189__D d_fabric_in[23] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_245 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_306 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0537__A1 _0526_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0514_ _0513_/X _0682_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1007__A _0981_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0915__B1_N _0914_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_186 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0846__A _0846_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1188__CLK _1201_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1099__D _1099_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0581__A _0581_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_201 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_245 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_278 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_12 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_66 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_245 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0491__A _0544_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_21 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0641__D _1117_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0767__A1 _1121_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_74 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_182 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_123 VGND VPWR sky130_fd_sc_hd__fill_1
X_0994_ _0948_/X _0956_/X _0954_/A _0940_/D _0995_/A VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0758__A1 _0668_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_342 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0930__A1 _1189_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_237 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_215 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_142 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0576__A _0587_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_292 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_307 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0726__D _0725_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0997__A1 _0968_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0742__C _0725_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0749__A1 _0663_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_68 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1203__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_11 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_66 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0921__A1 _0880_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_218 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_270 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0486__A reb VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_123 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0685__B1 _0550_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_104 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_98 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_8 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_215 VGND VPWR sky130_fd_sc_hd__fill_2
X_1193_ d_fabric_in[27] _1193_/Q _1221_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_36_145 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0546__D _0545_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1226__CLK _1226_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0977_ _0940_/C _0978_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_10_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_126_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_301 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_367 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_240 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_318 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_67 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_89 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_104_172 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0647__C _0641_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_145 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0658__B1 _0651_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0944__A _0968_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0900_ _0851_/A _0890_/X _0899_/X _0901_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_14_373 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_90 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1197__D d_fabric_in[31] VGND VPWR sky130_fd_sc_hd__diode_2
X_0831_ _1226_/Q _0841_/B _0835_/C _0831_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_127_220 VGND VPWR sky130_fd_sc_hd__decap_12
X_0762_ _0663_/A _0762_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0693_ _0676_/D _0627_/Y _0692_/X _0704_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_44_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_398 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0838__B _0838_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_207 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1015__A _1014_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0649__B1 _0648_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1176_ d_fabric_in[10] _0895_/D _1185_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0854__A _0854_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_262 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0821__B1 _1146_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_137_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_137_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_234 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_192 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0748__B _1086_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_56 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_240 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_159 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_265 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_276 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_354 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0812__B1 _0544_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_231 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_275 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_267 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_332 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_346 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_379 VGND VPWR sky130_fd_sc_hd__decap_12
X_1030_ _0945_/A _1025_/X _1029_/Y w_mask[12] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_46_262 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0674__A _0674_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0803__B1 _0487_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0814_ _0813_/X _1108_/Q _0676_/D _0808_/X d_fabric_out[25] VGND VPWR sky130_fd_sc_hd__o22a_4
X_0745_ _0550_/X _0745_/B _0744_/X _0745_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_115_245 VGND VPWR sky130_fd_sc_hd__decap_12
X_0676_ _0512_/X _0492_/C _0676_/C _0676_/D _0676_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_130_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_387 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_324 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0781__A2_N _0496_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_37_240 VGND VPWR sky130_fd_sc_hd__decap_4
X_1228_ conf[2] _0840_/A _1174_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_16_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0584__A _0505_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_210 VGND VPWR sky130_fd_sc_hd__fill_2
X_1159_ _1222_/Q _1159_/Q _1226_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1047__B1 _0958_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_304 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_162 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_106_256 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0573__A2 _0524_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_129 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1094__CLK _1142_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_66 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_335 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0730__C1 _0729_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_251 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0494__A _0493_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_349 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_265 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_98 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1038__B1 _1037_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0644__D _0720_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_80 VGND VPWR sky130_fd_sc_hd__decap_12
X_0530_ _0530_/A _0580_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0669__A _0740_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_198 VGND VPWR sky130_fd_sc_hd__fill_2
X_1013_ _0998_/X _1006_/X _1012_/X w_mask[8] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0835__C _0835_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_93 VGND VPWR sky130_fd_sc_hd__decap_12
X_0728_ _0721_/X _0728_/B _0723_/X _0728_/D _0728_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0579__A _0580_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0659_ _0659_/A _0658_/Y _0659_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_134_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_259 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_232 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0745__C _0744_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_265 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_224 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_8_0_clk clkbuf_4_8_0_clk/A _1114_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_43_79 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_156 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0794__A2 _0793_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0489__A _0503_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_270 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_397 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0952__A _0955_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_213 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_260 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_257 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_271 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_123 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_117_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0537__A2 _0532_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0513_ _0505_/A _0513_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_98_268 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_104_19 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0846__B _0852_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_146 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0581__B _0503_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_235 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_128 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_131_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_24 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_38_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_56 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1132__CLK _1116_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_13_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_290 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0767__A2 _0659_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_97 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_216 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0947__A _0940_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_179 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0682__A _0722_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0993_ _0968_/X _0992_/X _0989_/X w_mask[5] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_74_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0758__A2 _1128_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_354 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1018__A _1018_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0930__A2 _0926_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0857__A _1170_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1155__CLK _1174_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_290 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0576__B _0585_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_319 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0592__A _0579_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0997__A2 _0995_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_227 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0742__D _0695_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0749__A2 _0747_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_23 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_398 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0921__A2 _0833_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0486__B csb VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0685__A1 _0674_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_7 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1178__CLK _1187_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0929__B1_N _0870_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_335 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0677__A _0716_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1192_ d_fabric_in[26] _1192_/Q _1114_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_83_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_113 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_271 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_293 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_385 VGND VPWR sky130_fd_sc_hd__decap_12
X_0976_ _0968_/X _0974_/X _0975_/Y w_mask[2] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_99_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0587__A _0587_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_238 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_249 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_271 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_149 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_57 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_195 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0497__A _0497_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_76 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0647__D _0646_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0658__A1 _0501_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0658__B2 _0657_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_132_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_403 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_80 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_385 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0960__A _0988_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0830_ _0846_/A _0830_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_127_232 VGND VPWR sky130_fd_sc_hd__decap_12
X_0761_ _0675_/D _0750_/X _0759_/X _0760_/X _1088_/D VGND VPWR sky130_fd_sc_hd__o22a_4
X_0692_ _0739_/D _0558_/X _0692_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_37_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_154 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_1_0_clk clkbuf_0_clk/X clkbuf_2_3_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__0649__A1 _0626_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_19 VGND VPWR sky130_fd_sc_hd__decap_12
X_1175_ d_fabric_in[9] _0891_/D _1175_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_24_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_274 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1031__A _0981_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_160 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_32_193 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0821__B2 _0779_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0821__A1 _0663_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_27 VGND VPWR sky130_fd_sc_hd__decap_12
X_0959_ _0957_/X _0838_/B _0958_/X _0988_/C VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_118_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_176 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_403 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_222 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_288 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0812__A1 _0806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0812__B2 _0808_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_86 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1216__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0955__A _0955_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_241 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0674__B _0509_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0690__A _0544_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0803__B2 _0801_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0803__A1 _0799_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0813_ _0661_/Y _0813_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0744_ _0738_/X _0744_/B _0740_/X _0743_/X _0744_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_115_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_381 VGND VPWR sky130_fd_sc_hd__decap_12
X_0675_ _0740_/A _0677_/B _0676_/C _0675_/D _0684_/A VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_130_227 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1026__A _0985_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_185 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_399 VGND VPWR sky130_fd_sc_hd__decap_8
X_1227_ conf[1] _0841_/B _1142_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1158_ _1221_/Q _1158_/Q _1221_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_25_403 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0584__B _0585_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_406 VGND VPWR sky130_fd_sc_hd__fill_1
X_1089_ _1089_/D _1089_/Q _1114_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1047__A1 _1009_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0730__B1 _0719_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_347 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1038__A1 _0945_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_123 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_141 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_144 VGND VPWR sky130_fd_sc_hd__fill_2
X_1012_ _0985_/X _0983_/X _1011_/Y _1012_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_81_306 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_222 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_339 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_288 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0788__B1 _0739_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0727_ _0508_/A _0724_/X _0725_/X _0726_/X _0728_/D VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_103_238 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0579__B _0580_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0658_ _0501_/X _0551_/Y _0650_/X _0651_/Y _0657_/X _0658_/Y VGND VPWR sky130_fd_sc_hd__a32oi_4
X_0589_ _0579_/X _0580_/X _0583_/X _0588_/X _0589_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_69_141 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_111 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_336 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0595__A _1132_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0712__B1 _0487_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_277 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_269 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_138_168 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_134_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_282 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_339 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_169 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_158 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0952__B _0991_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_288 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_261 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_250 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_272 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_247 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0795__A2_N _0787_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_181 VGND VPWR sky130_fd_sc_hd__fill_2
X_0512_ _0722_/A _0512_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_100_208 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1084__CLK _1103_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_190 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_116_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_125 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_350 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_363 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_122_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_396 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_100 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_280 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0963__A _0950_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_361 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0682__B _0682_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_191 VGND VPWR sky130_fd_sc_hd__decap_3
X_0992_ _0991_/X _0992_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_8_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_206 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_4_7_0_clk clkbuf_4_7_0_clk/A _1201_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__1034__A _0948_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_261 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_306 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0576__C _0725_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_125 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_300 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_35 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0685__A2 _0684_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0783__A _0720_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_22 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_7 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_206 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0677__B _0677_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_239 VGND VPWR sky130_fd_sc_hd__decap_12
X_1191_ d_fabric_in[25] _1191_/Q _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_39_90 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0765__A1_N _0614_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_169 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_286 VGND VPWR sky130_fd_sc_hd__fill_2
X_0975_ _0946_/A _0966_/Y _0960_/X _0975_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
XANTENNA__1029__A _0988_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1122__CLK _1127_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0587__B _1153_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_250 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_147 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_253 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_117 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_59 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_150 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_109_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_136_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_272 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_158 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0658__A2 _0551_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_117 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_70 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0960__B _0955_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0760_ _0677_/D _0496_/A _0709_/X _0760_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__1145__CLK _1114_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_80 VGND VPWR sky130_fd_sc_hd__fill_1
X_0691_ _1142_/Q _0739_/D VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0688__A _0688_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_199 VGND VPWR sky130_fd_sc_hd__decap_12
X_1174_ d_fabric_in[8] _1174_/Q _1174_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0649__A2 _0632_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_117 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1031__B _1021_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_172 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0821__A2 _1114_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0958_ _0883_/A _0885_/A _0833_/A _0958_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_106_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_288 VGND VPWR sky130_fd_sc_hd__decap_12
X_0889_ _1174_/Q _0877_/X _0888_/Y d_sram_in[8] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_133_269 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0598__A _0579_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_323 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_264 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_275 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_286 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0928__B1_N _0867_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1168__CLK _1201_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0812__A2 _1107_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_247 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_301 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_98 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0955__B _0991_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_212 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_234 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_245 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0971__A _0940_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0690__B _0617_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0803__A2 _1100_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0812_ _0806_/X _1107_/Q _0544_/D _0808_/X d_fabric_out[24] VGND VPWR sky130_fd_sc_hd__o22a_4
X_0743_ _0616_/X _0509_/B _0741_/X _0743_/D _0743_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_6_393 VGND VPWR sky130_fd_sc_hd__decap_4
X_0674_ _0674_/A _0509_/B _0674_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_115_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_367 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1026__B _0995_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_337 VGND VPWR sky130_fd_sc_hd__decap_12
X_1226_ conf[0] _1226_/Q _1226_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_253 VGND VPWR sky130_fd_sc_hd__fill_1
X_1157_ _0840_/A _1157_/Q _1174_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0584__C _0585_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1042__A _0899_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1088_ _1088_/D _0763_/B _1114_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1047__A2 _0838_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0881__A _0835_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_79_109 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_239 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_57 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0730__A1 _1117_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_79 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_359 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_113_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_223 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_234 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_245 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1038__A2 _1035_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_289 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1102__D _0695_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_306 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_135 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_1_0_0_clk clkbuf_0_clk/X clkbuf_1_0_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_22_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_228 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0966__A _0966_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_315 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_220 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_66_337 VGND VPWR sky130_fd_sc_hd__decap_12
X_1011_ _1009_/X _1028_/A _0988_/C _1011_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_34_234 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0788__B2 _0787_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_128_361 VGND VPWR sky130_fd_sc_hd__decap_12
X_0726_ _0544_/A _0513_/X _1113_/D _0725_/C _0726_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_103_206 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_217 VGND VPWR sky130_fd_sc_hd__fill_1
X_0657_ _0716_/A _0502_/A _0655_/X _0656_/X _0657_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XANTENNA__0579__C _0579_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0588_ _0584_/X _0585_/X _0586_/X _0587_/X _0588_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0712__A1 _0750_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_175 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0876__A _0920_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0595__B _0583_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0712__B2 _0711_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1209_ addr_w[11] _0940_/C _1161_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_84_178 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_289 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_125 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1206__CLK _1221_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_311 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_250 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_366 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_304 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_337 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_359 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_123 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_156 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_251 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_240 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0952__C _1010_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_273 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_262 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_342 VGND VPWR sky130_fd_sc_hd__decap_12
X_0511_ _0544_/A _0722_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_98_226 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_39_304 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0696__A _0518_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0933__A1 _1191_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0709_ _0501_/X _0709_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_131_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_137 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_362 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_170 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_13 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_403 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0621__B1 _0620_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_312 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0924__A1 _1184_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_270 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_152 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0682__C _0682_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0991_ _0991_/A _0991_/B _0991_/C _0991_/D _0991_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0860__B1 _0880_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_263 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0915__A1 _0912_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_240 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0576__D _0505_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1034__B _0956_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_192 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1200__D addr_w[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0906__A1 _1178_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_389 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_47 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_240 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0783__B _0750_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_34 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_354 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1110__D _1142_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0677__C _0677_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1190_ d_fabric_in[24] _1190_/Q _1187_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0974__A _0973_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_137 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_398 VGND VPWR sky130_fd_sc_hd__decap_8
X_0974_ _0973_/X _0974_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1029__B _1029_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_315 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1045__A _0955_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0587__C _0587_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_19_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0884__A _0903_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_107 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_265 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1077__B1 _1076_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_129 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_354 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_173 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_195 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1097__CLK _1142_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_262 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_284 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1105__D _0723_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0658__A3 _0650_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_73_221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1068__B1 _1067_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_60 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_173 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_93 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0960__C _0988_/C VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_6_0_clk clkbuf_4_7_0_clk/A _1116_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_127_245 VGND VPWR sky130_fd_sc_hd__decap_12
X_0690_ _0544_/C _0617_/A _0690_/C _0679_/D _0690_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0969__A _0969_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0688__B _0687_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_240 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_178 VGND VPWR sky130_fd_sc_hd__decap_8
X_1173_ d_fabric_in[7] _1173_/Q _1187_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0649__A3 _0636_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_276 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_129 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1031__C _1024_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_192 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_140 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_324 VGND VPWR sky130_fd_sc_hd__decap_12
X_0957_ _0956_/X _0957_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_9_391 VGND VPWR sky130_fd_sc_hd__decap_12
X_0888_ _0880_/X _0887_/X _0861_/A _0888_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__0879__A _1010_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_140 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_184 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_221 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_32 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_268 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_278 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_11_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_127_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0955__C _0991_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_298 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1112__CLK _1103_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0690__C _0690_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0811_ _0806_/X _1106_/Q _1138_/Q _0808_/X d_fabric_out[23] VGND VPWR sky130_fd_sc_hd__o22a_4
X_0742_ _0725_/A _0544_/B _0725_/C _0695_/X _0743_/D VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_6_361 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0699__A _0699_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0673_ _0673_/A _0674_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_42_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_96_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_305 VGND VPWR sky130_fd_sc_hd__fill_2
X_1225_ addr_r[13] _1225_/Q _1185_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_84_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_232 VGND VPWR sky130_fd_sc_hd__fill_2
X_1156_ _0841_/B _1156_/Q _1174_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0584__D _0677_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_224 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1042__B _0899_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_268 VGND VPWR sky130_fd_sc_hd__fill_2
X_1087_ _0754_/X _0755_/B _1114_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_20_154 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_248 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_143 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0730__A2 _0548_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1135__CLK _1175_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_319 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_308 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_276 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_110 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_290 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_318 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_351 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_94 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_292 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_262 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_251 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_327 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_135 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_66_349 VGND VPWR sky130_fd_sc_hd__decap_12
X_1010_ _0948_/X _0956_/X _1010_/C _1028_/A VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_93_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_80 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0982__A _0991_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_246 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_373 VGND VPWR sky130_fd_sc_hd__decap_12
X_0725_ _0725_/A _0544_/B _0725_/C _0594_/A _0725_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0656_ _0544_/D _0656_/B _0656_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0579__D _1130_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_110 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1158__CLK _1221_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0927__B1_N _0862_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0587_ _0587_/A _1153_/Q _0587_/C _0720_/A _0587_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_69_121 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_69_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0712__A2 _0672_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1208_ addr_w[10] _0940_/A _1161_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_27_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_308 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1203__D addr_w[5] VGND VPWR sky130_fd_sc_hd__diode_2
X_1139_ d_sram_out[24] _0543_/A _1142_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_40_205 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_396 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_138_137 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_117 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_134_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_13 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_323 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_316 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_113 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_84_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1113__D _1113_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_363 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_252 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_241 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_230 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_274 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_263 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_159 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_354 VGND VPWR sky130_fd_sc_hd__decap_12
X_0510_ _1151_/Q _0544_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_3_161 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0977__A _0940_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0696__B _0701_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_179 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_74_190 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_62_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_227 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1048__A _1048_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0933__A2 _0932_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_205 VGND VPWR sky130_fd_sc_hd__decap_4
X_0708_ _0705_/X _0706_/Y _0707_/X _0708_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_0639_ _0723_/D _0639_/B _0639_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0887__A _0899_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_271 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_182 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0621__A1 _0591_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_343 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_324 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0924__A2 _0907_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_195 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_120 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1108__D _0602_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0797__A _1146_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_113 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_48_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_330 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_160 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_385 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0682__D _1128_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0990_ _0968_/X _0983_/X _0989_/X w_mask[4] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0860__A1 _0826_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_80 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_125_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_86 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0915__A2 _0907_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0500__A _0499_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_146 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1034__C _1024_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_296 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_190 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_333 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_131_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_335 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0906__A2 _0877_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_46 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_84 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_195 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_184 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_122_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_219 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1219__CLK _1124_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0677__D _0677_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_252 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_105 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_285 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_160 VGND VPWR sky130_fd_sc_hd__fill_2
X_0973_ _0978_/A _0982_/B _0973_/C _0991_/D _0973_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_72_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1029__C _1028_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_208 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_327 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1045__B _1009_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0587__D _0720_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_82_200 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_27_127 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_406 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1077__A1 _1025_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_160 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1211__D addr_w[13] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_176 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0760__B1 _0709_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_230 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_68 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_233 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_300 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1068__A1 _1006_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_50 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1121__D d_sram_out[6] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_94 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_127_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0751__B1 _0635_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0985__A _0985_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1191__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1172_ d_fabric_in[6] _1172_/Q _1114_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_64_200 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0649__A4 _0647_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_285 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_296 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_211 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_406 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1031__D _1003_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_118_202 VGND VPWR sky130_fd_sc_hd__decap_12
X_0956_ _0956_/A _0956_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0887_ _0899_/A _0899_/B _0903_/C _1174_/Q _0887_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0990__B1 _0989_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_163 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1056__A _1048_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_196 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_336 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1206__D addr_w[8] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_135 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0895__A _0899_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_44 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_247 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_174 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1116__D d_sram_out[1] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_403 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0955__D _0955_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_211 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_266 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_141 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0690__D _0679_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0810_ _0806_/X _1105_/Q _0723_/D _0808_/X d_fabric_out[22] VGND VPWR sky130_fd_sc_hd__o22a_4
X_0741_ _0544_/A _0513_/X _0724_/C _1130_/Q _0741_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_6_373 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0699__B _0699_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0672_ _0668_/X _0673_/A _0501_/X _0671_/X _0672_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_35_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_328 VGND VPWR sky130_fd_sc_hd__fill_2
X_1224_ addr_r[12] _1224_/Q _1161_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_92_361 VGND VPWR sky130_fd_sc_hd__decap_12
X_1155_ _1226_/Q _1155_/Q _1174_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1086_ _0747_/X _1086_/Q _1114_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1042__C _0835_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_247 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_258 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1087__CLK _1114_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0939_ _1197_/Q _0876_/X _0918_/Y d_sram_in[31] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_121_208 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0715__B1 _0714_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_15 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_5_0_clk clkbuf_3_2_0_clk/X _1175_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_16_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_113_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_288 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_363 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_271 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0706__B1 _0622_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_92 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0982__B _0982_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_394 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_385 VGND VPWR sky130_fd_sc_hd__decap_12
X_0724_ _0544_/A _0513_/X _0724_/C _0724_/D _0724_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0503__A _0503_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0655_ _1099_/D _0771_/B _0655_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0586_ _0585_/A _0585_/B _0587_/C _1117_/Q _0586_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_69_133 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_339 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0712__A3 _0710_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_188 VGND VPWR sky130_fd_sc_hd__fill_2
X_1207_ addr_w[9] _0956_/A _1221_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1138_ d_sram_out[23] _1138_/Q _1161_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_80_320 VGND VPWR sky130_fd_sc_hd__fill_2
X_1069_ _1015_/X _1059_/X _1067_/X w_mask[25] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_40_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_239 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0778__A1_N _0509_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_149 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_300 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1102__CLK _1116_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_335 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_328 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_331 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_191 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_217 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_242 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_231 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_220 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_275 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_264 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_253 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_173 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_306 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0696__C _0702_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_125 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_158 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0577__A2_N _0576_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_117 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_116_300 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1125__CLK _1103_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1048__B _1048_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0707_ _1116_/Q _0622_/Y _0550_/X _0707_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_89_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_239 VGND VPWR sky130_fd_sc_hd__decap_3
X_0638_ _0722_/D _0558_/X _0638_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0887__B _0899_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1064__A _1009_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0569_ _1153_/Q _0579_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_57_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1214__D addr_r[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_110_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_194 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0621__A2 _0619_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_355 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0909__B1 _0908_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0797__B _0659_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_261 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_187 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1124__D d_sram_out[9] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0911__B1_N _0910_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_172 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_93 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0860__A2 _0859_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1148__CLK _1174_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0988__A _0988_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1034__D _1003_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_54_128 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_19 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_301 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_108_108 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1059__A _1043_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_141 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1209__D addr_w[11] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_369 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_253 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_286 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_161 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_58 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1119__D d_sram_out[4] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_257 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0601__A _0583_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_242 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_128 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_312 VGND VPWR sky130_fd_sc_hd__decap_12
X_0972_ _0940_/D _0991_/D VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_118_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_301 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0511__A _0544_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_339 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1045__C _0973_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_275 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_223 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1077__A2 _1070_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_194 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_269 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_21 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_104_166 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0760__A1 _0677_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_361 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_161 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_40 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_312 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1068__A2 _1059_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_51 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_62 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_62 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_142 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_153 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_84 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_83 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0751__A1 _0668_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_1_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_44 VGND VPWR sky130_fd_sc_hd__decap_12
X_1171_ d_fabric_in[5] _1171_/Q _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_49_264 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_289 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0506__A _0505_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_197 VGND VPWR sky130_fd_sc_hd__fill_2
X_0955_ _0955_/A _0991_/B _0991_/C _0955_/D _0955_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0886_ _0908_/C _0903_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0990__A1 _0968_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1056__B _1056_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0895__B _0899_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1222__D addr_r[10] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_226 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_131 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_259 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1209__CLK _1161_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_269 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_124_239 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_11_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_191 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_180 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_204 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1132__D d_sram_out[17] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_93 VGND VPWR sky130_fd_sc_hd__decap_3
X_0740_ _0740_/A _0740_/B _0722_/C _1138_/Q _0740_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0699__C _0697_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0671_ _0512_/X _0677_/B _0676_/D _0487_/X _0771_/B _0671_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XFILLER_123_250 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_145 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_1223_ addr_r[11] _1223_/Q _1201_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_96_189 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_245 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_256 VGND VPWR sky130_fd_sc_hd__decap_12
X_1154_ _1162_/Q _1154_/Q _1185_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_92_373 VGND VPWR sky130_fd_sc_hd__decap_12
X_1085_ _1085_/D _1085_/Q _1114_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1042__D _1042_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0938_ _1196_/Q _0876_/X _0914_/Y d_sram_in[30] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_106_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_239 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_106_228 VGND VPWR sky130_fd_sc_hd__fill_2
X_0869_ _1172_/Q _0869_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1217__D addr_r[5] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0715__A1 _0663_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_59 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_3 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1181__CLK _1226_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_138_63 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_209 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1127__D d_sram_out[12] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0706__A1 _0674_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_145 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_148 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_245 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0982__C _0991_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_32 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0723_ _0740_/A _0740_/B _0722_/C _0723_/D _0723_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0654_ _0690_/C _0771_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_0585_ _0585_/A _0585_/B _0585_/C _1116_/Q _0585_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_69_123 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_111_231 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_318 VGND VPWR sky130_fd_sc_hd__decap_12
X_1206_ addr_w[8] baseaddr_w_sync[8] _1221_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA_clkbuf_4_7_0_clk_A clkbuf_4_7_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1137_ d_sram_out[22] _0723_/D _1124_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1068_ _1006_/X _1059_/X _1067_/X w_mask[24] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_33_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_106 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_323 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0936__A1 _1194_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_7 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_343 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_210 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_243 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_232 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_270 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_229 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_276 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_265 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_254 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_51 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0604__A _0557_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0927__A1 _1186_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_196 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0696__D _0695_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0863__B1 _0862_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_281 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0615__B1 _0678_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_251 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_4_0_clk clkbuf_3_2_0_clk/X _1142_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XANTENNA__0514__A _0513_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_312 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1048__C _1048_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0706_ _0674_/A _0629_/X _0622_/Y _0706_/Y VGND VPWR sky130_fd_sc_hd__a21oi_4
X_0637_ _1141_/Q _0722_/D VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0887__C _0903_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_240 VGND VPWR sky130_fd_sc_hd__fill_2
X_0568_ _0560_/Y _0562_/X _0567_/Y _0578_/B VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_97_295 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_284 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_262 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1064__B _1009_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0499_ _0620_/A _1147_/Q _0620_/C _0499_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_38_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_310 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_129 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_110_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_262 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0909__A1 _1171_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_367 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_122_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_144 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_135_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_284 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_192 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1140__D d_sram_out[25] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_93 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0988__B _0988_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_240 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_251 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_159 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_265 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0509__A _0509_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_313 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1013__B1 _1012_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_315 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1075__A _1066_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1225__D addr_r[13] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_45_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_3_4_0_clk_A clkbuf_3_5_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_302 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_64 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_269 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_15_0_clk_A clkbuf_3_7_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_307 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1135__D d_sram_out[20] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_91_235 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_170 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_354 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0818__B1 _0532_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_60 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1115__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_324 VGND VPWR sky130_fd_sc_hd__decap_12
X_0971_ _0940_/C _0973_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0999__A _0954_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_3 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1045__D _0987_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_254 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0809__B1 _0675_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_257 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_184 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0702__A _0724_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_2_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_189 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0760__A2 _0496_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_76_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1138__CLK _1161_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0925__B1_N _0855_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_276 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_132_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_129 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_30 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_279 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_52 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_324 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_63 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_74 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_85 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_198 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0612__A _0599_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0736__C1 _0735_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0751__A2 _1127_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_349 VGND VPWR sky130_fd_sc_hd__decap_12
X_1170_ d_fabric_in[4] _1170_/Q _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_2_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_154 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_80 VGND VPWR sky130_fd_sc_hd__decap_12
X_0954_ _0954_/A _0991_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_20_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_215 VGND VPWR sky130_fd_sc_hd__decap_12
X_0885_ _0885_/A _0908_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0522__A _1151_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0990__A2 _0983_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_110 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1056__C _1048_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0895__C _0903_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_268 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_279 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_110 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_154 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_198 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_305 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_279 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0607__A _1138_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_1_0_clk_A clkbuf_1_0_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_238 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_249 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_154 VGND VPWR sky130_fd_sc_hd__decap_12
X_0670_ _0602_/D _0676_/D VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0699__D _0698_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_273 VGND VPWR sky130_fd_sc_hd__fill_2
X_1222_ addr_r[10] _1222_/Q _1226_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_96_168 VGND VPWR sky130_fd_sc_hd__fill_2
X_1153_ _1161_/Q _1153_/Q _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_92_385 VGND VPWR sky130_fd_sc_hd__decap_12
X_1084_ _0712_/X _0714_/B _1103_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_268 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0517__A _0585_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_135 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0660__A1 _0487_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0937_ _1195_/Q _0932_/X _0910_/Y d_sram_in[29] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_20_179 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_3_0_clk_A clkbuf_4_3_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0868_ _0864_/Y _0833_/X _0867_/X d_sram_in[5] VGND VPWR sky130_fd_sc_hd__o21ai_4
X_0799_ _0661_/Y _0799_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_114_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_135 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0715__A2 _0712_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_87_168 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_87_146 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_319 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_113_45 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_330 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_341 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_227 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_238 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_271 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_135 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_125_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_75 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0706__A2 _0629_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_308 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_224 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1143__D d_sram_out[28] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_50 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_72 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_374 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0982__D _0991_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_190 VGND VPWR sky130_fd_sc_hd__decap_12
X_0722_ _0722_/A _0492_/C _0722_/C _0722_/D _0728_/B VGND VPWR sky130_fd_sc_hd__and4_4
X_0653_ _0740_/A _0716_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_40_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_0584_ _0505_/B _0585_/B _0585_/C _0677_/D _0584_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_111_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_113 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_105 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_84_149 VGND VPWR sky130_fd_sc_hd__fill_2
X_1205_ addr_w[7] baseaddr_w_sync[7] _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_65_330 VGND VPWR sky130_fd_sc_hd__decap_12
X_1136_ d_sram_out[21] _0675_/D _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_25_249 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_333 VGND VPWR sky130_fd_sc_hd__decap_3
X_1067_ _1044_/X _1025_/X _1066_/Y _1067_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_80_344 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_118 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_119_354 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0936__A2 _0932_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_335 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1228__D conf[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_16 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_232 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_124_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_287 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_102_276 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_127 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_330 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_149 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_182 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_200 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_355 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_233 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_222 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_277 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_266 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_255 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_244 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1138__D d_sram_out[23] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0927__A2 _0926_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_131 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0620__A _0620_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_105 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_93 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_333 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0863__A1 _0857_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_293 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0615__B2 _0558_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_324 VGND VPWR sky130_fd_sc_hd__decap_12
X_0705_ _0617_/X _0686_/X _0689_/X _0704_/X _0705_/X VGND VPWR sky130_fd_sc_hd__or4_4
XANTENNA__0530__A _0530_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0636_ _0676_/C _0686_/C _0635_/Y _0636_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XANTENNA__0887__D _1174_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0567_ _0583_/A _0580_/B _0530_/A _1118_/Q _0567_/Y VGND VPWR sky130_fd_sc_hd__nand4_4
XANTENNA__1064__C _0973_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_403 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0551__B1 _0550_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0498_ _1148_/Q _0620_/C VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1171__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_119 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_385 VGND VPWR sky130_fd_sc_hd__decap_12
X_1119_ d_sram_out[4] _0540_/D _1103_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_80_130 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_152 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0705__A _0617_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_119_184 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0909__A2 _0890_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_3_0_0_clk_A clkbuf_3_1_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0790__B1 _0532_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_122_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_241 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_156 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_11_0_clk_A clkbuf_3_5_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_73 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_110 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0988__C _0988_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0781__B1 _0676_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1194__CLK _1187_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_171 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0509__B _0509_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_141 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_325 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0525__A _1099_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1013__A1 _0998_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_327 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0772__B1 _0716_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1075__B _1074_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0619_ _0619_/A _0612_/Y _0618_/Y _0619_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_85_266 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_182 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_319 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_39_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_190 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_3_0_clk clkbuf_4_3_0_clk/A _1127_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_64_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_214 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_269 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_258 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0818__A1 _0813_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0818__B2 _0815_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1151__D _1159_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_185 VGND VPWR sky130_fd_sc_hd__fill_2
X_0970_ _0956_/A _0982_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0754__B1 _0752_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_200 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0809__A1 _0806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0809__B2 _0808_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_269 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_177 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0993__B1 _0989_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0702__B _0686_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_112_190 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_266 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_132_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_130 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_73_258 VGND VPWR sky130_fd_sc_hd__decap_6
XPHY_31 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_86 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_75 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_74 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0612__B _0612_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0736__B1 _0501_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_105 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1146__D d_sram_out[31] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_152 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_141 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_17_196 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_280 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0672__C1 _0671_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0953_ _0940_/C _0954_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_13_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_227 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0975__B1 _0960_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0884_ _0903_/B _0899_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_70_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_406 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0895__D _0895_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_46_19 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_225 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_236 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_216 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0713__A out_reg VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1105__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_328 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_203 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_258 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0607__B _0530_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_62 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_111_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_306 VGND VPWR sky130_fd_sc_hd__decap_12
X_1221_ addr_r[9] _1221_/Q _1221_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_96_158 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_309 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_236 VGND VPWR sky130_fd_sc_hd__fill_2
X_1152_ _1160_/Q _0504_/A _1201_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1083_ _0660_/X _0665_/A _1124_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_52_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_280 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_291 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0660__A2 _0496_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1128__CLK _1161_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0936_ _1194_/Q _0932_/X _0905_/Y d_sram_in[28] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__0533__A _0505_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0924__B1_N _0849_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0867_ _0864_/Y _0839_/X _0866_/Y _0867_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_0798_ _1130_/Q _0750_/X _0797_/X _0798_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0939__B1_N _0918_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_114_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_113_24 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_394 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_113_57 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_43_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_39 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_294 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_87 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_296 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_78_125 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_19_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_206 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0618__A _0552_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_386 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_261 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_94 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_283 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_300 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_56 VGND VPWR sky130_fd_sc_hd__decap_12
X_0721_ _0740_/A _0740_/B _0677_/C _1121_/Q _0721_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0652_ _0681_/A _0740_/A VGND VPWR sky130_fd_sc_hd__buf_1
X_0583_ _0583_/A _0579_/C _0583_/C _0673_/A _0583_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_88_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_158 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_128 VGND VPWR sky130_fd_sc_hd__decap_4
X_1204_ addr_w[6] baseaddr_w_sync[6] _1175_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1135_ d_sram_out[20] _0542_/D _1175_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0528__A _0527_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_301 VGND VPWR sky130_fd_sc_hd__fill_2
X_1066_ _1066_/A _1066_/B _1048_/C _1066_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_80_356 VGND VPWR sky130_fd_sc_hd__decap_12
X_0919_ _1181_/Q _0907_/X _0918_/Y d_sram_in[15] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_108_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_28 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_124_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_266 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_106 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_239 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_201 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_367 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_234 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_223 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_209 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_267 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_256 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_245 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_86 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0901__A _0854_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_110 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0620__B _1147_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1154__D _1162_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_342 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0863__A2 _0833_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_231 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_141 VGND VPWR sky130_fd_sc_hd__decap_12
X_0704_ _0690_/X _0704_/B _0699_/X _0704_/D _0704_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_131_306 VGND VPWR sky130_fd_sc_hd__decap_12
X_0635_ _0526_/X _0635_/B _0635_/C _0635_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_0566_ _0643_/B _0580_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1064__D _0955_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0497_ _0497_/A _0659_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0551__A1 _0509_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_139 VGND VPWR sky130_fd_sc_hd__fill_2
X_1118_ d_sram_out[3] _1118_/Q _1201_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1049_ _1044_/X _1006_/X _1048_/Y _1049_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_53_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0705__B _0686_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_196 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0721__A _0740_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_166 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0790__B2 _0787_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_220 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_168 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_139 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_97 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_52 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_80 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1149__D _1157_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0631__A _0700_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_306 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0781__B2 _0496_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_391 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_69_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_220 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_264 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_117 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_79_286 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_301 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_194 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0806__A _0661_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0525__B _0524_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1013__A2 _1006_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0541__A _0700_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_166 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0772__B2 _1130_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0772__A1 _0512_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_131_147 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1075__C _1048_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0618_ _0552_/Y _0613_/X _0615_/X _0617_/X _0618_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_112_361 VGND VPWR sky130_fd_sc_hd__decap_12
X_0549_ _0548_/X _0549_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_85_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_245 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0716__A _0716_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_199 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_41 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_372 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_234 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_289 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_131 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0818__A2 _1111_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_62 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0626__A _0682_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_73 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_84 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_50 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_280 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1161__CLK _1161_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0754__A1 _0542_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_147 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0754__B2 _0753_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_245 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_82_215 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_120 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0809__A2 _1104_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_164 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0536__A _0725_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_50_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_145 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0790__A2_N _0787_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0993__A1 _0968_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0702__C _0702_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_234 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_120 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_21 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_186 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_54 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_337 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_65 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_123 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_76 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1184__CLK _1187_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0612__C _0605_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0736__A1 _0668_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_110_117 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1162__D _1225_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_289 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_204 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0672__B1 _0501_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_93 VGND VPWR sky130_fd_sc_hd__decap_12
X_0952_ _0955_/A _0991_/B _1010_/C _0988_/A VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_9_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_239 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0975__A1 _0946_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0883_ _0883_/A _0903_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_63_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_123 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_204 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_218 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_123 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_318 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_2_0_clk clkbuf_4_3_0_clk/A _1163_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_87_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_270 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1157__D _0840_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_272 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_69_318 VGND VPWR sky130_fd_sc_hd__decap_12
X_1220_ addr_r[8] baseaddr_r_sync[8] _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_37_215 VGND VPWR sky130_fd_sc_hd__fill_2
X_1151_ _1159_/Q _1151_/Q _1116_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1082_ csb web _1163_/D VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_92_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_60_273 VGND VPWR sky130_fd_sc_hd__fill_2
X_0935_ _1193_/Q _0932_/X _0901_/Y d_sram_in[27] VGND VPWR sky130_fd_sc_hd__a21bo_4
X_0866_ _0866_/A _0866_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_9_171 VGND VPWR sky130_fd_sc_hd__decap_12
X_0797_ _1146_/Q _0659_/A _0797_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_28_204 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_270 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0724__A _0544_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_159 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0939__A1 _1197_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1061__B1 _1056_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1222__CLK _1226_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_242 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_85 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_96 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0618__B _0613_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_62 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0634__A _0542_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_295 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_312 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1052__B1 _1048_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_68 VGND VPWR sky130_fd_sc_hd__decap_12
X_0720_ _0720_/A _0506_/X _0720_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_6_141 VGND VPWR sky130_fd_sc_hd__decap_12
X_0651_ _0500_/X _0651_/Y VGND VPWR sky130_fd_sc_hd__inv_8
X_0582_ _0585_/C _0583_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_111_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_137 VGND VPWR sky130_fd_sc_hd__fill_2
X_1203_ addr_w[5] baseaddr_w_sync[5] _1171_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_26_3 VGND VPWR sky130_fd_sc_hd__fill_2
X_1134_ d_sram_out[19] _0695_/A _1201_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_65_354 VGND VPWR sky130_fd_sc_hd__decap_12
X_1065_ _1009_/A _0957_/X _1010_/C _1066_/B VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_80_368 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0544__A _0544_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_367 VGND VPWR sky130_fd_sc_hd__decap_12
X_0918_ _0854_/A _0918_/B _0918_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_134_337 VGND VPWR sky130_fd_sc_hd__decap_12
X_0849_ _0830_/Y _0839_/X _0848_/Y _0849_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_124_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0719__A _0651_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_140 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_302 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_83_184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_195 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_224 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_379 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_268 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_257 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_246 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_235 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_130_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_406 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_153 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_137_175 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0901__B _0901_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0620__C _0620_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0605__A1_N _0603_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1118__CLK _1201_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0629__A _0628_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_129 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1170__D d_fabric_in[4] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_313 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_151 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0938__B1_N _0914_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_276 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_337 VGND VPWR sky130_fd_sc_hd__decap_12
X_0703_ _0629_/X _0700_/X _0701_/X _0702_/X _0704_/D VGND VPWR sky130_fd_sc_hd__or4_4
X_0634_ _0542_/D _0690_/C _0635_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_131_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_232 VGND VPWR sky130_fd_sc_hd__fill_2
X_0565_ _0585_/B _0643_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_0496_ _0496_/A _0496_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0551__A2 _0546_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0539__A _0725_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_398 VGND VPWR sky130_fd_sc_hd__decap_8
X_1117_ d_sram_out[2] _1117_/Q _1187_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_110_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_1048_ _1048_/A _1048_/B _1048_/C _1048_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_53_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0705__C _0689_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1016__B1 _1012_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0721__B _0740_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_102_7 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_118 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_132 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_187 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0912__A _0903_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0631__B _0690_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1165__D _1165_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_257 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_151 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1090__CLK _1127_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0559__A1_N _0554_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_184 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0822__A d_sram_in[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_178 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0772__A2 _0677_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0617_ _0617_/A _0616_/X _0617_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_131_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_0548_ _0547_/X _0548_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_112_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_162 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_143 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0716__B _0720_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_56 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0732__A out_reg VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_53 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_162 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_44_121 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0907__A _0920_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_154 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0626__B _0686_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_32_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0642__A _0587_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_292 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0754__A2 _0750_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_213 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_293 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_271 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_260 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_198 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0552__A _1154_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0993__A2 _0992_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_281 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0702__D _1118_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_398 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0727__A _0508_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_154 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_22 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_198 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_165 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_22 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_44 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_349 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_66 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_157 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_179 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_99 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0612__D _0611_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_240 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0736__A2 _1126_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_235 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_268 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_110 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0637__A _1141_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_64_227 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0672__A1 _0668_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0951_ _0950_/Y _0991_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_32_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_342 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0975__A2 _0966_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0882_ _0903_/A _0899_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_56_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_99_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_319 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_330 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0547__A _0620_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_308 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_132_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1151__CLK _1116_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_208 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_312 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0920__A _1182_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_254 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_105 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0590__B1 _0578_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_138 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1173__D d_fabric_in[7] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_330 VGND VPWR sky130_fd_sc_hd__fill_2
X_1150_ _1158_/Q _0503_/A _1127_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1081_ _1040_/X _1043_/A _1079_/X w_mask[31] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_37_249 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_241 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_138 VGND VPWR sky130_fd_sc_hd__decap_12
X_0934_ _1192_/Q _0932_/X _0897_/Y d_sram_in[26] VGND VPWR sky130_fd_sc_hd__a21bo_4
X_0865_ _0827_/A _0859_/X _0844_/X _0866_/A VGND VPWR sky130_fd_sc_hd__a21o_4
XANTENNA__0830__A _0846_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0796_ _0713_/X _0795_/X _0785_/X _1097_/Q d_fabric_out[14] VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_114_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1083__D _0660_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1174__CLK _1174_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_374 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_300 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_227 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0724__B _0513_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_302 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1061__A1 _1044_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_56 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0939__A2 _0876_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_56 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_137_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0740__A _0740_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_311 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0618__C _0615_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_241 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_74 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0634__B _0690_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_324 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1052__A1 _1044_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1168__D d_fabric_in[2] VGND VPWR sky130_fd_sc_hd__diode_2
X_0650_ _0621_/Y _0623_/X _0549_/Y _0649_/X _0650_/X VGND VPWR sky130_fd_sc_hd__a211o_4
X_0581_ _0581_/A _0503_/A _0585_/C VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_97_403 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1197__CLK _1114_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_149 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_111_257 VGND VPWR sky130_fd_sc_hd__decap_12
X_1202_ addr_w[4] baseaddr_w_sync[4] _1124_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_19_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_300 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_130 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_1_0_clk clkbuf_4_0_0_clk/A _1103_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1133_ d_sram_out[18] _0594_/A _1116_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_92_185 VGND VPWR sky130_fd_sc_hd__fill_2
X_1064_ _1009_/A _1009_/B _0973_/C _0955_/D _1066_/A VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_25_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_314 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_325 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0825__A _0840_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_403 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0544__B _0544_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_302 VGND VPWR sky130_fd_sc_hd__decap_3
X_0917_ _1173_/Q _1046_/C _0916_/X _0918_/B VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_119_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0560__A _1127_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_108_15 VGND VPWR sky130_fd_sc_hd__decap_12
X_0848_ _0847_/X _0848_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_134_349 VGND VPWR sky130_fd_sc_hd__decap_12
X_0779_ _0776_/A _0779_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_307 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_102_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_246 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_174 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_225 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_258 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_247 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_236 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_274 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_269 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_137_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0793__B1 _0792_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_85 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_325 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0645__A _0583_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_288 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0784__B1 _0783_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0702_ _0724_/C _0686_/C _0702_/C _1118_/Q _0702_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_128_198 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_116_349 VGND VPWR sky130_fd_sc_hd__decap_12
X_0633_ _0594_/A _0702_/C _0635_/B VGND VPWR sky130_fd_sc_hd__and2_4
X_0564_ _0555_/Y _0585_/B VGND VPWR sky130_fd_sc_hd__buf_1
X_0495_ _0497_/A _0496_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_303 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_314 VGND VPWR sky130_fd_sc_hd__decap_12
X_1116_ d_sram_out[1] _1116_/Q _1116_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1212__CLK _1185_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1047_ _1009_/B _0838_/B _0958_/X _1048_/C VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0555__A _1153_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_200 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0705__D _0704_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_110 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1016__A1 _0998_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_266 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0721__C _0677_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0775__B1 _0773_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_266 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_130_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_299 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_163 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_56_196 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_20 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_100_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0912__B _0903_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0631__C _0686_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_97 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_125_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0766__B1 _0719_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_330 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1181__D d_fabric_in[15] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_94_269 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_111 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_281 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0772__A3 _1146_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0616_ _1151_/Q _0505_/A _1146_/Q _0580_/A _0616_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_124_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_406 VGND VPWR sky130_fd_sc_hd__fill_1
X_0547_ _0620_/A _0488_/Y _0620_/C _0547_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_112_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_236 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1091__D _1091_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_291 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_306 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0996__B1 _0988_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1108__CLK _1124_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_105 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0937__B1_N _0910_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_76 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_239 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_174 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0626__C _0626_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0642__B _0643_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_99_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_251 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1176__D d_fabric_in[10] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_144 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_125 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_50_158 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0833__A _0833_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_219 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_129_293 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1086__D _0747_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_104_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_217 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0727__B _0724_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_12 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_34 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_45 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_261 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_67 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_361 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0743__A _0616_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_203 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0918__A _0854_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_133 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0657__C1 _0656_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_291 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_125 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0672__A2 _0673_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0950_ _0956_/A _0950_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0653__A _0740_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_180 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0829__B1_N _0922_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_354 VGND VPWR sky130_fd_sc_hd__decap_12
X_0881_ _0835_/A _0903_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_99_136 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_342 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0828__A _0828_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0547__B _0488_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_261 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_283 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_158 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0563__A _0587_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_219 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_208 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_105_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_132_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_406 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0738__A _0681_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_174 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_230 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0920__B _0920_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_277 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_123_266 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_96_117 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0590__B2 _0589_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0590__A1 _0682_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_301 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_375 VGND VPWR sky130_fd_sc_hd__decap_3
X_1080_ _1035_/X _1070_/X _1079_/X w_mask[30] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_60_253 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_117 VGND VPWR sky130_fd_sc_hd__decap_12
X_0933_ _1191_/Q _0932_/X _0893_/Y d_sram_in[25] VGND VPWR sky130_fd_sc_hd__a21bo_4
X_0864_ _1171_/Q _0864_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_9_184 VGND VPWR sky130_fd_sc_hd__decap_12
X_0795_ _0575_/Y _0787_/X _1113_/D _0711_/X _0795_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_102_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_288 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0558__A _0505_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_172 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_386 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_334 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_345 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0724__C _0724_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_275 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_286 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1061__A2 _1022_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0740__B _0740_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_117 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_105_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_247 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_10 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_239 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_76 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_60 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0618__D _0617_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_86 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_97 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1052__A2 _1015_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_154 VGND VPWR sky130_fd_sc_hd__decap_12
X_0580_ _0580_/A _0580_/B _0580_/C _0580_/D _0580_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__1184__D d_fabric_in[18] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_117 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_214 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_269 VGND VPWR sky130_fd_sc_hd__decap_12
X_1201_ addr_w[3] baseaddr_w_sync[3] _1201_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_92_142 VGND VPWR sky130_fd_sc_hd__decap_4
X_1132_ d_sram_out[17] _1132_/Q _1116_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1063_ _1001_/X _1059_/X _1061_/X w_mask[23] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_65_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0544__C _0544_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0916_ _0903_/A _0903_/B _0908_/C _1181_/Q _0916_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__0841__A _1226_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0847_ _0880_/A _0946_/A _0844_/X _0846_/X _0847_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_127_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1141__CLK _1201_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0778_ _0509_/A _0496_/X _0544_/D _0496_/X _1091_/D VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XANTENNA__1094__D _0788_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_109 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_215 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_259 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_248 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_237 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_226 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_125_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_3 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0793__A1 _0679_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_20 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_301 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_97 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_172 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0926__A _0920_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0645__B _0643_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_80 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1179__D d_fabric_in[13] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0661__A out_reg VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1164__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0701_ _0724_/C _0701_/B _0628_/B _1132_/Q _0701_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_128_166 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0784__A1 _0722_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_391 VGND VPWR sky130_fd_sc_hd__decap_12
X_0632_ _0544_/D _0627_/Y _0629_/X _0631_/X _0632_/X VGND VPWR sky130_fd_sc_hd__a211o_4
XFILLER_124_361 VGND VPWR sky130_fd_sc_hd__decap_12
X_0563_ _0587_/A _0583_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_97_212 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_190 VGND VPWR sky130_fd_sc_hd__decap_8
X_0494_ _0493_/X _0497_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_38_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_153 VGND VPWR sky130_fd_sc_hd__fill_2
X_1115_ d_sram_out[0] _1115_/Q _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0836__A _0835_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_326 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_134 VGND VPWR sky130_fd_sc_hd__fill_2
X_1046_ _1009_/A _1009_/B _1046_/C _1048_/B VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_80_145 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_212 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_245 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1089__D _1089_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1016__A2 _1015_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_278 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0571__A _0571_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_107_306 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0775__A1 _1138_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0721__D _1121_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0775__B2 _0774_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_88_201 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_175 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_123 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_44_11 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_44 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1187__CLK _1187_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0912__C _0908_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0766__A1 _0609_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_147 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_0_0_clk clkbuf_4_0_0_clk/A _1124_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_5_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0631__D _1127_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_106_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_223 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_245 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_94_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_175 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0656__A _0544_/D VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_293 VGND VPWR sky130_fd_sc_hd__decap_12
X_0615_ _0614_/Y _0576_/X _0678_/A _0558_/X _0615_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
X_0546_ _0509_/B _0546_/B _0546_/C _0545_/X _0546_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_105_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_120 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0566__A _0643_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_101 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0693__B1 _0692_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1029_ _0988_/C _1029_/B _1028_/X _1029_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_41_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0996__A1 _0985_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_248 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_142 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_292 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_145 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0788__A1_N _0554_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_44_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_31 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0642__C _0587_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_8 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1202__CLK _1124_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_263 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1192__D d_fabric_in[26] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0911__A1 _1179_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_35_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_156 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_292 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1010__A _0948_/X VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_3_7_0_clk clkbuf_3_7_0_clk/A clkbuf_3_7_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_104_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_150 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0902__A1 _1177_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0529_ _0528_/X _0530_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_58_226 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_132_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_281 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_145 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0666__B1 _0665_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_13 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0727__C _0725_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_240 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_46 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_46 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_68 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_284 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0743__B _0509_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1225__CLK _1185_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_220 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_207 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0918__B _0918_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_123 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0657__B1 _0655_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_262 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_148 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_7 VGND VPWR sky130_fd_sc_hd__decap_6
X_0880_ _0880_/A _1046_/C _0880_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__1187__D d_fabric_in[21] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_253 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_354 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0896__B1 _0895_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0828__B _0826_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_270 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1005__A _0991_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0648__B1 _0622_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0547__C _0620_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0844__A d_sram_in[0] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0936__B1_N _0905_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1073__B1 _1071_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0820__B1 _1113_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1097__D _0795_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_127_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_127_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_321 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0738__B _0682_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_207 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_36_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_251 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_262 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_66 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_77 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_88 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0811__B1 _1138_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_108_264 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_123_245 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0590__A2 _0628_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_123_289 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_129 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_74 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_295 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0664__A out_reg VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_265 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_129 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_276 VGND VPWR sky130_fd_sc_hd__decap_12
X_0932_ _0920_/B _0932_/X VGND VPWR sky130_fd_sc_hd__buf_1
X_0863_ _0857_/Y _0833_/X _0862_/X d_sram_in[4] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0802__B1 _1099_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3 VGND VPWR sky130_fd_sc_hd__decap_12
X_0794_ _0713_/X _0793_/X _0785_/X _1096_/Q d_fabric_out[13] VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_5_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0839__A _0839_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_321 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0558__B _1153_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_28 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_184 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_68_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_357 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_379 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0574__A _0518_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_243 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_51_254 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_298 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0724__D _0724_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_306 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0740__C _0722_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_234 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_105_245 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_120_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_129 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_259 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_365 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_195 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_335 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1037__B1 _1036_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_265 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_128_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_204 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_361 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0659__A _0659_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_129 VGND VPWR sky130_fd_sc_hd__fill_1
X_1200_ addr_w[2] baseaddr_w_sync[2] _1163_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__1093__CLK _1103_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_1131_ d_sram_out[16] _1099_/D _1103_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_77_184 VGND VPWR sky130_fd_sc_hd__decap_12
X_1062_ _0995_/X _1059_/X _1061_/X w_mask[22] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_92_165 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_92_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_251 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0544__D _0544_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0915_ _0912_/D _0907_/X _0914_/Y d_sram_in[14] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__0841__B _0841_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0846_ _0846_/A _0852_/B _0846_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0777_ _0762_/X _1090_/D _0776_/X d_fabric_out[7] VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_102_204 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0569__A _1153_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_124_27 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_216 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_249 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_238 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_227 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1019__B1 _1011_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_125_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0793__A2 _0711_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_313 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_281 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_346 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_143 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_198 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0645__C _0530_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_202 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0942__A _0941_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0700_ _0700_/A _0700_/B _0656_/B _1130_/Q _0700_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_128_178 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0784__A2 _0711_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1195__D d_fabric_in[29] VGND VPWR sky130_fd_sc_hd__diode_2
X_0631_ _0700_/A _0690_/C _0686_/C _1127_/Q _0631_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0562_ _0561_/X _0562_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_124_373 VGND VPWR sky130_fd_sc_hd__decap_12
X_0493_ _0493_/A _0493_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_24_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_324 VGND VPWR sky130_fd_sc_hd__decap_12
X_1114_ _1146_/Q _1114_/Q _1114_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_65_143 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_338 VGND VPWR sky130_fd_sc_hd__decap_12
X_1045_ _0955_/A _1009_/B _0973_/C _0987_/D _1048_/A VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_0_94 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0852__A _0851_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_21_224 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_257 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_119_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_318 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0775__A2 _0750_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0829_ _0880_/A _0826_/X _0922_/A d_sram_in[1] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_135_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_257 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_130_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_102 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_202 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0762__A _0663_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_8_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0912__D _0912_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_88 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0766__A2 _0765_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_373 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_86 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0923__C1 _0922_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_268 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0656__B _0656_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1131__CLK _1103_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_62_135 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_70_190 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_0614_ _1113_/D _0614_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__1008__A _0950_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0545_ _0545_/A _0545_/B _0544_/X _0545_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_112_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_249 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_154 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_271 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_121_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0693__A1 _0676_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_135 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_157 VGND VPWR sky130_fd_sc_hd__fill_2
X_1028_ _1028_/A _1027_/X _1028_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_53_179 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0582__A _0585_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0996__A2 _0979_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_104 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_107_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_310 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_376 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0757__A _0679_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_290 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1154__CLK _1185_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_44 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_66 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_88 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_99 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0492__A _0620_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_385 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0642__D _0540_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_98 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_136_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_192 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_184 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0911__A2 _0907_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0667__A _0493_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_271 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_135 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_35_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_285 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1010__B _0956_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_129 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1177__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0528_ _0527_/X _0528_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_100_335 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_396 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0902__A2 _0877_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_27 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0666__A1 _0663_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0727__D _0726_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_47 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_58 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_138 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0743__C _0741_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_265 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_330 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_184 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0487__A _1132_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_66_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_271 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0657__A1 _0716_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_330 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0950__A _0956_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_265 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0896__A1 _0846_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_208 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_102_19 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1005__B _0982_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0648__A1 _0509_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_63_241 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0844__B _0826_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1021__A _0978_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1073__A1 _1022_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0820__A1 _0663_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0820__B2 _0815_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_202 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_127_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_213 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_311 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_193 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0738__C _0677_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_154 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_187 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_56 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0811__A1 _0806_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0811__B2 _0808_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0590__A3 _0509_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_97 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_6_0_clk clkbuf_3_7_0_clk/A clkbuf_3_6_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_37_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_399 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0945__A _0945_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_60_200 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_233 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_288 VGND VPWR sky130_fd_sc_hd__decap_12
X_0931_ _1190_/Q _0926_/X _0888_/Y d_sram_in[24] VGND VPWR sky130_fd_sc_hd__a21bo_4
XFILLER_13_171 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1198__D addr_w[0] VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0680__A _0544_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0802__A1 _0799_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0862_ _0857_/Y _0839_/X _0861_/Y _0862_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0802__B2 _0801_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0793_ _0679_/D _0711_/X _0792_/X _0793_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_114_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_141 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_333 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0558__C _0725_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1215__CLK _1142_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_230 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0574__B _0579_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_391 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_327 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0740__D _1138_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_105_213 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_120_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_300 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_86_174 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_241 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_103_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_403 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_233 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1037__A1 _0985_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_406 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0796__B1 _0785_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0659__B _0658_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0935__B1_N _0901_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_7 VGND VPWR sky130_fd_sc_hd__decap_12
X_1130_ d_sram_out[15] _1130_/Q _1201_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_77_141 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_163 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_196 VGND VPWR sky130_fd_sc_hd__decap_12
X_1061_ _1044_/X _1022_/X _1056_/Y _1061_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0675__A _0740_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_263 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_391 VGND VPWR sky130_fd_sc_hd__decap_12
X_0914_ _0847_/X _0913_/X _0914_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
XANTENNA__0841__C _0885_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0845_ _0835_/A _0943_/B _0885_/A _0852_/B VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_134_308 VGND VPWR sky130_fd_sc_hd__fill_2
X_0776_ _0776_/A _0776_/B _0776_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_88_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_163 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0585__A _0585_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_17_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_380 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_188 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_206 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_239 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_228 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1019__A1 _0985_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_12_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_137_135 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0778__B1 _0544_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_3_137 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_130 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_260 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_325 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0495__A _0497_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_47_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_200 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0645__D _1121_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_361 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_93 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_51 VGND VPWR sky130_fd_sc_hd__decap_8
X_0630_ _0594_/B _0690_/C VGND VPWR sky130_fd_sc_hd__buf_1
X_0561_ _0585_/A _0555_/Y _1151_/Q _0503_/A _0561_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_124_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_258 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_236 VGND VPWR sky130_fd_sc_hd__fill_2
X_0492_ _0620_/A _0488_/Y _0492_/C _1148_/Q _0493_/A VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_17_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0889__B1_N _0888_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_53_306 VGND VPWR sky130_fd_sc_hd__fill_2
X_1113_ _1113_/D _1113_/Q _1114_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1044_ _0843_/A _1044_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_80_125 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_158 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_236 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0852__B _0852_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_0828_ _0828_/A _0826_/X _0922_/A VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_115_330 VGND VPWR sky130_fd_sc_hd__decap_12
X_0759_ _0757_/X _0758_/X _0719_/X _0759_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_135_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_136 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1083__CLK _1124_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_98 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0923__B1 _0844_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_79_236 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_206 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_133 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_18_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_147 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0953__A _0940_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_116_105 VGND VPWR sky130_fd_sc_hd__decap_12
X_0613_ _0697_/A _0701_/B _0594_/B _1141_/Q _0613_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_112_300 VGND VPWR sky130_fd_sc_hd__decap_12
X_0544_ _0544_/A _0544_/B _0544_/C _0544_/D _0544_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__1024__A _0991_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_166 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_38_188 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_53_114 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0693__A2 _0627_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_1027_ _0981_/A _0956_/X _0954_/A _0955_/D _1027_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_34_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_30_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_115_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_322 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_141 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_388 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0757__B _0656_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_272 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_188 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_166 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_125 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_111_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0492__B _0488_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_230 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0948__A _0969_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_67_217 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_67_228 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_196 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0683__A _0509_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1010__C _1010_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_403 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0596__D1 _0595_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_132_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_116_29 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_98_364 VGND VPWR sky130_fd_sc_hd__decap_12
X_0527_ _0581_/A _0490_/A _0527_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_58_206 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0858__A _0852_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_369 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_209 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0666__A2 _0660_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_169 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_158 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_37 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0593__A _0587_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_264 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_48 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_106 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_297 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0743__D _0743_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_135_288 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1121__CLK _1201_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_11 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0657__A2 _0502_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_57_283 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_231 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_117 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_233 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_114_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_126_288 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0678__A _0678_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_301 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0896__A2 _0890_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1005__C _0978_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0648__A2 _0629_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1073__A2 _1070_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1021__B _1021_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0820__A2 _1113_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_11_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1144__CLK _1175_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_127_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0588__A _0584_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_172 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0738__D _0580_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_297 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_22_161 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_312 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0811__A2 _1106_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_288 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0498__A _1148_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_301 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_334 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_367 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_231 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_245 VGND VPWR sky130_fd_sc_hd__fill_2
X_0930_ _1189_/Q _0926_/X _0873_/X d_sram_in[23] VGND VPWR sky130_fd_sc_hd__a21bo_4
XANTENNA__1167__CLK _1175_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_110 VGND VPWR sky130_fd_sc_hd__decap_12
X_0861_ _0861_/A _0861_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XANTENNA__0802__A2 _1099_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0792_ _1128_/Q _0493_/X _0792_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_3_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0558__D _0505_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_315 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1032__A _1031_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0574__C _0573_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_137_306 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_138_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_137_339 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_120_239 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_315 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_68 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_212 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_223 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1037__A2 _1001_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0796__A1 _0713_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0796__B2 _1097_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_128_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_385 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0956__A _0956_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_153 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_77_175 VGND VPWR sky130_fd_sc_hd__decap_8
X_1060_ _0992_/X _1059_/X _1057_/X w_mask[21] VGND VPWR sky130_fd_sc_hd__o21ai_4
XANTENNA__0675__B _0677_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_92_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_201 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_329 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_245 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0691__A _1142_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_119_306 VGND VPWR sky130_fd_sc_hd__decap_12
X_0913_ _1172_/Q _1046_/C _0912_/X _0913_/X VGND VPWR sky130_fd_sc_hd__a21o_4
X_0844_ d_sram_in[0] _0826_/X _0844_/X VGND VPWR sky130_fd_sc_hd__and2_4
X_0775_ _1138_/Q _0750_/X _0773_/X _0774_/X _1090_/D VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_102_228 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1027__A _0981_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_272 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0866__A _0866_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_123 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_27 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0585__B _0585_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_1189_ d_fabric_in[23] _1189_/Q _1187_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_83_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_178 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_207 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_234 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_392 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_229 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_218 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_33_15 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1019__A2 _0992_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_59 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0778__B2 _0496_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_147 VGND VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_5_0_clk clkbuf_3_5_0_clk/A clkbuf_3_5_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_118_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_320 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_149 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_364 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_78 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_89 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_337 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_197 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0776__A _0776_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_212 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_215 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_395 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1205__CLK _1163_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0560_ _1127_/Q _0560_/Y VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_97_204 VGND VPWR sky130_fd_sc_hd__fill_2
X_0491_ _0544_/B _0492_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0686__A _0676_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_1112_ _0678_/A _1112_/Q _1103_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1043_ _1043_/A _1043_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_63 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_117 VGND VPWR sky130_fd_sc_hd__decap_12
X_0827_ _0827_/A _0828_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_115_342 VGND VPWR sky130_fd_sc_hd__decap_12
X_0758_ _0668_/X _1128_/Q _0687_/X _0758_/X VGND VPWR sky130_fd_sc_hd__a21o_4
XFILLER_88_215 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_135_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_237 VGND VPWR sky130_fd_sc_hd__fill_2
X_0689_ _0677_/C _0617_/A _0689_/C _0689_/X VGND VPWR sky130_fd_sc_hd__and3_4
XFILLER_28_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_112 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_292 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_56_123 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_148 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1228__CLK _1174_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0934__B1_N _0897_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_109_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_51 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0923__A1 _1183_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_121_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_123 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_85_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_156 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_115 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_80 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_117 VGND VPWR sky130_fd_sc_hd__decap_12
X_0612_ _0599_/X _0612_/B _0605_/X _0611_/Y _0612_/Y VGND VPWR sky130_fd_sc_hd__nor4_4
XFILLER_112_312 VGND VPWR sky130_fd_sc_hd__decap_12
X_0543_ _0543_/A _0544_/D VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_38_101 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_240 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_145 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1024__B _0982_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_295 VGND VPWR sky130_fd_sc_hd__fill_2
X_1026_ _0985_/A _0995_/X _1029_/B VGND VPWR sky130_fd_sc_hd__nor2_4
XFILLER_34_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1040__A _1039_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0850__B1 _0849_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_30_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_103_334 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_301 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_103_367 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_178 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_41 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0492__C _0492_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_34 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_242 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_398 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1100__D _1132_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_93 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0964__A _0981_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_243 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0683__B _0683_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_129 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_129_231 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0596__C1 _0526_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_332 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_112_142 VGND VPWR sky130_fd_sc_hd__decap_8
X_0526_ _0525_/X _0526_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_98_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_98_376 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_197 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1035__A _1034_/X VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_38 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VPWR sky130_fd_sc_hd__decap_3
X_1009_ _1009_/A _1009_/B _0991_/C _0987_/D _1009_/X VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__1076__B1 _1075_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_49 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_59 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_212 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_218 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_23 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_137 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1067__B1 _1066_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_72_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_354 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0814__B1 _0676_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_49_7 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1096__CLK _1103_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_262 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1005__D _1024_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0694__A _0700_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_221 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1058__B1 _1057_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_287 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1021__C _0978_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0805__B1 _0695_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_215 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0869__A _1172_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_151 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0588__B _0585_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_335 VGND VPWR sky130_fd_sc_hd__fill_1
X_0509_ _0509_/A _0509_/B _0509_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_100_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_276 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_7_0_clk_A clkbuf_3_7_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1049__B1 _1048_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_14_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_173 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_10_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_234 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0779__A _0776_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_117_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_11 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_346 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_265 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_276 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_287 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_80 VGND VPWR sky130_fd_sc_hd__decap_6
X_0860_ _0826_/X _0859_/X _0880_/A _0861_/A VGND VPWR sky130_fd_sc_hd__o21a_4
X_0791_ _0713_/X _0790_/X _0785_/X _1095_/Q d_fabric_out[12] VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_114_215 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0689__A _0677_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_176 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_91_360 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1111__CLK _1127_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_51_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_51_235 VGND VPWR sky130_fd_sc_hd__fill_2
X_0989_ _0985_/X _0974_/X _0988_/Y _0989_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__0599__A _0518_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_113_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_154 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_47_14 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_74_327 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_221 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_349 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_103_86 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_279 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0796__A2 _0795_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_10_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_146 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0675__C _0676_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1134__CLK _1201_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_18_276 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0972__A _0940_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_33_224 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_119_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_290 VGND VPWR sky130_fd_sc_hd__decap_12
X_0912_ _0903_/A _0903_/B _0908_/C _0912_/D _0912_/X VGND VPWR sky130_fd_sc_hd__and4_4
X_0843_ _0843_/A _0946_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_0774_ _0580_/D _0659_/A _0709_/X _0774_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XANTENNA__1027__B _0956_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_240 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_143 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_154 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_295 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1043__A _1043_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0585__C _0585_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_56_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_39 VGND VPWR sky130_fd_sc_hd__decap_12
X_1188_ d_fabric_in[22] _1188_/Q _1201_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_71_319 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0882__A _0903_/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_219 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_246 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_332 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_240 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_68 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1157__CLK _1174_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0776__B _0776_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_135 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_224 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0792__A _1128_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1103__D _0542_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_15_257 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_227 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_136_170 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_86 VGND VPWR sky130_fd_sc_hd__decap_12
X_0490_ _0490_/A _0544_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_124_398 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0686__B _0771_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_102 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_113 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_349 VGND VPWR sky130_fd_sc_hd__decap_12
X_1111_ _0532_/A _1111_/Q _1127_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
X_1042_ _0899_/A _0899_/B _0835_/C _1042_/D _1043_/A VGND VPWR sky130_fd_sc_hd__nand4_4
XFILLER_65_157 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_80_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_75 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_149 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_119_159 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_134_129 VGND VPWR sky130_fd_sc_hd__decap_12
X_0826_ _0835_/A _0943_/B _0835_/C _0826_/X VGND VPWR sky130_fd_sc_hd__o21a_4
X_0757_ _0679_/D _0656_/B _0757_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA_clkbuf_4_6_0_clk_A clkbuf_4_7_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_115_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_324 VGND VPWR sky130_fd_sc_hd__decap_12
X_0688_ _0688_/A _0687_/X _0689_/C VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__0877__A _0876_/X VGND VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_4_15_0_clk clkbuf_3_7_0_clk/X _1171_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_96_271 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_56_157 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_12_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_107_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_398 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0923__A2 _0876_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_51 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0787__A _0496_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_260 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_62_105 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_160 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_182 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_220 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_116_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_192 VGND VPWR sky130_fd_sc_hd__fill_2
X_0611_ _0724_/C _0617_/A _0610_/Y _0611_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
X_0542_ _0681_/A _0513_/X _0544_/C _0542_/D _0545_/B VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_112_324 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0697__A _0697_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_85_219 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_208 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_271 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1024__C _1024_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_81_403 VGND VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_4_0_clk clkbuf_3_5_0_clk/A clkbuf_4_8_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
X_1025_ _1024_/X _1025_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_46_190 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_160 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_182 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_193 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0850__A1 _0830_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_107 VGND VPWR sky130_fd_sc_hd__decap_12
X_0809_ _0806_/X _1104_/Q _0675_/D _0808_/X d_fabric_out[21] VGND VPWR sky130_fd_sc_hd__o22a_4
XFILLER_115_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_346 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_130_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_208 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_146 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_69 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_149 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_182 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0492__D _1148_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_138_276 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_121_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_92 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_75_241 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__0964__B _1021_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_138 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0683__C _0681_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_171 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_1_1_0_clk_A clkbuf_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_129_243 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0596__B1 _0718_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0525_ _1099_/D _0524_/X _0525_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_112_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_305 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_388 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0933__B1_N _0893_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1218__CLK _1124_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0615__A1_N _0614_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_26_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_285 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_28 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VPWR sky130_fd_sc_hd__decap_3
X_1008_ _0950_/Y _1009_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1076__A1 _0985_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_300 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_39 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_288 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0890__A _1046_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_34_182 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1201__D addr_w[3] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_135_224 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_135_257 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_3_3_0_clk_A clkbuf_3_3_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_165 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_263 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_149 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1067__A1 _1044_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_160 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_60_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_56 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0814__B2 _0808_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0814__A1 _0813_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_130 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1111__D _0532_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_14_0_clk_A clkbuf_3_7_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_126_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_241 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0694__B _0700_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_274 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_285 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_296 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1058__A1 _0983_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_16_171 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_299 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__1021__D _1024_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0805__A1 _0799_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0805__B2 _0801_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_163 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_227 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_205 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1046__A _1009_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0588__C _0586_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0508_ _0508_/A _0509_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_86_325 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_135 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_252 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1190__CLK _1187_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0885__A _0885_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_27_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_200 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_211 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1049__A1 _1044_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_42_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_255 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_266 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_246 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0980__B1 _0975_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_23 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_131_293 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1106__D _1138_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_133_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_93 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_299 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_9_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_196 VGND VPWR sky130_fd_sc_hd__decap_12
X_0790_ _0560_/Y _0787_/X _0532_/A _0787_/X _0790_/X VGND VPWR sky130_fd_sc_hd__a2bb2o_4
XFILLER_114_227 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0689__B _0617_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_133 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_3_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_199 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_24_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_36_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_258 VGND VPWR sky130_fd_sc_hd__fill_2
X_0988_ _0988_/A _0988_/B _0988_/C _0988_/Y VGND VPWR sky130_fd_sc_hd__nor3_4
XFILLER_105_238 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0599__B _0701_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_325 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_113_293 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_144 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_47_26 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_199 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_233 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_103_98 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_269 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1086__CLK _1114_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_137_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_166 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0650__C1 _0649_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_398 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_2_0_0_clk_A clkbuf_1_0_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_306 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0675__D _0675_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_58_380 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_169 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_73_361 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_288 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_236 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_269 VGND VPWR sky130_fd_sc_hd__decap_12
X_0911_ _1179_/Q _0907_/X _0910_/Y d_sram_in[13] VGND VPWR sky130_fd_sc_hd__a21bo_4
X_0842_ _0841_/X _0843_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_127_330 VGND VPWR sky130_fd_sc_hd__decap_12
X_0773_ _0771_/X _0772_/X _0719_/X _0773_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_52_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_102_208 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1027__C _0954_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_391 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0585__D _1116_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_83_136 VGND VPWR sky130_fd_sc_hd__fill_2
X_1187_ d_fabric_in[21] _1187_/Q _1187_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA_clkbuf_4_2_0_clk_A clkbuf_4_3_0_clk/A VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_209 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_258 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_39 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0632__C1 _0631_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_344 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_118_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_155 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0792__B _0493_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_320 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_236 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_56 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_105 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_228 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1101__CLK _1116_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_24_7 VGND VPWR sky130_fd_sc_hd__decap_12
X_1110_ _1142_/Q _1110_/Q _1103_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0686__C _0686_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_65_147 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0983__A _0982_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_1041_ _0945_/A _1040_/X _1037_/X w_mask[15] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_0_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_87 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_117 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_61_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_74 VGND VPWR sky130_fd_sc_hd__decap_12
X_0825_ _0840_/A _0835_/C VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_127_171 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0917__B1 _0916_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0756_ _0663_/X _0754_/X _0755_/X d_fabric_out[4] VGND VPWR sky130_fd_sc_hd__a21o_4
X_0687_ _0675_/D _0690_/C _0687_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_29_306 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1204__D addr_w[6] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_106 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0893__A _0866_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0853__C1 _0852_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_100_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_239 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_272 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1124__CLK _1124_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_109_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_24 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_196 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_103 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_294 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_114 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1114__D _1146_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_28_361 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_172 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_93 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_232 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_182 VGND VPWR sky130_fd_sc_hd__fill_1
X_0610_ _0675_/D _0583_/C _0688_/A _0608_/X _0609_/X _0610_/Y VGND VPWR sky130_fd_sc_hd__a2111oi_4
XFILLER_50_81 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_124_141 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0978__A _0978_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0541_ _0700_/A _0544_/C VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0697__B _0700_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_78_250 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_125 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_283 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1024__D _1024_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_169 VGND VPWR sky130_fd_sc_hd__fill_1
X_1024_ _0991_/A _0982_/B _1024_/C _1024_/D _1024_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_93_275 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_139 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0850__A2 _0833_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1147__CLK _1174_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_107_119 VGND VPWR sky130_fd_sc_hd__decap_3
X_0808_ _0776_/A _0808_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0888__A _0880_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0739_ _0722_/A _0492_/C _0722_/C _0739_/D _0744_/B VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_115_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_358 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_130_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_111_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_114 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_84_264 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_48 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_161 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_111_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_194 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_138_211 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_58 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_126_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_202 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_141 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1109__D _1141_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_96_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA_clkbuf_4_10_0_clk_A clkbuf_3_5_0_clk/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0964__C _0940_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_297 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_256 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_191 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_289 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_267 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_70 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_81 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_92 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0683__D _0683_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_312 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_334 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_367 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_14_0_clk clkbuf_3_7_0_clk/X _1226_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0596__A1 _0695_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0524_ _0581_/A _0544_/B _0524_/X VGND VPWR sky130_fd_sc_hd__and2_4
XANTENNA__0501__A _0500_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_166 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_317 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_117 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_212 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_29 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_223 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_245 VGND VPWR sky130_fd_sc_hd__decap_3
X_1007_ _0981_/A _1009_/A VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1076__A2 _1035_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_22_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_172 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_39 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_89_356 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_334 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_231 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_275 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__1067__A2 _1025_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_172 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_367 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0814__A2 _1108_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_197 VGND VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_3_0_clk clkbuf_3_3_0_clk/A clkbuf_4_7_0_clk/A VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_0_271 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0694__C _0583_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_201 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_245 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1058__A2 _1043_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0991__A _0991_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_142 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0805__A2 _1102_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_117_269 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_132_239 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1046__B _1009_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_86_304 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0588__D _0587_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0507_ _0506_/X _0508_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_86_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_234 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1049__A2 _1006_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1212__D addr_r[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_258 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0980__A1 _0968_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_117_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_35 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_197 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_175 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_315 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_133_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_204 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1122__D d_sram_out[7] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_237 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1208__CLK _1161_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_239 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0689__C _0689_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_123 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0986__A _0955_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_68_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_145 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_234 VGND VPWR sky130_fd_sc_hd__decap_4
X_0987_ _0955_/A _0957_/X _0991_/C _0987_/D _0988_/B VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_8_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_217 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0599__C _0628_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1207__D addr_w[9] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_59_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_178 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_38 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_340 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_204 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_215 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_237 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_59 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_105 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0650__B1 _0549_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_136_320 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_104_272 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_104_250 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1117__D d_sram_out[2] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_77_145 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_212 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_392 VGND VPWR sky130_fd_sc_hd__decap_4
X_0910_ _0866_/A _0910_/B _0910_/Y VGND VPWR sky130_fd_sc_hd__nor2_4
X_0841_ _1226_/Q _0841_/B _0885_/A _0841_/X VGND VPWR sky130_fd_sc_hd__or3_4
XFILLER_127_342 VGND VPWR sky130_fd_sc_hd__decap_12
X_0772_ _0512_/X _0677_/B _1146_/Q _0716_/A _1130_/Q _0772_/X VGND VPWR sky130_fd_sc_hd__a32o_4
XANTENNA__1180__CLK _1116_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_5_171 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1027__D _0955_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_110_220 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_110_264 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_167 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_189 VGND VPWR sky130_fd_sc_hd__fill_2
X_1186_ d_fabric_in[20] _1186_/Q _1226_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_32_270 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0632__B1 _0629_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_116_9 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_312 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0935__A1 _1193_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_356 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_101_220 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_134 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_114_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_264 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_178 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_297 VGND VPWR sky130_fd_sc_hd__fill_2
XPHY_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0871__B1 _0870_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_70_332 VGND VPWR sky130_fd_sc_hd__decap_4
XPHY_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_387 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_398 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_51 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0623__B1 _0622_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_312 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0686__D _1128_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_1040_ _1039_/X _1040_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_0_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_373 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0862__B1 _0861_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_61_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_80 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_192 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_86 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0504__A _0504_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0824_ _0841_/B _0943_/B VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0917__A1 _1173_/Q VGND VPWR sky130_fd_sc_hd__diode_2
X_0755_ _0733_/A _0755_/B _0755_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_115_367 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_207 VGND VPWR sky130_fd_sc_hd__decap_4
X_0686_ _0676_/C _0771_/B _0686_/C _1128_/Q _0686_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_130_337 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_318 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0893__B _0892_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_71_118 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_129 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1070__A _1043_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1169_ d_fabric_in[3] _0851_/A _1187_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0853__B1 _0844_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1220__D addr_r[8] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_138_404 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_100_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_240 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0605__B1 _1142_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_4_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_106_312 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_109_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_334 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1030__B1 _1029_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_36 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_304 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_229 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_240 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_273 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_170 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_181 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_43_354 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1130__D d_sram_out[15] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_109_150 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_93 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0978__B _0991_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0540_ _0681_/A _0682_/B _0682_/C _0540_/D _0545_/A VGND VPWR sky130_fd_sc_hd__and4_4
XANTENNA__1099__CLK _1116_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_337 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0697__C _0580_/C VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0994__A _0948_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_93_254 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_232 VGND VPWR sky130_fd_sc_hd__fill_2
X_1023_ _0998_/X _1022_/X _1019_/X w_mask[11] VGND VPWR sky130_fd_sc_hd__o21ai_4
XFILLER_53_118 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_34_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_61_173 VGND VPWR sky130_fd_sc_hd__decap_3
X_0807_ _0806_/X _1103_/Q _0542_/D _0801_/X d_fabric_out[20] VGND VPWR sky130_fd_sc_hd__o22a_4
XANTENNA__1012__B1 _1011_/Y VGND VPWR sky130_fd_sc_hd__diode_2
X_0738_ _0681_/A _0682_/B _0677_/C _0580_/D _0738_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_103_304 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0888__B _0887_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1065__A _1009_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_0669_ _0740_/B _0677_/B VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_130_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_240 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_262 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_84_210 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1215__D addr_r[3] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_243 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1079__B1 _1075_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_55_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_354 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0826__B1 _0835_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_40_324 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_112_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_121_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_56 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1125__D d_sram_out[10] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_75_221 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0964__D _0940_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0817__B1 _0739_/D VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_60 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_398 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_346 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_129_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_32 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0596__A2 _0580_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_98_302 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_335 VGND VPWR sky130_fd_sc_hd__fill_1
X_0523_ _0523_/A _0581_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_112_178 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_329 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_66_210 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_265 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_276 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_202 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__1114__CLK _1114_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_19 VGND VPWR sky130_fd_sc_hd__decap_3
X_1006_ _1005_/X _1006_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_81_257 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_268 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_324 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0899__A _0899_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_123 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_346 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_106_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_189 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_210 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_122_32 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_287 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_17_129 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_151 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_268 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_25_184 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_306 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_154 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_40_176 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_126_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_62 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0602__A _0697_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_48_210 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1137__CLK _1124_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0694__D _1126_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_63_213 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0991__B _0991_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_31_110 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_290 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_91 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_190 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_361 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0512__A _0722_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_125_281 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_154 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1046__C _1046_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0506_ _0505_/X _0506_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_98_176 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_276 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_198 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_108_215 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0980__A2 _0979_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_89_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_143 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_117_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_47 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_4_13_0_clk clkbuf_3_6_0_clk/X _1185_/CLK VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_133_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_235 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_249 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_147 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_342 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_319 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_382 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_290 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0507__A _0506_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0986_ _0955_/D _0987_/D VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__0599__D _0543_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_101_402 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_371 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_257 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1223__D addr_r[11] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_82_352 VGND VPWR sky130_fd_sc_hd__decap_12
Xclkbuf_3_2_0_clk clkbuf_3_3_0_clk/A clkbuf_3_2_0_clk/X VGND VPWR sky130_fd_sc_hd__clkbuf_1
XFILLER_63_27 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_396 VGND VPWR sky130_fd_sc_hd__fill_1
XPHY_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_293 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__0650__A1 _0621_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_6_117 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_136_332 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_136_398 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_2_312 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_149 VGND VPWR sky130_fd_sc_hd__fill_2
XANTENNA__1133__D d_sram_out[18] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_41_271 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_53_93 VGND VPWR sky130_fd_sc_hd__fill_2
X_0840_ _0840_/A _0885_/A VGND VPWR sky130_fd_sc_hd__inv_8
X_0771_ _1138_/Q _0771_/B _0771_/X VGND VPWR sky130_fd_sc_hd__and2_4
XFILLER_127_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_116 VGND VPWR sky130_fd_sc_hd__decap_4
X_1185_ d_fabric_in[19] _1185_/Q _1185_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_91_193 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_64_396 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0632__A1 _0544_/D VGND VPWR sky130_fd_sc_hd__diode_2
X_0969_ _0969_/A _0978_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_118_398 VGND VPWR sky130_fd_sc_hd__decap_8
XANTENNA__0935__A2 _0932_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1218__D addr_r[6] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_133_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0700__A _0700_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_105 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0931__B1_N _0888_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_74_15 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_300 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_130_32 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0871__A1 _0869_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_293 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0623__A1 _1115_/Q VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_128_129 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_74 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_354 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_124_324 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1128__D d_sram_out[13] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_97_208 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_65_105 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_93 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_300 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0862__A1 _0857_/Y VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_9_98 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_80 VGND VPWR sky130_fd_sc_hd__decap_4
X_0823_ _1226_/Q _0835_/A VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_127_184 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0917__A2 _1046_/C VGND VPWR sky130_fd_sc_hd__diode_2
X_0754_ _0542_/D _0750_/X _0752_/X _0753_/X _0754_/X VGND VPWR sky130_fd_sc_hd__o22a_4
X_0685_ _0674_/X _0684_/Y _0550_/X _0685_/X VGND VPWR sky130_fd_sc_hd__o21a_4
XFILLER_115_379 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0520__A _0682_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_130_349 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_241 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_127 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_149 VGND VPWR sky130_fd_sc_hd__fill_2
X_1168_ d_fabric_in[2] _0846_/A _1201_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XANTENNA__0853__A1 _0827_/A VGND VPWR sky130_fd_sc_hd__diode_2
X_1099_ _1099_/D _1099_/Q _1116_/CLK VGND VPWR sky130_fd_sc_hd__dfxtp_4
XFILLER_100_68 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0605__B2 _0639_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_60_28 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_252 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_133_110 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_114_7 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1030__A1 _0945_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_69_48 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_379 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_208 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_125_98 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1170__CLK _1171_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_90_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_28_385 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_130 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_70_141 VGND VPWR sky130_fd_sc_hd__decap_12
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_245 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_162 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_109_184 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_124_154 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0978__C _0978_/C VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_112_349 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0697__D _0580_/D VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0780__B1 _0762_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0994__B _0956_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_38_116 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_330 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_149 VGND VPWR sky130_fd_sc_hd__fill_2
X_1022_ _1021_/X _1022_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_34_300 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_299 VGND VPWR sky130_fd_sc_hd__decap_6
XANTENNA__0515__A _0682_/B VGND VPWR sky130_fd_sc_hd__diode_2
X_0806_ _0661_/Y _0806_/X VGND VPWR sky130_fd_sc_hd__buf_1
XFILLER_115_110 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1012__A1 _0985_/X VGND VPWR sky130_fd_sc_hd__diode_2
X_0737_ _1126_/Q _0506_/X _0745_/B VGND VPWR sky130_fd_sc_hd__or2_4
XANTENNA__0888__C _0861_/A VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1065__B _0957_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_39_29 VGND VPWR sky130_fd_sc_hd__decap_12
X_0668_ _0716_/A _0668_/X VGND VPWR sky130_fd_sc_hd__buf_1
XANTENNA__1193__CLK _1221_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
X_0599_ _0518_/X _0701_/B _0628_/B _0543_/A _0599_/X VGND VPWR sky130_fd_sc_hd__and4_4
XFILLER_57_403 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__1079__A1 _0985_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_84_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_39 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_111_45 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0826__A1 _0835_/A VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_52_174 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_27 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_71_38 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_138_268 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_215 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_105_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_154 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_121_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_68 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_62 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_51 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_233 VGND VPWR sky130_fd_sc_hd__decap_8
XFILLER_35_108 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_288 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_16_300 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0817__A1 _0813_/X VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__0817__B2 _0815_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_43_130 VGND VPWR sky130_fd_sc_hd__decap_3
XANTENNA__1141__D d_sram_out[26] VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_358 VGND VPWR sky130_fd_sc_hd__decap_8
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_129_257 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_7 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_44 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_314 VGND VPWR sky130_fd_sc_hd__decap_12
X_0522_ _1151_/Q _0523_/A VGND VPWR sky130_fd_sc_hd__inv_8
XFILLER_3_281 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0753__B1 _0709_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_20_3 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_403 VGND VPWR sky130_fd_sc_hd__decap_4
XFILLER_120_190 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_222 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_19_171 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_81_236 VGND VPWR sky130_fd_sc_hd__fill_2
X_1005_ _0991_/A _0982_/B _0978_/C _1024_/D _1005_/X VGND VPWR sky130_fd_sc_hd__or4_4
XFILLER_34_152 VGND VPWR sky130_fd_sc_hd__fill_1
XANTENNA__0899__B _0899_/B VGND VPWR sky130_fd_sc_hd__diode_2
XANTENNA__1226__D conf[0] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_103_135 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_106_56 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_103_179 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_103_168 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_122_44 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1089__CLK _1114_/CLK VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_25_196 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_280 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_86 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_318 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_391 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_126_227 VGND VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_74 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0602__B _0701_/B VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_134_271 VGND VPWR sky130_fd_sc_hd__decap_4
XANTENNA__0735__B1 _0695_/X VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_95_306 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__1136__D d_sram_out[21] VGND VPWR sky130_fd_sc_hd__diode_2
XFILLER_36_406 VGND VPWR sky130_fd_sc_hd__fill_1
XFILLER_48_266 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_225 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_141 VGND VPWR sky130_fd_sc_hd__decap_12
XANTENNA__0991__C _0991_/C VGND VPWR sky130_fd_sc_hd__diode_2
XPHY_191 VGND VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_188 VGND VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_373 VGND VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3 VGND VPWR sky130_fd_sc_hd__fill_2
XFILLER_125_293 VGND VPWR sky130_fd_sc_hd__decap_12
X_0505_ _0505_/A _0505_/B _0505_/X VGND VPWR sky130_fd_sc_hd__or2_4
XFILLER_100_105 VGND VPWR sky130_fd_sc_hd__decap_12
.ends

