magic
tech sky130A
magscale 1 2
timestamp 1607364296
<< checkpaint >>
rect -3932 -3932 33932 83932
<< locali >>
rect 15761 56219 15795 56389
rect 15301 55063 15335 55233
rect 17693 55131 17727 55301
rect 15393 54587 15427 54757
rect 15117 51255 15151 51425
rect 20913 50711 20947 50881
rect 23765 50711 23799 50813
rect 21557 49147 21591 49317
rect 20177 47991 20211 48229
rect 21833 46495 21867 46597
rect 23765 46359 23799 46461
rect 22477 43095 22511 43401
rect 11897 39831 11931 40069
rect 21649 38811 21683 38981
rect 15577 38199 15611 38505
rect 15301 37655 15335 37893
rect 15761 36635 15795 36805
rect 8861 35547 8895 35717
rect 10057 35479 10091 35649
rect 10425 35479 10459 35717
rect 18889 35683 18923 35785
rect 14197 34935 14231 35241
rect 6009 34391 6043 34629
rect 22661 33303 22695 33609
rect 14657 32963 14691 33065
rect 9413 32827 9447 32929
rect 8493 31739 8527 31977
rect 9689 31875 9723 31977
rect 15117 31807 15151 31977
rect 7757 31331 7791 31433
rect 9689 28475 9723 28713
rect 11621 27999 11655 28101
rect 16221 27999 16255 28169
rect 16037 26911 16071 27013
rect 12173 26231 12207 26537
rect 10793 24599 10827 24905
rect 15577 22423 15611 22525
rect 10701 21335 10735 21437
rect 17693 21335 17727 21641
rect 14749 19159 14783 19261
rect 12633 18683 12667 18921
rect 13829 14943 13863 15113
<< viali >>
rect 13829 77333 13863 77367
rect 19165 77129 19199 77163
rect 13737 76993 13771 77027
rect 14105 76993 14139 77027
rect 19625 76993 19659 77027
rect 13829 76925 13863 76959
rect 19349 76925 19383 76959
rect 21005 76857 21039 76891
rect 15209 76789 15243 76823
rect 9965 76449 9999 76483
rect 21189 76449 21223 76483
rect 9689 76381 9723 76415
rect 12173 76381 12207 76415
rect 12449 76381 12483 76415
rect 19441 76381 19475 76415
rect 20913 76381 20947 76415
rect 13737 76313 13771 76347
rect 11253 76245 11287 76279
rect 22477 76245 22511 76279
rect 9781 76041 9815 76075
rect 20913 76041 20947 76075
rect 12173 75837 12207 75871
rect 13553 75837 13587 75871
rect 13829 75837 13863 75871
rect 10149 75701 10183 75735
rect 12633 75701 12667 75735
rect 13369 75701 13403 75735
rect 15117 75701 15151 75735
rect 21373 75701 21407 75735
rect 25053 75497 25087 75531
rect 10701 75361 10735 75395
rect 10425 75293 10459 75327
rect 23673 75293 23707 75327
rect 23949 75293 23983 75327
rect 11989 75157 12023 75191
rect 13553 75157 13587 75191
rect 10517 74953 10551 74987
rect 18889 74953 18923 74987
rect 24225 74953 24259 74987
rect 19349 74817 19383 74851
rect 19073 74749 19107 74783
rect 10793 74613 10827 74647
rect 20453 74613 20487 74647
rect 23949 74613 23983 74647
rect 19165 74409 19199 74443
rect 12449 74273 12483 74307
rect 12173 74205 12207 74239
rect 13553 74069 13587 74103
rect 12173 73865 12207 73899
rect 12633 73525 12667 73559
rect 14381 73253 14415 73287
rect 13001 73185 13035 73219
rect 12725 73117 12759 73151
rect 12817 72777 12851 72811
rect 13093 72437 13127 72471
rect 22569 72165 22603 72199
rect 21189 72097 21223 72131
rect 20913 72029 20947 72063
rect 20913 71349 20947 71383
rect 21373 71349 21407 71383
rect 22569 71077 22603 71111
rect 21189 71009 21223 71043
rect 20913 70941 20947 70975
rect 20913 70533 20947 70567
rect 26065 70465 26099 70499
rect 26433 70465 26467 70499
rect 21373 70397 21407 70431
rect 26157 70397 26191 70431
rect 27537 70261 27571 70295
rect 2789 70057 2823 70091
rect 26157 70057 26191 70091
rect 1409 69921 1443 69955
rect 1685 69853 1719 69887
rect 11345 69445 11379 69479
rect 2053 69377 2087 69411
rect 26065 69377 26099 69411
rect 26433 69377 26467 69411
rect 1685 69309 1719 69343
rect 11529 69309 11563 69343
rect 11805 69309 11839 69343
rect 26157 69309 26191 69343
rect 27721 69173 27755 69207
rect 26249 68969 26283 69003
rect 9137 68425 9171 68459
rect 9689 68425 9723 68459
rect 9321 68221 9355 68255
rect 10701 67337 10735 67371
rect 10885 67133 10919 67167
rect 11253 66997 11287 67031
rect 21649 66793 21683 66827
rect 17233 66657 17267 66691
rect 17693 66657 17727 66691
rect 21833 66657 21867 66691
rect 16957 66589 16991 66623
rect 17601 66521 17635 66555
rect 18245 66453 18279 66487
rect 21741 66249 21775 66283
rect 18061 66113 18095 66147
rect 18337 66045 18371 66079
rect 16865 65977 16899 66011
rect 17785 65977 17819 66011
rect 19717 65977 19751 66011
rect 16405 65909 16439 65943
rect 17233 65909 17267 65943
rect 18613 65637 18647 65671
rect 15301 65569 15335 65603
rect 15669 65569 15703 65603
rect 16129 65569 16163 65603
rect 17877 65569 17911 65603
rect 18337 65569 18371 65603
rect 17601 65501 17635 65535
rect 16129 65433 16163 65467
rect 17141 65161 17175 65195
rect 21649 65161 21683 65195
rect 24409 65161 24443 65195
rect 16037 65093 16071 65127
rect 14657 65025 14691 65059
rect 15117 65025 15151 65059
rect 15301 65025 15335 65059
rect 24869 65025 24903 65059
rect 15577 64957 15611 64991
rect 16037 64957 16071 64991
rect 16589 64957 16623 64991
rect 21833 64957 21867 64991
rect 24593 64957 24627 64991
rect 14381 64889 14415 64923
rect 17601 64889 17635 64923
rect 18245 64889 18279 64923
rect 22201 64889 22235 64923
rect 21741 64481 21775 64515
rect 21465 64413 21499 64447
rect 15117 64345 15151 64379
rect 15577 64277 15611 64311
rect 15945 64277 15979 64311
rect 23029 64277 23063 64311
rect 21557 64073 21591 64107
rect 21833 64073 21867 64107
rect 17049 63937 17083 63971
rect 18613 63937 18647 63971
rect 19073 63937 19107 63971
rect 15853 63869 15887 63903
rect 16129 63869 16163 63903
rect 16313 63869 16347 63903
rect 16773 63869 16807 63903
rect 18797 63869 18831 63903
rect 20453 63801 20487 63835
rect 15485 63733 15519 63767
rect 18889 63529 18923 63563
rect 23673 63461 23707 63495
rect 15669 63393 15703 63427
rect 16129 63393 16163 63427
rect 23581 63393 23615 63427
rect 24409 63393 24443 63427
rect 15485 63325 15519 63359
rect 24501 63325 24535 63359
rect 16129 63257 16163 63291
rect 23489 62985 23523 63019
rect 26065 62849 26099 62883
rect 26433 62849 26467 62883
rect 15669 62781 15703 62815
rect 23949 62781 23983 62815
rect 26157 62781 26191 62815
rect 16037 62713 16071 62747
rect 27813 62713 27847 62747
rect 15393 62645 15427 62679
rect 24225 62645 24259 62679
rect 26157 62441 26191 62475
rect 15945 62373 15979 62407
rect 16773 62305 16807 62339
rect 16497 62237 16531 62271
rect 16957 62237 16991 62271
rect 19073 62101 19107 62135
rect 13829 61897 13863 61931
rect 12449 61761 12483 61795
rect 20085 61761 20119 61795
rect 26065 61761 26099 61795
rect 26433 61761 26467 61795
rect 12173 61693 12207 61727
rect 12725 61693 12759 61727
rect 18981 61693 19015 61727
rect 19349 61693 19383 61727
rect 19809 61693 19843 61727
rect 26157 61693 26191 61727
rect 27813 61625 27847 61659
rect 15945 61557 15979 61591
rect 16313 61557 16347 61591
rect 16681 61557 16715 61591
rect 17325 61557 17359 61591
rect 18797 61557 18831 61591
rect 1593 61353 1627 61387
rect 12449 61353 12483 61387
rect 20729 61353 20763 61387
rect 26157 61353 26191 61387
rect 21465 61285 21499 61319
rect 26709 61285 26743 61319
rect 17141 61217 17175 61251
rect 17785 61217 17819 61251
rect 18061 61217 18095 61251
rect 19165 61217 19199 61251
rect 21189 61217 21223 61251
rect 22201 61217 22235 61251
rect 27445 61217 27479 61251
rect 17417 61149 17451 61183
rect 21373 61149 21407 61183
rect 22293 61149 22327 61183
rect 26617 61149 26651 61183
rect 27537 61149 27571 61183
rect 18061 61081 18095 61115
rect 19073 61081 19107 61115
rect 16221 61013 16255 61047
rect 18613 61013 18647 61047
rect 19349 61013 19383 61047
rect 2789 60809 2823 60843
rect 22017 60809 22051 60843
rect 22937 60809 22971 60843
rect 26893 60809 26927 60843
rect 27353 60809 27387 60843
rect 18889 60741 18923 60775
rect 1409 60673 1443 60707
rect 16129 60673 16163 60707
rect 16819 60673 16853 60707
rect 17509 60673 17543 60707
rect 19441 60673 19475 60707
rect 20637 60673 20671 60707
rect 22569 60673 22603 60707
rect 26525 60673 26559 60707
rect 1685 60605 1719 60639
rect 16037 60605 16071 60639
rect 16681 60605 16715 60639
rect 16957 60605 16991 60639
rect 17877 60605 17911 60639
rect 18245 60605 18279 60639
rect 18613 60605 18647 60639
rect 18889 60605 18923 60639
rect 20545 60605 20579 60639
rect 20913 60605 20947 60639
rect 16221 60265 16255 60299
rect 18245 60265 18279 60299
rect 16865 60197 16899 60231
rect 18797 60197 18831 60231
rect 17693 60129 17727 60163
rect 19441 60129 19475 60163
rect 19717 60129 19751 60163
rect 20637 60129 20671 60163
rect 21465 60129 21499 60163
rect 21741 60129 21775 60163
rect 22937 60129 22971 60163
rect 17417 60061 17451 60095
rect 17877 60061 17911 60095
rect 18981 60061 19015 60095
rect 21097 60061 21131 60095
rect 21833 60061 21867 60095
rect 22845 60061 22879 60095
rect 19717 59993 19751 60027
rect 1685 59925 1719 59959
rect 15853 59925 15887 59959
rect 16773 59925 16807 59959
rect 17785 59721 17819 59755
rect 15301 59653 15335 59687
rect 17509 59585 17543 59619
rect 20269 59585 20303 59619
rect 20913 59585 20947 59619
rect 21833 59585 21867 59619
rect 14933 59517 14967 59551
rect 16313 59517 16347 59551
rect 16589 59517 16623 59551
rect 16773 59517 16807 59551
rect 18613 59517 18647 59551
rect 18797 59517 18831 59551
rect 19073 59517 19107 59551
rect 19533 59517 19567 59551
rect 20637 59517 20671 59551
rect 21281 59517 21315 59551
rect 21557 59517 21591 59551
rect 22477 59517 22511 59551
rect 15761 59449 15795 59483
rect 19809 59449 19843 59483
rect 15577 59381 15611 59415
rect 17049 59381 17083 59415
rect 22201 59381 22235 59415
rect 22845 59381 22879 59415
rect 19809 59177 19843 59211
rect 15761 59109 15795 59143
rect 17601 59109 17635 59143
rect 21189 59109 21223 59143
rect 21465 59109 21499 59143
rect 15117 59041 15151 59075
rect 16221 59041 16255 59075
rect 16773 59041 16807 59075
rect 18613 59041 18647 59075
rect 19625 59041 19659 59075
rect 20085 59041 20119 59075
rect 22293 59041 22327 59075
rect 22477 59041 22511 59075
rect 23489 59041 23523 59075
rect 15945 58973 15979 59007
rect 17785 58973 17819 59007
rect 18337 58973 18371 59007
rect 18797 58973 18831 59007
rect 22017 58973 22051 59007
rect 23305 58973 23339 59007
rect 16681 58905 16715 58939
rect 17325 58905 17359 58939
rect 20453 58905 20487 58939
rect 14657 58837 14691 58871
rect 19073 58837 19107 58871
rect 19533 58837 19567 58871
rect 24317 58837 24351 58871
rect 2973 58633 3007 58667
rect 14473 58633 14507 58667
rect 16681 58633 16715 58667
rect 20269 58633 20303 58667
rect 21833 58633 21867 58667
rect 22201 58633 22235 58667
rect 23121 58633 23155 58667
rect 22477 58565 22511 58599
rect 3433 58497 3467 58531
rect 16405 58497 16439 58531
rect 18613 58497 18647 58531
rect 19165 58497 19199 58531
rect 19901 58497 19935 58531
rect 23673 58497 23707 58531
rect 24685 58497 24719 58531
rect 3157 58429 3191 58463
rect 14289 58429 14323 58463
rect 15301 58429 15335 58463
rect 15669 58429 15703 58463
rect 16221 58429 16255 58463
rect 19441 58429 19475 58463
rect 19625 58429 19659 58463
rect 21005 58429 21039 58463
rect 21281 58429 21315 58463
rect 21465 58429 21499 58463
rect 22293 58429 22327 58463
rect 24225 58429 24259 58463
rect 24501 58429 24535 58463
rect 4813 58361 4847 58395
rect 14197 58361 14231 58395
rect 18429 58361 18463 58395
rect 20453 58361 20487 58395
rect 14841 58293 14875 58327
rect 15209 58293 15243 58327
rect 17233 58293 17267 58327
rect 17877 58293 17911 58327
rect 23397 58293 23431 58327
rect 11989 58089 12023 58123
rect 14381 58089 14415 58123
rect 23397 58089 23431 58123
rect 20913 58021 20947 58055
rect 12173 57953 12207 57987
rect 14197 57953 14231 57987
rect 15761 57953 15795 57987
rect 16129 57953 16163 57987
rect 17233 57953 17267 57987
rect 19349 57953 19383 57987
rect 19717 57953 19751 57987
rect 21741 57953 21775 57987
rect 23765 57953 23799 57987
rect 23949 57953 23983 57987
rect 24501 57953 24535 57987
rect 3249 57885 3283 57919
rect 15393 57885 15427 57919
rect 16773 57885 16807 57919
rect 17601 57885 17635 57919
rect 17785 57885 17819 57919
rect 18981 57885 19015 57919
rect 21465 57885 21499 57919
rect 21925 57885 21959 57919
rect 22201 57885 22235 57919
rect 2697 57817 2731 57851
rect 14105 57817 14139 57851
rect 16129 57817 16163 57851
rect 17398 57817 17432 57851
rect 19717 57817 19751 57851
rect 24409 57817 24443 57851
rect 13553 57749 13587 57783
rect 14749 57749 14783 57783
rect 15025 57749 15059 57783
rect 17049 57749 17083 57783
rect 17509 57749 17543 57783
rect 18337 57749 18371 57783
rect 18613 57749 18647 57783
rect 20453 57749 20487 57783
rect 22569 57749 22603 57783
rect 23029 57749 23063 57783
rect 6561 57545 6595 57579
rect 13461 57545 13495 57579
rect 17141 57545 17175 57579
rect 18705 57545 18739 57579
rect 19533 57545 19567 57579
rect 22201 57545 22235 57579
rect 22753 57545 22787 57579
rect 23489 57545 23523 57579
rect 24225 57545 24259 57579
rect 18337 57477 18371 57511
rect 23949 57477 23983 57511
rect 2513 57409 2547 57443
rect 2697 57409 2731 57443
rect 2789 57409 2823 57443
rect 7297 57409 7331 57443
rect 14013 57409 14047 57443
rect 14657 57409 14691 57443
rect 18429 57409 18463 57443
rect 19809 57409 19843 57443
rect 3513 57341 3547 57375
rect 3617 57341 3651 57375
rect 7021 57341 7055 57375
rect 13553 57341 13587 57375
rect 14933 57341 14967 57375
rect 15485 57341 15519 57375
rect 16957 57341 16991 57375
rect 18208 57341 18242 57375
rect 20269 57341 20303 57375
rect 20545 57341 20579 57375
rect 21097 57341 21131 57375
rect 21649 57341 21683 57375
rect 22385 57341 22419 57375
rect 8677 57273 8711 57307
rect 15669 57273 15703 57307
rect 18061 57273 18095 57307
rect 20821 57273 20855 57307
rect 2145 57205 2179 57239
rect 12081 57205 12115 57239
rect 13737 57205 13771 57239
rect 14381 57205 14415 57239
rect 16221 57205 16255 57239
rect 16865 57205 16899 57239
rect 17417 57205 17451 57239
rect 17785 57205 17819 57239
rect 19073 57205 19107 57239
rect 2789 57001 2823 57035
rect 7021 57001 7055 57035
rect 13369 57001 13403 57035
rect 13737 57001 13771 57035
rect 14381 57001 14415 57035
rect 17877 57001 17911 57035
rect 20729 57001 20763 57035
rect 21097 57001 21131 57035
rect 21741 57001 21775 57035
rect 22109 57001 22143 57035
rect 23213 57001 23247 57035
rect 14105 56933 14139 56967
rect 17233 56933 17267 56967
rect 20269 56933 20303 56967
rect 21373 56933 21407 56967
rect 1685 56865 1719 56899
rect 13185 56865 13219 56899
rect 14197 56865 14231 56899
rect 15669 56865 15703 56899
rect 16221 56865 16255 56899
rect 18889 56865 18923 56899
rect 19349 56865 19383 56899
rect 19809 56865 19843 56899
rect 20913 56865 20947 56899
rect 22845 56865 22879 56899
rect 1409 56797 1443 56831
rect 15393 56797 15427 56831
rect 17601 56797 17635 56831
rect 19993 56797 20027 56831
rect 22477 56797 22511 56831
rect 16129 56729 16163 56763
rect 17049 56729 17083 56763
rect 18613 56729 18647 56763
rect 14749 56661 14783 56695
rect 15117 56661 15151 56695
rect 17371 56661 17405 56695
rect 17509 56661 17543 56695
rect 18245 56661 18279 56695
rect 1685 56457 1719 56491
rect 2053 56457 2087 56491
rect 15209 56457 15243 56491
rect 18521 56457 18555 56491
rect 19717 56457 19751 56491
rect 21741 56457 21775 56491
rect 23121 56457 23155 56491
rect 26065 56457 26099 56491
rect 13737 56389 13771 56423
rect 14841 56389 14875 56423
rect 15761 56389 15795 56423
rect 16405 56389 16439 56423
rect 16589 56389 16623 56423
rect 18337 56389 18371 56423
rect 21373 56389 21407 56423
rect 14933 56321 14967 56355
rect 14712 56253 14746 56287
rect 15945 56321 15979 56355
rect 16497 56321 16531 56355
rect 18429 56321 18463 56355
rect 19625 56321 19659 56355
rect 20085 56321 20119 56355
rect 26157 56321 26191 56355
rect 16276 56253 16310 56287
rect 18208 56253 18242 56287
rect 19073 56253 19107 56287
rect 19901 56253 19935 56287
rect 20361 56253 20395 56287
rect 20821 56253 20855 56287
rect 21925 56253 21959 56287
rect 22385 56253 22419 56287
rect 26433 56253 26467 56287
rect 14565 56185 14599 56219
rect 15761 56185 15795 56219
rect 16129 56185 16163 56219
rect 18061 56185 18095 56219
rect 21097 56185 21131 56219
rect 13277 56117 13311 56151
rect 14105 56117 14139 56151
rect 14473 56117 14507 56151
rect 15577 56117 15611 56151
rect 17233 56117 17267 56151
rect 17785 56117 17819 56151
rect 22109 56117 22143 56151
rect 22753 56117 22787 56151
rect 27721 56117 27755 56151
rect 14013 55913 14047 55947
rect 14381 55913 14415 55947
rect 17601 55913 17635 55947
rect 18429 55913 18463 55947
rect 20085 55913 20119 55947
rect 20453 55913 20487 55947
rect 22937 55913 22971 55947
rect 26157 55913 26191 55947
rect 17325 55845 17359 55879
rect 18797 55845 18831 55879
rect 10793 55777 10827 55811
rect 13185 55777 13219 55811
rect 14197 55777 14231 55811
rect 15577 55777 15611 55811
rect 16589 55777 16623 55811
rect 19625 55777 19659 55811
rect 20913 55777 20947 55811
rect 21373 55777 21407 55811
rect 21925 55777 21959 55811
rect 22385 55777 22419 55811
rect 23765 55777 23799 55811
rect 10517 55709 10551 55743
rect 16957 55709 16991 55743
rect 18061 55709 18095 55743
rect 19349 55709 19383 55743
rect 19809 55709 19843 55743
rect 22661 55709 22695 55743
rect 23397 55709 23431 55743
rect 23489 55709 23523 55743
rect 13369 55641 13403 55675
rect 14749 55641 14783 55675
rect 16865 55641 16899 55675
rect 12081 55573 12115 55607
rect 13645 55573 13679 55607
rect 15117 55573 15151 55607
rect 15761 55573 15795 55607
rect 16129 55573 16163 55607
rect 16497 55573 16531 55607
rect 16754 55573 16788 55607
rect 21097 55573 21131 55607
rect 21833 55573 21867 55607
rect 24869 55573 24903 55607
rect 10609 55369 10643 55403
rect 10885 55369 10919 55403
rect 13001 55369 13035 55403
rect 14933 55369 14967 55403
rect 16202 55369 16236 55403
rect 16681 55369 16715 55403
rect 17417 55369 17451 55403
rect 18226 55369 18260 55403
rect 19441 55369 19475 55403
rect 23121 55369 23155 55403
rect 23857 55369 23891 55403
rect 14749 55301 14783 55335
rect 16313 55301 16347 55335
rect 17049 55301 17083 55335
rect 17693 55301 17727 55335
rect 18337 55301 18371 55335
rect 22017 55301 22051 55335
rect 14620 55233 14654 55267
rect 14841 55233 14875 55267
rect 15301 55233 15335 55267
rect 16405 55233 16439 55267
rect 13461 55165 13495 55199
rect 14473 55165 14507 55199
rect 16037 55165 16071 55199
rect 18429 55233 18463 55267
rect 22661 55233 22695 55267
rect 25237 55233 25271 55267
rect 26065 55233 26099 55267
rect 26433 55233 26467 55267
rect 18061 55165 18095 55199
rect 19073 55165 19107 55199
rect 19993 55165 20027 55199
rect 20637 55165 20671 55199
rect 21281 55165 21315 55199
rect 22201 55165 22235 55199
rect 22569 55165 22603 55199
rect 24317 55165 24351 55199
rect 24409 55165 24443 55199
rect 25145 55165 25179 55199
rect 26157 55165 26191 55199
rect 17693 55097 17727 55131
rect 17785 55097 17819 55131
rect 18797 55097 18831 55131
rect 20085 55097 20119 55131
rect 13277 55029 13311 55063
rect 13645 55029 13679 55063
rect 14197 55029 14231 55063
rect 15301 55029 15335 55063
rect 15485 55029 15519 55063
rect 15945 55029 15979 55063
rect 21649 55029 21683 55063
rect 23489 55029 23523 55063
rect 27721 55029 27755 55063
rect 14105 54825 14139 54859
rect 17141 54825 17175 54859
rect 18153 54825 18187 54859
rect 19349 54825 19383 54859
rect 19625 54825 19659 54859
rect 20729 54825 20763 54859
rect 22385 54825 22419 54859
rect 24225 54825 24259 54859
rect 24685 54825 24719 54859
rect 12081 54757 12115 54791
rect 12725 54757 12759 54791
rect 15117 54757 15151 54791
rect 15393 54757 15427 54791
rect 16681 54757 16715 54791
rect 18245 54757 18279 54791
rect 23029 54757 23063 54791
rect 12173 54689 12207 54723
rect 13185 54689 13219 54723
rect 14197 54689 14231 54723
rect 14657 54621 14691 54655
rect 15669 54689 15703 54723
rect 18061 54689 18095 54723
rect 19441 54689 19475 54723
rect 19901 54689 19935 54723
rect 21097 54689 21131 54723
rect 21833 54689 21867 54723
rect 21925 54689 21959 54723
rect 22753 54689 22787 54723
rect 23765 54689 23799 54723
rect 27445 54689 27479 54723
rect 16037 54621 16071 54655
rect 17693 54621 17727 54655
rect 17877 54621 17911 54655
rect 18613 54621 18647 54655
rect 21005 54621 21039 54655
rect 22937 54621 22971 54655
rect 23857 54621 23891 54655
rect 26617 54621 26651 54655
rect 26709 54621 26743 54655
rect 27537 54621 27571 54655
rect 13001 54553 13035 54587
rect 13369 54553 13403 54587
rect 14381 54553 14415 54587
rect 15393 54553 15427 54587
rect 15945 54553 15979 54587
rect 18889 54553 18923 54587
rect 12357 54485 12391 54519
rect 13737 54485 13771 54519
rect 15485 54485 15519 54519
rect 15807 54485 15841 54519
rect 16313 54485 16347 54519
rect 20361 54485 20395 54519
rect 26249 54485 26283 54519
rect 12265 54281 12299 54315
rect 15853 54281 15887 54315
rect 16589 54281 16623 54315
rect 18521 54281 18555 54315
rect 19533 54281 19567 54315
rect 20913 54281 20947 54315
rect 27905 54281 27939 54315
rect 13185 54213 13219 54247
rect 16037 54213 16071 54247
rect 22017 54213 22051 54247
rect 11897 54145 11931 54179
rect 12909 54145 12943 54179
rect 15945 54145 15979 54179
rect 17141 54145 17175 54179
rect 18061 54145 18095 54179
rect 25881 54145 25915 54179
rect 26249 54145 26283 54179
rect 11345 54077 11379 54111
rect 13001 54077 13035 54111
rect 13461 54077 13495 54111
rect 14657 54077 14691 54111
rect 15724 54077 15758 54111
rect 18337 54077 18371 54111
rect 19809 54077 19843 54111
rect 21281 54077 21315 54111
rect 22201 54077 22235 54111
rect 22523 54077 22557 54111
rect 22661 54077 22695 54111
rect 23029 54077 23063 54111
rect 23673 54077 23707 54111
rect 24133 54077 24167 54111
rect 24685 54077 24719 54111
rect 25973 54077 26007 54111
rect 14013 54009 14047 54043
rect 15025 54009 15059 54043
rect 15393 54009 15427 54043
rect 15577 54009 15611 54043
rect 18245 54009 18279 54043
rect 20453 54009 20487 54043
rect 21649 54009 21683 54043
rect 11529 53941 11563 53975
rect 13829 53941 13863 53975
rect 17417 53941 17451 53975
rect 17785 53941 17819 53975
rect 19073 53941 19107 53975
rect 23489 53941 23523 53975
rect 23765 53941 23799 53975
rect 27353 53941 27387 53975
rect 11805 53737 11839 53771
rect 18061 53737 18095 53771
rect 20269 53737 20303 53771
rect 20729 53737 20763 53771
rect 21925 53737 21959 53771
rect 22385 53737 22419 53771
rect 26709 53737 26743 53771
rect 13921 53669 13955 53703
rect 16957 53669 16991 53703
rect 19257 53669 19291 53703
rect 27077 53669 27111 53703
rect 11253 53601 11287 53635
rect 12541 53601 12575 53635
rect 16221 53601 16255 53635
rect 18061 53601 18095 53635
rect 18245 53601 18279 53635
rect 18613 53601 18647 53635
rect 19533 53601 19567 53635
rect 19717 53601 19751 53635
rect 20913 53601 20947 53635
rect 21005 53601 21039 53635
rect 21189 53601 21223 53635
rect 22937 53601 22971 53635
rect 23121 53601 23155 53635
rect 23949 53601 23983 53635
rect 24041 53601 24075 53635
rect 12265 53533 12299 53567
rect 16589 53533 16623 53567
rect 17601 53533 17635 53567
rect 21373 53533 21407 53567
rect 23213 53533 23247 53567
rect 25973 53533 26007 53567
rect 16037 53465 16071 53499
rect 16359 53465 16393 53499
rect 19901 53465 19935 53499
rect 11437 53397 11471 53431
rect 12081 53397 12115 53431
rect 14289 53397 14323 53431
rect 14657 53397 14691 53431
rect 15025 53397 15059 53431
rect 15669 53397 15703 53431
rect 16497 53397 16531 53431
rect 17325 53397 17359 53431
rect 24501 53397 24535 53431
rect 10517 53193 10551 53227
rect 10885 53193 10919 53227
rect 11897 53193 11931 53227
rect 14473 53193 14507 53227
rect 16221 53193 16255 53227
rect 16681 53193 16715 53227
rect 17049 53193 17083 53227
rect 21465 53193 21499 53227
rect 23121 53193 23155 53227
rect 23489 53193 23523 53227
rect 17877 53125 17911 53159
rect 12449 53057 12483 53091
rect 18061 53057 18095 53091
rect 20637 53057 20671 53091
rect 24133 53057 24167 53091
rect 24501 53057 24535 53091
rect 11345 52989 11379 53023
rect 12725 52989 12759 53023
rect 15025 52989 15059 53023
rect 16497 52989 16531 53023
rect 18337 52989 18371 53023
rect 18797 52989 18831 53023
rect 19717 52989 19751 53023
rect 20085 52989 20119 53023
rect 20545 52989 20579 53023
rect 21649 52989 21683 53023
rect 21741 52989 21775 53023
rect 24225 52989 24259 53023
rect 11253 52921 11287 52955
rect 18429 52921 18463 52955
rect 21097 52921 21131 52955
rect 22201 52921 22235 52955
rect 11529 52853 11563 52887
rect 12173 52853 12207 52887
rect 14013 52853 14047 52887
rect 14841 52853 14875 52887
rect 15209 52853 15243 52887
rect 17417 52853 17451 52887
rect 18245 52853 18279 52887
rect 19165 52853 19199 52887
rect 19625 52853 19659 52887
rect 22477 52853 22511 52887
rect 25605 52853 25639 52887
rect 10793 52649 10827 52683
rect 11805 52649 11839 52683
rect 13829 52649 13863 52683
rect 16497 52649 16531 52683
rect 18153 52649 18187 52683
rect 19165 52649 19199 52683
rect 19717 52649 19751 52683
rect 20085 52649 20119 52683
rect 21005 52649 21039 52683
rect 22845 52649 22879 52683
rect 11529 52581 11563 52615
rect 13185 52581 13219 52615
rect 14013 52581 14047 52615
rect 14381 52581 14415 52615
rect 14749 52581 14783 52615
rect 15025 52581 15059 52615
rect 22293 52581 22327 52615
rect 1685 52513 1719 52547
rect 3065 52513 3099 52547
rect 10609 52513 10643 52547
rect 11621 52513 11655 52547
rect 12633 52513 12667 52547
rect 13553 52513 13587 52547
rect 13921 52513 13955 52547
rect 15945 52513 15979 52547
rect 16865 52513 16899 52547
rect 17049 52513 17083 52547
rect 18245 52513 18279 52547
rect 18705 52513 18739 52547
rect 19073 52513 19107 52547
rect 21097 52513 21131 52547
rect 21465 52513 21499 52547
rect 23305 52513 23339 52547
rect 23857 52513 23891 52547
rect 1409 52445 1443 52479
rect 12449 52445 12483 52479
rect 13645 52445 13679 52479
rect 15301 52445 15335 52479
rect 17325 52445 17359 52479
rect 21741 52445 21775 52479
rect 23121 52445 23155 52479
rect 23765 52377 23799 52411
rect 12081 52309 12115 52343
rect 12817 52309 12851 52343
rect 17693 52309 17727 52343
rect 20361 52309 20395 52343
rect 24317 52309 24351 52343
rect 1685 52105 1719 52139
rect 8401 52105 8435 52139
rect 10885 52105 10919 52139
rect 11253 52105 11287 52139
rect 11897 52105 11931 52139
rect 12265 52105 12299 52139
rect 14841 52105 14875 52139
rect 15209 52105 15243 52139
rect 18337 52105 18371 52139
rect 20269 52105 20303 52139
rect 21833 52105 21867 52139
rect 22569 52105 22603 52139
rect 23305 52105 23339 52139
rect 25053 52105 25087 52139
rect 17049 52037 17083 52071
rect 19257 52037 19291 52071
rect 14197 51969 14231 52003
rect 15301 51969 15335 52003
rect 17509 51969 17543 52003
rect 19165 51969 19199 52003
rect 19901 51969 19935 52003
rect 23029 51969 23063 52003
rect 24409 51969 24443 52003
rect 8033 51901 8067 51935
rect 10333 51901 10367 51935
rect 11345 51901 11379 51935
rect 12817 51901 12851 51935
rect 13093 51901 13127 51935
rect 15393 51901 15427 51935
rect 16865 51901 16899 51935
rect 17877 51901 17911 51935
rect 18521 51901 18555 51935
rect 19257 51901 19291 51935
rect 20361 51901 20395 51935
rect 21005 51901 21039 51935
rect 21097 51901 21131 51935
rect 21373 51901 21407 51935
rect 21557 51901 21591 51935
rect 22385 51901 22419 51935
rect 24685 51901 24719 51935
rect 16773 51833 16807 51867
rect 23673 51833 23707 51867
rect 23857 51833 23891 51867
rect 24041 51833 24075 51867
rect 1961 51765 1995 51799
rect 7849 51765 7883 51799
rect 10517 51765 10551 51799
rect 11529 51765 11563 51799
rect 12633 51765 12667 51799
rect 16313 51765 16347 51799
rect 22201 51765 22235 51799
rect 23949 51765 23983 51799
rect 10425 51561 10459 51595
rect 11069 51561 11103 51595
rect 11529 51561 11563 51595
rect 13093 51561 13127 51595
rect 14841 51561 14875 51595
rect 16681 51561 16715 51595
rect 17877 51561 17911 51595
rect 19073 51561 19107 51595
rect 20453 51561 20487 51595
rect 24501 51561 24535 51595
rect 12173 51493 12207 51527
rect 13645 51493 13679 51527
rect 15945 51493 15979 51527
rect 6101 51425 6135 51459
rect 10609 51425 10643 51459
rect 11621 51425 11655 51459
rect 12633 51425 12667 51459
rect 13792 51425 13826 51459
rect 15117 51425 15151 51459
rect 16037 51425 16071 51459
rect 16184 51425 16218 51459
rect 17509 51425 17543 51459
rect 17785 51425 17819 51459
rect 18061 51425 18095 51459
rect 18429 51425 18463 51459
rect 19533 51425 19567 51459
rect 20085 51425 20119 51459
rect 21557 51425 21591 51459
rect 21925 51425 21959 51459
rect 22017 51425 22051 51459
rect 22385 51425 22419 51459
rect 23029 51425 23063 51459
rect 23213 51425 23247 51459
rect 24041 51425 24075 51459
rect 24225 51425 24259 51459
rect 12541 51357 12575 51391
rect 14013 51357 14047 51391
rect 13553 51289 13587 51323
rect 13921 51289 13955 51323
rect 16405 51357 16439 51391
rect 21465 51357 21499 51391
rect 23765 51357 23799 51391
rect 19717 51289 19751 51323
rect 5917 51221 5951 51255
rect 11805 51221 11839 51255
rect 12817 51221 12851 51255
rect 14289 51221 14323 51255
rect 15117 51221 15151 51255
rect 15485 51221 15519 51255
rect 16313 51221 16347 51255
rect 17141 51221 17175 51255
rect 19441 51221 19475 51255
rect 21005 51221 21039 51255
rect 24961 51221 24995 51255
rect 6009 51017 6043 51051
rect 10425 51017 10459 51051
rect 11253 51017 11287 51051
rect 12265 51017 12299 51051
rect 14289 51017 14323 51051
rect 14749 51017 14783 51051
rect 14979 51017 15013 51051
rect 18337 51017 18371 51051
rect 22201 51017 22235 51051
rect 22937 51017 22971 51051
rect 24317 51017 24351 51051
rect 11529 50949 11563 50983
rect 15117 50949 15151 50983
rect 16405 50949 16439 50983
rect 23305 50949 23339 50983
rect 13277 50881 13311 50915
rect 15209 50881 15243 50915
rect 15853 50881 15887 50915
rect 16221 50881 16255 50915
rect 17141 50881 17175 50915
rect 20361 50881 20395 50915
rect 20913 50881 20947 50915
rect 21925 50881 21959 50915
rect 24409 50881 24443 50915
rect 11345 50813 11379 50847
rect 11805 50813 11839 50847
rect 12817 50813 12851 50847
rect 13553 50813 13587 50847
rect 14841 50813 14875 50847
rect 16589 50813 16623 50847
rect 16681 50813 16715 50847
rect 19441 50813 19475 50847
rect 19717 50813 19751 50847
rect 19901 50813 19935 50847
rect 13461 50745 13495 50779
rect 13645 50745 13679 50779
rect 14013 50745 14047 50779
rect 17417 50745 17451 50779
rect 17785 50745 17819 50779
rect 18889 50745 18923 50779
rect 21373 50813 21407 50847
rect 23765 50813 23799 50847
rect 24685 50813 24719 50847
rect 21005 50745 21039 50779
rect 21189 50745 21223 50779
rect 21557 50745 21591 50779
rect 13185 50677 13219 50711
rect 15485 50677 15519 50711
rect 18797 50677 18831 50711
rect 20637 50677 20671 50711
rect 20913 50677 20947 50711
rect 21465 50677 21499 50711
rect 23765 50677 23799 50711
rect 23949 50677 23983 50711
rect 25789 50677 25823 50711
rect 12633 50473 12667 50507
rect 13001 50473 13035 50507
rect 13369 50473 13403 50507
rect 14841 50473 14875 50507
rect 16497 50473 16531 50507
rect 16865 50473 16899 50507
rect 18521 50473 18555 50507
rect 20361 50473 20395 50507
rect 20729 50473 20763 50507
rect 21189 50473 21223 50507
rect 23489 50473 23523 50507
rect 24317 50473 24351 50507
rect 16221 50405 16255 50439
rect 17417 50405 17451 50439
rect 17785 50405 17819 50439
rect 22477 50405 22511 50439
rect 22845 50405 22879 50439
rect 23213 50405 23247 50439
rect 10425 50337 10459 50371
rect 13921 50337 13955 50371
rect 14197 50337 14231 50371
rect 15669 50337 15703 50371
rect 15761 50337 15795 50371
rect 17233 50337 17267 50371
rect 17325 50337 17359 50371
rect 18981 50337 19015 50371
rect 19441 50337 19475 50371
rect 21557 50337 21591 50371
rect 22661 50337 22695 50371
rect 22753 50337 22787 50371
rect 24317 50337 24351 50371
rect 10701 50269 10735 50303
rect 14381 50269 14415 50303
rect 17049 50269 17083 50303
rect 18797 50269 18831 50303
rect 19717 50269 19751 50303
rect 11805 50133 11839 50167
rect 15485 50133 15519 50167
rect 18153 50133 18187 50167
rect 21925 50133 21959 50167
rect 22293 50133 22327 50167
rect 8953 49929 8987 49963
rect 9873 49929 9907 49963
rect 12265 49929 12299 49963
rect 12909 49929 12943 49963
rect 15393 49929 15427 49963
rect 17509 49929 17543 49963
rect 17877 49929 17911 49963
rect 18429 49929 18463 49963
rect 20269 49929 20303 49963
rect 22201 49929 22235 49963
rect 22477 49929 22511 49963
rect 22845 49929 22879 49963
rect 23489 49929 23523 49963
rect 10241 49861 10275 49895
rect 16405 49861 16439 49895
rect 17049 49861 17083 49895
rect 25421 49861 25455 49895
rect 7389 49793 7423 49827
rect 10333 49793 10367 49827
rect 11253 49793 11287 49827
rect 13001 49793 13035 49827
rect 13277 49793 13311 49827
rect 14381 49793 14415 49827
rect 24409 49793 24443 49827
rect 7665 49725 7699 49759
rect 10793 49725 10827 49759
rect 11161 49725 11195 49759
rect 14933 49725 14967 49759
rect 15485 49725 15519 49759
rect 16037 49725 16071 49759
rect 16405 49725 16439 49759
rect 18705 49725 18739 49759
rect 18981 49725 19015 49759
rect 19441 49725 19475 49759
rect 20545 49725 20579 49759
rect 21281 49725 21315 49759
rect 23765 49725 23799 49759
rect 24685 49725 24719 49759
rect 25237 49725 25271 49759
rect 19625 49657 19659 49691
rect 20913 49657 20947 49691
rect 21097 49657 21131 49691
rect 21465 49657 21499 49691
rect 21833 49657 21867 49691
rect 7205 49589 7239 49623
rect 11805 49589 11839 49623
rect 21373 49589 21407 49623
rect 25697 49589 25731 49623
rect 7389 49385 7423 49419
rect 10793 49385 10827 49419
rect 12633 49385 12667 49419
rect 14749 49385 14783 49419
rect 16497 49385 16531 49419
rect 17785 49385 17819 49419
rect 18153 49385 18187 49419
rect 19993 49385 20027 49419
rect 21373 49385 21407 49419
rect 15025 49317 15059 49351
rect 15853 49317 15887 49351
rect 16221 49317 16255 49351
rect 21557 49317 21591 49351
rect 11437 49249 11471 49283
rect 13001 49249 13035 49283
rect 15393 49249 15427 49283
rect 16681 49249 16715 49283
rect 16865 49249 16899 49283
rect 17233 49249 17267 49283
rect 18889 49249 18923 49283
rect 19165 49249 19199 49283
rect 19625 49249 19659 49283
rect 20913 49249 20947 49283
rect 11345 49181 11379 49215
rect 12725 49181 12759 49215
rect 18337 49181 18371 49215
rect 19349 49181 19383 49215
rect 22385 49249 22419 49283
rect 22569 49249 22603 49283
rect 22753 49249 22787 49283
rect 23673 49249 23707 49283
rect 24777 49249 24811 49283
rect 10425 49113 10459 49147
rect 21097 49113 21131 49147
rect 21557 49113 21591 49147
rect 21741 49113 21775 49147
rect 22201 49113 22235 49147
rect 11161 49045 11195 49079
rect 11621 49045 11655 49079
rect 14105 49045 14139 49079
rect 15577 49045 15611 49079
rect 20637 49045 20671 49079
rect 23213 49045 23247 49079
rect 23949 49045 23983 49079
rect 24409 49045 24443 49079
rect 11805 48841 11839 48875
rect 12265 48841 12299 48875
rect 13093 48841 13127 48875
rect 13553 48841 13587 48875
rect 16037 48841 16071 48875
rect 17877 48841 17911 48875
rect 19441 48841 19475 48875
rect 21097 48841 21131 48875
rect 22937 48841 22971 48875
rect 24777 48841 24811 48875
rect 25421 48841 25455 48875
rect 15485 48773 15519 48807
rect 16497 48773 16531 48807
rect 21465 48773 21499 48807
rect 14197 48705 14231 48739
rect 16773 48705 16807 48739
rect 19993 48705 20027 48739
rect 20729 48705 20763 48739
rect 22661 48705 22695 48739
rect 23673 48705 23707 48739
rect 12633 48637 12667 48671
rect 13645 48637 13679 48671
rect 14565 48637 14599 48671
rect 14657 48637 14691 48671
rect 15025 48637 15059 48671
rect 15577 48637 15611 48671
rect 16957 48637 16991 48671
rect 18061 48637 18095 48671
rect 18889 48637 18923 48671
rect 19073 48637 19107 48671
rect 20269 48637 20303 48671
rect 22201 48637 22235 48671
rect 22477 48637 22511 48671
rect 23489 48637 23523 48671
rect 23765 48637 23799 48671
rect 25237 48637 25271 48671
rect 25697 48637 25731 48671
rect 20177 48569 20211 48603
rect 20361 48569 20395 48603
rect 21833 48569 21867 48603
rect 11437 48501 11471 48535
rect 12817 48501 12851 48535
rect 13829 48501 13863 48535
rect 17141 48501 17175 48535
rect 17509 48501 17543 48535
rect 18337 48501 18371 48535
rect 19809 48501 19843 48535
rect 12449 48297 12483 48331
rect 13277 48297 13311 48331
rect 14749 48297 14783 48331
rect 17509 48297 17543 48331
rect 20269 48297 20303 48331
rect 21189 48297 21223 48331
rect 12909 48229 12943 48263
rect 13369 48229 13403 48263
rect 16957 48229 16991 48263
rect 18889 48229 18923 48263
rect 20177 48229 20211 48263
rect 22385 48229 22419 48263
rect 25145 48229 25179 48263
rect 14197 48161 14231 48195
rect 16129 48161 16163 48195
rect 16405 48161 16439 48195
rect 17693 48161 17727 48195
rect 18061 48161 18095 48195
rect 18245 48161 18279 48195
rect 19533 48161 19567 48195
rect 13921 48093 13955 48127
rect 14381 48093 14415 48127
rect 15577 48093 15611 48127
rect 16589 48093 16623 48127
rect 17233 48093 17267 48127
rect 19441 48093 19475 48127
rect 19993 48093 20027 48127
rect 15025 48025 15059 48059
rect 20913 48161 20947 48195
rect 21097 48161 21131 48195
rect 21265 48161 21299 48195
rect 22661 48161 22695 48195
rect 22845 48161 22879 48195
rect 23673 48161 23707 48195
rect 24133 48161 24167 48195
rect 24501 48161 24535 48195
rect 24685 48161 24719 48195
rect 21649 48093 21683 48127
rect 22937 48093 22971 48127
rect 23765 48093 23799 48127
rect 20729 48025 20763 48059
rect 19165 47957 19199 47991
rect 20177 47957 20211 47991
rect 21925 47957 21959 47991
rect 22477 47957 22511 47991
rect 24869 47957 24903 47991
rect 26249 47957 26283 47991
rect 8033 47753 8067 47787
rect 13093 47753 13127 47787
rect 13461 47753 13495 47787
rect 14289 47753 14323 47787
rect 14657 47753 14691 47787
rect 15301 47753 15335 47787
rect 16865 47753 16899 47787
rect 17417 47753 17451 47787
rect 19809 47753 19843 47787
rect 20177 47753 20211 47787
rect 23121 47753 23155 47787
rect 24961 47753 24995 47787
rect 27721 47753 27755 47787
rect 12725 47685 12759 47719
rect 8493 47617 8527 47651
rect 13829 47617 13863 47651
rect 15577 47617 15611 47651
rect 16497 47617 16531 47651
rect 18337 47617 18371 47651
rect 19533 47617 19567 47651
rect 22845 47617 22879 47651
rect 24685 47617 24719 47651
rect 26157 47617 26191 47651
rect 8217 47549 8251 47583
rect 14473 47549 14507 47583
rect 16037 47549 16071 47583
rect 16313 47549 16347 47583
rect 17601 47549 17635 47583
rect 18613 47549 18647 47583
rect 18981 47549 19015 47583
rect 19257 47549 19291 47583
rect 20453 47549 20487 47583
rect 20913 47549 20947 47583
rect 21373 47549 21407 47583
rect 21465 47549 21499 47583
rect 21925 47549 21959 47583
rect 23489 47549 23523 47583
rect 24225 47549 24259 47583
rect 24501 47549 24535 47583
rect 25421 47549 25455 47583
rect 26433 47549 26467 47583
rect 17233 47481 17267 47515
rect 23673 47481 23707 47515
rect 9781 47413 9815 47447
rect 12173 47413 12207 47447
rect 15025 47413 15059 47447
rect 20637 47413 20671 47447
rect 21557 47413 21591 47447
rect 23305 47413 23339 47447
rect 25973 47413 26007 47447
rect 8217 47209 8251 47243
rect 13737 47209 13771 47243
rect 14013 47209 14047 47243
rect 14381 47209 14415 47243
rect 14749 47209 14783 47243
rect 16957 47209 16991 47243
rect 20729 47209 20763 47243
rect 22385 47209 22419 47243
rect 23765 47209 23799 47243
rect 24133 47209 24167 47243
rect 26709 47209 26743 47243
rect 15117 47141 15151 47175
rect 17233 47141 17267 47175
rect 18153 47141 18187 47175
rect 20913 47141 20947 47175
rect 22477 47141 22511 47175
rect 12541 47073 12575 47107
rect 13277 47073 13311 47107
rect 14197 47073 14231 47107
rect 15669 47073 15703 47107
rect 16221 47073 16255 47107
rect 17417 47073 17451 47107
rect 18981 47073 19015 47107
rect 19257 47073 19291 47107
rect 20177 47073 20211 47107
rect 21005 47073 21039 47107
rect 22937 47073 22971 47107
rect 23121 47073 23155 47107
rect 23305 47073 23339 47107
rect 24501 47073 24535 47107
rect 25329 47073 25363 47107
rect 26525 47073 26559 47107
rect 12633 47005 12667 47039
rect 15393 47005 15427 47039
rect 18521 47005 18555 47039
rect 24593 47005 24627 47039
rect 25421 47005 25455 47039
rect 16129 46937 16163 46971
rect 17601 46937 17635 46971
rect 19257 46937 19291 46971
rect 25789 46937 25823 46971
rect 19901 46869 19935 46903
rect 22017 46869 22051 46903
rect 26157 46869 26191 46903
rect 13553 46665 13587 46699
rect 14473 46665 14507 46699
rect 14933 46665 14967 46699
rect 15209 46665 15243 46699
rect 17417 46665 17451 46699
rect 17877 46665 17911 46699
rect 26801 46665 26835 46699
rect 12541 46597 12575 46631
rect 19625 46597 19659 46631
rect 21557 46597 21591 46631
rect 21833 46597 21867 46631
rect 23397 46597 23431 46631
rect 27169 46597 27203 46631
rect 15853 46529 15887 46563
rect 18061 46529 18095 46563
rect 18797 46529 18831 46563
rect 19717 46529 19751 46563
rect 20269 46529 20303 46563
rect 20729 46529 20763 46563
rect 24225 46529 24259 46563
rect 12265 46461 12299 46495
rect 12449 46461 12483 46495
rect 12725 46461 12759 46495
rect 15025 46461 15059 46495
rect 16221 46461 16255 46495
rect 16405 46461 16439 46495
rect 16865 46461 16899 46495
rect 18337 46461 18371 46495
rect 20545 46461 20579 46495
rect 21741 46461 21775 46495
rect 21833 46461 21867 46495
rect 22201 46461 22235 46495
rect 23765 46461 23799 46495
rect 24409 46461 24443 46495
rect 24869 46461 24903 46495
rect 25421 46461 25455 46495
rect 25973 46461 26007 46495
rect 26065 46461 26099 46495
rect 17141 46393 17175 46427
rect 18245 46393 18279 46427
rect 21005 46393 21039 46427
rect 22017 46393 22051 46427
rect 22385 46393 22419 46427
rect 22753 46393 22787 46427
rect 25145 46393 25179 46427
rect 26525 46393 26559 46427
rect 11897 46325 11931 46359
rect 12909 46325 12943 46359
rect 14197 46325 14231 46359
rect 15577 46325 15611 46359
rect 19165 46325 19199 46359
rect 21373 46325 21407 46359
rect 22293 46325 22327 46359
rect 23029 46325 23063 46359
rect 23765 46325 23799 46359
rect 23857 46325 23891 46359
rect 25881 46325 25915 46359
rect 11897 46121 11931 46155
rect 12265 46121 12299 46155
rect 15025 46121 15059 46155
rect 16681 46121 16715 46155
rect 17509 46121 17543 46155
rect 18705 46121 18739 46155
rect 19717 46121 19751 46155
rect 24133 46121 24167 46155
rect 24593 46121 24627 46155
rect 25973 46121 26007 46155
rect 20637 46053 20671 46087
rect 25605 46053 25639 46087
rect 12449 45985 12483 46019
rect 12725 45985 12759 46019
rect 15485 45985 15519 46019
rect 15669 45985 15703 46019
rect 16129 45985 16163 46019
rect 17233 45985 17267 46019
rect 17693 45985 17727 46019
rect 19257 45985 19291 46019
rect 19533 45985 19567 46019
rect 20913 45985 20947 46019
rect 21097 45985 21131 46019
rect 22937 45985 22971 46019
rect 23305 45985 23339 46019
rect 23397 45985 23431 46019
rect 24317 45985 24351 46019
rect 24869 45985 24903 46019
rect 13185 45917 13219 45951
rect 19165 45917 19199 45951
rect 19349 45917 19383 45951
rect 12541 45849 12575 45883
rect 16129 45849 16163 45883
rect 17049 45849 17083 45883
rect 22753 45849 22787 45883
rect 1593 45781 1627 45815
rect 14473 45781 14507 45815
rect 18337 45781 18371 45815
rect 20269 45781 20303 45815
rect 22017 45781 22051 45815
rect 12541 45577 12575 45611
rect 14933 45577 14967 45611
rect 15485 45577 15519 45611
rect 19717 45577 19751 45611
rect 21373 45577 21407 45611
rect 23029 45577 23063 45611
rect 25053 45577 25087 45611
rect 11253 45509 11287 45543
rect 16497 45509 16531 45543
rect 17141 45509 17175 45543
rect 17877 45509 17911 45543
rect 18153 45509 18187 45543
rect 1409 45441 1443 45475
rect 1685 45441 1719 45475
rect 14013 45441 14047 45475
rect 14381 45441 14415 45475
rect 18797 45441 18831 45475
rect 23489 45441 23523 45475
rect 23765 45441 23799 45475
rect 11345 45373 11379 45407
rect 11897 45373 11931 45407
rect 12541 45373 12575 45407
rect 12817 45373 12851 45407
rect 13461 45373 13495 45407
rect 14473 45373 14507 45407
rect 14749 45373 14783 45407
rect 15945 45373 15979 45407
rect 16865 45373 16899 45407
rect 16957 45373 16991 45407
rect 18061 45373 18095 45407
rect 18337 45373 18371 45407
rect 19625 45373 19659 45407
rect 19993 45373 20027 45407
rect 20361 45373 20395 45407
rect 20913 45373 20947 45407
rect 21925 45373 21959 45407
rect 22385 45373 22419 45407
rect 24593 45373 24627 45407
rect 24685 45373 24719 45407
rect 25881 45373 25915 45407
rect 26985 45373 27019 45407
rect 27353 45373 27387 45407
rect 3065 45305 3099 45339
rect 12265 45305 12299 45339
rect 14657 45305 14691 45339
rect 17509 45305 17543 45339
rect 22661 45305 22695 45339
rect 23857 45305 23891 45339
rect 25421 45305 25455 45339
rect 25605 45305 25639 45339
rect 25973 45305 26007 45339
rect 26341 45305 26375 45339
rect 11529 45237 11563 45271
rect 19349 45237 19383 45271
rect 21741 45237 21775 45271
rect 25789 45237 25823 45271
rect 26617 45237 26651 45271
rect 1685 45033 1719 45067
rect 1961 45033 1995 45067
rect 12541 45033 12575 45067
rect 14565 45033 14599 45067
rect 15577 45033 15611 45067
rect 16037 45033 16071 45067
rect 16865 45033 16899 45067
rect 17233 45033 17267 45067
rect 18153 45033 18187 45067
rect 18797 45033 18831 45067
rect 23305 45033 23339 45067
rect 23673 45033 23707 45067
rect 24869 45033 24903 45067
rect 25605 45033 25639 45067
rect 26709 45033 26743 45067
rect 13645 44965 13679 44999
rect 19165 44965 19199 44999
rect 21833 44965 21867 44999
rect 25237 44965 25271 44999
rect 26249 44965 26283 44999
rect 26893 44965 26927 44999
rect 11805 44897 11839 44931
rect 13461 44897 13495 44931
rect 16681 44897 16715 44931
rect 17693 44897 17727 44931
rect 17969 44897 18003 44931
rect 19257 44897 19291 44931
rect 22477 44897 22511 44931
rect 22845 44897 22879 44931
rect 23949 44897 23983 44931
rect 25421 44897 25455 44931
rect 25973 44897 26007 44931
rect 26801 44897 26835 44931
rect 11897 44829 11931 44863
rect 19625 44829 19659 44863
rect 19717 44829 19751 44863
rect 20637 44829 20671 44863
rect 21189 44829 21223 44863
rect 22385 44829 22419 44863
rect 22937 44829 22971 44863
rect 23857 44829 23891 44863
rect 26525 44829 26559 44863
rect 27261 44829 27295 44863
rect 16589 44761 16623 44795
rect 17785 44761 17819 44795
rect 19533 44761 19567 44795
rect 2329 44693 2363 44727
rect 19395 44693 19429 44727
rect 20269 44693 20303 44727
rect 21741 44693 21775 44727
rect 27537 44693 27571 44727
rect 2973 44489 3007 44523
rect 14197 44489 14231 44523
rect 15761 44489 15795 44523
rect 19717 44489 19751 44523
rect 21649 44489 21683 44523
rect 23121 44489 23155 44523
rect 25605 44489 25639 44523
rect 12265 44421 12299 44455
rect 12725 44421 12759 44455
rect 17141 44421 17175 44455
rect 1409 44353 1443 44387
rect 12817 44353 12851 44387
rect 16773 44353 16807 44387
rect 18613 44353 18647 44387
rect 19993 44353 20027 44387
rect 20177 44353 20211 44387
rect 24869 44353 24903 44387
rect 25237 44353 25271 44387
rect 26065 44353 26099 44387
rect 26433 44353 26467 44387
rect 1685 44285 1719 44319
rect 10241 44285 10275 44319
rect 10977 44285 11011 44319
rect 12596 44285 12630 44319
rect 14013 44285 14047 44319
rect 14473 44285 14507 44319
rect 15945 44285 15979 44319
rect 16957 44285 16991 44319
rect 18521 44285 18555 44319
rect 19257 44285 19291 44319
rect 20361 44285 20395 44319
rect 20913 44285 20947 44319
rect 21281 44285 21315 44319
rect 22201 44285 22235 44319
rect 22385 44285 22419 44319
rect 22569 44285 22603 44319
rect 23949 44285 23983 44319
rect 24777 44285 24811 44319
rect 26157 44285 26191 44319
rect 28089 44285 28123 44319
rect 11897 44217 11931 44251
rect 12449 44217 12483 44251
rect 20545 44217 20579 44251
rect 21741 44217 21775 44251
rect 24041 44217 24075 44251
rect 10793 44149 10827 44183
rect 11437 44149 11471 44183
rect 13093 44149 13127 44183
rect 13461 44149 13495 44183
rect 13921 44149 13955 44183
rect 16129 44149 16163 44183
rect 17509 44149 17543 44183
rect 17785 44149 17819 44183
rect 20453 44149 20487 44183
rect 23489 44149 23523 44183
rect 27721 44149 27755 44183
rect 17141 43945 17175 43979
rect 19073 43945 19107 43979
rect 19717 43945 19751 43979
rect 21281 43945 21315 43979
rect 23857 43945 23891 43979
rect 25881 43945 25915 43979
rect 26709 43945 26743 43979
rect 26801 43945 26835 43979
rect 16865 43877 16899 43911
rect 26525 43877 26559 43911
rect 26893 43877 26927 43911
rect 1501 43809 1535 43843
rect 7849 43809 7883 43843
rect 8585 43809 8619 43843
rect 8677 43809 8711 43843
rect 11805 43809 11839 43843
rect 12081 43809 12115 43843
rect 13093 43809 13127 43843
rect 16313 43809 16347 43843
rect 16405 43809 16439 43843
rect 17693 43809 17727 43843
rect 17785 43809 17819 43843
rect 17969 43809 18003 43843
rect 19901 43809 19935 43843
rect 21097 43809 21131 43843
rect 22569 43809 22603 43843
rect 22753 43809 22787 43843
rect 22937 43809 22971 43843
rect 26341 43809 26375 43843
rect 1777 43741 1811 43775
rect 3157 43741 3191 43775
rect 7757 43741 7791 43775
rect 11253 43741 11287 43775
rect 12265 43741 12299 43775
rect 12633 43741 12667 43775
rect 18429 43741 18463 43775
rect 23949 43741 23983 43775
rect 24225 43741 24259 43775
rect 25605 43741 25639 43775
rect 27261 43741 27295 43775
rect 13001 43673 13035 43707
rect 16129 43673 16163 43707
rect 22385 43673 22419 43707
rect 13277 43605 13311 43639
rect 17601 43605 17635 43639
rect 18705 43605 18739 43639
rect 20545 43605 20579 43639
rect 21833 43605 21867 43639
rect 23489 43605 23523 43639
rect 27537 43605 27571 43639
rect 7757 43401 7791 43435
rect 8493 43401 8527 43435
rect 11345 43401 11379 43435
rect 12817 43401 12851 43435
rect 16129 43401 16163 43435
rect 16589 43401 16623 43435
rect 17141 43401 17175 43435
rect 17693 43401 17727 43435
rect 19441 43401 19475 43435
rect 21833 43401 21867 43435
rect 22477 43401 22511 43435
rect 22753 43401 22787 43435
rect 23121 43401 23155 43435
rect 24041 43401 24075 43435
rect 25973 43401 26007 43435
rect 26525 43401 26559 43435
rect 26985 43401 27019 43435
rect 27353 43401 27387 43435
rect 8125 43333 8159 43367
rect 10977 43333 11011 43367
rect 15853 43333 15887 43367
rect 20085 43333 20119 43367
rect 1777 43265 1811 43299
rect 13829 43265 13863 43299
rect 18061 43265 18095 43299
rect 22293 43265 22327 43299
rect 1501 43197 1535 43231
rect 3157 43197 3191 43231
rect 10793 43197 10827 43231
rect 11713 43197 11747 43231
rect 12173 43197 12207 43231
rect 13001 43197 13035 43231
rect 13369 43197 13403 43231
rect 13737 43197 13771 43231
rect 16957 43197 16991 43231
rect 18337 43197 18371 43231
rect 21097 43197 21131 43231
rect 21373 43197 21407 43231
rect 21557 43197 21591 43231
rect 20361 43129 20395 43163
rect 20545 43129 20579 43163
rect 23489 43333 23523 43367
rect 28273 43333 28307 43367
rect 24501 43265 24535 43299
rect 27077 43265 27111 43299
rect 22569 43197 22603 43231
rect 24593 43197 24627 43231
rect 24869 43197 24903 43231
rect 27169 43197 27203 43231
rect 27905 43197 27939 43231
rect 10609 43061 10643 43095
rect 22477 43061 22511 43095
rect 1685 42857 1719 42891
rect 17049 42857 17083 42891
rect 17509 42857 17543 42891
rect 20637 42857 20671 42891
rect 27353 42857 27387 42891
rect 2329 42789 2363 42823
rect 11437 42789 11471 42823
rect 21649 42789 21683 42823
rect 11345 42721 11379 42755
rect 12081 42721 12115 42755
rect 12449 42721 12483 42755
rect 17601 42721 17635 42755
rect 19809 42721 19843 42755
rect 21557 42721 21591 42755
rect 22293 42721 22327 42755
rect 22661 42721 22695 42755
rect 22753 42721 22787 42755
rect 23949 42721 23983 42755
rect 24225 42721 24259 42755
rect 26525 42721 26559 42755
rect 26617 42721 26651 42755
rect 11989 42653 12023 42687
rect 12541 42653 12575 42687
rect 17877 42653 17911 42687
rect 21189 42653 21223 42687
rect 22385 42653 22419 42687
rect 25881 42653 25915 42687
rect 26249 42653 26283 42687
rect 20177 42585 20211 42619
rect 2053 42517 2087 42551
rect 8677 42517 8711 42551
rect 13001 42517 13035 42551
rect 18981 42517 19015 42551
rect 23121 42517 23155 42551
rect 23765 42517 23799 42551
rect 25329 42517 25363 42551
rect 26801 42517 26835 42551
rect 1593 42313 1627 42347
rect 10885 42313 10919 42347
rect 11897 42313 11931 42347
rect 12173 42313 12207 42347
rect 14473 42313 14507 42347
rect 17785 42313 17819 42347
rect 18337 42313 18371 42347
rect 21005 42313 21039 42347
rect 25053 42313 25087 42347
rect 17417 42245 17451 42279
rect 18889 42245 18923 42279
rect 19625 42245 19659 42279
rect 19993 42245 20027 42279
rect 23949 42245 23983 42279
rect 25605 42245 25639 42279
rect 25973 42245 26007 42279
rect 8493 42177 8527 42211
rect 14197 42177 14231 42211
rect 22569 42177 22603 42211
rect 26433 42177 26467 42211
rect 8769 42109 8803 42143
rect 8953 42109 8987 42143
rect 9229 42109 9263 42143
rect 9597 42109 9631 42143
rect 10057 42109 10091 42143
rect 10241 42109 10275 42143
rect 11345 42109 11379 42143
rect 14289 42109 14323 42143
rect 18705 42109 18739 42143
rect 19165 42109 19199 42143
rect 20177 42109 20211 42143
rect 20361 42109 20395 42143
rect 20545 42109 20579 42143
rect 21465 42109 21499 42143
rect 22109 42109 22143 42143
rect 22385 42109 22419 42143
rect 24133 42109 24167 42143
rect 24317 42109 24351 42143
rect 24501 42109 24535 42143
rect 26157 42109 26191 42143
rect 11253 42041 11287 42075
rect 15117 42041 15151 42075
rect 21557 42041 21591 42075
rect 23489 42041 23523 42075
rect 8125 41973 8159 42007
rect 11529 41973 11563 42007
rect 12633 41973 12667 42007
rect 14013 41973 14047 42007
rect 22937 41973 22971 42007
rect 27537 41973 27571 42007
rect 8677 41769 8711 41803
rect 17693 41769 17727 41803
rect 18153 41769 18187 41803
rect 19625 41769 19659 41803
rect 20361 41769 20395 41803
rect 21833 41769 21867 41803
rect 22201 41769 22235 41803
rect 24041 41769 24075 41803
rect 25697 41769 25731 41803
rect 26249 41769 26283 41803
rect 27537 41769 27571 41803
rect 10793 41701 10827 41735
rect 20729 41701 20763 41735
rect 21465 41701 21499 41735
rect 26525 41701 26559 41735
rect 11529 41633 11563 41667
rect 11897 41633 11931 41667
rect 19809 41633 19843 41667
rect 20913 41633 20947 41667
rect 21097 41633 21131 41667
rect 22569 41633 22603 41667
rect 23121 41633 23155 41667
rect 25145 41633 25179 41667
rect 27169 41633 27203 41667
rect 11437 41565 11471 41599
rect 11989 41565 12023 41599
rect 23213 41565 23247 41599
rect 24317 41565 24351 41599
rect 24409 41565 24443 41599
rect 25237 41565 25271 41599
rect 10425 41497 10459 41531
rect 19993 41497 20027 41531
rect 9045 41429 9079 41463
rect 10977 41429 11011 41463
rect 16129 41429 16163 41463
rect 23397 41429 23431 41463
rect 11805 41225 11839 41259
rect 19809 41225 19843 41259
rect 20085 41225 20119 41259
rect 22477 41225 22511 41259
rect 22845 41225 22879 41259
rect 26341 41225 26375 41259
rect 11161 41157 11195 41191
rect 16405 41157 16439 41191
rect 19533 41157 19567 41191
rect 20545 41157 20579 41191
rect 26801 41157 26835 41191
rect 9873 41089 9907 41123
rect 21189 41089 21223 41123
rect 22017 41089 22051 41123
rect 24685 41089 24719 41123
rect 10333 41021 10367 41055
rect 10701 41021 10735 41055
rect 11253 41021 11287 41055
rect 16589 41021 16623 41055
rect 16773 41021 16807 41055
rect 16957 41021 16991 41055
rect 19625 41021 19659 41055
rect 21097 41021 21131 41055
rect 21925 41021 21959 41055
rect 23765 41021 23799 41055
rect 24225 41021 24259 41055
rect 24777 41021 24811 41055
rect 25053 41021 25087 41055
rect 16037 40953 16071 40987
rect 20913 40953 20947 40987
rect 23489 40953 23523 40987
rect 10149 40885 10183 40919
rect 12081 40885 12115 40919
rect 12725 40885 12759 40919
rect 13093 40885 13127 40919
rect 23949 40885 23983 40919
rect 10885 40681 10919 40715
rect 20729 40681 20763 40715
rect 21557 40681 21591 40715
rect 21925 40681 21959 40715
rect 23397 40681 23431 40715
rect 25053 40681 25087 40715
rect 25513 40681 25547 40715
rect 22569 40613 22603 40647
rect 22845 40613 22879 40647
rect 10425 40545 10459 40579
rect 12081 40545 12115 40579
rect 12449 40545 12483 40579
rect 14013 40545 14047 40579
rect 16589 40545 16623 40579
rect 17049 40545 17083 40579
rect 21005 40545 21039 40579
rect 22017 40545 22051 40579
rect 22109 40545 22143 40579
rect 24225 40545 24259 40579
rect 24593 40545 24627 40579
rect 10057 40477 10091 40511
rect 11989 40477 12023 40511
rect 12541 40477 12575 40511
rect 16773 40477 16807 40511
rect 24133 40477 24167 40511
rect 24685 40477 24719 40511
rect 11345 40409 11379 40443
rect 16221 40409 16255 40443
rect 21189 40409 21223 40443
rect 1593 40341 1627 40375
rect 10609 40341 10643 40375
rect 11529 40341 11563 40375
rect 12909 40341 12943 40375
rect 13277 40341 13311 40375
rect 14197 40341 14231 40375
rect 15669 40341 15703 40375
rect 18153 40341 18187 40375
rect 23673 40341 23707 40375
rect 11805 40137 11839 40171
rect 15117 40137 15151 40171
rect 17601 40137 17635 40171
rect 22385 40137 22419 40171
rect 11897 40069 11931 40103
rect 12081 40069 12115 40103
rect 25421 40069 25455 40103
rect 1777 40001 1811 40035
rect 9965 40001 9999 40035
rect 11253 40001 11287 40035
rect 1501 39933 1535 39967
rect 9137 39933 9171 39967
rect 10517 39933 10551 39967
rect 10609 39933 10643 39967
rect 10885 39933 10919 39967
rect 11437 39933 11471 39967
rect 3157 39865 3191 39899
rect 9505 39865 9539 39899
rect 15945 40001 15979 40035
rect 25145 40001 25179 40035
rect 13369 39933 13403 39967
rect 15669 39933 15703 39967
rect 22017 39933 22051 39967
rect 23673 39933 23707 39967
rect 24225 39933 24259 39967
rect 25237 39933 25271 39967
rect 25697 39933 25731 39967
rect 13829 39865 13863 39899
rect 21097 39865 21131 39899
rect 23489 39865 23523 39899
rect 24409 39865 24443 39899
rect 9873 39797 9907 39831
rect 11897 39797 11931 39831
rect 12633 39797 12667 39831
rect 13645 39797 13679 39831
rect 17049 39797 17083 39831
rect 21833 39797 21867 39831
rect 23029 39797 23063 39831
rect 24685 39797 24719 39831
rect 1685 39593 1719 39627
rect 10517 39593 10551 39627
rect 16589 39593 16623 39627
rect 19441 39593 19475 39627
rect 21833 39593 21867 39627
rect 22385 39593 22419 39627
rect 24501 39593 24535 39627
rect 24777 39593 24811 39627
rect 11161 39525 11195 39559
rect 9505 39457 9539 39491
rect 11621 39457 11655 39491
rect 11805 39457 11839 39491
rect 11989 39457 12023 39491
rect 12909 39457 12943 39491
rect 13001 39457 13035 39491
rect 13553 39457 13587 39491
rect 13737 39457 13771 39491
rect 14749 39457 14783 39491
rect 15301 39457 15335 39491
rect 16773 39457 16807 39491
rect 21557 39457 21591 39491
rect 21741 39457 21775 39491
rect 23581 39457 23615 39491
rect 24593 39457 24627 39491
rect 12265 39389 12299 39423
rect 12541 39389 12575 39423
rect 14105 39389 14139 39423
rect 16681 39389 16715 39423
rect 17601 39389 17635 39423
rect 18061 39389 18095 39423
rect 18337 39389 18371 39423
rect 9137 39321 9171 39355
rect 10057 39253 10091 39287
rect 10793 39253 10827 39287
rect 12725 39253 12759 39287
rect 13185 39253 13219 39287
rect 14381 39253 14415 39287
rect 15485 39253 15519 39287
rect 15761 39253 15795 39287
rect 16221 39253 16255 39287
rect 16957 39253 16991 39287
rect 21465 39253 21499 39287
rect 23765 39253 23799 39287
rect 24041 39253 24075 39287
rect 3157 39049 3191 39083
rect 12909 39049 12943 39083
rect 15209 39049 15243 39083
rect 17049 39049 17083 39083
rect 19441 39049 19475 39083
rect 21189 39049 21223 39083
rect 23857 39049 23891 39083
rect 27537 39049 27571 39083
rect 10425 38981 10459 39015
rect 21557 38981 21591 39015
rect 21649 38981 21683 39015
rect 21833 38981 21867 39015
rect 1593 38913 1627 38947
rect 10149 38913 10183 38947
rect 11529 38913 11563 38947
rect 17877 38913 17911 38947
rect 1869 38845 1903 38879
rect 9597 38845 9631 38879
rect 9689 38845 9723 38879
rect 11161 38845 11195 38879
rect 12449 38845 12483 38879
rect 12633 38845 12667 38879
rect 12725 38845 12759 38879
rect 13553 38845 13587 38879
rect 13921 38845 13955 38879
rect 14013 38845 14047 38879
rect 14197 38845 14231 38879
rect 15393 38845 15427 38879
rect 17509 38845 17543 38879
rect 18061 38845 18095 38879
rect 18337 38845 18371 38879
rect 22845 38913 22879 38947
rect 26065 38913 26099 38947
rect 22017 38845 22051 38879
rect 22109 38845 22143 38879
rect 22569 38845 22603 38879
rect 26157 38845 26191 38879
rect 26433 38845 26467 38879
rect 9137 38777 9171 38811
rect 10977 38777 11011 38811
rect 11805 38777 11839 38811
rect 14565 38777 14599 38811
rect 16221 38777 16255 38811
rect 21649 38777 21683 38811
rect 8769 38709 8803 38743
rect 9505 38709 9539 38743
rect 10793 38709 10827 38743
rect 12173 38709 12207 38743
rect 14841 38709 14875 38743
rect 15577 38709 15611 38743
rect 15853 38709 15887 38743
rect 16773 38709 16807 38743
rect 24593 38709 24627 38743
rect 8769 38505 8803 38539
rect 9505 38505 9539 38539
rect 15577 38505 15611 38539
rect 16497 38505 16531 38539
rect 18153 38505 18187 38539
rect 20269 38505 20303 38539
rect 26157 38505 26191 38539
rect 8125 38437 8159 38471
rect 9689 38437 9723 38471
rect 12081 38437 12115 38471
rect 8585 38369 8619 38403
rect 10333 38369 10367 38403
rect 10701 38369 10735 38403
rect 10885 38369 10919 38403
rect 13185 38369 13219 38403
rect 14197 38369 14231 38403
rect 14657 38369 14691 38403
rect 15301 38369 15335 38403
rect 8493 38301 8527 38335
rect 10425 38301 10459 38335
rect 12541 38301 12575 38335
rect 1961 38233 1995 38267
rect 9045 38233 9079 38267
rect 11253 38233 11287 38267
rect 14105 38233 14139 38267
rect 18429 38437 18463 38471
rect 16313 38369 16347 38403
rect 23673 38369 23707 38403
rect 15853 38233 15887 38267
rect 1593 38165 1627 38199
rect 11529 38165 11563 38199
rect 12449 38165 12483 38199
rect 13553 38165 13587 38199
rect 14381 38165 14415 38199
rect 15025 38165 15059 38199
rect 15485 38165 15519 38199
rect 15577 38165 15611 38199
rect 16221 38165 16255 38199
rect 16773 38165 16807 38199
rect 17233 38165 17267 38199
rect 17601 38165 17635 38199
rect 8953 37961 8987 37995
rect 9689 37961 9723 37995
rect 11069 37961 11103 37995
rect 15025 37961 15059 37995
rect 16589 37961 16623 37995
rect 18613 37961 18647 37995
rect 18981 37961 19015 37995
rect 23489 37961 23523 37995
rect 25973 37961 26007 37995
rect 10931 37893 10965 37927
rect 15301 37893 15335 37927
rect 7573 37825 7607 37859
rect 11161 37825 11195 37859
rect 11529 37825 11563 37859
rect 11897 37825 11931 37859
rect 12449 37825 12483 37859
rect 14749 37825 14783 37859
rect 7941 37757 7975 37791
rect 8401 37757 8435 37791
rect 9413 37757 9447 37791
rect 9505 37757 9539 37791
rect 10793 37757 10827 37791
rect 12265 37757 12299 37791
rect 12633 37757 12667 37791
rect 14289 37757 14323 37791
rect 8309 37689 8343 37723
rect 9229 37689 9263 37723
rect 12817 37689 12851 37723
rect 13185 37689 13219 37723
rect 14013 37689 14047 37723
rect 14381 37689 14415 37723
rect 17417 37825 17451 37859
rect 20085 37825 20119 37859
rect 21189 37825 21223 37859
rect 26433 37825 26467 37859
rect 16313 37757 16347 37791
rect 17693 37757 17727 37791
rect 20269 37757 20303 37791
rect 21097 37757 21131 37791
rect 23765 37757 23799 37791
rect 24593 37757 24627 37791
rect 24685 37757 24719 37791
rect 26157 37757 26191 37791
rect 15577 37689 15611 37723
rect 15761 37689 15795 37723
rect 15945 37689 15979 37723
rect 17049 37689 17083 37723
rect 20361 37689 20395 37723
rect 23857 37689 23891 37723
rect 7205 37621 7239 37655
rect 8585 37621 8619 37655
rect 10241 37621 10275 37655
rect 10609 37621 10643 37655
rect 12725 37621 12759 37655
rect 13461 37621 13495 37655
rect 13921 37621 13955 37655
rect 14197 37621 14231 37655
rect 15301 37621 15335 37655
rect 15393 37621 15427 37655
rect 15853 37621 15887 37655
rect 18337 37621 18371 37655
rect 27537 37621 27571 37655
rect 6929 37417 6963 37451
rect 9413 37417 9447 37451
rect 12633 37417 12667 37451
rect 14197 37417 14231 37451
rect 15945 37417 15979 37451
rect 19625 37417 19659 37451
rect 20269 37417 20303 37451
rect 25513 37417 25547 37451
rect 26249 37417 26283 37451
rect 3065 37349 3099 37383
rect 8677 37349 8711 37383
rect 10333 37349 10367 37383
rect 10885 37349 10919 37383
rect 11529 37349 11563 37383
rect 13369 37349 13403 37383
rect 13461 37349 13495 37383
rect 13829 37349 13863 37383
rect 15117 37349 15151 37383
rect 1685 37281 1719 37315
rect 7297 37281 7331 37315
rect 9781 37281 9815 37315
rect 9873 37281 9907 37315
rect 11345 37281 11379 37315
rect 11437 37281 11471 37315
rect 12173 37281 12207 37315
rect 13277 37281 13311 37315
rect 15301 37281 15335 37315
rect 16681 37281 16715 37315
rect 16865 37281 16899 37315
rect 17601 37281 17635 37315
rect 18245 37281 18279 37315
rect 18429 37281 18463 37315
rect 21925 37281 21959 37315
rect 22017 37281 22051 37315
rect 22753 37281 22787 37315
rect 23673 37281 23707 37315
rect 24225 37281 24259 37315
rect 1409 37213 1443 37247
rect 7021 37213 7055 37247
rect 11161 37213 11195 37247
rect 11897 37213 11931 37247
rect 13093 37213 13127 37247
rect 15669 37213 15703 37247
rect 17233 37213 17267 37247
rect 22845 37213 22879 37247
rect 23949 37213 23983 37247
rect 15466 37145 15500 37179
rect 16405 37145 16439 37179
rect 18613 37145 18647 37179
rect 6193 37077 6227 37111
rect 6469 37077 6503 37111
rect 9045 37077 9079 37111
rect 12909 37077 12943 37111
rect 14473 37077 14507 37111
rect 15577 37077 15611 37111
rect 17003 37077 17037 37111
rect 17141 37077 17175 37111
rect 17969 37077 18003 37111
rect 18981 37077 19015 37111
rect 19349 37077 19383 37111
rect 1685 36873 1719 36907
rect 6285 36873 6319 36907
rect 8953 36873 8987 36907
rect 10931 36873 10965 36907
rect 11069 36873 11103 36907
rect 11805 36873 11839 36907
rect 12725 36873 12759 36907
rect 13074 36873 13108 36907
rect 17417 36873 17451 36907
rect 18521 36873 18555 36907
rect 22201 36873 22235 36907
rect 22661 36873 22695 36907
rect 23949 36873 23983 36907
rect 24409 36873 24443 36907
rect 6561 36805 6595 36839
rect 10609 36805 10643 36839
rect 13185 36805 13219 36839
rect 15761 36805 15795 36839
rect 15945 36805 15979 36839
rect 18245 36805 18279 36839
rect 19257 36805 19291 36839
rect 2145 36737 2179 36771
rect 7113 36737 7147 36771
rect 10241 36737 10275 36771
rect 11161 36737 11195 36771
rect 11529 36737 11563 36771
rect 13277 36737 13311 36771
rect 14473 36737 14507 36771
rect 15209 36737 15243 36771
rect 1869 36669 1903 36703
rect 5549 36669 5583 36703
rect 6837 36669 6871 36703
rect 9413 36669 9447 36703
rect 9597 36669 9631 36703
rect 10793 36669 10827 36703
rect 12909 36669 12943 36703
rect 14381 36669 14415 36703
rect 16773 36737 16807 36771
rect 17141 36737 17175 36771
rect 20545 36737 20579 36771
rect 26065 36737 26099 36771
rect 26157 36737 26191 36771
rect 16313 36669 16347 36703
rect 18061 36669 18095 36703
rect 18889 36669 18923 36703
rect 19073 36669 19107 36703
rect 19533 36669 19567 36703
rect 19901 36669 19935 36703
rect 20637 36669 20671 36703
rect 21097 36669 21131 36703
rect 26433 36669 26467 36703
rect 8493 36601 8527 36635
rect 12265 36601 12299 36635
rect 14749 36601 14783 36635
rect 14841 36601 14875 36635
rect 15761 36601 15795 36635
rect 16037 36601 16071 36635
rect 16405 36601 16439 36635
rect 17785 36601 17819 36635
rect 21373 36601 21407 36635
rect 21925 36601 21959 36635
rect 3249 36533 3283 36567
rect 5917 36533 5951 36567
rect 9229 36533 9263 36567
rect 9689 36533 9723 36567
rect 13553 36533 13587 36567
rect 14013 36533 14047 36567
rect 14657 36533 14691 36567
rect 15577 36533 15611 36567
rect 16221 36533 16255 36567
rect 27721 36533 27755 36567
rect 1961 36329 1995 36363
rect 6929 36329 6963 36363
rect 7573 36329 7607 36363
rect 8309 36329 8343 36363
rect 10149 36329 10183 36363
rect 14565 36329 14599 36363
rect 19625 36329 19659 36363
rect 19993 36329 20027 36363
rect 20729 36329 20763 36363
rect 8401 36261 8435 36295
rect 8769 36261 8803 36295
rect 13277 36261 13311 36295
rect 14013 36261 14047 36295
rect 17141 36261 17175 36295
rect 17233 36261 17267 36295
rect 17601 36261 17635 36295
rect 21833 36261 21867 36295
rect 4905 36193 4939 36227
rect 8217 36193 8251 36227
rect 10149 36193 10183 36227
rect 10609 36193 10643 36227
rect 10701 36193 10735 36227
rect 11253 36193 11287 36227
rect 13093 36193 13127 36227
rect 13185 36193 13219 36227
rect 15945 36193 15979 36227
rect 17049 36193 17083 36227
rect 18521 36193 18555 36227
rect 19809 36193 19843 36227
rect 22569 36193 22603 36227
rect 4629 36125 4663 36159
rect 8033 36125 8067 36159
rect 9505 36125 9539 36159
rect 12909 36125 12943 36159
rect 13645 36125 13679 36159
rect 16037 36125 16071 36159
rect 16865 36125 16899 36159
rect 18429 36125 18463 36159
rect 21741 36125 21775 36159
rect 22661 36125 22695 36159
rect 12173 36057 12207 36091
rect 16773 36057 16807 36091
rect 20269 36057 20303 36091
rect 2329 35989 2363 36023
rect 6009 35989 6043 36023
rect 7849 35989 7883 36023
rect 9045 35989 9079 36023
rect 11713 35989 11747 36023
rect 12541 35989 12575 36023
rect 14841 35989 14875 36023
rect 16405 35989 16439 36023
rect 18061 35989 18095 36023
rect 18705 35989 18739 36023
rect 19349 35989 19383 36023
rect 21189 35989 21223 36023
rect 23673 35989 23707 36023
rect 26249 35989 26283 36023
rect 4629 35785 4663 35819
rect 4905 35785 4939 35819
rect 5181 35785 5215 35819
rect 8585 35785 8619 35819
rect 17233 35785 17267 35819
rect 18889 35785 18923 35819
rect 19625 35785 19659 35819
rect 21281 35785 21315 35819
rect 22477 35785 22511 35819
rect 4169 35717 4203 35751
rect 8861 35717 8895 35751
rect 8953 35717 8987 35751
rect 10425 35717 10459 35751
rect 10517 35717 10551 35751
rect 13553 35717 13587 35751
rect 15853 35717 15887 35751
rect 2881 35649 2915 35683
rect 8309 35649 8343 35683
rect 2513 35581 2547 35615
rect 3157 35581 3191 35615
rect 4721 35581 4755 35615
rect 5733 35581 5767 35615
rect 6193 35581 6227 35615
rect 7113 35581 7147 35615
rect 7849 35581 7883 35615
rect 9873 35649 9907 35683
rect 10057 35649 10091 35683
rect 9137 35581 9171 35615
rect 2329 35513 2363 35547
rect 5641 35513 5675 35547
rect 6653 35513 6687 35547
rect 7573 35513 7607 35547
rect 7941 35513 7975 35547
rect 8861 35513 8895 35547
rect 9321 35513 9355 35547
rect 9505 35513 9539 35547
rect 10241 35581 10275 35615
rect 1593 35445 1627 35479
rect 2145 35445 2179 35479
rect 5917 35445 5951 35479
rect 7389 35445 7423 35479
rect 7757 35445 7791 35479
rect 9413 35445 9447 35479
rect 10057 35445 10091 35479
rect 19073 35717 19107 35751
rect 13185 35649 13219 35683
rect 14013 35649 14047 35683
rect 15485 35649 15519 35683
rect 15945 35649 15979 35683
rect 16957 35649 16991 35683
rect 17877 35649 17911 35683
rect 18061 35649 18095 35683
rect 18797 35649 18831 35683
rect 18889 35649 18923 35683
rect 23489 35649 23523 35683
rect 23949 35649 23983 35683
rect 26157 35649 26191 35683
rect 26433 35649 26467 35683
rect 11897 35581 11931 35615
rect 14289 35581 14323 35615
rect 15724 35581 15758 35615
rect 18245 35581 18279 35615
rect 19901 35581 19935 35615
rect 21649 35581 21683 35615
rect 23673 35581 23707 35615
rect 26065 35581 26099 35615
rect 10701 35513 10735 35547
rect 11069 35513 11103 35547
rect 11437 35513 11471 35547
rect 12265 35513 12299 35547
rect 12449 35513 12483 35547
rect 12817 35513 12851 35547
rect 14381 35513 14415 35547
rect 14749 35513 14783 35547
rect 15577 35513 15611 35547
rect 18429 35513 18463 35547
rect 20545 35513 20579 35547
rect 22109 35513 22143 35547
rect 25329 35513 25363 35547
rect 27813 35513 27847 35547
rect 10425 35445 10459 35479
rect 10885 35445 10919 35479
rect 10977 35445 11011 35479
rect 12633 35445 12667 35479
rect 12725 35445 12759 35479
rect 13921 35445 13955 35479
rect 14197 35445 14231 35479
rect 15025 35445 15059 35479
rect 16221 35445 16255 35479
rect 18337 35445 18371 35479
rect 20821 35445 20855 35479
rect 22845 35445 22879 35479
rect 4629 35241 4663 35275
rect 5641 35241 5675 35275
rect 9965 35241 9999 35275
rect 10701 35241 10735 35275
rect 11069 35241 11103 35275
rect 13461 35241 13495 35275
rect 14197 35241 14231 35275
rect 16405 35241 16439 35275
rect 18153 35241 18187 35275
rect 19441 35241 19475 35275
rect 19901 35241 19935 35275
rect 20545 35241 20579 35275
rect 9137 35173 9171 35207
rect 11253 35173 11287 35207
rect 11989 35173 12023 35207
rect 12541 35173 12575 35207
rect 5089 35105 5123 35139
rect 6101 35105 6135 35139
rect 7113 35105 7147 35139
rect 9873 35105 9907 35139
rect 10041 35105 10075 35139
rect 10425 35105 10459 35139
rect 11483 35105 11517 35139
rect 12817 35105 12851 35139
rect 12964 35105 12998 35139
rect 6009 35037 6043 35071
rect 7389 35037 7423 35071
rect 9689 35037 9723 35071
rect 11621 35037 11655 35071
rect 13185 35037 13219 35071
rect 3893 34969 3927 35003
rect 15301 35173 15335 35207
rect 15669 35173 15703 35207
rect 17233 35173 17267 35207
rect 17601 35173 17635 35207
rect 18429 35173 18463 35207
rect 14473 35105 14507 35139
rect 15485 35105 15519 35139
rect 15577 35105 15611 35139
rect 17049 35105 17083 35139
rect 17141 35105 17175 35139
rect 19073 35105 19107 35139
rect 21741 35105 21775 35139
rect 22017 35105 22051 35139
rect 23397 35105 23431 35139
rect 16037 35037 16071 35071
rect 16865 35037 16899 35071
rect 21189 35037 21223 35071
rect 22201 35037 22235 35071
rect 23121 35037 23155 35071
rect 1593 34901 1627 34935
rect 3433 34901 3467 34935
rect 4997 34901 5031 34935
rect 5273 34901 5307 34935
rect 6285 34901 6319 34935
rect 6561 34901 6595 34935
rect 7021 34901 7055 34935
rect 8677 34901 8711 34935
rect 9413 34901 9447 34935
rect 11418 34901 11452 34935
rect 13093 34901 13127 34935
rect 14013 34901 14047 34935
rect 14197 34901 14231 34935
rect 15117 34901 15151 34935
rect 16681 34901 16715 34935
rect 22477 34901 22511 34935
rect 23029 34901 23063 34935
rect 24501 34901 24535 34935
rect 26249 34901 26283 34935
rect 4537 34697 4571 34731
rect 12173 34697 12207 34731
rect 15301 34697 15335 34731
rect 16773 34697 16807 34731
rect 17141 34697 17175 34731
rect 17877 34697 17911 34731
rect 19441 34697 19475 34731
rect 20269 34697 20303 34731
rect 21925 34697 21959 34731
rect 22569 34697 22603 34731
rect 23121 34697 23155 34731
rect 25973 34697 26007 34731
rect 27721 34697 27755 34731
rect 5089 34629 5123 34663
rect 6009 34629 6043 34663
rect 6653 34629 6687 34663
rect 9781 34629 9815 34663
rect 18337 34629 18371 34663
rect 19993 34629 20027 34663
rect 22293 34629 22327 34663
rect 3893 34561 3927 34595
rect 5365 34561 5399 34595
rect 5917 34561 5951 34595
rect 1409 34493 1443 34527
rect 1685 34493 1719 34527
rect 3525 34493 3559 34527
rect 4261 34493 4295 34527
rect 4353 34493 4387 34527
rect 5457 34493 5491 34527
rect 7849 34561 7883 34595
rect 8125 34561 8159 34595
rect 8953 34561 8987 34595
rect 13277 34561 13311 34595
rect 14105 34561 14139 34595
rect 14197 34561 14231 34595
rect 18429 34561 18463 34595
rect 19073 34561 19107 34595
rect 20545 34561 20579 34595
rect 21557 34561 21591 34595
rect 23489 34561 23523 34595
rect 25053 34561 25087 34595
rect 26433 34561 26467 34595
rect 7021 34493 7055 34527
rect 7573 34493 7607 34527
rect 8493 34493 8527 34527
rect 8677 34493 8711 34527
rect 9045 34493 9079 34527
rect 10057 34493 10091 34527
rect 10517 34493 10551 34527
rect 10701 34493 10735 34527
rect 10885 34493 10919 34527
rect 12541 34493 12575 34527
rect 12725 34493 12759 34527
rect 12893 34493 12927 34527
rect 14381 34493 14415 34527
rect 14933 34493 14967 34527
rect 15761 34493 15795 34527
rect 18208 34493 18242 34527
rect 20821 34493 20855 34527
rect 21373 34493 21407 34527
rect 23673 34493 23707 34527
rect 23949 34493 23983 34527
rect 26157 34493 26191 34527
rect 13553 34425 13587 34459
rect 14565 34425 14599 34459
rect 16129 34425 16163 34459
rect 16497 34425 16531 34459
rect 18061 34425 18095 34459
rect 2789 34357 2823 34391
rect 6009 34357 6043 34391
rect 6285 34357 6319 34391
rect 7205 34357 7239 34391
rect 11345 34357 11379 34391
rect 11897 34357 11931 34391
rect 12817 34357 12851 34391
rect 14473 34357 14507 34391
rect 15945 34357 15979 34391
rect 16037 34357 16071 34391
rect 18705 34357 18739 34391
rect 1685 34153 1719 34187
rect 3433 34153 3467 34187
rect 4353 34153 4387 34187
rect 4629 34153 4663 34187
rect 4997 34153 5031 34187
rect 5641 34153 5675 34187
rect 6561 34153 6595 34187
rect 12173 34153 12207 34187
rect 13921 34153 13955 34187
rect 16773 34153 16807 34187
rect 17693 34153 17727 34187
rect 18061 34153 18095 34187
rect 20269 34153 20303 34187
rect 22385 34153 22419 34187
rect 5365 34085 5399 34119
rect 5733 34085 5767 34119
rect 5825 34085 5859 34119
rect 9689 34085 9723 34119
rect 12357 34085 12391 34119
rect 13645 34085 13679 34119
rect 14013 34085 14047 34119
rect 14657 34085 14691 34119
rect 15025 34085 15059 34119
rect 21281 34085 21315 34119
rect 4445 34017 4479 34051
rect 5457 34017 5491 34051
rect 10149 34017 10183 34051
rect 10333 34017 10367 34051
rect 10609 34017 10643 34051
rect 10793 34017 10827 34051
rect 12265 34017 12299 34051
rect 13553 34017 13587 34051
rect 13829 34017 13863 34051
rect 15301 34017 15335 34051
rect 15448 34017 15482 34051
rect 16865 34017 16899 34051
rect 17049 34017 17083 34051
rect 18521 34017 18555 34051
rect 21097 34017 21131 34051
rect 21189 34017 21223 34051
rect 23397 34017 23431 34051
rect 23489 34017 23523 34051
rect 25237 34017 25271 34051
rect 6193 33949 6227 33983
rect 7021 33949 7055 33983
rect 7297 33949 7331 33983
rect 9505 33949 9539 33983
rect 11069 33949 11103 33983
rect 11897 33949 11931 33983
rect 11989 33949 12023 33983
rect 12725 33949 12759 33983
rect 14381 33949 14415 33983
rect 15669 33949 15703 33983
rect 17325 33949 17359 33983
rect 18245 33949 18279 33983
rect 20913 33949 20947 33983
rect 21649 33949 21683 33983
rect 22569 33949 22603 33983
rect 22661 33949 22695 33983
rect 24409 33949 24443 33983
rect 24961 33949 24995 33983
rect 25421 33949 25455 33983
rect 11529 33881 11563 33915
rect 21925 33881 21959 33915
rect 3801 33813 3835 33847
rect 6929 33813 6963 33847
rect 8401 33813 8435 33847
rect 9045 33813 9079 33847
rect 13093 33813 13127 33847
rect 15577 33813 15611 33847
rect 15761 33813 15795 33847
rect 16405 33813 16439 33847
rect 19809 33813 19843 33847
rect 20729 33813 20763 33847
rect 23857 33813 23891 33847
rect 24317 33813 24351 33847
rect 26249 33813 26283 33847
rect 4537 33609 4571 33643
rect 6285 33609 6319 33643
rect 6653 33609 6687 33643
rect 7113 33609 7147 33643
rect 9045 33609 9079 33643
rect 11713 33609 11747 33643
rect 13645 33609 13679 33643
rect 17601 33609 17635 33643
rect 19165 33609 19199 33643
rect 22661 33609 22695 33643
rect 22937 33609 22971 33643
rect 23213 33609 23247 33643
rect 23857 33609 23891 33643
rect 24501 33609 24535 33643
rect 25973 33609 26007 33643
rect 3525 33541 3559 33575
rect 10977 33541 11011 33575
rect 2789 33473 2823 33507
rect 3157 33473 3191 33507
rect 5365 33473 5399 33507
rect 7297 33473 7331 33507
rect 7941 33473 7975 33507
rect 8125 33473 8159 33507
rect 20913 33473 20947 33507
rect 22569 33473 22603 33507
rect 4261 33405 4295 33439
rect 4353 33405 4387 33439
rect 5457 33405 5491 33439
rect 7849 33405 7883 33439
rect 8217 33405 8251 33439
rect 9689 33405 9723 33439
rect 9965 33405 9999 33439
rect 10149 33405 10183 33439
rect 10333 33405 10367 33439
rect 10701 33405 10735 33439
rect 12449 33405 12483 33439
rect 12633 33405 12667 33439
rect 13185 33405 13219 33439
rect 15117 33405 15151 33439
rect 15577 33405 15611 33439
rect 15853 33405 15887 33439
rect 16129 33405 16163 33439
rect 18705 33405 18739 33439
rect 19993 33405 20027 33439
rect 20821 33405 20855 33439
rect 22109 33405 22143 33439
rect 3893 33337 3927 33371
rect 4905 33337 4939 33371
rect 5917 33337 5951 33371
rect 9229 33337 9263 33371
rect 12817 33337 12851 33371
rect 14013 33337 14047 33371
rect 16957 33337 16991 33371
rect 18797 33337 18831 33371
rect 20085 33337 20119 33371
rect 21833 33337 21867 33371
rect 22201 33337 22235 33371
rect 25145 33541 25179 33575
rect 24869 33473 24903 33507
rect 26157 33473 26191 33507
rect 26433 33405 26467 33439
rect 5273 33269 5307 33303
rect 8677 33269 8711 33303
rect 11989 33269 12023 33303
rect 12725 33269 12759 33303
rect 14381 33269 14415 33303
rect 14933 33269 14967 33303
rect 17325 33269 17359 33303
rect 19441 33269 19475 33303
rect 21373 33269 21407 33303
rect 21649 33269 21683 33303
rect 22017 33269 22051 33303
rect 22661 33269 22695 33303
rect 27537 33269 27571 33303
rect 4629 33065 4663 33099
rect 4905 33065 4939 33099
rect 7757 33065 7791 33099
rect 9229 33065 9263 33099
rect 11621 33065 11655 33099
rect 14565 33065 14599 33099
rect 14657 33065 14691 33099
rect 14933 33065 14967 33099
rect 15485 33065 15519 33099
rect 16313 33065 16347 33099
rect 17049 33065 17083 33099
rect 18613 33065 18647 33099
rect 19625 33065 19659 33099
rect 20729 33065 20763 33099
rect 22937 33065 22971 33099
rect 23673 33065 23707 33099
rect 25145 33065 25179 33099
rect 8033 32997 8067 33031
rect 9689 32997 9723 33031
rect 12449 32997 12483 33031
rect 12725 32997 12759 33031
rect 15669 32997 15703 33031
rect 16037 32997 16071 33031
rect 23305 32997 23339 33031
rect 4721 32929 4755 32963
rect 8309 32929 8343 32963
rect 9413 32929 9447 32963
rect 10333 32929 10367 32963
rect 10701 32929 10735 32963
rect 11713 32929 11747 32963
rect 13185 32929 13219 32963
rect 13461 32929 13495 32963
rect 13553 32929 13587 32963
rect 14197 32929 14231 32963
rect 14657 32929 14691 32963
rect 15577 32929 15611 32963
rect 17233 32929 17267 32963
rect 19717 32929 19751 32963
rect 20913 32929 20947 32963
rect 3525 32861 3559 32895
rect 5733 32861 5767 32895
rect 6009 32861 6043 32895
rect 7389 32861 7423 32895
rect 8217 32861 8251 32895
rect 8769 32861 8803 32895
rect 10241 32861 10275 32895
rect 10793 32861 10827 32895
rect 13829 32861 13863 32895
rect 15301 32861 15335 32895
rect 17509 32861 17543 32895
rect 21189 32861 21223 32895
rect 22293 32861 22327 32895
rect 23765 32861 23799 32895
rect 24041 32861 24075 32895
rect 9413 32793 9447 32827
rect 3893 32725 3927 32759
rect 5457 32725 5491 32759
rect 11161 32725 11195 32759
rect 11897 32725 11931 32759
rect 16681 32725 16715 32759
rect 19165 32725 19199 32759
rect 19901 32725 19935 32759
rect 20269 32725 20303 32759
rect 26249 32725 26283 32759
rect 3433 32521 3467 32555
rect 4905 32521 4939 32555
rect 5181 32521 5215 32555
rect 6193 32521 6227 32555
rect 7941 32521 7975 32555
rect 9689 32521 9723 32555
rect 11897 32521 11931 32555
rect 12909 32521 12943 32555
rect 13829 32521 13863 32555
rect 17785 32521 17819 32555
rect 21189 32521 21223 32555
rect 23489 32521 23523 32555
rect 4261 32453 4295 32487
rect 7389 32453 7423 32487
rect 12725 32453 12759 32487
rect 18245 32453 18279 32487
rect 22477 32453 22511 32487
rect 23029 32453 23063 32487
rect 4629 32385 4663 32419
rect 8493 32385 8527 32419
rect 12596 32385 12630 32419
rect 14013 32385 14047 32419
rect 15761 32385 15795 32419
rect 15945 32385 15979 32419
rect 19073 32385 19107 32419
rect 19441 32385 19475 32419
rect 4721 32317 4755 32351
rect 5733 32317 5767 32351
rect 7573 32317 7607 32351
rect 8401 32317 8435 32351
rect 8769 32317 8803 32351
rect 9229 32317 9263 32351
rect 10149 32317 10183 32351
rect 10517 32317 10551 32351
rect 10885 32317 10919 32351
rect 11253 32317 11287 32351
rect 12788 32317 12822 32351
rect 16405 32317 16439 32351
rect 16589 32317 16623 32351
rect 16957 32317 16991 32351
rect 17141 32317 17175 32351
rect 18061 32317 18095 32351
rect 19165 32317 19199 32351
rect 21557 32317 21591 32351
rect 21649 32317 21683 32351
rect 22017 32317 22051 32351
rect 22569 32317 22603 32351
rect 5641 32249 5675 32283
rect 8861 32249 8895 32283
rect 12449 32249 12483 32283
rect 14289 32249 14323 32283
rect 14381 32249 14415 32283
rect 14749 32249 14783 32283
rect 18521 32249 18555 32283
rect 20821 32249 20855 32283
rect 3893 32181 3927 32215
rect 5917 32181 5951 32215
rect 6561 32181 6595 32215
rect 8677 32181 8711 32215
rect 10149 32181 10183 32215
rect 12265 32181 12299 32215
rect 13461 32181 13495 32215
rect 14197 32181 14231 32215
rect 15393 32181 15427 32215
rect 17417 32181 17451 32215
rect 23949 32181 23983 32215
rect 24317 32181 24351 32215
rect 24593 32181 24627 32215
rect 2881 31977 2915 32011
rect 4997 31977 5031 32011
rect 5273 31977 5307 32011
rect 8309 31977 8343 32011
rect 8493 31977 8527 32011
rect 9137 31977 9171 32011
rect 9413 31977 9447 32011
rect 9689 31977 9723 32011
rect 10057 31977 10091 32011
rect 10793 31977 10827 32011
rect 11253 31977 11287 32011
rect 13645 31977 13679 32011
rect 14197 31977 14231 32011
rect 14933 31977 14967 32011
rect 15117 31977 15151 32011
rect 15485 31977 15519 32011
rect 18245 31977 18279 32011
rect 20637 31977 20671 32011
rect 21741 31977 21775 32011
rect 22201 31977 22235 32011
rect 23489 31977 23523 32011
rect 4629 31909 4663 31943
rect 5733 31909 5767 31943
rect 7481 31909 7515 31943
rect 1501 31841 1535 31875
rect 6101 31841 6135 31875
rect 1777 31773 1811 31807
rect 5825 31773 5859 31807
rect 10149 31909 10183 31943
rect 8585 31841 8619 31875
rect 9689 31841 9723 31875
rect 9781 31841 9815 31875
rect 9965 31841 9999 31875
rect 10517 31841 10551 31875
rect 11805 31841 11839 31875
rect 12173 31841 12207 31875
rect 12265 31841 12299 31875
rect 13185 31841 13219 31875
rect 13461 31841 13495 31875
rect 17969 31909 18003 31943
rect 23121 31909 23155 31943
rect 15301 31841 15335 31875
rect 18613 31841 18647 31875
rect 19441 31841 19475 31875
rect 19809 31841 19843 31875
rect 20269 31841 20303 31875
rect 21005 31841 21039 31875
rect 22937 31841 22971 31875
rect 11345 31773 11379 31807
rect 12817 31773 12851 31807
rect 13277 31773 13311 31807
rect 15117 31773 15151 31807
rect 16129 31773 16163 31807
rect 16313 31773 16347 31807
rect 16589 31773 16623 31807
rect 18981 31773 19015 31807
rect 19349 31773 19383 31807
rect 19717 31773 19751 31807
rect 20913 31773 20947 31807
rect 8493 31705 8527 31739
rect 8769 31705 8803 31739
rect 15761 31705 15795 31739
rect 7849 31637 7883 31671
rect 21189 31637 21223 31671
rect 6653 31433 6687 31467
rect 7757 31433 7791 31467
rect 7941 31433 7975 31467
rect 8861 31433 8895 31467
rect 11437 31433 11471 31467
rect 11897 31433 11931 31467
rect 12725 31433 12759 31467
rect 13921 31433 13955 31467
rect 14289 31433 14323 31467
rect 15393 31433 15427 31467
rect 16405 31433 16439 31467
rect 17325 31433 17359 31467
rect 19625 31433 19659 31467
rect 21741 31433 21775 31467
rect 5549 31365 5583 31399
rect 6285 31365 6319 31399
rect 7573 31365 7607 31399
rect 16957 31365 16991 31399
rect 7757 31297 7791 31331
rect 8033 31297 8067 31331
rect 9321 31297 9355 31331
rect 10701 31297 10735 31331
rect 12817 31297 12851 31331
rect 15761 31297 15795 31331
rect 18061 31297 18095 31331
rect 21373 31297 21407 31331
rect 23489 31297 23523 31331
rect 23949 31297 23983 31331
rect 26065 31297 26099 31331
rect 27629 31297 27663 31331
rect 7021 31229 7055 31263
rect 8125 31229 8159 31263
rect 9873 31229 9907 31263
rect 10057 31229 10091 31263
rect 10333 31229 10367 31263
rect 10793 31229 10827 31263
rect 14565 31229 14599 31263
rect 16497 31229 16531 31263
rect 17693 31229 17727 31263
rect 18337 31229 18371 31263
rect 20545 31229 20579 31263
rect 20729 31229 20763 31263
rect 21925 31229 21959 31263
rect 22385 31229 22419 31263
rect 22845 31229 22879 31263
rect 23673 31229 23707 31263
rect 26157 31229 26191 31263
rect 26433 31229 26467 31263
rect 1961 31161 1995 31195
rect 8585 31161 8619 31195
rect 9413 31161 9447 31195
rect 13185 31161 13219 31195
rect 13553 31161 13587 31195
rect 14381 31161 14415 31195
rect 14657 31161 14691 31195
rect 14749 31161 14783 31195
rect 15117 31161 15151 31195
rect 21097 31161 21131 31195
rect 1685 31093 1719 31127
rect 4813 31093 4847 31127
rect 5181 31093 5215 31127
rect 5825 31093 5859 31127
rect 7205 31093 7239 31127
rect 12265 31093 12299 31127
rect 13001 31093 13035 31127
rect 13093 31093 13127 31127
rect 19993 31093 20027 31127
rect 20361 31093 20395 31127
rect 22109 31093 22143 31127
rect 25053 31093 25087 31127
rect 6009 30889 6043 30923
rect 9965 30889 9999 30923
rect 10517 30889 10551 30923
rect 11713 30889 11747 30923
rect 13461 30889 13495 30923
rect 13829 30889 13863 30923
rect 16681 30889 16715 30923
rect 23765 30889 23799 30923
rect 9413 30821 9447 30855
rect 10333 30821 10367 30855
rect 10701 30821 10735 30855
rect 11069 30821 11103 30855
rect 12725 30821 12759 30855
rect 12817 30821 12851 30855
rect 16313 30821 16347 30855
rect 21465 30821 21499 30855
rect 6101 30753 6135 30787
rect 8585 30753 8619 30787
rect 9137 30753 9171 30787
rect 10609 30753 10643 30787
rect 12357 30753 12391 30787
rect 12449 30753 12483 30787
rect 12633 30753 12667 30787
rect 13185 30753 13219 30787
rect 14197 30753 14231 30787
rect 15301 30753 15335 30787
rect 15577 30753 15611 30787
rect 17693 30753 17727 30787
rect 20913 30753 20947 30787
rect 6377 30685 6411 30719
rect 8125 30685 8159 30719
rect 12081 30685 12115 30719
rect 14749 30685 14783 30719
rect 16037 30685 16071 30719
rect 17049 30685 17083 30719
rect 17969 30685 18003 30719
rect 20361 30685 20395 30719
rect 21833 30685 21867 30719
rect 22201 30685 22235 30719
rect 8769 30617 8803 30651
rect 14381 30617 14415 30651
rect 15393 30617 15427 30651
rect 19993 30617 20027 30651
rect 21097 30617 21131 30651
rect 5549 30549 5583 30583
rect 7481 30549 7515 30583
rect 8493 30549 8527 30583
rect 12173 30549 12207 30583
rect 15025 30549 15059 30583
rect 17601 30549 17635 30583
rect 19073 30549 19107 30583
rect 19625 30549 19659 30583
rect 26157 30549 26191 30583
rect 8677 30345 8711 30379
rect 10609 30345 10643 30379
rect 11529 30345 11563 30379
rect 11897 30345 11931 30379
rect 16681 30345 16715 30379
rect 20913 30345 20947 30379
rect 5273 30277 5307 30311
rect 6009 30277 6043 30311
rect 14289 30277 14323 30311
rect 14749 30277 14783 30311
rect 17049 30277 17083 30311
rect 18337 30277 18371 30311
rect 20269 30277 20303 30311
rect 5641 30209 5675 30243
rect 7113 30209 7147 30243
rect 10241 30209 10275 30243
rect 10885 30209 10919 30243
rect 12909 30209 12943 30243
rect 13645 30209 13679 30243
rect 17417 30209 17451 30243
rect 17785 30209 17819 30243
rect 18521 30209 18555 30243
rect 19901 30209 19935 30243
rect 4445 30141 4479 30175
rect 4813 30141 4847 30175
rect 6653 30141 6687 30175
rect 7297 30141 7331 30175
rect 7481 30141 7515 30175
rect 7849 30141 7883 30175
rect 7941 30141 7975 30175
rect 9137 30141 9171 30175
rect 9781 30141 9815 30175
rect 10057 30141 10091 30175
rect 11345 30141 11379 30175
rect 14749 30141 14783 30175
rect 14933 30141 14967 30175
rect 15301 30141 15335 30175
rect 15945 30141 15979 30175
rect 16405 30141 16439 30175
rect 18705 30141 18739 30175
rect 19073 30141 19107 30175
rect 19165 30141 19199 30175
rect 20085 30141 20119 30175
rect 20545 30141 20579 30175
rect 6377 30073 6411 30107
rect 9229 30073 9263 30107
rect 13093 30073 13127 30107
rect 13277 30073 13311 30107
rect 21281 30073 21315 30107
rect 21649 30073 21683 30107
rect 4261 30005 4295 30039
rect 6469 30005 6503 30039
rect 12173 30005 12207 30039
rect 12817 30005 12851 30039
rect 13185 30005 13219 30039
rect 19533 30005 19567 30039
rect 6561 29801 6595 29835
rect 8309 29801 8343 29835
rect 9045 29801 9079 29835
rect 9413 29801 9447 29835
rect 13461 29801 13495 29835
rect 16405 29801 16439 29835
rect 17877 29801 17911 29835
rect 19901 29801 19935 29835
rect 20453 29801 20487 29835
rect 21649 29801 21683 29835
rect 6193 29733 6227 29767
rect 6929 29733 6963 29767
rect 7941 29733 7975 29767
rect 12357 29733 12391 29767
rect 12449 29733 12483 29767
rect 15117 29733 15151 29767
rect 17049 29733 17083 29767
rect 17601 29733 17635 29767
rect 18705 29733 18739 29767
rect 19165 29733 19199 29767
rect 21189 29733 21223 29767
rect 7021 29665 7055 29699
rect 8125 29665 8159 29699
rect 10517 29665 10551 29699
rect 12265 29665 12299 29699
rect 13645 29665 13679 29699
rect 13792 29665 13826 29699
rect 15301 29665 15335 29699
rect 16865 29665 16899 29699
rect 17141 29665 17175 29699
rect 18613 29665 18647 29699
rect 18781 29665 18815 29699
rect 19533 29665 19567 29699
rect 20177 29665 20211 29699
rect 21833 29665 21867 29699
rect 5457 29597 5491 29631
rect 7573 29597 7607 29631
rect 9689 29597 9723 29631
rect 10241 29597 10275 29631
rect 10701 29597 10735 29631
rect 12081 29597 12115 29631
rect 12817 29597 12851 29631
rect 14013 29597 14047 29631
rect 14657 29597 14691 29631
rect 15669 29597 15703 29631
rect 18429 29597 18463 29631
rect 7205 29529 7239 29563
rect 11529 29529 11563 29563
rect 13093 29529 13127 29563
rect 15577 29529 15611 29563
rect 18245 29529 18279 29563
rect 19993 29529 20027 29563
rect 5825 29461 5859 29495
rect 11069 29461 11103 29495
rect 11989 29461 12023 29495
rect 13921 29461 13955 29495
rect 14289 29461 14323 29495
rect 15439 29461 15473 29495
rect 15761 29461 15795 29495
rect 16681 29461 16715 29495
rect 6653 29257 6687 29291
rect 7113 29257 7147 29291
rect 9137 29257 9171 29291
rect 11437 29257 11471 29291
rect 11713 29257 11747 29291
rect 12633 29257 12667 29291
rect 14657 29257 14691 29291
rect 15761 29257 15795 29291
rect 16451 29257 16485 29291
rect 16589 29257 16623 29291
rect 17325 29257 17359 29291
rect 18337 29257 18371 29291
rect 19625 29257 19659 29291
rect 19901 29257 19935 29291
rect 21005 29257 21039 29291
rect 21741 29257 21775 29291
rect 9413 29189 9447 29223
rect 9689 29189 9723 29223
rect 12173 29189 12207 29223
rect 17877 29189 17911 29223
rect 18889 29189 18923 29223
rect 19349 29189 19383 29223
rect 7757 29121 7791 29155
rect 8769 29121 8803 29155
rect 13093 29121 13127 29155
rect 15485 29121 15519 29155
rect 16681 29121 16715 29155
rect 18061 29121 18095 29155
rect 20269 29121 20303 29155
rect 5549 29053 5583 29087
rect 6285 29053 6319 29087
rect 8217 29053 8251 29087
rect 8309 29053 8343 29087
rect 10241 29053 10275 29087
rect 10333 29053 10367 29087
rect 10609 29053 10643 29087
rect 10793 29053 10827 29087
rect 13185 29053 13219 29087
rect 13461 29053 13495 29087
rect 14289 29053 14323 29087
rect 14933 29053 14967 29087
rect 16313 29053 16347 29087
rect 18153 29053 18187 29087
rect 19441 29053 19475 29087
rect 20637 29053 20671 29087
rect 5825 28985 5859 29019
rect 8125 28985 8159 29019
rect 13545 28985 13579 29019
rect 13921 28985 13955 29019
rect 14749 28985 14783 29019
rect 15117 28985 15151 29019
rect 17049 28985 17083 29019
rect 13369 28917 13403 28951
rect 15025 28917 15059 28951
rect 16129 28917 16163 28951
rect 5549 28713 5583 28747
rect 6193 28713 6227 28747
rect 6561 28713 6595 28747
rect 9413 28713 9447 28747
rect 9689 28713 9723 28747
rect 14013 28713 14047 28747
rect 15577 28713 15611 28747
rect 16313 28713 16347 28747
rect 17509 28713 17543 28747
rect 18153 28713 18187 28747
rect 18889 28713 18923 28747
rect 19349 28713 19383 28747
rect 19993 28713 20027 28747
rect 20361 28713 20395 28747
rect 9137 28645 9171 28679
rect 1409 28577 1443 28611
rect 5733 28577 5767 28611
rect 8585 28577 8619 28611
rect 1685 28509 1719 28543
rect 6929 28509 6963 28543
rect 7757 28509 7791 28543
rect 8309 28509 8343 28543
rect 8769 28509 8803 28543
rect 12817 28645 12851 28679
rect 12909 28645 12943 28679
rect 13645 28645 13679 28679
rect 15485 28645 15519 28679
rect 15669 28645 15703 28679
rect 16865 28645 16899 28679
rect 10793 28577 10827 28611
rect 11345 28577 11379 28611
rect 12081 28577 12115 28611
rect 12449 28577 12483 28611
rect 12725 28577 12759 28611
rect 14105 28577 14139 28611
rect 14933 28577 14967 28611
rect 18429 28577 18463 28611
rect 19441 28577 19475 28611
rect 11437 28509 11471 28543
rect 12541 28509 12575 28543
rect 13277 28509 13311 28543
rect 15301 28509 15335 28543
rect 16037 28509 16071 28543
rect 17012 28509 17046 28543
rect 17233 28509 17267 28543
rect 7297 28441 7331 28475
rect 9689 28441 9723 28475
rect 10333 28441 10367 28475
rect 10701 28441 10735 28475
rect 14289 28441 14323 28475
rect 14565 28441 14599 28475
rect 2973 28373 3007 28407
rect 7665 28373 7699 28407
rect 9873 28373 9907 28407
rect 16681 28373 16715 28407
rect 17141 28373 17175 28407
rect 18613 28373 18647 28407
rect 19625 28373 19659 28407
rect 21741 28373 21775 28407
rect 3157 28169 3191 28203
rect 8953 28169 8987 28203
rect 11253 28169 11287 28203
rect 13737 28169 13771 28203
rect 16221 28169 16255 28203
rect 16405 28169 16439 28203
rect 16773 28169 16807 28203
rect 17693 28169 17727 28203
rect 19441 28169 19475 28203
rect 20913 28169 20947 28203
rect 21557 28169 21591 28203
rect 7205 28101 7239 28135
rect 9321 28101 9355 28135
rect 11621 28101 11655 28135
rect 11897 28101 11931 28135
rect 1593 28033 1627 28067
rect 9965 28033 9999 28067
rect 12173 28033 12207 28067
rect 14289 28033 14323 28067
rect 18337 28101 18371 28135
rect 20729 28101 20763 28135
rect 16497 28033 16531 28067
rect 17417 28033 17451 28067
rect 20361 28033 20395 28067
rect 21741 28033 21775 28067
rect 22661 28033 22695 28067
rect 1869 27965 1903 27999
rect 6653 27965 6687 27999
rect 7021 27965 7055 27999
rect 8033 27965 8067 27999
rect 8585 27965 8619 27999
rect 9505 27965 9539 27999
rect 9689 27965 9723 27999
rect 10057 27965 10091 27999
rect 11345 27965 11379 27999
rect 11621 27965 11655 27999
rect 12449 27965 12483 27999
rect 12633 27965 12667 27999
rect 12725 27965 12759 27999
rect 13185 27965 13219 27999
rect 14197 27965 14231 27999
rect 14565 27965 14599 27999
rect 14933 27965 14967 27999
rect 15669 27965 15703 27999
rect 16221 27965 16255 27999
rect 16589 27965 16623 27999
rect 18521 27965 18555 27999
rect 18705 27965 18739 27999
rect 18889 27965 18923 27999
rect 19901 27965 19935 27999
rect 21097 27965 21131 27999
rect 22569 27965 22603 27999
rect 5641 27897 5675 27931
rect 7849 27897 7883 27931
rect 10885 27897 10919 27931
rect 16037 27897 16071 27931
rect 21833 27897 21867 27931
rect 6285 27829 6319 27863
rect 8217 27829 8251 27863
rect 11529 27829 11563 27863
rect 14105 27829 14139 27863
rect 20085 27829 20119 27863
rect 2329 27625 2363 27659
rect 7389 27625 7423 27659
rect 13369 27625 13403 27659
rect 14473 27625 14507 27659
rect 15853 27625 15887 27659
rect 18521 27625 18555 27659
rect 4629 27557 4663 27591
rect 7205 27557 7239 27591
rect 9873 27557 9907 27591
rect 11529 27557 11563 27591
rect 14841 27557 14875 27591
rect 19349 27557 19383 27591
rect 21741 27557 21775 27591
rect 4813 27489 4847 27523
rect 6837 27489 6871 27523
rect 7941 27489 7975 27523
rect 8309 27489 8343 27523
rect 10057 27489 10091 27523
rect 10425 27489 10459 27523
rect 10885 27489 10919 27523
rect 12081 27489 12115 27523
rect 12541 27489 12575 27523
rect 13921 27489 13955 27523
rect 15393 27489 15427 27523
rect 16681 27489 16715 27523
rect 18889 27489 18923 27523
rect 20085 27489 20119 27523
rect 5089 27421 5123 27455
rect 7757 27421 7791 27455
rect 8217 27421 8251 27455
rect 9137 27421 9171 27455
rect 13001 27421 13035 27455
rect 16405 27421 16439 27455
rect 19717 27421 19751 27455
rect 10885 27353 10919 27387
rect 12081 27353 12115 27387
rect 14105 27353 14139 27387
rect 19073 27353 19107 27387
rect 1593 27285 1627 27319
rect 1961 27285 1995 27319
rect 6193 27285 6227 27319
rect 9413 27285 9447 27319
rect 11805 27285 11839 27319
rect 13737 27285 13771 27319
rect 15577 27285 15611 27319
rect 16313 27285 16347 27319
rect 17785 27285 17819 27319
rect 21097 27285 21131 27319
rect 1593 27081 1627 27115
rect 6653 27081 6687 27115
rect 8309 27081 8343 27115
rect 8953 27081 8987 27115
rect 11069 27081 11103 27115
rect 11897 27081 11931 27115
rect 15945 27081 15979 27115
rect 19625 27081 19659 27115
rect 20085 27081 20119 27115
rect 10517 27013 10551 27047
rect 13921 27013 13955 27047
rect 16037 27013 16071 27047
rect 16221 27013 16255 27047
rect 4261 26945 4295 26979
rect 6285 26945 6319 26979
rect 7205 26945 7239 26979
rect 13185 26945 13219 26979
rect 15577 26945 15611 26979
rect 17877 26945 17911 26979
rect 18337 26945 18371 26979
rect 4721 26877 4755 26911
rect 5181 26877 5215 26911
rect 5365 26877 5399 26911
rect 5733 26877 5767 26911
rect 5917 26877 5951 26911
rect 6929 26877 6963 26911
rect 9413 26877 9447 26911
rect 9582 26877 9616 26911
rect 10237 26877 10271 26911
rect 10333 26877 10367 26911
rect 12633 26877 12667 26911
rect 14105 26877 14139 26911
rect 14565 26877 14599 26911
rect 15025 26877 15059 26911
rect 15485 26877 15519 26911
rect 16037 26877 16071 26911
rect 16405 26877 16439 26911
rect 16497 26877 16531 26911
rect 17233 26877 17267 26911
rect 18061 26877 18095 26911
rect 4629 26809 4663 26843
rect 12449 26809 12483 26843
rect 12817 26809 12851 26843
rect 13645 26809 13679 26843
rect 16957 26809 16991 26843
rect 3801 26741 3835 26775
rect 9229 26741 9263 26775
rect 11529 26741 11563 26775
rect 12265 26741 12299 26775
rect 12725 26741 12759 26775
rect 8125 26537 8159 26571
rect 8769 26537 8803 26571
rect 9137 26537 9171 26571
rect 11897 26537 11931 26571
rect 12173 26537 12207 26571
rect 14105 26537 14139 26571
rect 14841 26537 14875 26571
rect 16221 26537 16255 26571
rect 16865 26537 16899 26571
rect 18889 26537 18923 26571
rect 3065 26469 3099 26503
rect 1409 26401 1443 26435
rect 5273 26401 5307 26435
rect 8585 26401 8619 26435
rect 10333 26401 10367 26435
rect 10517 26401 10551 26435
rect 10701 26401 10735 26435
rect 1685 26333 1719 26367
rect 5549 26333 5583 26367
rect 7757 26333 7791 26367
rect 9873 26333 9907 26367
rect 11069 26333 11103 26367
rect 11253 26333 11287 26367
rect 5089 26265 5123 26299
rect 7297 26265 7331 26299
rect 15853 26469 15887 26503
rect 17877 26469 17911 26503
rect 18153 26469 18187 26503
rect 18521 26469 18555 26503
rect 13093 26401 13127 26435
rect 13185 26401 13219 26435
rect 13461 26401 13495 26435
rect 15393 26401 15427 26435
rect 17417 26401 17451 26435
rect 13553 26333 13587 26367
rect 15301 26333 15335 26367
rect 17325 26333 17359 26367
rect 12541 26265 12575 26299
rect 4813 26197 4847 26231
rect 6653 26197 6687 26231
rect 8493 26197 8527 26231
rect 9413 26197 9447 26231
rect 12173 26197 12207 26231
rect 12265 26197 12299 26231
rect 14565 26197 14599 26231
rect 16589 26197 16623 26231
rect 1685 25993 1719 26027
rect 2053 25993 2087 26027
rect 6653 25993 6687 26027
rect 7205 25993 7239 26027
rect 8309 25993 8343 26027
rect 10701 25993 10735 26027
rect 11805 25993 11839 26027
rect 15761 25993 15795 26027
rect 17785 25993 17819 26027
rect 18337 25993 18371 26027
rect 18705 25993 18739 26027
rect 10149 25925 10183 25959
rect 12541 25925 12575 25959
rect 14289 25925 14323 25959
rect 4261 25857 4295 25891
rect 8493 25857 8527 25891
rect 10793 25857 10827 25891
rect 11529 25857 11563 25891
rect 13277 25857 13311 25891
rect 14381 25857 14415 25891
rect 15117 25857 15151 25891
rect 16405 25857 16439 25891
rect 4721 25789 4755 25823
rect 5181 25789 5215 25823
rect 5365 25789 5399 25823
rect 5733 25789 5767 25823
rect 5917 25789 5951 25823
rect 7941 25789 7975 25823
rect 8585 25789 8619 25823
rect 9137 25789 9171 25823
rect 9321 25789 9355 25823
rect 12173 25789 12207 25823
rect 12449 25789 12483 25823
rect 13001 25789 13035 25823
rect 16589 25789 16623 25823
rect 16957 25789 16991 25823
rect 17049 25789 17083 25823
rect 3893 25721 3927 25755
rect 7573 25721 7607 25755
rect 11069 25721 11103 25755
rect 11161 25721 11195 25755
rect 13921 25721 13955 25755
rect 14565 25721 14599 25755
rect 14749 25721 14783 25755
rect 4629 25653 4663 25687
rect 9597 25653 9631 25687
rect 10977 25653 11011 25687
rect 14657 25653 14691 25687
rect 15485 25653 15519 25687
rect 16221 25653 16255 25687
rect 17509 25653 17543 25687
rect 1685 25449 1719 25483
rect 5641 25449 5675 25483
rect 7021 25449 7055 25483
rect 9137 25449 9171 25483
rect 9505 25449 9539 25483
rect 9965 25449 9999 25483
rect 10885 25449 10919 25483
rect 11253 25449 11287 25483
rect 12909 25449 12943 25483
rect 14933 25449 14967 25483
rect 15577 25449 15611 25483
rect 16037 25449 16071 25483
rect 13461 25381 13495 25415
rect 14473 25381 14507 25415
rect 1409 25313 1443 25347
rect 1593 25313 1627 25347
rect 7113 25313 7147 25347
rect 10149 25313 10183 25347
rect 11713 25313 11747 25347
rect 11897 25313 11931 25347
rect 12081 25313 12115 25347
rect 12265 25313 12299 25347
rect 12633 25313 12667 25347
rect 16129 25313 16163 25347
rect 7389 25245 7423 25279
rect 13829 25245 13863 25279
rect 13921 25245 13955 25279
rect 16405 25245 16439 25279
rect 5273 25177 5307 25211
rect 4813 25109 4847 25143
rect 8493 25109 8527 25143
rect 10333 25109 10367 25143
rect 13369 25109 13403 25143
rect 13599 25109 13633 25143
rect 13737 25109 13771 25143
rect 17509 25109 17543 25143
rect 10793 24905 10827 24939
rect 11897 24905 11931 24939
rect 16221 24905 16255 24939
rect 16589 24905 16623 24939
rect 17325 24905 17359 24939
rect 17693 24905 17727 24939
rect 9137 24837 9171 24871
rect 6653 24769 6687 24803
rect 8125 24769 8159 24803
rect 9689 24769 9723 24803
rect 10609 24769 10643 24803
rect 7389 24701 7423 24735
rect 8033 24701 8067 24735
rect 8401 24701 8435 24735
rect 8585 24701 8619 24735
rect 9505 24701 9539 24735
rect 10517 24701 10551 24735
rect 1685 24633 1719 24667
rect 7297 24633 7331 24667
rect 9781 24633 9815 24667
rect 12265 24769 12299 24803
rect 13369 24769 13403 24803
rect 14289 24769 14323 24803
rect 11437 24701 11471 24735
rect 12909 24701 12943 24735
rect 13277 24701 13311 24735
rect 14197 24701 14231 24735
rect 14933 24701 14967 24735
rect 16037 24701 16071 24735
rect 18061 24701 18095 24735
rect 18521 24701 18555 24735
rect 12449 24633 12483 24667
rect 15669 24633 15703 24667
rect 1961 24565 1995 24599
rect 6285 24565 6319 24599
rect 10793 24565 10827 24599
rect 11069 24565 11103 24599
rect 13737 24565 13771 24599
rect 15393 24565 15427 24599
rect 16865 24565 16899 24599
rect 18245 24565 18279 24599
rect 7113 24361 7147 24395
rect 7849 24361 7883 24395
rect 9873 24361 9907 24395
rect 10517 24361 10551 24395
rect 11253 24361 11287 24395
rect 12541 24361 12575 24395
rect 12817 24361 12851 24395
rect 14933 24361 14967 24395
rect 15485 24361 15519 24395
rect 17049 24361 17083 24395
rect 18061 24361 18095 24395
rect 7481 24293 7515 24327
rect 11897 24293 11931 24327
rect 15577 24293 15611 24327
rect 15669 24293 15703 24327
rect 11437 24225 11471 24259
rect 13001 24225 13035 24259
rect 13185 24225 13219 24259
rect 13553 24225 13587 24259
rect 16865 24225 16899 24259
rect 17877 24225 17911 24259
rect 11345 24157 11379 24191
rect 15301 24157 15335 24191
rect 16037 24157 16071 24191
rect 9505 24089 9539 24123
rect 16405 24089 16439 24123
rect 16773 24089 16807 24123
rect 10885 24021 10919 24055
rect 14197 24021 14231 24055
rect 14565 24021 14599 24055
rect 7113 23817 7147 23851
rect 8585 23817 8619 23851
rect 10333 23817 10367 23851
rect 10701 23817 10735 23851
rect 13369 23817 13403 23851
rect 15853 23817 15887 23851
rect 16957 23817 16991 23851
rect 18337 23817 18371 23851
rect 11069 23749 11103 23783
rect 16497 23749 16531 23783
rect 13001 23681 13035 23715
rect 8769 23613 8803 23647
rect 11437 23613 11471 23647
rect 12265 23613 12299 23647
rect 12449 23613 12483 23647
rect 12541 23613 12575 23647
rect 13921 23613 13955 23647
rect 14289 23613 14323 23647
rect 14657 23613 14691 23647
rect 14841 23613 14875 23647
rect 15209 23613 15243 23647
rect 16313 23613 16347 23647
rect 8677 23545 8711 23579
rect 11805 23477 11839 23511
rect 14289 23477 14323 23511
rect 16221 23477 16255 23511
rect 8769 23273 8803 23307
rect 11437 23273 11471 23307
rect 11897 23273 11931 23307
rect 12081 23273 12115 23307
rect 14473 23273 14507 23307
rect 15117 23273 15151 23307
rect 18153 23273 18187 23307
rect 10149 23205 10183 23239
rect 15485 23205 15519 23239
rect 15669 23205 15703 23239
rect 16037 23205 16071 23239
rect 6837 23137 6871 23171
rect 7205 23137 7239 23171
rect 7389 23137 7423 23171
rect 8585 23137 8619 23171
rect 10977 23137 11011 23171
rect 11989 23137 12023 23171
rect 12817 23137 12851 23171
rect 13001 23137 13035 23171
rect 13921 23137 13955 23171
rect 15577 23137 15611 23171
rect 6193 23069 6227 23103
rect 6929 23069 6963 23103
rect 10701 23069 10735 23103
rect 11161 23069 11195 23103
rect 15301 23069 15335 23103
rect 13829 23001 13863 23035
rect 7757 22933 7791 22967
rect 13369 22933 13403 22967
rect 14105 22933 14139 22967
rect 16405 22933 16439 22967
rect 5917 22729 5951 22763
rect 8217 22729 8251 22763
rect 9873 22729 9907 22763
rect 10241 22729 10275 22763
rect 11713 22729 11747 22763
rect 13369 22729 13403 22763
rect 15301 22729 15335 22763
rect 6285 22661 6319 22695
rect 6653 22661 6687 22695
rect 11989 22661 12023 22695
rect 13737 22661 13771 22695
rect 16129 22661 16163 22695
rect 6837 22593 6871 22627
rect 7113 22593 7147 22627
rect 12449 22593 12483 22627
rect 14933 22593 14967 22627
rect 17877 22593 17911 22627
rect 18337 22593 18371 22627
rect 26065 22593 26099 22627
rect 26433 22593 26467 22627
rect 8861 22525 8895 22559
rect 9229 22525 9263 22559
rect 9321 22525 9355 22559
rect 10333 22525 10367 22559
rect 11161 22525 11195 22559
rect 12541 22525 12575 22559
rect 14105 22525 14139 22559
rect 14289 22525 14323 22559
rect 14657 22525 14691 22559
rect 15577 22525 15611 22559
rect 16405 22525 16439 22559
rect 18061 22525 18095 22559
rect 26157 22525 26191 22559
rect 10885 22457 10919 22491
rect 13001 22457 13035 22491
rect 5549 22389 5583 22423
rect 9505 22389 9539 22423
rect 10517 22389 10551 22423
rect 15577 22389 15611 22423
rect 15669 22389 15703 22423
rect 16773 22389 16807 22423
rect 19441 22389 19475 22423
rect 27721 22389 27755 22423
rect 13001 22185 13035 22219
rect 14105 22185 14139 22219
rect 14473 22185 14507 22219
rect 17049 22185 17083 22219
rect 26157 22185 26191 22219
rect 6101 22049 6135 22083
rect 8585 22049 8619 22083
rect 12173 22049 12207 22083
rect 13277 22049 13311 22083
rect 15393 22049 15427 22083
rect 16865 22049 16899 22083
rect 18981 22049 19015 22083
rect 19349 22049 19383 22083
rect 6377 21981 6411 22015
rect 9505 21981 9539 22015
rect 9689 21981 9723 22015
rect 9965 21981 9999 22015
rect 13185 21981 13219 22015
rect 15301 21981 15335 22015
rect 16129 21981 16163 22015
rect 18429 21981 18463 22015
rect 19073 21981 19107 22015
rect 19257 21981 19291 22015
rect 12357 21913 12391 21947
rect 7665 21845 7699 21879
rect 8769 21845 8803 21879
rect 11253 21845 11287 21879
rect 12081 21845 12115 21879
rect 12725 21845 12759 21879
rect 13461 21845 13495 21879
rect 15577 21845 15611 21879
rect 16681 21845 16715 21879
rect 18153 21845 18187 21879
rect 8585 21641 8619 21675
rect 9781 21641 9815 21675
rect 10793 21641 10827 21675
rect 11897 21641 11931 21675
rect 13829 21641 13863 21675
rect 17417 21641 17451 21675
rect 17693 21641 17727 21675
rect 19349 21641 19383 21675
rect 5917 21573 5951 21607
rect 9137 21573 9171 21607
rect 6653 21505 6687 21539
rect 7389 21505 7423 21539
rect 12265 21505 12299 21539
rect 14565 21505 14599 21539
rect 16221 21505 16255 21539
rect 16589 21505 16623 21539
rect 7573 21437 7607 21471
rect 7941 21437 7975 21471
rect 8033 21437 8067 21471
rect 8953 21437 8987 21471
rect 10149 21437 10183 21471
rect 10701 21437 10735 21471
rect 10977 21437 11011 21471
rect 11069 21437 11103 21471
rect 12541 21437 12575 21471
rect 13277 21437 13311 21471
rect 13461 21437 13495 21471
rect 14657 21437 14691 21471
rect 16497 21437 16531 21471
rect 16681 21437 16715 21471
rect 17141 21437 17175 21471
rect 6929 21369 6963 21403
rect 11529 21369 11563 21403
rect 14473 21369 14507 21403
rect 17877 21505 17911 21539
rect 18061 21505 18095 21539
rect 18521 21437 18555 21471
rect 18705 21437 18739 21471
rect 18889 21437 18923 21471
rect 19717 21369 19751 21403
rect 6285 21301 6319 21335
rect 9965 21301 9999 21335
rect 10517 21301 10551 21335
rect 10701 21301 10735 21335
rect 12541 21301 12575 21335
rect 15577 21301 15611 21335
rect 16313 21301 16347 21335
rect 17693 21301 17727 21335
rect 6193 21097 6227 21131
rect 6929 21097 6963 21131
rect 7389 21097 7423 21131
rect 8953 21097 8987 21131
rect 9505 21097 9539 21131
rect 9873 21097 9907 21131
rect 10885 21097 10919 21131
rect 13093 21097 13127 21131
rect 14381 21097 14415 21131
rect 15945 21097 15979 21131
rect 17785 21097 17819 21131
rect 18429 21097 18463 21131
rect 3157 21029 3191 21063
rect 12541 21029 12575 21063
rect 14105 21029 14139 21063
rect 18705 21029 18739 21063
rect 1777 20961 1811 20995
rect 9689 20961 9723 20995
rect 11069 20961 11103 20995
rect 11161 20961 11195 20995
rect 12817 20961 12851 20995
rect 13001 20961 13035 20995
rect 14197 20961 14231 20995
rect 15393 20961 15427 20995
rect 22661 20961 22695 20995
rect 1501 20893 1535 20927
rect 16405 20893 16439 20927
rect 16681 20893 16715 20927
rect 22385 20893 22419 20927
rect 10425 20825 10459 20859
rect 12081 20825 12115 20859
rect 14749 20825 14783 20859
rect 11345 20757 11379 20791
rect 13645 20757 13679 20791
rect 15025 20757 15059 20791
rect 15577 20757 15611 20791
rect 16313 20757 16347 20791
rect 19165 20757 19199 20791
rect 23765 20757 23799 20791
rect 2053 20553 2087 20587
rect 9413 20553 9447 20587
rect 10149 20553 10183 20587
rect 11621 20553 11655 20587
rect 12265 20553 12299 20587
rect 15485 20553 15519 20587
rect 17785 20553 17819 20587
rect 22845 20553 22879 20587
rect 12817 20485 12851 20519
rect 13277 20485 13311 20519
rect 18337 20485 18371 20519
rect 10885 20417 10919 20451
rect 16405 20417 16439 20451
rect 16773 20417 16807 20451
rect 11161 20349 11195 20383
rect 11345 20349 11379 20383
rect 13277 20349 13311 20383
rect 13645 20349 13679 20383
rect 13829 20349 13863 20383
rect 14197 20349 14231 20383
rect 14565 20349 14599 20383
rect 16497 20349 16531 20383
rect 16865 20349 16899 20383
rect 17509 20349 17543 20383
rect 18521 20349 18555 20383
rect 18705 20349 18739 20383
rect 18889 20349 18923 20383
rect 10333 20281 10367 20315
rect 15853 20281 15887 20315
rect 1593 20213 1627 20247
rect 9781 20213 9815 20247
rect 22385 20213 22419 20247
rect 7481 20009 7515 20043
rect 9965 20009 9999 20043
rect 10425 20009 10459 20043
rect 14197 20009 14231 20043
rect 14473 20009 14507 20043
rect 15485 20009 15519 20043
rect 15945 20009 15979 20043
rect 8769 19941 8803 19975
rect 10793 19941 10827 19975
rect 12081 19941 12115 19975
rect 13185 19941 13219 19975
rect 19533 19941 19567 19975
rect 8217 19873 8251 19907
rect 8309 19873 8343 19907
rect 11253 19873 11287 19907
rect 11621 19873 11655 19907
rect 12725 19873 12759 19907
rect 13461 19873 13495 19907
rect 14013 19873 14047 19907
rect 15301 19873 15335 19907
rect 19073 19873 19107 19907
rect 11713 19805 11747 19839
rect 12633 19805 12667 19839
rect 16497 19805 16531 19839
rect 16773 19805 16807 19839
rect 18429 19805 18463 19839
rect 18981 19805 19015 19839
rect 12541 19737 12575 19771
rect 7849 19669 7883 19703
rect 13829 19669 13863 19703
rect 14841 19669 14875 19703
rect 16313 19669 16347 19703
rect 18061 19669 18095 19703
rect 8953 19465 8987 19499
rect 11437 19465 11471 19499
rect 11897 19465 11931 19499
rect 14013 19465 14047 19499
rect 15393 19465 15427 19499
rect 16865 19465 16899 19499
rect 18337 19465 18371 19499
rect 18981 19465 19015 19499
rect 11069 19397 11103 19431
rect 8125 19329 8159 19363
rect 10057 19329 10091 19363
rect 12449 19329 12483 19363
rect 15485 19329 15519 19363
rect 7297 19261 7331 19295
rect 8033 19261 8067 19295
rect 8401 19261 8435 19295
rect 8585 19261 8619 19295
rect 9321 19261 9355 19295
rect 10149 19261 10183 19295
rect 10517 19261 10551 19295
rect 10609 19261 10643 19295
rect 12909 19261 12943 19295
rect 13093 19261 13127 19295
rect 13277 19261 13311 19295
rect 14473 19261 14507 19295
rect 14749 19261 14783 19295
rect 15761 19261 15795 19295
rect 18061 19261 18095 19295
rect 18153 19261 18187 19295
rect 19349 19261 19383 19295
rect 12265 19193 12299 19227
rect 6653 19125 6687 19159
rect 7665 19125 7699 19159
rect 9781 19125 9815 19159
rect 14657 19125 14691 19159
rect 14749 19125 14783 19159
rect 15025 19125 15059 19159
rect 17417 19125 17451 19159
rect 17785 19125 17819 19159
rect 8493 18921 8527 18955
rect 9965 18921 9999 18955
rect 10793 18921 10827 18955
rect 12633 18921 12667 18955
rect 14013 18921 14047 18955
rect 14841 18921 14875 18955
rect 15761 18921 15795 18955
rect 16313 18921 16347 18955
rect 18153 18921 18187 18955
rect 12541 18853 12575 18887
rect 7389 18785 7423 18819
rect 11345 18785 11379 18819
rect 11713 18785 11747 18819
rect 7113 18717 7147 18751
rect 11437 18717 11471 18751
rect 11621 18717 11655 18751
rect 13553 18785 13587 18819
rect 15945 18785 15979 18819
rect 16957 18785 16991 18819
rect 12725 18717 12759 18751
rect 13277 18717 13311 18751
rect 13737 18717 13771 18751
rect 16865 18717 16899 18751
rect 12633 18649 12667 18683
rect 14381 18649 14415 18683
rect 9413 18581 9447 18615
rect 10241 18581 10275 18615
rect 16681 18581 16715 18615
rect 17141 18581 17175 18615
rect 17693 18581 17727 18615
rect 3249 18377 3283 18411
rect 7573 18377 7607 18411
rect 9229 18377 9263 18411
rect 11069 18377 11103 18411
rect 12173 18377 12207 18411
rect 14381 18377 14415 18411
rect 16313 18377 16347 18411
rect 17049 18377 17083 18411
rect 17325 18377 17359 18411
rect 17693 18377 17727 18411
rect 7205 18309 7239 18343
rect 11805 18309 11839 18343
rect 16681 18309 16715 18343
rect 9781 18241 9815 18275
rect 10333 18241 10367 18275
rect 10793 18241 10827 18275
rect 13001 18241 13035 18275
rect 13737 18241 13771 18275
rect 15025 18241 15059 18275
rect 1869 18173 1903 18207
rect 2145 18173 2179 18207
rect 8953 18173 8987 18207
rect 10609 18173 10643 18207
rect 12449 18173 12483 18207
rect 13277 18173 13311 18207
rect 13461 18173 13495 18207
rect 14841 18173 14875 18207
rect 15209 18173 15243 18207
rect 15393 18173 15427 18207
rect 15761 18173 15795 18207
rect 16865 18173 16899 18207
rect 11529 18105 11563 18139
rect 1685 18037 1719 18071
rect 9689 18037 9723 18071
rect 8309 17833 8343 17867
rect 9137 17833 9171 17867
rect 11621 17833 11655 17867
rect 12265 17833 12299 17867
rect 13553 17833 13587 17867
rect 14657 17833 14691 17867
rect 15577 17833 15611 17867
rect 16773 17833 16807 17867
rect 18705 17833 18739 17867
rect 10333 17765 10367 17799
rect 11161 17697 11195 17731
rect 12541 17697 12575 17731
rect 13093 17697 13127 17731
rect 13277 17697 13311 17731
rect 15117 17697 15151 17731
rect 15945 17697 15979 17731
rect 16313 17697 16347 17731
rect 17601 17697 17635 17731
rect 9413 17629 9447 17663
rect 10885 17629 10919 17663
rect 11345 17629 11379 17663
rect 12357 17629 12391 17663
rect 14197 17629 14231 17663
rect 15761 17629 15795 17663
rect 16221 17629 16255 17663
rect 17325 17629 17359 17663
rect 10241 17561 10275 17595
rect 1961 17493 1995 17527
rect 17233 17493 17267 17527
rect 2789 17289 2823 17323
rect 8493 17289 8527 17323
rect 9873 17289 9907 17323
rect 11897 17289 11931 17323
rect 12265 17289 12299 17323
rect 14013 17289 14047 17323
rect 15301 17289 15335 17323
rect 15761 17289 15795 17323
rect 16221 17289 16255 17323
rect 10149 17221 10183 17255
rect 1685 17153 1719 17187
rect 8953 17153 8987 17187
rect 9137 17153 9171 17187
rect 10793 17153 10827 17187
rect 11253 17153 11287 17187
rect 14197 17153 14231 17187
rect 16313 17153 16347 17187
rect 16865 17153 16899 17187
rect 1409 17085 1443 17119
rect 8861 17085 8895 17119
rect 9229 17085 9263 17119
rect 10977 17085 11011 17119
rect 11345 17085 11379 17119
rect 12725 17085 12759 17119
rect 13645 17085 13679 17119
rect 14289 17085 14323 17119
rect 14841 17085 14875 17119
rect 15025 17085 15059 17119
rect 16405 17085 16439 17119
rect 17417 17085 17451 17119
rect 7757 17017 7791 17051
rect 13277 17017 13311 17051
rect 8125 16949 8159 16983
rect 10609 16949 10643 16983
rect 17785 16949 17819 16983
rect 1685 16745 1719 16779
rect 8309 16745 8343 16779
rect 9505 16745 9539 16779
rect 10333 16745 10367 16779
rect 12449 16745 12483 16779
rect 14749 16745 14783 16779
rect 15577 16745 15611 16779
rect 16681 16745 16715 16779
rect 23673 16745 23707 16779
rect 7757 16677 7791 16711
rect 10057 16677 10091 16711
rect 10701 16677 10735 16711
rect 12081 16677 12115 16711
rect 13185 16677 13219 16711
rect 15025 16677 15059 16711
rect 6377 16609 6411 16643
rect 11253 16609 11287 16643
rect 11529 16609 11563 16643
rect 12817 16609 12851 16643
rect 13829 16609 13863 16643
rect 14105 16609 14139 16643
rect 15485 16609 15519 16643
rect 15853 16609 15887 16643
rect 16129 16609 16163 16643
rect 17233 16609 17267 16643
rect 22293 16609 22327 16643
rect 6101 16541 6135 16575
rect 11713 16541 11747 16575
rect 13461 16541 13495 16575
rect 14381 16541 14415 16575
rect 22569 16541 22603 16575
rect 2053 16405 2087 16439
rect 17417 16405 17451 16439
rect 4997 16201 5031 16235
rect 6561 16201 6595 16235
rect 7849 16201 7883 16235
rect 9689 16201 9723 16235
rect 10977 16201 11011 16235
rect 14013 16201 14047 16235
rect 16405 16201 16439 16235
rect 16773 16201 16807 16235
rect 17325 16201 17359 16235
rect 19625 16201 19659 16235
rect 10609 16133 10643 16167
rect 16037 16133 16071 16167
rect 3341 16065 3375 16099
rect 8217 16065 8251 16099
rect 3433 15997 3467 16031
rect 3709 15997 3743 16031
rect 8309 15997 8343 16031
rect 8585 15997 8619 16031
rect 10793 15997 10827 16031
rect 11621 15997 11655 16031
rect 12265 15997 12299 16031
rect 12909 15997 12943 16031
rect 14657 15997 14691 16031
rect 15117 15997 15151 16031
rect 15577 15997 15611 16031
rect 15853 15997 15887 16031
rect 18061 15997 18095 16031
rect 18337 15997 18371 16031
rect 10333 15929 10367 15963
rect 13369 15929 13403 15963
rect 13645 15929 13679 15963
rect 14473 15929 14507 15963
rect 6101 15861 6135 15895
rect 11345 15861 11379 15895
rect 17785 15861 17819 15895
rect 22385 15861 22419 15895
rect 22753 15861 22787 15895
rect 3525 15657 3559 15691
rect 6653 15657 6687 15691
rect 10057 15657 10091 15691
rect 10425 15657 10459 15691
rect 12541 15657 12575 15691
rect 14197 15657 14231 15691
rect 15117 15657 15151 15691
rect 8677 15589 8711 15623
rect 14657 15589 14691 15623
rect 15485 15589 15519 15623
rect 6837 15521 6871 15555
rect 7297 15521 7331 15555
rect 9873 15521 9907 15555
rect 13185 15521 13219 15555
rect 13277 15521 13311 15555
rect 13645 15521 13679 15555
rect 13737 15521 13771 15555
rect 16221 15521 16255 15555
rect 7021 15453 7055 15487
rect 15945 15453 15979 15487
rect 18061 15453 18095 15487
rect 12909 15317 12943 15351
rect 17325 15317 17359 15351
rect 6653 15113 6687 15147
rect 7113 15113 7147 15147
rect 7849 15113 7883 15147
rect 10333 15113 10367 15147
rect 12265 15113 12299 15147
rect 13553 15113 13587 15147
rect 13829 15113 13863 15147
rect 13921 15113 13955 15147
rect 16037 15113 16071 15147
rect 8217 14977 8251 15011
rect 8585 14977 8619 15011
rect 13277 14977 13311 15011
rect 15209 15045 15243 15079
rect 16497 14977 16531 15011
rect 8309 14909 8343 14943
rect 10793 14909 10827 14943
rect 11253 14909 11287 14943
rect 11897 14909 11931 14943
rect 12633 14909 12667 14943
rect 13829 14909 13863 14943
rect 14289 14909 14323 14943
rect 14381 14909 14415 14943
rect 14749 14909 14783 14943
rect 14841 14909 14875 14943
rect 16589 14909 16623 14943
rect 16681 14909 16715 14943
rect 17141 14841 17175 14875
rect 7389 14773 7423 14807
rect 9689 14773 9723 14807
rect 10977 14773 11011 14807
rect 17417 14773 17451 14807
rect 7481 14569 7515 14603
rect 10149 14569 10183 14603
rect 11161 14569 11195 14603
rect 14473 14569 14507 14603
rect 7573 14501 7607 14535
rect 12265 14501 12299 14535
rect 13737 14501 13771 14535
rect 14197 14501 14231 14535
rect 8217 14433 8251 14467
rect 8585 14433 8619 14467
rect 9965 14433 9999 14467
rect 10977 14433 11011 14467
rect 12633 14433 12667 14467
rect 13093 14433 13127 14467
rect 13185 14433 13219 14467
rect 17141 14433 17175 14467
rect 17325 14433 17359 14467
rect 17509 14433 17543 14467
rect 8125 14365 8159 14399
rect 8493 14365 8527 14399
rect 12449 14365 12483 14399
rect 14933 14365 14967 14399
rect 16957 14297 16991 14331
rect 9137 14229 9171 14263
rect 15945 14229 15979 14263
rect 7297 14025 7331 14059
rect 9965 14025 9999 14059
rect 10701 14025 10735 14059
rect 11345 14025 11379 14059
rect 12909 14025 12943 14059
rect 13553 14025 13587 14059
rect 14289 14025 14323 14059
rect 15393 14025 15427 14059
rect 17141 14025 17175 14059
rect 17417 14025 17451 14059
rect 7665 13957 7699 13991
rect 16773 13957 16807 13991
rect 9321 13889 9355 13923
rect 11897 13889 11931 13923
rect 15577 13889 15611 13923
rect 26065 13889 26099 13923
rect 27629 13889 27663 13923
rect 8401 13821 8435 13855
rect 8861 13821 8895 13855
rect 9045 13821 9079 13855
rect 9413 13821 9447 13855
rect 10517 13821 10551 13855
rect 12173 13821 12207 13855
rect 12817 13821 12851 13855
rect 13921 13821 13955 13855
rect 14657 13821 14691 13855
rect 15669 13821 15703 13855
rect 26157 13821 26191 13855
rect 26433 13821 26467 13855
rect 8309 13753 8343 13787
rect 10977 13685 11011 13719
rect 7849 13481 7883 13515
rect 8769 13481 8803 13515
rect 13001 13481 13035 13515
rect 22569 13481 22603 13515
rect 26249 13481 26283 13515
rect 8493 13413 8527 13447
rect 7481 13345 7515 13379
rect 10701 13345 10735 13379
rect 12265 13345 12299 13379
rect 13553 13345 13587 13379
rect 21189 13345 21223 13379
rect 12173 13277 12207 13311
rect 21465 13277 21499 13311
rect 13737 13209 13771 13243
rect 7297 13141 7331 13175
rect 11069 13141 11103 13175
rect 12449 13141 12483 13175
rect 7389 12937 7423 12971
rect 10057 12937 10091 12971
rect 10701 12937 10735 12971
rect 12173 12937 12207 12971
rect 13921 12937 13955 12971
rect 21281 12937 21315 12971
rect 21649 12937 21683 12971
rect 13553 12869 13587 12903
rect 8585 12801 8619 12835
rect 8953 12801 8987 12835
rect 8677 12733 8711 12767
rect 11161 12733 11195 12767
rect 11621 12733 11655 12767
rect 12449 12733 12483 12767
rect 12909 12733 12943 12767
rect 11345 12597 11379 12631
rect 12633 12597 12667 12631
rect 12541 12393 12575 12427
rect 12817 12393 12851 12427
rect 9781 12257 9815 12291
rect 11621 12257 11655 12291
rect 11805 12257 11839 12291
rect 11989 12257 12023 12291
rect 13185 12257 13219 12291
rect 13277 12257 13311 12291
rect 13645 12257 13679 12291
rect 13737 12257 13771 12291
rect 16221 12257 16255 12291
rect 11437 12121 11471 12155
rect 16037 12121 16071 12155
rect 8677 12053 8711 12087
rect 9965 12053 9999 12087
rect 10425 12053 10459 12087
rect 14197 12053 14231 12087
rect 15577 12053 15611 12087
rect 15853 12053 15887 12087
rect 9137 11849 9171 11883
rect 9505 11849 9539 11883
rect 9873 11849 9907 11883
rect 11713 11849 11747 11883
rect 14105 11849 14139 11883
rect 14933 11849 14967 11883
rect 15393 11849 15427 11883
rect 16957 11849 16991 11883
rect 10149 11781 10183 11815
rect 14473 11781 14507 11815
rect 12173 11713 12207 11747
rect 15577 11713 15611 11747
rect 16037 11713 16071 11747
rect 9321 11645 9355 11679
rect 10793 11645 10827 11679
rect 10977 11645 11011 11679
rect 11161 11645 11195 11679
rect 12449 11645 12483 11679
rect 12633 11645 12667 11679
rect 13093 11645 13127 11679
rect 13185 11645 13219 11679
rect 15761 11645 15795 11679
rect 16129 11645 16163 11679
rect 10333 11577 10367 11611
rect 13737 11577 13771 11611
rect 16589 11577 16623 11611
rect 10425 11305 10459 11339
rect 11621 11305 11655 11339
rect 12081 11305 12115 11339
rect 12449 11305 12483 11339
rect 12817 11305 12851 11339
rect 14657 11305 14691 11339
rect 16681 11305 16715 11339
rect 17785 11305 17819 11339
rect 11345 11237 11379 11271
rect 8033 11169 8067 11203
rect 10885 11169 10919 11203
rect 13185 11169 13219 11203
rect 13645 11169 13679 11203
rect 13737 11169 13771 11203
rect 15577 11169 15611 11203
rect 17969 11169 18003 11203
rect 10793 11101 10827 11135
rect 13001 11101 13035 11135
rect 14289 11101 14323 11135
rect 15301 11101 15335 11135
rect 7849 11033 7883 11067
rect 7849 10761 7883 10795
rect 10793 10761 10827 10795
rect 11253 10761 11287 10795
rect 13093 10761 13127 10795
rect 15393 10761 15427 10795
rect 17877 10761 17911 10795
rect 20821 10761 20855 10795
rect 13369 10693 13403 10727
rect 13737 10693 13771 10727
rect 19257 10625 19291 10659
rect 19533 10557 19567 10591
rect 19073 10489 19107 10523
rect 12725 10421 12759 10455
rect 15669 10421 15703 10455
rect 18797 10217 18831 10251
rect 19257 10217 19291 10251
rect 16405 10081 16439 10115
rect 18981 10081 19015 10115
rect 16313 10013 16347 10047
rect 16589 9877 16623 9911
rect 12817 9673 12851 9707
rect 18797 9673 18831 9707
rect 15025 9537 15059 9571
rect 15485 9537 15519 9571
rect 16865 9537 16899 9571
rect 17509 9537 17543 9571
rect 12265 9469 12299 9503
rect 12541 9469 12575 9503
rect 12633 9469 12667 9503
rect 13461 9469 13495 9503
rect 13921 9469 13955 9503
rect 14473 9469 14507 9503
rect 15209 9469 15243 9503
rect 17141 9469 17175 9503
rect 14105 9333 14139 9367
rect 3065 9061 3099 9095
rect 1409 8993 1443 9027
rect 9689 8993 9723 9027
rect 9965 8993 9999 9027
rect 12633 8993 12667 9027
rect 13001 8993 13035 9027
rect 13093 8993 13127 9027
rect 16681 8993 16715 9027
rect 16865 8993 16899 9027
rect 17049 8993 17083 9027
rect 1685 8925 1719 8959
rect 12173 8925 12207 8959
rect 16497 8857 16531 8891
rect 9137 8789 9171 8823
rect 11069 8789 11103 8823
rect 13553 8789 13587 8823
rect 15485 8789 15519 8823
rect 2053 8585 2087 8619
rect 8861 8585 8895 8619
rect 10517 8585 10551 8619
rect 12173 8585 12207 8619
rect 12633 8585 12667 8619
rect 16589 8585 16623 8619
rect 16957 8585 16991 8619
rect 8585 8517 8619 8551
rect 11805 8517 11839 8551
rect 16313 8517 16347 8551
rect 13737 8449 13771 8483
rect 14013 8449 14047 8483
rect 14381 8449 14415 8483
rect 9505 8381 9539 8415
rect 9689 8381 9723 8415
rect 10028 8381 10062 8415
rect 10241 8381 10275 8415
rect 13277 8381 13311 8415
rect 14105 8381 14139 8415
rect 14473 8381 14507 8415
rect 1593 8313 1627 8347
rect 9045 8313 9079 8347
rect 9137 8041 9171 8075
rect 9873 8041 9907 8075
rect 12449 8041 12483 8075
rect 13829 8041 13863 8075
rect 18153 8041 18187 8075
rect 13553 7973 13587 8007
rect 11069 7905 11103 7939
rect 11345 7905 11379 7939
rect 16865 7905 16899 7939
rect 16589 7837 16623 7871
rect 11161 7497 11195 7531
rect 14473 7497 14507 7531
rect 16681 7497 16715 7531
rect 17049 7497 17083 7531
rect 11437 7429 11471 7463
rect 13001 7361 13035 7395
rect 13369 7361 13403 7395
rect 13093 7293 13127 7327
rect 13093 6613 13127 6647
rect 14565 6613 14599 6647
rect 14381 6409 14415 6443
rect 14841 6273 14875 6307
rect 14565 6205 14599 6239
rect 15945 6069 15979 6103
rect 13829 5729 13863 5763
rect 14197 5729 14231 5763
rect 14381 5729 14415 5763
rect 15945 5729 15979 5763
rect 16313 5729 16347 5763
rect 16405 5729 16439 5763
rect 13921 5661 13955 5695
rect 15761 5661 15795 5695
rect 13093 5525 13127 5559
rect 13461 5525 13495 5559
rect 15577 5525 15611 5559
rect 12173 5321 12207 5355
rect 13001 5321 13035 5355
rect 15301 5321 15335 5355
rect 15669 5321 15703 5355
rect 16037 5321 16071 5355
rect 13093 5117 13127 5151
rect 13369 5117 13403 5151
rect 14473 4981 14507 5015
rect 13645 4777 13679 4811
rect 14013 4777 14047 4811
rect 15577 4777 15611 4811
rect 12633 4709 12667 4743
rect 10977 4641 11011 4675
rect 11253 4641 11287 4675
rect 13277 4641 13311 4675
rect 11345 4097 11379 4131
rect 11069 3961 11103 3995
rect 9965 3689 9999 3723
rect 11805 3689 11839 3723
rect 19441 3689 19475 3723
rect 10425 3553 10459 3587
rect 17877 3553 17911 3587
rect 10701 3485 10735 3519
rect 18153 3485 18187 3519
rect 11437 3145 11471 3179
rect 18245 3145 18279 3179
rect 18613 3077 18647 3111
rect 9781 3009 9815 3043
rect 10149 3009 10183 3043
rect 9873 2941 9907 2975
rect 10793 2601 10827 2635
rect 14013 2601 14047 2635
rect 17785 2601 17819 2635
rect 20545 2601 20579 2635
rect 12909 2465 12943 2499
rect 18153 2465 18187 2499
rect 21741 2465 21775 2499
rect 12081 2397 12115 2431
rect 12633 2397 12667 2431
rect 18337 2397 18371 2431
rect 18613 2397 18647 2431
rect 21465 2397 21499 2431
rect 20913 2329 20947 2363
rect 10517 2261 10551 2295
rect 12449 2261 12483 2295
rect 19717 2261 19751 2295
rect 23029 2261 23063 2295
<< metal1 >>
rect 1104 77818 28888 77840
rect 1104 77766 10982 77818
rect 11034 77766 11046 77818
rect 11098 77766 11110 77818
rect 11162 77766 11174 77818
rect 11226 77766 20982 77818
rect 21034 77766 21046 77818
rect 21098 77766 21110 77818
rect 21162 77766 21174 77818
rect 21226 77766 28888 77818
rect 1104 77744 28888 77766
rect 3326 77324 3332 77376
rect 3384 77364 3390 77376
rect 10318 77364 10324 77376
rect 3384 77336 10324 77364
rect 3384 77324 3390 77336
rect 10318 77324 10324 77336
rect 10376 77324 10382 77376
rect 13814 77364 13820 77376
rect 13775 77336 13820 77364
rect 13814 77324 13820 77336
rect 13872 77324 13878 77376
rect 23842 77324 23848 77376
rect 23900 77364 23906 77376
rect 25866 77364 25872 77376
rect 23900 77336 25872 77364
rect 23900 77324 23906 77336
rect 25866 77324 25872 77336
rect 25924 77324 25930 77376
rect 1104 77274 28888 77296
rect 1104 77222 5982 77274
rect 6034 77222 6046 77274
rect 6098 77222 6110 77274
rect 6162 77222 6174 77274
rect 6226 77222 15982 77274
rect 16034 77222 16046 77274
rect 16098 77222 16110 77274
rect 16162 77222 16174 77274
rect 16226 77222 25982 77274
rect 26034 77222 26046 77274
rect 26098 77222 26110 77274
rect 26162 77222 26174 77274
rect 26226 77222 28888 77274
rect 1104 77200 28888 77222
rect 17494 77120 17500 77172
rect 17552 77160 17558 77172
rect 19153 77163 19211 77169
rect 19153 77160 19165 77163
rect 17552 77132 19165 77160
rect 17552 77120 17558 77132
rect 19153 77129 19165 77132
rect 19199 77129 19211 77163
rect 19153 77123 19211 77129
rect 13725 77027 13783 77033
rect 13725 76993 13737 77027
rect 13771 77024 13783 77027
rect 14093 77027 14151 77033
rect 14093 77024 14105 77027
rect 13771 76996 14105 77024
rect 13771 76993 13783 76996
rect 13725 76987 13783 76993
rect 14093 76993 14105 76996
rect 14139 77024 14151 77027
rect 14274 77024 14280 77036
rect 14139 76996 14280 77024
rect 14139 76993 14151 76996
rect 14093 76987 14151 76993
rect 14274 76984 14280 76996
rect 14332 76984 14338 77036
rect 19168 77024 19196 77123
rect 19613 77027 19671 77033
rect 19613 77024 19625 77027
rect 19168 76996 19625 77024
rect 19613 76993 19625 76996
rect 19659 76993 19671 77027
rect 19613 76987 19671 76993
rect 13814 76956 13820 76968
rect 13775 76928 13820 76956
rect 13814 76916 13820 76928
rect 13872 76916 13878 76968
rect 19334 76956 19340 76968
rect 19295 76928 19340 76956
rect 19334 76916 19340 76928
rect 19392 76916 19398 76968
rect 20993 76891 21051 76897
rect 20993 76857 21005 76891
rect 21039 76888 21051 76891
rect 22738 76888 22744 76900
rect 21039 76860 22744 76888
rect 21039 76857 21051 76860
rect 20993 76851 21051 76857
rect 22738 76848 22744 76860
rect 22796 76848 22802 76900
rect 15197 76823 15255 76829
rect 15197 76789 15209 76823
rect 15243 76820 15255 76823
rect 15286 76820 15292 76832
rect 15243 76792 15292 76820
rect 15243 76789 15255 76792
rect 15197 76783 15255 76789
rect 15286 76780 15292 76792
rect 15344 76780 15350 76832
rect 1104 76730 28888 76752
rect 1104 76678 10982 76730
rect 11034 76678 11046 76730
rect 11098 76678 11110 76730
rect 11162 76678 11174 76730
rect 11226 76678 20982 76730
rect 21034 76678 21046 76730
rect 21098 76678 21110 76730
rect 21162 76678 21174 76730
rect 21226 76678 28888 76730
rect 1104 76656 28888 76678
rect 8754 76440 8760 76492
rect 8812 76480 8818 76492
rect 9766 76480 9772 76492
rect 8812 76452 9772 76480
rect 8812 76440 8818 76452
rect 9766 76440 9772 76452
rect 9824 76480 9830 76492
rect 9953 76483 10011 76489
rect 9953 76480 9965 76483
rect 9824 76452 9965 76480
rect 9824 76440 9830 76452
rect 9953 76449 9965 76452
rect 9999 76449 10011 76483
rect 9953 76443 10011 76449
rect 20806 76440 20812 76492
rect 20864 76480 20870 76492
rect 21177 76483 21235 76489
rect 21177 76480 21189 76483
rect 20864 76452 21189 76480
rect 20864 76440 20870 76452
rect 21177 76449 21189 76452
rect 21223 76449 21235 76483
rect 21177 76443 21235 76449
rect 9677 76415 9735 76421
rect 9677 76381 9689 76415
rect 9723 76412 9735 76415
rect 10042 76412 10048 76424
rect 9723 76384 10048 76412
rect 9723 76381 9735 76384
rect 9677 76375 9735 76381
rect 10042 76372 10048 76384
rect 10100 76372 10106 76424
rect 12161 76415 12219 76421
rect 12161 76381 12173 76415
rect 12207 76412 12219 76415
rect 12342 76412 12348 76424
rect 12207 76384 12348 76412
rect 12207 76381 12219 76384
rect 12161 76375 12219 76381
rect 12342 76372 12348 76384
rect 12400 76372 12406 76424
rect 12434 76372 12440 76424
rect 12492 76412 12498 76424
rect 12492 76384 12537 76412
rect 12492 76372 12498 76384
rect 19242 76372 19248 76424
rect 19300 76412 19306 76424
rect 19429 76415 19487 76421
rect 19429 76412 19441 76415
rect 19300 76384 19441 76412
rect 19300 76372 19306 76384
rect 19429 76381 19441 76384
rect 19475 76412 19487 76415
rect 20901 76415 20959 76421
rect 20901 76412 20913 76415
rect 19475 76384 20913 76412
rect 19475 76381 19487 76384
rect 19429 76375 19487 76381
rect 20901 76381 20913 76384
rect 20947 76412 20959 76415
rect 21358 76412 21364 76424
rect 20947 76384 21364 76412
rect 20947 76381 20959 76384
rect 20901 76375 20959 76381
rect 21358 76372 21364 76384
rect 21416 76372 21422 76424
rect 13722 76344 13728 76356
rect 13683 76316 13728 76344
rect 13722 76304 13728 76316
rect 13780 76304 13786 76356
rect 11241 76279 11299 76285
rect 11241 76245 11253 76279
rect 11287 76276 11299 76279
rect 11606 76276 11612 76288
rect 11287 76248 11612 76276
rect 11287 76245 11299 76248
rect 11241 76239 11299 76245
rect 11606 76236 11612 76248
rect 11664 76236 11670 76288
rect 22465 76279 22523 76285
rect 22465 76245 22477 76279
rect 22511 76276 22523 76279
rect 22646 76276 22652 76288
rect 22511 76248 22652 76276
rect 22511 76245 22523 76248
rect 22465 76239 22523 76245
rect 22646 76236 22652 76248
rect 22704 76236 22710 76288
rect 1104 76186 28888 76208
rect 1104 76134 5982 76186
rect 6034 76134 6046 76186
rect 6098 76134 6110 76186
rect 6162 76134 6174 76186
rect 6226 76134 15982 76186
rect 16034 76134 16046 76186
rect 16098 76134 16110 76186
rect 16162 76134 16174 76186
rect 16226 76134 25982 76186
rect 26034 76134 26046 76186
rect 26098 76134 26110 76186
rect 26162 76134 26174 76186
rect 26226 76134 28888 76186
rect 1104 76112 28888 76134
rect 9766 76072 9772 76084
rect 9727 76044 9772 76072
rect 9766 76032 9772 76044
rect 9824 76032 9830 76084
rect 20806 76032 20812 76084
rect 20864 76072 20870 76084
rect 20901 76075 20959 76081
rect 20901 76072 20913 76075
rect 20864 76044 20913 76072
rect 20864 76032 20870 76044
rect 20901 76041 20913 76044
rect 20947 76041 20959 76075
rect 20901 76035 20959 76041
rect 12434 75896 12440 75948
rect 12492 75896 12498 75948
rect 1394 75828 1400 75880
rect 1452 75868 1458 75880
rect 1854 75868 1860 75880
rect 1452 75840 1860 75868
rect 1452 75828 1458 75840
rect 1854 75828 1860 75840
rect 1912 75828 1918 75880
rect 12158 75868 12164 75880
rect 12119 75840 12164 75868
rect 12158 75828 12164 75840
rect 12216 75868 12222 75880
rect 12452 75868 12480 75896
rect 13538 75868 13544 75880
rect 12216 75840 12480 75868
rect 12636 75840 13544 75868
rect 12216 75828 12222 75840
rect 10134 75732 10140 75744
rect 10095 75704 10140 75732
rect 10134 75692 10140 75704
rect 10192 75692 10198 75744
rect 12342 75692 12348 75744
rect 12400 75732 12406 75744
rect 12434 75732 12440 75744
rect 12400 75704 12440 75732
rect 12400 75692 12406 75704
rect 12434 75692 12440 75704
rect 12492 75732 12498 75744
rect 12636 75741 12664 75840
rect 13538 75828 13544 75840
rect 13596 75828 13602 75880
rect 13817 75871 13875 75877
rect 13817 75868 13829 75871
rect 13648 75840 13829 75868
rect 12621 75735 12679 75741
rect 12621 75732 12633 75735
rect 12492 75704 12633 75732
rect 12492 75692 12498 75704
rect 12621 75701 12633 75704
rect 12667 75701 12679 75735
rect 13354 75732 13360 75744
rect 13315 75704 13360 75732
rect 12621 75695 12679 75701
rect 13354 75692 13360 75704
rect 13412 75732 13418 75744
rect 13648 75732 13676 75840
rect 13817 75837 13829 75840
rect 13863 75837 13875 75871
rect 13817 75831 13875 75837
rect 15102 75732 15108 75744
rect 13412 75704 13676 75732
rect 15063 75704 15108 75732
rect 13412 75692 13418 75704
rect 15102 75692 15108 75704
rect 15160 75692 15166 75744
rect 21358 75732 21364 75744
rect 21319 75704 21364 75732
rect 21358 75692 21364 75704
rect 21416 75692 21422 75744
rect 1104 75642 28888 75664
rect 1104 75590 10982 75642
rect 11034 75590 11046 75642
rect 11098 75590 11110 75642
rect 11162 75590 11174 75642
rect 11226 75590 20982 75642
rect 21034 75590 21046 75642
rect 21098 75590 21110 75642
rect 21162 75590 21174 75642
rect 21226 75590 28888 75642
rect 1104 75568 28888 75590
rect 25038 75528 25044 75540
rect 24999 75500 25044 75528
rect 25038 75488 25044 75500
rect 25096 75488 25102 75540
rect 10502 75352 10508 75404
rect 10560 75392 10566 75404
rect 10689 75395 10747 75401
rect 10689 75392 10701 75395
rect 10560 75364 10701 75392
rect 10560 75352 10566 75364
rect 10689 75361 10701 75364
rect 10735 75392 10747 75395
rect 11330 75392 11336 75404
rect 10735 75364 11336 75392
rect 10735 75361 10747 75364
rect 10689 75355 10747 75361
rect 11330 75352 11336 75364
rect 11388 75352 11394 75404
rect 10134 75284 10140 75336
rect 10192 75324 10198 75336
rect 10413 75327 10471 75333
rect 10413 75324 10425 75327
rect 10192 75296 10425 75324
rect 10192 75284 10198 75296
rect 10413 75293 10425 75296
rect 10459 75324 10471 75327
rect 10778 75324 10784 75336
rect 10459 75296 10784 75324
rect 10459 75293 10471 75296
rect 10413 75287 10471 75293
rect 10778 75284 10784 75296
rect 10836 75284 10842 75336
rect 23658 75324 23664 75336
rect 23619 75296 23664 75324
rect 23658 75284 23664 75296
rect 23716 75284 23722 75336
rect 23934 75324 23940 75336
rect 23895 75296 23940 75324
rect 23934 75284 23940 75296
rect 23992 75284 23998 75336
rect 11974 75188 11980 75200
rect 11935 75160 11980 75188
rect 11974 75148 11980 75160
rect 12032 75148 12038 75200
rect 12434 75148 12440 75200
rect 12492 75188 12498 75200
rect 13541 75191 13599 75197
rect 13541 75188 13553 75191
rect 12492 75160 13553 75188
rect 12492 75148 12498 75160
rect 13541 75157 13553 75160
rect 13587 75157 13599 75191
rect 13541 75151 13599 75157
rect 1104 75098 28888 75120
rect 1104 75046 5982 75098
rect 6034 75046 6046 75098
rect 6098 75046 6110 75098
rect 6162 75046 6174 75098
rect 6226 75046 15982 75098
rect 16034 75046 16046 75098
rect 16098 75046 16110 75098
rect 16162 75046 16174 75098
rect 16226 75046 25982 75098
rect 26034 75046 26046 75098
rect 26098 75046 26110 75098
rect 26162 75046 26174 75098
rect 26226 75046 28888 75098
rect 1104 75024 28888 75046
rect 10502 74984 10508 74996
rect 10463 74956 10508 74984
rect 10502 74944 10508 74956
rect 10560 74944 10566 74996
rect 17954 74944 17960 74996
rect 18012 74984 18018 74996
rect 18877 74987 18935 74993
rect 18877 74984 18889 74987
rect 18012 74956 18889 74984
rect 18012 74944 18018 74956
rect 18877 74953 18889 74956
rect 18923 74953 18935 74987
rect 18877 74947 18935 74953
rect 18892 74848 18920 74947
rect 23658 74944 23664 74996
rect 23716 74984 23722 74996
rect 24213 74987 24271 74993
rect 24213 74984 24225 74987
rect 23716 74956 24225 74984
rect 23716 74944 23722 74956
rect 24213 74953 24225 74956
rect 24259 74984 24271 74987
rect 24762 74984 24768 74996
rect 24259 74956 24768 74984
rect 24259 74953 24271 74956
rect 24213 74947 24271 74953
rect 24762 74944 24768 74956
rect 24820 74944 24826 74996
rect 19337 74851 19395 74857
rect 19337 74848 19349 74851
rect 18892 74820 19349 74848
rect 19337 74817 19349 74820
rect 19383 74817 19395 74851
rect 19337 74811 19395 74817
rect 4154 74740 4160 74792
rect 4212 74780 4218 74792
rect 5442 74780 5448 74792
rect 4212 74752 5448 74780
rect 4212 74740 4218 74752
rect 5442 74740 5448 74752
rect 5500 74740 5506 74792
rect 12526 74740 12532 74792
rect 12584 74780 12590 74792
rect 13722 74780 13728 74792
rect 12584 74752 13728 74780
rect 12584 74740 12590 74752
rect 13722 74740 13728 74752
rect 13780 74740 13786 74792
rect 13814 74740 13820 74792
rect 13872 74780 13878 74792
rect 14734 74780 14740 74792
rect 13872 74752 14740 74780
rect 13872 74740 13878 74752
rect 14734 74740 14740 74752
rect 14792 74740 14798 74792
rect 15654 74740 15660 74792
rect 15712 74780 15718 74792
rect 16482 74780 16488 74792
rect 15712 74752 16488 74780
rect 15712 74740 15718 74752
rect 16482 74740 16488 74752
rect 16540 74740 16546 74792
rect 19061 74783 19119 74789
rect 19061 74749 19073 74783
rect 19107 74780 19119 74783
rect 19150 74780 19156 74792
rect 19107 74752 19156 74780
rect 19107 74749 19119 74752
rect 19061 74743 19119 74749
rect 19150 74740 19156 74752
rect 19208 74740 19214 74792
rect 4614 74604 4620 74656
rect 4672 74644 4678 74656
rect 5534 74644 5540 74656
rect 4672 74616 5540 74644
rect 4672 74604 4678 74616
rect 5534 74604 5540 74616
rect 5592 74604 5598 74656
rect 6454 74604 6460 74656
rect 6512 74644 6518 74656
rect 6914 74644 6920 74656
rect 6512 74616 6920 74644
rect 6512 74604 6518 74616
rect 6914 74604 6920 74616
rect 6972 74604 6978 74656
rect 10778 74644 10784 74656
rect 10739 74616 10784 74644
rect 10778 74604 10784 74616
rect 10836 74604 10842 74656
rect 20346 74604 20352 74656
rect 20404 74644 20410 74656
rect 20441 74647 20499 74653
rect 20441 74644 20453 74647
rect 20404 74616 20453 74644
rect 20404 74604 20410 74616
rect 20441 74613 20453 74616
rect 20487 74613 20499 74647
rect 20441 74607 20499 74613
rect 22094 74604 22100 74656
rect 22152 74644 22158 74656
rect 22554 74644 22560 74656
rect 22152 74616 22560 74644
rect 22152 74604 22158 74616
rect 22554 74604 22560 74616
rect 22612 74604 22618 74656
rect 23934 74644 23940 74656
rect 23895 74616 23940 74644
rect 23934 74604 23940 74616
rect 23992 74604 23998 74656
rect 27614 74604 27620 74656
rect 27672 74644 27678 74656
rect 28994 74644 29000 74656
rect 27672 74616 29000 74644
rect 27672 74604 27678 74616
rect 28994 74604 29000 74616
rect 29052 74604 29058 74656
rect 1104 74554 28888 74576
rect 1104 74502 10982 74554
rect 11034 74502 11046 74554
rect 11098 74502 11110 74554
rect 11162 74502 11174 74554
rect 11226 74502 20982 74554
rect 21034 74502 21046 74554
rect 21098 74502 21110 74554
rect 21162 74502 21174 74554
rect 21226 74502 28888 74554
rect 1104 74480 28888 74502
rect 19153 74443 19211 74449
rect 19153 74409 19165 74443
rect 19199 74440 19211 74443
rect 19242 74440 19248 74452
rect 19199 74412 19248 74440
rect 19199 74409 19211 74412
rect 19153 74403 19211 74409
rect 19242 74400 19248 74412
rect 19300 74400 19306 74452
rect 11974 74264 11980 74316
rect 12032 74304 12038 74316
rect 12437 74307 12495 74313
rect 12437 74304 12449 74307
rect 12032 74276 12449 74304
rect 12032 74264 12038 74276
rect 12437 74273 12449 74276
rect 12483 74273 12495 74307
rect 12437 74267 12495 74273
rect 12161 74239 12219 74245
rect 12161 74205 12173 74239
rect 12207 74236 12219 74239
rect 12342 74236 12348 74248
rect 12207 74208 12348 74236
rect 12207 74205 12219 74208
rect 12161 74199 12219 74205
rect 12342 74196 12348 74208
rect 12400 74196 12406 74248
rect 13078 74060 13084 74112
rect 13136 74100 13142 74112
rect 13541 74103 13599 74109
rect 13541 74100 13553 74103
rect 13136 74072 13553 74100
rect 13136 74060 13142 74072
rect 13541 74069 13553 74072
rect 13587 74069 13599 74103
rect 13541 74063 13599 74069
rect 1104 74010 28888 74032
rect 1104 73958 5982 74010
rect 6034 73958 6046 74010
rect 6098 73958 6110 74010
rect 6162 73958 6174 74010
rect 6226 73958 15982 74010
rect 16034 73958 16046 74010
rect 16098 73958 16110 74010
rect 16162 73958 16174 74010
rect 16226 73958 25982 74010
rect 26034 73958 26046 74010
rect 26098 73958 26110 74010
rect 26162 73958 26174 74010
rect 26226 73958 28888 74010
rect 1104 73936 28888 73958
rect 11974 73856 11980 73908
rect 12032 73896 12038 73908
rect 12161 73899 12219 73905
rect 12161 73896 12173 73899
rect 12032 73868 12173 73896
rect 12032 73856 12038 73868
rect 12161 73865 12173 73868
rect 12207 73865 12219 73899
rect 12161 73859 12219 73865
rect 12434 73516 12440 73568
rect 12492 73556 12498 73568
rect 12621 73559 12679 73565
rect 12621 73556 12633 73559
rect 12492 73528 12633 73556
rect 12492 73516 12498 73528
rect 12621 73525 12633 73528
rect 12667 73525 12679 73559
rect 12621 73519 12679 73525
rect 1104 73466 28888 73488
rect 1104 73414 10982 73466
rect 11034 73414 11046 73466
rect 11098 73414 11110 73466
rect 11162 73414 11174 73466
rect 11226 73414 20982 73466
rect 21034 73414 21046 73466
rect 21098 73414 21110 73466
rect 21162 73414 21174 73466
rect 21226 73414 28888 73466
rect 1104 73392 28888 73414
rect 14366 73284 14372 73296
rect 14327 73256 14372 73284
rect 14366 73244 14372 73256
rect 14424 73244 14430 73296
rect 12989 73219 13047 73225
rect 12989 73185 13001 73219
rect 13035 73216 13047 73219
rect 13078 73216 13084 73228
rect 13035 73188 13084 73216
rect 13035 73185 13047 73188
rect 12989 73179 13047 73185
rect 13078 73176 13084 73188
rect 13136 73176 13142 73228
rect 12434 73108 12440 73160
rect 12492 73148 12498 73160
rect 12713 73151 12771 73157
rect 12713 73148 12725 73151
rect 12492 73120 12725 73148
rect 12492 73108 12498 73120
rect 12713 73117 12725 73120
rect 12759 73117 12771 73151
rect 12713 73111 12771 73117
rect 1104 72922 28888 72944
rect 1104 72870 5982 72922
rect 6034 72870 6046 72922
rect 6098 72870 6110 72922
rect 6162 72870 6174 72922
rect 6226 72870 15982 72922
rect 16034 72870 16046 72922
rect 16098 72870 16110 72922
rect 16162 72870 16174 72922
rect 16226 72870 25982 72922
rect 26034 72870 26046 72922
rect 26098 72870 26110 72922
rect 26162 72870 26174 72922
rect 26226 72870 28888 72922
rect 1104 72848 28888 72870
rect 12805 72811 12863 72817
rect 12805 72777 12817 72811
rect 12851 72808 12863 72811
rect 13078 72808 13084 72820
rect 12851 72780 13084 72808
rect 12851 72777 12863 72780
rect 12805 72771 12863 72777
rect 13078 72768 13084 72780
rect 13136 72768 13142 72820
rect 12434 72428 12440 72480
rect 12492 72468 12498 72480
rect 13081 72471 13139 72477
rect 13081 72468 13093 72471
rect 12492 72440 13093 72468
rect 12492 72428 12498 72440
rect 13081 72437 13093 72440
rect 13127 72437 13139 72471
rect 13081 72431 13139 72437
rect 1104 72378 28888 72400
rect 1104 72326 10982 72378
rect 11034 72326 11046 72378
rect 11098 72326 11110 72378
rect 11162 72326 11174 72378
rect 11226 72326 20982 72378
rect 21034 72326 21046 72378
rect 21098 72326 21110 72378
rect 21162 72326 21174 72378
rect 21226 72326 28888 72378
rect 1104 72304 28888 72326
rect 22554 72196 22560 72208
rect 22515 72168 22560 72196
rect 22554 72156 22560 72168
rect 22612 72156 22618 72208
rect 20806 72088 20812 72140
rect 20864 72128 20870 72140
rect 21177 72131 21235 72137
rect 21177 72128 21189 72131
rect 20864 72100 21189 72128
rect 20864 72088 20870 72100
rect 21177 72097 21189 72100
rect 21223 72097 21235 72131
rect 21177 72091 21235 72097
rect 20901 72063 20959 72069
rect 20901 72029 20913 72063
rect 20947 72060 20959 72063
rect 21358 72060 21364 72072
rect 20947 72032 21364 72060
rect 20947 72029 20959 72032
rect 20901 72023 20959 72029
rect 21358 72020 21364 72032
rect 21416 72020 21422 72072
rect 1104 71834 28888 71856
rect 1104 71782 5982 71834
rect 6034 71782 6046 71834
rect 6098 71782 6110 71834
rect 6162 71782 6174 71834
rect 6226 71782 15982 71834
rect 16034 71782 16046 71834
rect 16098 71782 16110 71834
rect 16162 71782 16174 71834
rect 16226 71782 25982 71834
rect 26034 71782 26046 71834
rect 26098 71782 26110 71834
rect 26162 71782 26174 71834
rect 26226 71782 28888 71834
rect 1104 71760 28888 71782
rect 20806 71340 20812 71392
rect 20864 71380 20870 71392
rect 20901 71383 20959 71389
rect 20901 71380 20913 71383
rect 20864 71352 20913 71380
rect 20864 71340 20870 71352
rect 20901 71349 20913 71352
rect 20947 71349 20959 71383
rect 21358 71380 21364 71392
rect 21319 71352 21364 71380
rect 20901 71343 20959 71349
rect 21358 71340 21364 71352
rect 21416 71340 21422 71392
rect 1104 71290 28888 71312
rect 1104 71238 10982 71290
rect 11034 71238 11046 71290
rect 11098 71238 11110 71290
rect 11162 71238 11174 71290
rect 11226 71238 20982 71290
rect 21034 71238 21046 71290
rect 21098 71238 21110 71290
rect 21162 71238 21174 71290
rect 21226 71238 28888 71290
rect 1104 71216 28888 71238
rect 7558 71068 7564 71120
rect 7616 71108 7622 71120
rect 8018 71108 8024 71120
rect 7616 71080 8024 71108
rect 7616 71068 7622 71080
rect 8018 71068 8024 71080
rect 8076 71068 8082 71120
rect 22557 71111 22615 71117
rect 22557 71077 22569 71111
rect 22603 71108 22615 71111
rect 23382 71108 23388 71120
rect 22603 71080 23388 71108
rect 22603 71077 22615 71080
rect 22557 71071 22615 71077
rect 23382 71068 23388 71080
rect 23440 71068 23446 71120
rect 20990 71000 20996 71052
rect 21048 71040 21054 71052
rect 21177 71043 21235 71049
rect 21177 71040 21189 71043
rect 21048 71012 21189 71040
rect 21048 71000 21054 71012
rect 21177 71009 21189 71012
rect 21223 71009 21235 71043
rect 21177 71003 21235 71009
rect 20901 70975 20959 70981
rect 20901 70941 20913 70975
rect 20947 70972 20959 70975
rect 21358 70972 21364 70984
rect 20947 70944 21364 70972
rect 20947 70941 20959 70944
rect 20901 70935 20959 70941
rect 21358 70932 21364 70944
rect 21416 70932 21422 70984
rect 23106 70932 23112 70984
rect 23164 70972 23170 70984
rect 23382 70972 23388 70984
rect 23164 70944 23388 70972
rect 23164 70932 23170 70944
rect 23382 70932 23388 70944
rect 23440 70932 23446 70984
rect 1104 70746 28888 70768
rect 1104 70694 5982 70746
rect 6034 70694 6046 70746
rect 6098 70694 6110 70746
rect 6162 70694 6174 70746
rect 6226 70694 15982 70746
rect 16034 70694 16046 70746
rect 16098 70694 16110 70746
rect 16162 70694 16174 70746
rect 16226 70694 25982 70746
rect 26034 70694 26046 70746
rect 26098 70694 26110 70746
rect 26162 70694 26174 70746
rect 26226 70694 28888 70746
rect 1104 70672 28888 70694
rect 20898 70564 20904 70576
rect 20859 70536 20904 70564
rect 20898 70524 20904 70536
rect 20956 70524 20962 70576
rect 26053 70499 26111 70505
rect 26053 70465 26065 70499
rect 26099 70496 26111 70499
rect 26418 70496 26424 70508
rect 26099 70468 26424 70496
rect 26099 70465 26111 70468
rect 26053 70459 26111 70465
rect 26418 70456 26424 70468
rect 26476 70456 26482 70508
rect 21358 70428 21364 70440
rect 21271 70400 21364 70428
rect 21358 70388 21364 70400
rect 21416 70428 21422 70440
rect 21726 70428 21732 70440
rect 21416 70400 21732 70428
rect 21416 70388 21422 70400
rect 21726 70388 21732 70400
rect 21784 70388 21790 70440
rect 24854 70388 24860 70440
rect 24912 70428 24918 70440
rect 26142 70428 26148 70440
rect 24912 70400 26148 70428
rect 24912 70388 24918 70400
rect 26142 70388 26148 70400
rect 26200 70388 26206 70440
rect 27706 70320 27712 70372
rect 27764 70360 27770 70372
rect 27890 70360 27896 70372
rect 27764 70332 27896 70360
rect 27764 70320 27770 70332
rect 27890 70320 27896 70332
rect 27948 70320 27954 70372
rect 26418 70252 26424 70304
rect 26476 70292 26482 70304
rect 27525 70295 27583 70301
rect 27525 70292 27537 70295
rect 26476 70264 27537 70292
rect 26476 70252 26482 70264
rect 27525 70261 27537 70264
rect 27571 70261 27583 70295
rect 27525 70255 27583 70261
rect 1104 70202 28888 70224
rect 1104 70150 10982 70202
rect 11034 70150 11046 70202
rect 11098 70150 11110 70202
rect 11162 70150 11174 70202
rect 11226 70150 20982 70202
rect 21034 70150 21046 70202
rect 21098 70150 21110 70202
rect 21162 70150 21174 70202
rect 21226 70150 28888 70202
rect 1104 70128 28888 70150
rect 2774 70048 2780 70100
rect 2832 70088 2838 70100
rect 2832 70060 2877 70088
rect 2832 70048 2838 70060
rect 25866 70048 25872 70100
rect 25924 70088 25930 70100
rect 26142 70088 26148 70100
rect 25924 70060 26148 70088
rect 25924 70048 25930 70060
rect 26142 70048 26148 70060
rect 26200 70048 26206 70100
rect 1397 69955 1455 69961
rect 1397 69921 1409 69955
rect 1443 69952 1455 69955
rect 2038 69952 2044 69964
rect 1443 69924 2044 69952
rect 1443 69921 1455 69924
rect 1397 69915 1455 69921
rect 2038 69912 2044 69924
rect 2096 69912 2102 69964
rect 1670 69884 1676 69896
rect 1631 69856 1676 69884
rect 1670 69844 1676 69856
rect 1728 69844 1734 69896
rect 1104 69658 28888 69680
rect 1104 69606 5982 69658
rect 6034 69606 6046 69658
rect 6098 69606 6110 69658
rect 6162 69606 6174 69658
rect 6226 69606 15982 69658
rect 16034 69606 16046 69658
rect 16098 69606 16110 69658
rect 16162 69606 16174 69658
rect 16226 69606 25982 69658
rect 26034 69606 26046 69658
rect 26098 69606 26110 69658
rect 26162 69606 26174 69658
rect 26226 69606 28888 69658
rect 1104 69584 28888 69606
rect 11333 69479 11391 69485
rect 11333 69445 11345 69479
rect 11379 69476 11391 69479
rect 12342 69476 12348 69488
rect 11379 69448 12348 69476
rect 11379 69445 11391 69448
rect 11333 69439 11391 69445
rect 12342 69436 12348 69448
rect 12400 69436 12406 69488
rect 1578 69368 1584 69420
rect 1636 69408 1642 69420
rect 2038 69408 2044 69420
rect 1636 69380 2044 69408
rect 1636 69368 1642 69380
rect 2038 69368 2044 69380
rect 2096 69368 2102 69420
rect 26053 69411 26111 69417
rect 26053 69377 26065 69411
rect 26099 69408 26111 69411
rect 26418 69408 26424 69420
rect 26099 69380 26424 69408
rect 26099 69377 26111 69380
rect 26053 69371 26111 69377
rect 26418 69368 26424 69380
rect 26476 69368 26482 69420
rect 1670 69340 1676 69352
rect 1631 69312 1676 69340
rect 1670 69300 1676 69312
rect 1728 69300 1734 69352
rect 11330 69300 11336 69352
rect 11388 69340 11394 69352
rect 11517 69343 11575 69349
rect 11517 69340 11529 69343
rect 11388 69312 11529 69340
rect 11388 69300 11394 69312
rect 11517 69309 11529 69312
rect 11563 69340 11575 69343
rect 11793 69343 11851 69349
rect 11793 69340 11805 69343
rect 11563 69312 11805 69340
rect 11563 69309 11575 69312
rect 11517 69303 11575 69309
rect 11793 69309 11805 69312
rect 11839 69309 11851 69343
rect 11793 69303 11851 69309
rect 24854 69300 24860 69352
rect 24912 69340 24918 69352
rect 25866 69340 25872 69352
rect 24912 69312 25872 69340
rect 24912 69300 24918 69312
rect 25866 69300 25872 69312
rect 25924 69340 25930 69352
rect 26145 69343 26203 69349
rect 26145 69340 26157 69343
rect 25924 69312 26157 69340
rect 25924 69300 25930 69312
rect 26145 69309 26157 69312
rect 26191 69340 26203 69343
rect 26234 69340 26240 69352
rect 26191 69312 26240 69340
rect 26191 69309 26203 69312
rect 26145 69303 26203 69309
rect 26234 69300 26240 69312
rect 26292 69300 26298 69352
rect 27706 69204 27712 69216
rect 27667 69176 27712 69204
rect 27706 69164 27712 69176
rect 27764 69164 27770 69216
rect 1104 69114 28888 69136
rect 1104 69062 10982 69114
rect 11034 69062 11046 69114
rect 11098 69062 11110 69114
rect 11162 69062 11174 69114
rect 11226 69062 20982 69114
rect 21034 69062 21046 69114
rect 21098 69062 21110 69114
rect 21162 69062 21174 69114
rect 21226 69062 28888 69114
rect 1104 69040 28888 69062
rect 26234 69000 26240 69012
rect 26195 68972 26240 69000
rect 26234 68960 26240 68972
rect 26292 68960 26298 69012
rect 1104 68570 28888 68592
rect 1104 68518 5982 68570
rect 6034 68518 6046 68570
rect 6098 68518 6110 68570
rect 6162 68518 6174 68570
rect 6226 68518 15982 68570
rect 16034 68518 16046 68570
rect 16098 68518 16110 68570
rect 16162 68518 16174 68570
rect 16226 68518 25982 68570
rect 26034 68518 26046 68570
rect 26098 68518 26110 68570
rect 26162 68518 26174 68570
rect 26226 68518 28888 68570
rect 1104 68496 28888 68518
rect 9122 68456 9128 68468
rect 9083 68428 9128 68456
rect 9122 68416 9128 68428
rect 9180 68416 9186 68468
rect 9677 68459 9735 68465
rect 9677 68425 9689 68459
rect 9723 68456 9735 68459
rect 10686 68456 10692 68468
rect 9723 68428 10692 68456
rect 9723 68425 9735 68428
rect 9677 68419 9735 68425
rect 9309 68255 9367 68261
rect 9309 68221 9321 68255
rect 9355 68252 9367 68255
rect 9692 68252 9720 68419
rect 10686 68416 10692 68428
rect 10744 68456 10750 68468
rect 11330 68456 11336 68468
rect 10744 68428 11336 68456
rect 10744 68416 10750 68428
rect 11330 68416 11336 68428
rect 11388 68416 11394 68468
rect 9355 68224 9720 68252
rect 9355 68221 9367 68224
rect 9309 68215 9367 68221
rect 1104 68026 28888 68048
rect 1104 67974 10982 68026
rect 11034 67974 11046 68026
rect 11098 67974 11110 68026
rect 11162 67974 11174 68026
rect 11226 67974 20982 68026
rect 21034 67974 21046 68026
rect 21098 67974 21110 68026
rect 21162 67974 21174 68026
rect 21226 67974 28888 68026
rect 1104 67952 28888 67974
rect 11238 67600 11244 67652
rect 11296 67640 11302 67652
rect 11974 67640 11980 67652
rect 11296 67612 11980 67640
rect 11296 67600 11302 67612
rect 11974 67600 11980 67612
rect 12032 67600 12038 67652
rect 16390 67600 16396 67652
rect 16448 67640 16454 67652
rect 16574 67640 16580 67652
rect 16448 67612 16580 67640
rect 16448 67600 16454 67612
rect 16574 67600 16580 67612
rect 16632 67600 16638 67652
rect 1104 67482 28888 67504
rect 1104 67430 5982 67482
rect 6034 67430 6046 67482
rect 6098 67430 6110 67482
rect 6162 67430 6174 67482
rect 6226 67430 15982 67482
rect 16034 67430 16046 67482
rect 16098 67430 16110 67482
rect 16162 67430 16174 67482
rect 16226 67430 25982 67482
rect 26034 67430 26046 67482
rect 26098 67430 26110 67482
rect 26162 67430 26174 67482
rect 26226 67430 28888 67482
rect 1104 67408 28888 67430
rect 10686 67368 10692 67380
rect 10647 67340 10692 67368
rect 10686 67328 10692 67340
rect 10744 67328 10750 67380
rect 10873 67167 10931 67173
rect 10873 67133 10885 67167
rect 10919 67164 10931 67167
rect 10919 67136 11284 67164
rect 10919 67133 10931 67136
rect 10873 67127 10931 67133
rect 11256 67037 11284 67136
rect 11241 67031 11299 67037
rect 11241 66997 11253 67031
rect 11287 67028 11299 67031
rect 11974 67028 11980 67040
rect 11287 67000 11980 67028
rect 11287 66997 11299 67000
rect 11241 66991 11299 66997
rect 11974 66988 11980 67000
rect 12032 66988 12038 67040
rect 1104 66938 28888 66960
rect 1104 66886 10982 66938
rect 11034 66886 11046 66938
rect 11098 66886 11110 66938
rect 11162 66886 11174 66938
rect 11226 66886 20982 66938
rect 21034 66886 21046 66938
rect 21098 66886 21110 66938
rect 21162 66886 21174 66938
rect 21226 66886 28888 66938
rect 1104 66864 28888 66886
rect 21637 66827 21695 66833
rect 21637 66793 21649 66827
rect 21683 66824 21695 66827
rect 21726 66824 21732 66836
rect 21683 66796 21732 66824
rect 21683 66793 21695 66796
rect 21637 66787 21695 66793
rect 21726 66784 21732 66796
rect 21784 66784 21790 66836
rect 17218 66688 17224 66700
rect 17179 66660 17224 66688
rect 17218 66648 17224 66660
rect 17276 66648 17282 66700
rect 17681 66691 17739 66697
rect 17681 66657 17693 66691
rect 17727 66688 17739 66691
rect 17862 66688 17868 66700
rect 17727 66660 17868 66688
rect 17727 66657 17739 66660
rect 17681 66651 17739 66657
rect 17862 66648 17868 66660
rect 17920 66648 17926 66700
rect 21818 66688 21824 66700
rect 21779 66660 21824 66688
rect 21818 66648 21824 66660
rect 21876 66648 21882 66700
rect 16942 66620 16948 66632
rect 16903 66592 16948 66620
rect 16942 66580 16948 66592
rect 17000 66580 17006 66632
rect 17586 66552 17592 66564
rect 17547 66524 17592 66552
rect 17586 66512 17592 66524
rect 17644 66512 17650 66564
rect 18046 66444 18052 66496
rect 18104 66484 18110 66496
rect 18233 66487 18291 66493
rect 18233 66484 18245 66487
rect 18104 66456 18245 66484
rect 18104 66444 18110 66456
rect 18233 66453 18245 66456
rect 18279 66484 18291 66487
rect 18874 66484 18880 66496
rect 18279 66456 18880 66484
rect 18279 66453 18291 66456
rect 18233 66447 18291 66453
rect 18874 66444 18880 66456
rect 18932 66444 18938 66496
rect 1104 66394 28888 66416
rect 1104 66342 5982 66394
rect 6034 66342 6046 66394
rect 6098 66342 6110 66394
rect 6162 66342 6174 66394
rect 6226 66342 15982 66394
rect 16034 66342 16046 66394
rect 16098 66342 16110 66394
rect 16162 66342 16174 66394
rect 16226 66342 25982 66394
rect 26034 66342 26046 66394
rect 26098 66342 26110 66394
rect 26162 66342 26174 66394
rect 26226 66342 28888 66394
rect 1104 66320 28888 66342
rect 21729 66283 21787 66289
rect 21729 66249 21741 66283
rect 21775 66280 21787 66283
rect 21818 66280 21824 66292
rect 21775 66252 21824 66280
rect 21775 66249 21787 66252
rect 21729 66243 21787 66249
rect 21818 66240 21824 66252
rect 21876 66240 21882 66292
rect 27706 66240 27712 66292
rect 27764 66280 27770 66292
rect 27982 66280 27988 66292
rect 27764 66252 27988 66280
rect 27764 66240 27770 66252
rect 27982 66240 27988 66252
rect 28040 66240 28046 66292
rect 18046 66144 18052 66156
rect 18007 66116 18052 66144
rect 18046 66104 18052 66116
rect 18104 66104 18110 66156
rect 18325 66079 18383 66085
rect 18325 66076 18337 66079
rect 18156 66048 18337 66076
rect 16853 66011 16911 66017
rect 16853 65977 16865 66011
rect 16899 66008 16911 66011
rect 16942 66008 16948 66020
rect 16899 65980 16948 66008
rect 16899 65977 16911 65980
rect 16853 65971 16911 65977
rect 16942 65968 16948 65980
rect 17000 66008 17006 66020
rect 17586 66008 17592 66020
rect 17000 65980 17592 66008
rect 17000 65968 17006 65980
rect 17586 65968 17592 65980
rect 17644 65968 17650 66020
rect 17770 66008 17776 66020
rect 17731 65980 17776 66008
rect 17770 65968 17776 65980
rect 17828 66008 17834 66020
rect 18156 66008 18184 66048
rect 18325 66045 18337 66048
rect 18371 66045 18383 66079
rect 18325 66039 18383 66045
rect 17828 65980 18184 66008
rect 19705 66011 19763 66017
rect 17828 65968 17834 65980
rect 19705 65977 19717 66011
rect 19751 66008 19763 66011
rect 20530 66008 20536 66020
rect 19751 65980 20536 66008
rect 19751 65977 19763 65980
rect 19705 65971 19763 65977
rect 20530 65968 20536 65980
rect 20588 65968 20594 66020
rect 15470 65900 15476 65952
rect 15528 65940 15534 65952
rect 16393 65943 16451 65949
rect 16393 65940 16405 65943
rect 15528 65912 16405 65940
rect 15528 65900 15534 65912
rect 16393 65909 16405 65912
rect 16439 65909 16451 65943
rect 17218 65940 17224 65952
rect 17179 65912 17224 65940
rect 16393 65903 16451 65909
rect 17218 65900 17224 65912
rect 17276 65900 17282 65952
rect 1104 65850 28888 65872
rect 1104 65798 10982 65850
rect 11034 65798 11046 65850
rect 11098 65798 11110 65850
rect 11162 65798 11174 65850
rect 11226 65798 20982 65850
rect 21034 65798 21046 65850
rect 21098 65798 21110 65850
rect 21162 65798 21174 65850
rect 21226 65798 28888 65850
rect 1104 65776 28888 65798
rect 18598 65668 18604 65680
rect 18559 65640 18604 65668
rect 18598 65628 18604 65640
rect 18656 65628 18662 65680
rect 14366 65560 14372 65612
rect 14424 65600 14430 65612
rect 15289 65603 15347 65609
rect 15289 65600 15301 65603
rect 14424 65572 15301 65600
rect 14424 65560 14430 65572
rect 15289 65569 15301 65572
rect 15335 65569 15347 65603
rect 15654 65600 15660 65612
rect 15615 65572 15660 65600
rect 15289 65563 15347 65569
rect 15654 65560 15660 65572
rect 15712 65560 15718 65612
rect 15838 65560 15844 65612
rect 15896 65600 15902 65612
rect 16117 65603 16175 65609
rect 16117 65600 16129 65603
rect 15896 65572 16129 65600
rect 15896 65560 15902 65572
rect 16117 65569 16129 65572
rect 16163 65569 16175 65603
rect 17862 65600 17868 65612
rect 17823 65572 17868 65600
rect 16117 65563 16175 65569
rect 17862 65560 17868 65572
rect 17920 65560 17926 65612
rect 17954 65560 17960 65612
rect 18012 65600 18018 65612
rect 18230 65600 18236 65612
rect 18012 65572 18236 65600
rect 18012 65560 18018 65572
rect 18230 65560 18236 65572
rect 18288 65600 18294 65612
rect 18325 65603 18383 65609
rect 18325 65600 18337 65603
rect 18288 65572 18337 65600
rect 18288 65560 18294 65572
rect 18325 65569 18337 65572
rect 18371 65569 18383 65603
rect 18325 65563 18383 65569
rect 17586 65532 17592 65544
rect 17547 65504 17592 65532
rect 17586 65492 17592 65504
rect 17644 65492 17650 65544
rect 24946 65492 24952 65544
rect 25004 65532 25010 65544
rect 25774 65532 25780 65544
rect 25004 65504 25780 65532
rect 25004 65492 25010 65504
rect 25774 65492 25780 65504
rect 25832 65492 25838 65544
rect 15194 65424 15200 65476
rect 15252 65464 15258 65476
rect 16117 65467 16175 65473
rect 16117 65464 16129 65467
rect 15252 65436 16129 65464
rect 15252 65424 15258 65436
rect 16117 65433 16129 65436
rect 16163 65433 16175 65467
rect 16117 65427 16175 65433
rect 1104 65306 28888 65328
rect 1104 65254 5982 65306
rect 6034 65254 6046 65306
rect 6098 65254 6110 65306
rect 6162 65254 6174 65306
rect 6226 65254 15982 65306
rect 16034 65254 16046 65306
rect 16098 65254 16110 65306
rect 16162 65254 16174 65306
rect 16226 65254 25982 65306
rect 26034 65254 26046 65306
rect 26098 65254 26110 65306
rect 26162 65254 26174 65306
rect 26226 65254 28888 65306
rect 1104 65232 28888 65254
rect 17129 65195 17187 65201
rect 17129 65192 17141 65195
rect 14660 65164 17141 65192
rect 14366 65016 14372 65068
rect 14424 65056 14430 65068
rect 14660 65065 14688 65164
rect 17129 65161 17141 65164
rect 17175 65192 17187 65195
rect 17862 65192 17868 65204
rect 17175 65164 17868 65192
rect 17175 65161 17187 65164
rect 17129 65155 17187 65161
rect 17862 65152 17868 65164
rect 17920 65152 17926 65204
rect 21637 65195 21695 65201
rect 21637 65161 21649 65195
rect 21683 65192 21695 65195
rect 21818 65192 21824 65204
rect 21683 65164 21824 65192
rect 21683 65161 21695 65164
rect 21637 65155 21695 65161
rect 21818 65152 21824 65164
rect 21876 65152 21882 65204
rect 24397 65195 24455 65201
rect 24397 65161 24409 65195
rect 24443 65192 24455 65195
rect 24762 65192 24768 65204
rect 24443 65164 24768 65192
rect 24443 65161 24455 65164
rect 24397 65155 24455 65161
rect 24762 65152 24768 65164
rect 24820 65152 24826 65204
rect 15378 65084 15384 65136
rect 15436 65124 15442 65136
rect 16025 65127 16083 65133
rect 16025 65124 16037 65127
rect 15436 65096 16037 65124
rect 15436 65084 15442 65096
rect 16025 65093 16037 65096
rect 16071 65093 16083 65127
rect 16025 65087 16083 65093
rect 14645 65059 14703 65065
rect 14645 65056 14657 65059
rect 14424 65028 14657 65056
rect 14424 65016 14430 65028
rect 14645 65025 14657 65028
rect 14691 65025 14703 65059
rect 14645 65019 14703 65025
rect 15105 65059 15163 65065
rect 15105 65025 15117 65059
rect 15151 65056 15163 65059
rect 15289 65059 15347 65065
rect 15289 65056 15301 65059
rect 15151 65028 15301 65056
rect 15151 65025 15163 65028
rect 15105 65019 15163 65025
rect 15289 65025 15301 65028
rect 15335 65056 15347 65059
rect 17218 65056 17224 65068
rect 15335 65028 17224 65056
rect 15335 65025 15347 65028
rect 15289 65019 15347 65025
rect 17218 65016 17224 65028
rect 17276 65016 17282 65068
rect 21836 65056 21864 65152
rect 24857 65059 24915 65065
rect 24857 65056 24869 65059
rect 21836 65028 24869 65056
rect 15565 64991 15623 64997
rect 15565 64957 15577 64991
rect 15611 64988 15623 64991
rect 15611 64960 15645 64988
rect 15611 64957 15623 64960
rect 15565 64951 15623 64957
rect 14369 64923 14427 64929
rect 14369 64889 14381 64923
rect 14415 64920 14427 64923
rect 15580 64920 15608 64951
rect 15838 64948 15844 65000
rect 15896 64988 15902 65000
rect 24596 64997 24624 65028
rect 24857 65025 24869 65028
rect 24903 65025 24915 65059
rect 24857 65019 24915 65025
rect 16025 64991 16083 64997
rect 16025 64988 16037 64991
rect 15896 64960 16037 64988
rect 15896 64948 15902 64960
rect 16025 64957 16037 64960
rect 16071 64988 16083 64991
rect 16577 64991 16635 64997
rect 16577 64988 16589 64991
rect 16071 64960 16589 64988
rect 16071 64957 16083 64960
rect 16025 64951 16083 64957
rect 16577 64957 16589 64960
rect 16623 64957 16635 64991
rect 16577 64951 16635 64957
rect 21821 64991 21879 64997
rect 21821 64957 21833 64991
rect 21867 64957 21879 64991
rect 21821 64951 21879 64957
rect 24581 64991 24639 64997
rect 24581 64957 24593 64991
rect 24627 64957 24639 64991
rect 24581 64951 24639 64957
rect 15654 64920 15660 64932
rect 14415 64892 15660 64920
rect 14415 64889 14427 64892
rect 14369 64883 14427 64889
rect 15654 64880 15660 64892
rect 15712 64880 15718 64932
rect 17586 64920 17592 64932
rect 17547 64892 17592 64920
rect 17586 64880 17592 64892
rect 17644 64880 17650 64932
rect 18230 64920 18236 64932
rect 18191 64892 18236 64920
rect 18230 64880 18236 64892
rect 18288 64880 18294 64932
rect 21836 64920 21864 64951
rect 22189 64923 22247 64929
rect 22189 64920 22201 64923
rect 21836 64892 22201 64920
rect 22189 64889 22201 64892
rect 22235 64920 22247 64923
rect 22462 64920 22468 64932
rect 22235 64892 22468 64920
rect 22235 64889 22247 64892
rect 22189 64883 22247 64889
rect 22462 64880 22468 64892
rect 22520 64880 22526 64932
rect 1104 64762 28888 64784
rect 1104 64710 10982 64762
rect 11034 64710 11046 64762
rect 11098 64710 11110 64762
rect 11162 64710 11174 64762
rect 11226 64710 20982 64762
rect 21034 64710 21046 64762
rect 21098 64710 21110 64762
rect 21162 64710 21174 64762
rect 21226 64710 28888 64762
rect 1104 64688 28888 64710
rect 20714 64472 20720 64524
rect 20772 64512 20778 64524
rect 21542 64512 21548 64524
rect 20772 64484 21548 64512
rect 20772 64472 20778 64484
rect 21542 64472 21548 64484
rect 21600 64512 21606 64524
rect 21729 64515 21787 64521
rect 21729 64512 21741 64515
rect 21600 64484 21741 64512
rect 21600 64472 21606 64484
rect 21729 64481 21741 64484
rect 21775 64481 21787 64515
rect 21729 64475 21787 64481
rect 21453 64447 21511 64453
rect 21453 64413 21465 64447
rect 21499 64444 21511 64447
rect 21634 64444 21640 64456
rect 21499 64416 21640 64444
rect 21499 64413 21511 64416
rect 21453 64407 21511 64413
rect 21634 64404 21640 64416
rect 21692 64404 21698 64456
rect 15105 64379 15163 64385
rect 15105 64345 15117 64379
rect 15151 64376 15163 64379
rect 15838 64376 15844 64388
rect 15151 64348 15844 64376
rect 15151 64345 15163 64348
rect 15105 64339 15163 64345
rect 15838 64336 15844 64348
rect 15896 64336 15902 64388
rect 15565 64311 15623 64317
rect 15565 64277 15577 64311
rect 15611 64308 15623 64311
rect 15654 64308 15660 64320
rect 15611 64280 15660 64308
rect 15611 64277 15623 64280
rect 15565 64271 15623 64277
rect 15654 64268 15660 64280
rect 15712 64308 15718 64320
rect 15933 64311 15991 64317
rect 15933 64308 15945 64311
rect 15712 64280 15945 64308
rect 15712 64268 15718 64280
rect 15933 64277 15945 64280
rect 15979 64277 15991 64311
rect 15933 64271 15991 64277
rect 23017 64311 23075 64317
rect 23017 64277 23029 64311
rect 23063 64308 23075 64311
rect 23474 64308 23480 64320
rect 23063 64280 23480 64308
rect 23063 64277 23075 64280
rect 23017 64271 23075 64277
rect 23474 64268 23480 64280
rect 23532 64268 23538 64320
rect 1104 64218 28888 64240
rect 1104 64166 5982 64218
rect 6034 64166 6046 64218
rect 6098 64166 6110 64218
rect 6162 64166 6174 64218
rect 6226 64166 15982 64218
rect 16034 64166 16046 64218
rect 16098 64166 16110 64218
rect 16162 64166 16174 64218
rect 16226 64166 25982 64218
rect 26034 64166 26046 64218
rect 26098 64166 26110 64218
rect 26162 64166 26174 64218
rect 26226 64166 28888 64218
rect 1104 64144 28888 64166
rect 21542 64104 21548 64116
rect 21503 64076 21548 64104
rect 21542 64064 21548 64076
rect 21600 64064 21606 64116
rect 21634 64064 21640 64116
rect 21692 64104 21698 64116
rect 21821 64107 21879 64113
rect 21821 64104 21833 64107
rect 21692 64076 21833 64104
rect 21692 64064 21698 64076
rect 21821 64073 21833 64076
rect 21867 64073 21879 64107
rect 21821 64067 21879 64073
rect 15654 63928 15660 63980
rect 15712 63968 15718 63980
rect 17034 63968 17040 63980
rect 15712 63940 16344 63968
rect 16995 63940 17040 63968
rect 15712 63928 15718 63940
rect 15841 63903 15899 63909
rect 15841 63869 15853 63903
rect 15887 63900 15899 63903
rect 16117 63903 16175 63909
rect 16117 63900 16129 63903
rect 15887 63872 16129 63900
rect 15887 63869 15899 63872
rect 15841 63863 15899 63869
rect 16117 63869 16129 63872
rect 16163 63900 16175 63903
rect 16206 63900 16212 63912
rect 16163 63872 16212 63900
rect 16163 63869 16175 63872
rect 16117 63863 16175 63869
rect 16206 63860 16212 63872
rect 16264 63860 16270 63912
rect 16316 63909 16344 63940
rect 17034 63928 17040 63940
rect 17092 63928 17098 63980
rect 18598 63968 18604 63980
rect 18559 63940 18604 63968
rect 18598 63928 18604 63940
rect 18656 63968 18662 63980
rect 19061 63971 19119 63977
rect 19061 63968 19073 63971
rect 18656 63940 19073 63968
rect 18656 63928 18662 63940
rect 19061 63937 19073 63940
rect 19107 63937 19119 63971
rect 19061 63931 19119 63937
rect 16301 63903 16359 63909
rect 16301 63869 16313 63903
rect 16347 63869 16359 63903
rect 16301 63863 16359 63869
rect 16761 63903 16819 63909
rect 16761 63869 16773 63903
rect 16807 63869 16819 63903
rect 16761 63863 16819 63869
rect 18785 63903 18843 63909
rect 18785 63869 18797 63903
rect 18831 63900 18843 63903
rect 18874 63900 18880 63912
rect 18831 63872 18880 63900
rect 18831 63869 18843 63872
rect 18785 63863 18843 63869
rect 16776 63832 16804 63863
rect 18874 63860 18880 63872
rect 18932 63860 18938 63912
rect 20438 63832 20444 63844
rect 15764 63804 16804 63832
rect 20399 63804 20444 63832
rect 15764 63776 15792 63804
rect 20438 63792 20444 63804
rect 20496 63792 20502 63844
rect 15473 63767 15531 63773
rect 15473 63733 15485 63767
rect 15519 63764 15531 63767
rect 15746 63764 15752 63776
rect 15519 63736 15752 63764
rect 15519 63733 15531 63736
rect 15473 63727 15531 63733
rect 15746 63724 15752 63736
rect 15804 63724 15810 63776
rect 1104 63674 28888 63696
rect 1104 63622 10982 63674
rect 11034 63622 11046 63674
rect 11098 63622 11110 63674
rect 11162 63622 11174 63674
rect 11226 63622 20982 63674
rect 21034 63622 21046 63674
rect 21098 63622 21110 63674
rect 21162 63622 21174 63674
rect 21226 63622 28888 63674
rect 1104 63600 28888 63622
rect 18874 63560 18880 63572
rect 18835 63532 18880 63560
rect 18874 63520 18880 63532
rect 18932 63520 18938 63572
rect 23658 63492 23664 63504
rect 23619 63464 23664 63492
rect 23658 63452 23664 63464
rect 23716 63452 23722 63504
rect 15654 63424 15660 63436
rect 15615 63396 15660 63424
rect 15654 63384 15660 63396
rect 15712 63384 15718 63436
rect 15746 63384 15752 63436
rect 15804 63424 15810 63436
rect 16117 63427 16175 63433
rect 16117 63424 16129 63427
rect 15804 63396 16129 63424
rect 15804 63384 15810 63396
rect 16117 63393 16129 63396
rect 16163 63393 16175 63427
rect 16117 63387 16175 63393
rect 23569 63427 23627 63433
rect 23569 63393 23581 63427
rect 23615 63424 23627 63427
rect 24210 63424 24216 63436
rect 23615 63396 24216 63424
rect 23615 63393 23627 63396
rect 23569 63387 23627 63393
rect 24210 63384 24216 63396
rect 24268 63384 24274 63436
rect 24394 63424 24400 63436
rect 24355 63396 24400 63424
rect 24394 63384 24400 63396
rect 24452 63384 24458 63436
rect 15473 63359 15531 63365
rect 15473 63325 15485 63359
rect 15519 63356 15531 63359
rect 15562 63356 15568 63368
rect 15519 63328 15568 63356
rect 15519 63325 15531 63328
rect 15473 63319 15531 63325
rect 15562 63316 15568 63328
rect 15620 63316 15626 63368
rect 24026 63316 24032 63368
rect 24084 63356 24090 63368
rect 24489 63359 24547 63365
rect 24489 63356 24501 63359
rect 24084 63328 24501 63356
rect 24084 63316 24090 63328
rect 24489 63325 24501 63328
rect 24535 63325 24547 63359
rect 24489 63319 24547 63325
rect 15102 63248 15108 63300
rect 15160 63288 15166 63300
rect 16117 63291 16175 63297
rect 16117 63288 16129 63291
rect 15160 63260 16129 63288
rect 15160 63248 15166 63260
rect 16117 63257 16129 63260
rect 16163 63257 16175 63291
rect 16117 63251 16175 63257
rect 1104 63130 28888 63152
rect 1104 63078 5982 63130
rect 6034 63078 6046 63130
rect 6098 63078 6110 63130
rect 6162 63078 6174 63130
rect 6226 63078 15982 63130
rect 16034 63078 16046 63130
rect 16098 63078 16110 63130
rect 16162 63078 16174 63130
rect 16226 63078 25982 63130
rect 26034 63078 26046 63130
rect 26098 63078 26110 63130
rect 26162 63078 26174 63130
rect 26226 63078 28888 63130
rect 1104 63056 28888 63078
rect 23474 63016 23480 63028
rect 23435 62988 23480 63016
rect 23474 62976 23480 62988
rect 23532 63016 23538 63028
rect 24394 63016 24400 63028
rect 23532 62988 24400 63016
rect 23532 62976 23538 62988
rect 24394 62976 24400 62988
rect 24452 62976 24458 63028
rect 25866 62840 25872 62892
rect 25924 62880 25930 62892
rect 26053 62883 26111 62889
rect 26053 62880 26065 62883
rect 25924 62852 26065 62880
rect 25924 62840 25930 62852
rect 26053 62849 26065 62852
rect 26099 62880 26111 62883
rect 26421 62883 26479 62889
rect 26421 62880 26433 62883
rect 26099 62852 26433 62880
rect 26099 62849 26111 62852
rect 26053 62843 26111 62849
rect 26421 62849 26433 62852
rect 26467 62849 26479 62883
rect 26421 62843 26479 62849
rect 27614 62840 27620 62892
rect 27672 62880 27678 62892
rect 27798 62880 27804 62892
rect 27672 62852 27804 62880
rect 27672 62840 27678 62852
rect 27798 62840 27804 62852
rect 27856 62840 27862 62892
rect 14090 62772 14096 62824
rect 14148 62812 14154 62824
rect 15654 62812 15660 62824
rect 14148 62784 15660 62812
rect 14148 62772 14154 62784
rect 15654 62772 15660 62784
rect 15712 62772 15718 62824
rect 23937 62815 23995 62821
rect 23937 62781 23949 62815
rect 23983 62812 23995 62815
rect 24210 62812 24216 62824
rect 23983 62784 24216 62812
rect 23983 62781 23995 62784
rect 23937 62775 23995 62781
rect 24210 62772 24216 62784
rect 24268 62772 24274 62824
rect 24854 62772 24860 62824
rect 24912 62812 24918 62824
rect 26142 62812 26148 62824
rect 24912 62784 26148 62812
rect 24912 62772 24918 62784
rect 26142 62772 26148 62784
rect 26200 62772 26206 62824
rect 13354 62704 13360 62756
rect 13412 62744 13418 62756
rect 15746 62744 15752 62756
rect 13412 62716 15752 62744
rect 13412 62704 13418 62716
rect 15746 62704 15752 62716
rect 15804 62744 15810 62756
rect 16025 62747 16083 62753
rect 16025 62744 16037 62747
rect 15804 62716 16037 62744
rect 15804 62704 15810 62716
rect 16025 62713 16037 62716
rect 16071 62713 16083 62747
rect 27798 62744 27804 62756
rect 27759 62716 27804 62744
rect 16025 62707 16083 62713
rect 27798 62704 27804 62716
rect 27856 62704 27862 62756
rect 15381 62679 15439 62685
rect 15381 62645 15393 62679
rect 15427 62676 15439 62679
rect 15562 62676 15568 62688
rect 15427 62648 15568 62676
rect 15427 62645 15439 62648
rect 15381 62639 15439 62645
rect 15562 62636 15568 62648
rect 15620 62636 15626 62688
rect 24026 62636 24032 62688
rect 24084 62676 24090 62688
rect 24213 62679 24271 62685
rect 24213 62676 24225 62679
rect 24084 62648 24225 62676
rect 24084 62636 24090 62648
rect 24213 62645 24225 62648
rect 24259 62645 24271 62679
rect 24213 62639 24271 62645
rect 1104 62586 28888 62608
rect 1104 62534 10982 62586
rect 11034 62534 11046 62586
rect 11098 62534 11110 62586
rect 11162 62534 11174 62586
rect 11226 62534 20982 62586
rect 21034 62534 21046 62586
rect 21098 62534 21110 62586
rect 21162 62534 21174 62586
rect 21226 62534 28888 62586
rect 1104 62512 28888 62534
rect 15470 62432 15476 62484
rect 15528 62472 15534 62484
rect 15654 62472 15660 62484
rect 15528 62444 15660 62472
rect 15528 62432 15534 62444
rect 15654 62432 15660 62444
rect 15712 62432 15718 62484
rect 25866 62432 25872 62484
rect 25924 62472 25930 62484
rect 26142 62472 26148 62484
rect 25924 62444 26148 62472
rect 25924 62432 25930 62444
rect 26142 62432 26148 62444
rect 26200 62432 26206 62484
rect 15838 62364 15844 62416
rect 15896 62404 15902 62416
rect 15933 62407 15991 62413
rect 15933 62404 15945 62407
rect 15896 62376 15945 62404
rect 15896 62364 15902 62376
rect 15933 62373 15945 62376
rect 15979 62373 15991 62407
rect 15933 62367 15991 62373
rect 13722 62296 13728 62348
rect 13780 62336 13786 62348
rect 15470 62336 15476 62348
rect 13780 62308 15476 62336
rect 13780 62296 13786 62308
rect 15470 62296 15476 62308
rect 15528 62296 15534 62348
rect 16298 62296 16304 62348
rect 16356 62336 16362 62348
rect 16761 62339 16819 62345
rect 16761 62336 16773 62339
rect 16356 62308 16773 62336
rect 16356 62296 16362 62308
rect 16761 62305 16773 62308
rect 16807 62305 16819 62339
rect 16761 62299 16819 62305
rect 16485 62271 16543 62277
rect 16485 62237 16497 62271
rect 16531 62268 16543 62271
rect 16666 62268 16672 62280
rect 16531 62240 16672 62268
rect 16531 62237 16543 62240
rect 16485 62231 16543 62237
rect 16666 62228 16672 62240
rect 16724 62228 16730 62280
rect 16945 62271 17003 62277
rect 16945 62237 16957 62271
rect 16991 62237 17003 62271
rect 16945 62231 17003 62237
rect 16574 62160 16580 62212
rect 16632 62200 16638 62212
rect 16960 62200 16988 62231
rect 17862 62200 17868 62212
rect 16632 62172 17868 62200
rect 16632 62160 16638 62172
rect 17862 62160 17868 62172
rect 17920 62160 17926 62212
rect 19061 62135 19119 62141
rect 19061 62101 19073 62135
rect 19107 62132 19119 62135
rect 19242 62132 19248 62144
rect 19107 62104 19248 62132
rect 19107 62101 19119 62104
rect 19061 62095 19119 62101
rect 19242 62092 19248 62104
rect 19300 62092 19306 62144
rect 1104 62042 28888 62064
rect 1104 61990 5982 62042
rect 6034 61990 6046 62042
rect 6098 61990 6110 62042
rect 6162 61990 6174 62042
rect 6226 61990 15982 62042
rect 16034 61990 16046 62042
rect 16098 61990 16110 62042
rect 16162 61990 16174 62042
rect 16226 61990 25982 62042
rect 26034 61990 26046 62042
rect 26098 61990 26110 62042
rect 26162 61990 26174 62042
rect 26226 61990 28888 62042
rect 1104 61968 28888 61990
rect 13814 61928 13820 61940
rect 13775 61900 13820 61928
rect 13814 61888 13820 61900
rect 13872 61888 13878 61940
rect 12434 61752 12440 61804
rect 12492 61792 12498 61804
rect 20070 61792 20076 61804
rect 12492 61764 12537 61792
rect 20031 61764 20076 61792
rect 12492 61752 12498 61764
rect 20070 61752 20076 61764
rect 20128 61752 20134 61804
rect 25774 61752 25780 61804
rect 25832 61792 25838 61804
rect 26053 61795 26111 61801
rect 26053 61792 26065 61795
rect 25832 61764 26065 61792
rect 25832 61752 25838 61764
rect 26053 61761 26065 61764
rect 26099 61792 26111 61795
rect 26421 61795 26479 61801
rect 26421 61792 26433 61795
rect 26099 61764 26433 61792
rect 26099 61761 26111 61764
rect 26053 61755 26111 61761
rect 26421 61761 26433 61764
rect 26467 61761 26479 61795
rect 26421 61755 26479 61761
rect 12158 61724 12164 61736
rect 12119 61696 12164 61724
rect 12158 61684 12164 61696
rect 12216 61724 12222 61736
rect 12713 61727 12771 61733
rect 12713 61724 12725 61727
rect 12216 61696 12725 61724
rect 12216 61684 12222 61696
rect 12713 61693 12725 61696
rect 12759 61693 12771 61727
rect 18969 61727 19027 61733
rect 18969 61724 18981 61727
rect 12713 61687 12771 61693
rect 18800 61696 18981 61724
rect 16574 61656 16580 61668
rect 15948 61628 16580 61656
rect 15838 61548 15844 61600
rect 15896 61588 15902 61600
rect 15948 61597 15976 61628
rect 16574 61616 16580 61628
rect 16632 61616 16638 61668
rect 18800 61600 18828 61696
rect 18969 61693 18981 61696
rect 19015 61693 19027 61727
rect 18969 61687 19027 61693
rect 19242 61684 19248 61736
rect 19300 61724 19306 61736
rect 19337 61727 19395 61733
rect 19337 61724 19349 61727
rect 19300 61696 19349 61724
rect 19300 61684 19306 61696
rect 19337 61693 19349 61696
rect 19383 61693 19395 61727
rect 19337 61687 19395 61693
rect 19426 61684 19432 61736
rect 19484 61724 19490 61736
rect 19794 61724 19800 61736
rect 19484 61696 19800 61724
rect 19484 61684 19490 61696
rect 19794 61684 19800 61696
rect 19852 61684 19858 61736
rect 25866 61684 25872 61736
rect 25924 61724 25930 61736
rect 26145 61727 26203 61733
rect 26145 61724 26157 61727
rect 25924 61696 26157 61724
rect 25924 61684 25930 61696
rect 26145 61693 26157 61696
rect 26191 61693 26203 61727
rect 26145 61687 26203 61693
rect 27801 61659 27859 61665
rect 27801 61625 27813 61659
rect 27847 61656 27859 61659
rect 28074 61656 28080 61668
rect 27847 61628 28080 61656
rect 27847 61625 27859 61628
rect 27801 61619 27859 61625
rect 28074 61616 28080 61628
rect 28132 61616 28138 61668
rect 15933 61591 15991 61597
rect 15933 61588 15945 61591
rect 15896 61560 15945 61588
rect 15896 61548 15902 61560
rect 15933 61557 15945 61560
rect 15979 61557 15991 61591
rect 16298 61588 16304 61600
rect 16259 61560 16304 61588
rect 15933 61551 15991 61557
rect 16298 61548 16304 61560
rect 16356 61548 16362 61600
rect 16666 61588 16672 61600
rect 16627 61560 16672 61588
rect 16666 61548 16672 61560
rect 16724 61548 16730 61600
rect 17313 61591 17371 61597
rect 17313 61557 17325 61591
rect 17359 61588 17371 61591
rect 17678 61588 17684 61600
rect 17359 61560 17684 61588
rect 17359 61557 17371 61560
rect 17313 61551 17371 61557
rect 17678 61548 17684 61560
rect 17736 61588 17742 61600
rect 18046 61588 18052 61600
rect 17736 61560 18052 61588
rect 17736 61548 17742 61560
rect 18046 61548 18052 61560
rect 18104 61548 18110 61600
rect 18782 61588 18788 61600
rect 18743 61560 18788 61588
rect 18782 61548 18788 61560
rect 18840 61548 18846 61600
rect 1104 61498 28888 61520
rect 1104 61446 10982 61498
rect 11034 61446 11046 61498
rect 11098 61446 11110 61498
rect 11162 61446 11174 61498
rect 11226 61446 20982 61498
rect 21034 61446 21046 61498
rect 21098 61446 21110 61498
rect 21162 61446 21174 61498
rect 21226 61446 28888 61498
rect 1104 61424 28888 61446
rect 1578 61384 1584 61396
rect 1539 61356 1584 61384
rect 1578 61344 1584 61356
rect 1636 61344 1642 61396
rect 12434 61344 12440 61396
rect 12492 61384 12498 61396
rect 20714 61384 20720 61396
rect 12492 61356 12537 61384
rect 20675 61356 20720 61384
rect 12492 61344 12498 61356
rect 20714 61344 20720 61356
rect 20772 61344 20778 61396
rect 25866 61344 25872 61396
rect 25924 61384 25930 61396
rect 26145 61387 26203 61393
rect 26145 61384 26157 61387
rect 25924 61356 26157 61384
rect 25924 61344 25930 61356
rect 26145 61353 26157 61356
rect 26191 61353 26203 61387
rect 26145 61347 26203 61353
rect 17862 61276 17868 61328
rect 17920 61316 17926 61328
rect 21450 61316 21456 61328
rect 17920 61288 19196 61316
rect 21411 61288 21456 61316
rect 17920 61276 17926 61288
rect 19168 61260 19196 61288
rect 21450 61276 21456 61288
rect 21508 61276 21514 61328
rect 26694 61316 26700 61328
rect 26655 61288 26700 61316
rect 26694 61276 26700 61288
rect 26752 61276 26758 61328
rect 17129 61251 17187 61257
rect 17129 61217 17141 61251
rect 17175 61248 17187 61251
rect 17773 61251 17831 61257
rect 17773 61248 17785 61251
rect 17175 61220 17785 61248
rect 17175 61217 17187 61220
rect 17129 61211 17187 61217
rect 17773 61217 17785 61220
rect 17819 61217 17831 61251
rect 18046 61248 18052 61260
rect 18007 61220 18052 61248
rect 17773 61211 17831 61217
rect 17405 61183 17463 61189
rect 17405 61149 17417 61183
rect 17451 61180 17463 61183
rect 17494 61180 17500 61192
rect 17451 61152 17500 61180
rect 17451 61149 17463 61152
rect 17405 61143 17463 61149
rect 17494 61140 17500 61152
rect 17552 61140 17558 61192
rect 17788 61180 17816 61211
rect 18046 61208 18052 61220
rect 18104 61208 18110 61260
rect 19150 61248 19156 61260
rect 19063 61220 19156 61248
rect 19150 61208 19156 61220
rect 19208 61208 19214 61260
rect 21177 61251 21235 61257
rect 21177 61217 21189 61251
rect 21223 61248 21235 61251
rect 22002 61248 22008 61260
rect 21223 61220 22008 61248
rect 21223 61217 21235 61220
rect 21177 61211 21235 61217
rect 22002 61208 22008 61220
rect 22060 61248 22066 61260
rect 22189 61251 22247 61257
rect 22189 61248 22201 61251
rect 22060 61220 22201 61248
rect 22060 61208 22066 61220
rect 22189 61217 22201 61220
rect 22235 61217 22247 61251
rect 22189 61211 22247 61217
rect 27338 61208 27344 61260
rect 27396 61248 27402 61260
rect 27433 61251 27491 61257
rect 27433 61248 27445 61251
rect 27396 61220 27445 61248
rect 27396 61208 27402 61220
rect 27433 61217 27445 61220
rect 27479 61248 27491 61251
rect 27798 61248 27804 61260
rect 27479 61220 27804 61248
rect 27479 61217 27491 61220
rect 27433 61211 27491 61217
rect 27798 61208 27804 61220
rect 27856 61208 27862 61260
rect 21358 61180 21364 61192
rect 17788 61152 19104 61180
rect 21319 61152 21364 61180
rect 17954 61072 17960 61124
rect 18012 61112 18018 61124
rect 19076 61121 19104 61152
rect 21358 61140 21364 61152
rect 21416 61140 21422 61192
rect 22281 61183 22339 61189
rect 22281 61149 22293 61183
rect 22327 61180 22339 61183
rect 22830 61180 22836 61192
rect 22327 61152 22836 61180
rect 22327 61149 22339 61152
rect 22281 61143 22339 61149
rect 22830 61140 22836 61152
rect 22888 61140 22894 61192
rect 26510 61140 26516 61192
rect 26568 61180 26574 61192
rect 26605 61183 26663 61189
rect 26605 61180 26617 61183
rect 26568 61152 26617 61180
rect 26568 61140 26574 61152
rect 26605 61149 26617 61152
rect 26651 61149 26663 61183
rect 26605 61143 26663 61149
rect 26878 61140 26884 61192
rect 26936 61180 26942 61192
rect 27525 61183 27583 61189
rect 27525 61180 27537 61183
rect 26936 61152 27537 61180
rect 26936 61140 26942 61152
rect 27525 61149 27537 61152
rect 27571 61149 27583 61183
rect 27525 61143 27583 61149
rect 18049 61115 18107 61121
rect 18049 61112 18061 61115
rect 18012 61084 18061 61112
rect 18012 61072 18018 61084
rect 18049 61081 18061 61084
rect 18095 61081 18107 61115
rect 18049 61075 18107 61081
rect 19061 61115 19119 61121
rect 19061 61081 19073 61115
rect 19107 61112 19119 61115
rect 19242 61112 19248 61124
rect 19107 61084 19248 61112
rect 19107 61081 19119 61084
rect 19061 61075 19119 61081
rect 19242 61072 19248 61084
rect 19300 61112 19306 61124
rect 21266 61112 21272 61124
rect 19300 61084 21272 61112
rect 19300 61072 19306 61084
rect 21266 61072 21272 61084
rect 21324 61072 21330 61124
rect 16209 61047 16267 61053
rect 16209 61013 16221 61047
rect 16255 61044 16267 61047
rect 16574 61044 16580 61056
rect 16255 61016 16580 61044
rect 16255 61013 16267 61016
rect 16209 61007 16267 61013
rect 16574 61004 16580 61016
rect 16632 61004 16638 61056
rect 18598 61044 18604 61056
rect 18559 61016 18604 61044
rect 18598 61004 18604 61016
rect 18656 61004 18662 61056
rect 19337 61047 19395 61053
rect 19337 61013 19349 61047
rect 19383 61044 19395 61047
rect 19610 61044 19616 61056
rect 19383 61016 19616 61044
rect 19383 61013 19395 61016
rect 19337 61007 19395 61013
rect 19610 61004 19616 61016
rect 19668 61004 19674 61056
rect 20806 61004 20812 61056
rect 20864 61044 20870 61056
rect 21450 61044 21456 61056
rect 20864 61016 21456 61044
rect 20864 61004 20870 61016
rect 21450 61004 21456 61016
rect 21508 61004 21514 61056
rect 1104 60954 28888 60976
rect 1104 60902 5982 60954
rect 6034 60902 6046 60954
rect 6098 60902 6110 60954
rect 6162 60902 6174 60954
rect 6226 60902 15982 60954
rect 16034 60902 16046 60954
rect 16098 60902 16110 60954
rect 16162 60902 16174 60954
rect 16226 60902 25982 60954
rect 26034 60902 26046 60954
rect 26098 60902 26110 60954
rect 26162 60902 26174 60954
rect 26226 60902 28888 60954
rect 1104 60880 28888 60902
rect 2774 60800 2780 60852
rect 2832 60840 2838 60852
rect 2832 60812 2877 60840
rect 2832 60800 2838 60812
rect 19058 60800 19064 60852
rect 19116 60840 19122 60852
rect 19242 60840 19248 60852
rect 19116 60812 19248 60840
rect 19116 60800 19122 60812
rect 19242 60800 19248 60812
rect 19300 60800 19306 60852
rect 22002 60840 22008 60852
rect 21963 60812 22008 60840
rect 22002 60800 22008 60812
rect 22060 60800 22066 60852
rect 22830 60800 22836 60852
rect 22888 60840 22894 60852
rect 22925 60843 22983 60849
rect 22925 60840 22937 60843
rect 22888 60812 22937 60840
rect 22888 60800 22894 60812
rect 22925 60809 22937 60812
rect 22971 60840 22983 60843
rect 25498 60840 25504 60852
rect 22971 60812 25504 60840
rect 22971 60809 22983 60812
rect 22925 60803 22983 60809
rect 25498 60800 25504 60812
rect 25556 60840 25562 60852
rect 26878 60840 26884 60852
rect 25556 60812 26884 60840
rect 25556 60800 25562 60812
rect 26878 60800 26884 60812
rect 26936 60800 26942 60852
rect 27338 60840 27344 60852
rect 27299 60812 27344 60840
rect 27338 60800 27344 60812
rect 27396 60800 27402 60852
rect 18874 60772 18880 60784
rect 18835 60744 18880 60772
rect 18874 60732 18880 60744
rect 18932 60732 18938 60784
rect 19150 60732 19156 60784
rect 19208 60772 19214 60784
rect 19208 60744 19288 60772
rect 19208 60732 19214 60744
rect 1397 60707 1455 60713
rect 1397 60673 1409 60707
rect 1443 60704 1455 60707
rect 1578 60704 1584 60716
rect 1443 60676 1584 60704
rect 1443 60673 1455 60676
rect 1397 60667 1455 60673
rect 1578 60664 1584 60676
rect 1636 60664 1642 60716
rect 15654 60664 15660 60716
rect 15712 60704 15718 60716
rect 16117 60707 16175 60713
rect 16117 60704 16129 60707
rect 15712 60676 16129 60704
rect 15712 60664 15718 60676
rect 16117 60673 16129 60676
rect 16163 60673 16175 60707
rect 16807 60707 16865 60713
rect 16807 60704 16819 60707
rect 16117 60667 16175 60673
rect 16500 60676 16819 60704
rect 1670 60636 1676 60648
rect 1631 60608 1676 60636
rect 1670 60596 1676 60608
rect 1728 60596 1734 60648
rect 16025 60639 16083 60645
rect 16025 60605 16037 60639
rect 16071 60636 16083 60639
rect 16500 60636 16528 60676
rect 16807 60673 16819 60676
rect 16853 60704 16865 60707
rect 17034 60704 17040 60716
rect 16853 60676 17040 60704
rect 16853 60673 16865 60676
rect 16807 60667 16865 60673
rect 17034 60664 17040 60676
rect 17092 60664 17098 60716
rect 17494 60704 17500 60716
rect 17455 60676 17500 60704
rect 17494 60664 17500 60676
rect 17552 60664 17558 60716
rect 19260 60704 19288 60744
rect 19429 60707 19487 60713
rect 19429 60704 19441 60707
rect 19260 60676 19441 60704
rect 19429 60673 19441 60676
rect 19475 60673 19487 60707
rect 20622 60704 20628 60716
rect 20583 60676 20628 60704
rect 19429 60667 19487 60673
rect 20622 60664 20628 60676
rect 20680 60664 20686 60716
rect 21266 60664 21272 60716
rect 21324 60664 21330 60716
rect 21358 60664 21364 60716
rect 21416 60704 21422 60716
rect 22557 60707 22615 60713
rect 22557 60704 22569 60707
rect 21416 60676 22569 60704
rect 21416 60664 21422 60676
rect 22557 60673 22569 60676
rect 22603 60673 22615 60707
rect 26510 60704 26516 60716
rect 26471 60676 26516 60704
rect 22557 60667 22615 60673
rect 26510 60664 26516 60676
rect 26568 60664 26574 60716
rect 16071 60608 16528 60636
rect 16071 60605 16083 60608
rect 16025 60599 16083 60605
rect 16574 60596 16580 60648
rect 16632 60636 16638 60648
rect 16669 60639 16727 60645
rect 16669 60636 16681 60639
rect 16632 60608 16681 60636
rect 16632 60596 16638 60608
rect 16669 60605 16681 60608
rect 16715 60605 16727 60639
rect 16669 60599 16727 60605
rect 16945 60639 17003 60645
rect 16945 60605 16957 60639
rect 16991 60605 17003 60639
rect 16945 60599 17003 60605
rect 17865 60639 17923 60645
rect 17865 60605 17877 60639
rect 17911 60636 17923 60639
rect 18230 60636 18236 60648
rect 17911 60608 18236 60636
rect 17911 60605 17923 60608
rect 17865 60599 17923 60605
rect 16206 60528 16212 60580
rect 16264 60568 16270 60580
rect 16960 60568 16988 60599
rect 18230 60596 18236 60608
rect 18288 60596 18294 60648
rect 18598 60636 18604 60648
rect 18559 60608 18604 60636
rect 18598 60596 18604 60608
rect 18656 60596 18662 60648
rect 18874 60636 18880 60648
rect 18835 60608 18880 60636
rect 18874 60596 18880 60608
rect 18932 60596 18938 60648
rect 20533 60639 20591 60645
rect 20533 60605 20545 60639
rect 20579 60636 20591 60639
rect 20714 60636 20720 60648
rect 20579 60608 20720 60636
rect 20579 60605 20591 60608
rect 20533 60599 20591 60605
rect 20714 60596 20720 60608
rect 20772 60636 20778 60648
rect 20901 60639 20959 60645
rect 20901 60636 20913 60639
rect 20772 60608 20913 60636
rect 20772 60596 20778 60608
rect 20901 60605 20913 60608
rect 20947 60605 20959 60639
rect 21284 60636 21312 60664
rect 21542 60636 21548 60648
rect 21284 60608 21548 60636
rect 20901 60599 20959 60605
rect 21542 60596 21548 60608
rect 21600 60596 21606 60648
rect 18616 60568 18644 60596
rect 19334 60568 19340 60580
rect 16264 60540 19340 60568
rect 16264 60528 16270 60540
rect 19334 60528 19340 60540
rect 19392 60528 19398 60580
rect 1104 60410 28888 60432
rect 1104 60358 10982 60410
rect 11034 60358 11046 60410
rect 11098 60358 11110 60410
rect 11162 60358 11174 60410
rect 11226 60358 20982 60410
rect 21034 60358 21046 60410
rect 21098 60358 21110 60410
rect 21162 60358 21174 60410
rect 21226 60358 28888 60410
rect 1104 60336 28888 60358
rect 15654 60256 15660 60308
rect 15712 60296 15718 60308
rect 16206 60296 16212 60308
rect 15712 60268 16212 60296
rect 15712 60256 15718 60268
rect 16206 60256 16212 60268
rect 16264 60256 16270 60308
rect 17678 60296 17684 60308
rect 16868 60268 17684 60296
rect 16868 60240 16896 60268
rect 17678 60256 17684 60268
rect 17736 60256 17742 60308
rect 18233 60299 18291 60305
rect 18233 60265 18245 60299
rect 18279 60296 18291 60299
rect 18874 60296 18880 60308
rect 18279 60268 18880 60296
rect 18279 60265 18291 60268
rect 18233 60259 18291 60265
rect 18874 60256 18880 60268
rect 18932 60256 18938 60308
rect 19426 60256 19432 60308
rect 19484 60256 19490 60308
rect 16850 60228 16856 60240
rect 16763 60200 16856 60228
rect 16850 60188 16856 60200
rect 16908 60188 16914 60240
rect 18785 60231 18843 60237
rect 18785 60197 18797 60231
rect 18831 60228 18843 60231
rect 19444 60228 19472 60256
rect 18831 60200 19748 60228
rect 18831 60197 18843 60200
rect 18785 60191 18843 60197
rect 17034 60120 17040 60172
rect 17092 60160 17098 60172
rect 17218 60160 17224 60172
rect 17092 60132 17224 60160
rect 17092 60120 17098 60132
rect 17218 60120 17224 60132
rect 17276 60160 17282 60172
rect 17681 60163 17739 60169
rect 17681 60160 17693 60163
rect 17276 60132 17693 60160
rect 17276 60120 17282 60132
rect 17681 60129 17693 60132
rect 17727 60129 17739 60163
rect 17681 60123 17739 60129
rect 19429 60163 19487 60169
rect 19429 60129 19441 60163
rect 19475 60160 19487 60163
rect 19518 60160 19524 60172
rect 19475 60132 19524 60160
rect 19475 60129 19487 60132
rect 19429 60123 19487 60129
rect 19518 60120 19524 60132
rect 19576 60120 19582 60172
rect 19720 60169 19748 60200
rect 20732 60200 21772 60228
rect 19705 60163 19763 60169
rect 19705 60129 19717 60163
rect 19751 60129 19763 60163
rect 19705 60123 19763 60129
rect 19794 60120 19800 60172
rect 19852 60160 19858 60172
rect 20622 60160 20628 60172
rect 19852 60132 20628 60160
rect 19852 60120 19858 60132
rect 20622 60120 20628 60132
rect 20680 60160 20686 60172
rect 20732 60160 20760 60200
rect 20680 60132 20760 60160
rect 21453 60163 21511 60169
rect 20680 60120 20686 60132
rect 21453 60129 21465 60163
rect 21499 60160 21511 60163
rect 21542 60160 21548 60172
rect 21499 60132 21548 60160
rect 21499 60129 21511 60132
rect 21453 60123 21511 60129
rect 21542 60120 21548 60132
rect 21600 60120 21606 60172
rect 21744 60169 21772 60200
rect 21729 60163 21787 60169
rect 21729 60129 21741 60163
rect 21775 60129 21787 60163
rect 21729 60123 21787 60129
rect 22738 60120 22744 60172
rect 22796 60160 22802 60172
rect 22922 60160 22928 60172
rect 22796 60132 22928 60160
rect 22796 60120 22802 60132
rect 22922 60120 22928 60132
rect 22980 60120 22986 60172
rect 17405 60095 17463 60101
rect 17405 60061 17417 60095
rect 17451 60061 17463 60095
rect 17405 60055 17463 60061
rect 17865 60095 17923 60101
rect 17865 60061 17877 60095
rect 17911 60061 17923 60095
rect 17865 60055 17923 60061
rect 17420 60024 17448 60055
rect 17678 60024 17684 60036
rect 17420 59996 17684 60024
rect 17678 59984 17684 59996
rect 17736 59984 17742 60036
rect 1670 59956 1676 59968
rect 1583 59928 1676 59956
rect 1670 59916 1676 59928
rect 1728 59956 1734 59968
rect 2038 59956 2044 59968
rect 1728 59928 2044 59956
rect 1728 59916 1734 59928
rect 2038 59916 2044 59928
rect 2096 59916 2102 59968
rect 15841 59959 15899 59965
rect 15841 59925 15853 59959
rect 15887 59956 15899 59959
rect 16761 59959 16819 59965
rect 16761 59956 16773 59959
rect 15887 59928 16773 59956
rect 15887 59925 15899 59928
rect 15841 59919 15899 59925
rect 16761 59925 16773 59928
rect 16807 59956 16819 59959
rect 17310 59956 17316 59968
rect 16807 59928 17316 59956
rect 16807 59925 16819 59928
rect 16761 59919 16819 59925
rect 17310 59916 17316 59928
rect 17368 59956 17374 59968
rect 17880 59956 17908 60055
rect 18230 60052 18236 60104
rect 18288 60092 18294 60104
rect 18782 60092 18788 60104
rect 18288 60064 18788 60092
rect 18288 60052 18294 60064
rect 18782 60052 18788 60064
rect 18840 60092 18846 60104
rect 18969 60095 19027 60101
rect 18969 60092 18981 60095
rect 18840 60064 18981 60092
rect 18840 60052 18846 60064
rect 18969 60061 18981 60064
rect 19015 60061 19027 60095
rect 18969 60055 19027 60061
rect 21085 60095 21143 60101
rect 21085 60061 21097 60095
rect 21131 60061 21143 60095
rect 21818 60092 21824 60104
rect 21779 60064 21824 60092
rect 21085 60055 21143 60061
rect 19702 60024 19708 60036
rect 19663 59996 19708 60024
rect 19702 59984 19708 59996
rect 19760 59984 19766 60036
rect 21100 60024 21128 60055
rect 21818 60052 21824 60064
rect 21876 60052 21882 60104
rect 22830 60092 22836 60104
rect 22791 60064 22836 60092
rect 22830 60052 22836 60064
rect 22888 60052 22894 60104
rect 22186 60024 22192 60036
rect 21100 59996 22192 60024
rect 22186 59984 22192 59996
rect 22244 59984 22250 60036
rect 17368 59928 17908 59956
rect 17368 59916 17374 59928
rect 1104 59866 28888 59888
rect 1104 59814 5982 59866
rect 6034 59814 6046 59866
rect 6098 59814 6110 59866
rect 6162 59814 6174 59866
rect 6226 59814 15982 59866
rect 16034 59814 16046 59866
rect 16098 59814 16110 59866
rect 16162 59814 16174 59866
rect 16226 59814 25982 59866
rect 26034 59814 26046 59866
rect 26098 59814 26110 59866
rect 26162 59814 26174 59866
rect 26226 59814 28888 59866
rect 1104 59792 28888 59814
rect 17494 59712 17500 59764
rect 17552 59752 17558 59764
rect 17773 59755 17831 59761
rect 17773 59752 17785 59755
rect 17552 59724 17785 59752
rect 17552 59712 17558 59724
rect 17773 59721 17785 59724
rect 17819 59752 17831 59755
rect 19058 59752 19064 59764
rect 17819 59724 19064 59752
rect 17819 59721 17831 59724
rect 17773 59715 17831 59721
rect 19058 59712 19064 59724
rect 19116 59712 19122 59764
rect 15289 59687 15347 59693
rect 15289 59653 15301 59687
rect 15335 59684 15347 59687
rect 17678 59684 17684 59696
rect 15335 59656 17684 59684
rect 15335 59653 15347 59656
rect 15289 59647 15347 59653
rect 17678 59644 17684 59656
rect 17736 59644 17742 59696
rect 22830 59684 22836 59696
rect 20916 59656 22836 59684
rect 17497 59619 17555 59625
rect 17497 59585 17509 59619
rect 17543 59616 17555 59619
rect 18874 59616 18880 59628
rect 17543 59588 18880 59616
rect 17543 59585 17555 59588
rect 17497 59579 17555 59585
rect 18874 59576 18880 59588
rect 18932 59616 18938 59628
rect 20916 59625 20944 59656
rect 22830 59644 22836 59656
rect 22888 59644 22894 59696
rect 20257 59619 20315 59625
rect 18932 59588 19564 59616
rect 18932 59576 18938 59588
rect 14921 59551 14979 59557
rect 14921 59517 14933 59551
rect 14967 59548 14979 59551
rect 16206 59548 16212 59560
rect 14967 59520 16212 59548
rect 14967 59517 14979 59520
rect 14921 59511 14979 59517
rect 16206 59508 16212 59520
rect 16264 59548 16270 59560
rect 16301 59551 16359 59557
rect 16301 59548 16313 59551
rect 16264 59520 16313 59548
rect 16264 59508 16270 59520
rect 16301 59517 16313 59520
rect 16347 59517 16359 59551
rect 16301 59511 16359 59517
rect 16577 59551 16635 59557
rect 16577 59517 16589 59551
rect 16623 59517 16635 59551
rect 16577 59511 16635 59517
rect 16761 59551 16819 59557
rect 16761 59517 16773 59551
rect 16807 59548 16819 59551
rect 17310 59548 17316 59560
rect 16807 59520 17316 59548
rect 16807 59517 16819 59520
rect 16761 59511 16819 59517
rect 15746 59480 15752 59492
rect 15707 59452 15752 59480
rect 15746 59440 15752 59452
rect 15804 59440 15810 59492
rect 14550 59372 14556 59424
rect 14608 59412 14614 59424
rect 15562 59412 15568 59424
rect 14608 59384 15568 59412
rect 14608 59372 14614 59384
rect 15562 59372 15568 59384
rect 15620 59412 15626 59424
rect 16592 59412 16620 59511
rect 17310 59508 17316 59520
rect 17368 59508 17374 59560
rect 18601 59551 18659 59557
rect 18601 59517 18613 59551
rect 18647 59548 18659 59551
rect 18782 59548 18788 59560
rect 18647 59520 18788 59548
rect 18647 59517 18659 59520
rect 18601 59511 18659 59517
rect 18782 59508 18788 59520
rect 18840 59508 18846 59560
rect 19058 59548 19064 59560
rect 19019 59520 19064 59548
rect 19058 59508 19064 59520
rect 19116 59508 19122 59560
rect 19536 59557 19564 59588
rect 20257 59585 20269 59619
rect 20303 59616 20315 59619
rect 20901 59619 20959 59625
rect 20901 59616 20913 59619
rect 20303 59588 20913 59616
rect 20303 59585 20315 59588
rect 20257 59579 20315 59585
rect 20901 59585 20913 59588
rect 20947 59585 20959 59619
rect 20901 59579 20959 59585
rect 21821 59619 21879 59625
rect 21821 59585 21833 59619
rect 21867 59616 21879 59619
rect 21910 59616 21916 59628
rect 21867 59588 21916 59616
rect 21867 59585 21879 59588
rect 21821 59579 21879 59585
rect 21910 59576 21916 59588
rect 21968 59576 21974 59628
rect 19521 59551 19579 59557
rect 19521 59517 19533 59551
rect 19567 59517 19579 59551
rect 19521 59511 19579 59517
rect 20625 59551 20683 59557
rect 20625 59517 20637 59551
rect 20671 59548 20683 59551
rect 21266 59548 21272 59560
rect 20671 59520 21272 59548
rect 20671 59517 20683 59520
rect 20625 59511 20683 59517
rect 21266 59508 21272 59520
rect 21324 59508 21330 59560
rect 21358 59508 21364 59560
rect 21416 59548 21422 59560
rect 21545 59551 21603 59557
rect 21545 59548 21557 59551
rect 21416 59520 21557 59548
rect 21416 59508 21422 59520
rect 21545 59517 21557 59520
rect 21591 59517 21603 59551
rect 21545 59511 21603 59517
rect 21634 59508 21640 59560
rect 21692 59548 21698 59560
rect 22465 59551 22523 59557
rect 22465 59548 22477 59551
rect 21692 59520 22477 59548
rect 21692 59508 21698 59520
rect 22465 59517 22477 59520
rect 22511 59517 22523 59551
rect 22465 59511 22523 59517
rect 19794 59480 19800 59492
rect 19755 59452 19800 59480
rect 19794 59440 19800 59452
rect 19852 59440 19858 59492
rect 17034 59412 17040 59424
rect 15620 59384 16620 59412
rect 16995 59384 17040 59412
rect 15620 59372 15626 59384
rect 17034 59372 17040 59384
rect 17092 59372 17098 59424
rect 22186 59412 22192 59424
rect 22147 59384 22192 59412
rect 22186 59372 22192 59384
rect 22244 59372 22250 59424
rect 22738 59372 22744 59424
rect 22796 59412 22802 59424
rect 22833 59415 22891 59421
rect 22833 59412 22845 59415
rect 22796 59384 22845 59412
rect 22796 59372 22802 59384
rect 22833 59381 22845 59384
rect 22879 59381 22891 59415
rect 22833 59375 22891 59381
rect 1104 59322 28888 59344
rect 1104 59270 10982 59322
rect 11034 59270 11046 59322
rect 11098 59270 11110 59322
rect 11162 59270 11174 59322
rect 11226 59270 20982 59322
rect 21034 59270 21046 59322
rect 21098 59270 21110 59322
rect 21162 59270 21174 59322
rect 21226 59270 28888 59322
rect 1104 59248 28888 59270
rect 19334 59168 19340 59220
rect 19392 59208 19398 59220
rect 19797 59211 19855 59217
rect 19797 59208 19809 59211
rect 19392 59180 19809 59208
rect 19392 59168 19398 59180
rect 19797 59177 19809 59180
rect 19843 59177 19855 59211
rect 19797 59171 19855 59177
rect 15749 59143 15807 59149
rect 15749 59109 15761 59143
rect 15795 59140 15807 59143
rect 17586 59140 17592 59152
rect 15795 59112 16804 59140
rect 17547 59112 17592 59140
rect 15795 59109 15807 59112
rect 15749 59103 15807 59109
rect 14734 59032 14740 59084
rect 14792 59072 14798 59084
rect 15105 59075 15163 59081
rect 15105 59072 15117 59075
rect 14792 59044 15117 59072
rect 14792 59032 14798 59044
rect 15105 59041 15117 59044
rect 15151 59072 15163 59075
rect 15654 59072 15660 59084
rect 15151 59044 15660 59072
rect 15151 59041 15163 59044
rect 15105 59035 15163 59041
rect 15654 59032 15660 59044
rect 15712 59072 15718 59084
rect 16776 59081 16804 59112
rect 17586 59100 17592 59112
rect 17644 59140 17650 59152
rect 21177 59143 21235 59149
rect 17644 59112 18644 59140
rect 17644 59100 17650 59112
rect 16209 59075 16267 59081
rect 16209 59072 16221 59075
rect 15712 59044 16221 59072
rect 15712 59032 15718 59044
rect 16209 59041 16221 59044
rect 16255 59041 16267 59075
rect 16209 59035 16267 59041
rect 16761 59075 16819 59081
rect 16761 59041 16773 59075
rect 16807 59072 16819 59075
rect 16850 59072 16856 59084
rect 16807 59044 16856 59072
rect 16807 59041 16819 59044
rect 16761 59035 16819 59041
rect 16850 59032 16856 59044
rect 16908 59032 16914 59084
rect 17678 59032 17684 59084
rect 17736 59072 17742 59084
rect 18616 59081 18644 59112
rect 21177 59109 21189 59143
rect 21223 59140 21235 59143
rect 21358 59140 21364 59152
rect 21223 59112 21364 59140
rect 21223 59109 21235 59112
rect 21177 59103 21235 59109
rect 21358 59100 21364 59112
rect 21416 59140 21422 59152
rect 21453 59143 21511 59149
rect 21453 59140 21465 59143
rect 21416 59112 21465 59140
rect 21416 59100 21422 59112
rect 21453 59109 21465 59112
rect 21499 59109 21511 59143
rect 21453 59103 21511 59109
rect 18601 59075 18659 59081
rect 17736 59044 18184 59072
rect 17736 59032 17742 59044
rect 18156 59016 18184 59044
rect 18601 59041 18613 59075
rect 18647 59041 18659 59075
rect 19610 59072 19616 59084
rect 19571 59044 19616 59072
rect 18601 59035 18659 59041
rect 19610 59032 19616 59044
rect 19668 59072 19674 59084
rect 20073 59075 20131 59081
rect 20073 59072 20085 59075
rect 19668 59044 20085 59072
rect 19668 59032 19674 59044
rect 20073 59041 20085 59044
rect 20119 59041 20131 59075
rect 20073 59035 20131 59041
rect 21818 59032 21824 59084
rect 21876 59072 21882 59084
rect 22281 59075 22339 59081
rect 22281 59072 22293 59075
rect 21876 59044 22293 59072
rect 21876 59032 21882 59044
rect 22281 59041 22293 59044
rect 22327 59041 22339 59075
rect 22281 59035 22339 59041
rect 22465 59075 22523 59081
rect 22465 59041 22477 59075
rect 22511 59072 22523 59075
rect 22830 59072 22836 59084
rect 22511 59044 22836 59072
rect 22511 59041 22523 59044
rect 22465 59035 22523 59041
rect 22830 59032 22836 59044
rect 22888 59032 22894 59084
rect 23474 59072 23480 59084
rect 23435 59044 23480 59072
rect 23474 59032 23480 59044
rect 23532 59032 23538 59084
rect 15562 58964 15568 59016
rect 15620 59004 15626 59016
rect 15933 59007 15991 59013
rect 15933 59004 15945 59007
rect 15620 58976 15945 59004
rect 15620 58964 15626 58976
rect 15933 58973 15945 58976
rect 15979 58973 15991 59007
rect 15933 58967 15991 58973
rect 17773 59007 17831 59013
rect 17773 58973 17785 59007
rect 17819 59004 17831 59007
rect 17954 59004 17960 59016
rect 17819 58976 17960 59004
rect 17819 58973 17831 58976
rect 17773 58967 17831 58973
rect 17954 58964 17960 58976
rect 18012 58964 18018 59016
rect 18138 58964 18144 59016
rect 18196 59004 18202 59016
rect 18325 59007 18383 59013
rect 18325 59004 18337 59007
rect 18196 58976 18337 59004
rect 18196 58964 18202 58976
rect 18325 58973 18337 58976
rect 18371 58973 18383 59007
rect 18325 58967 18383 58973
rect 18785 59007 18843 59013
rect 18785 58973 18797 59007
rect 18831 59004 18843 59007
rect 18966 59004 18972 59016
rect 18831 58976 18972 59004
rect 18831 58973 18843 58976
rect 18785 58967 18843 58973
rect 16666 58936 16672 58948
rect 16627 58908 16672 58936
rect 16666 58896 16672 58908
rect 16724 58896 16730 58948
rect 17310 58936 17316 58948
rect 17223 58908 17316 58936
rect 17310 58896 17316 58908
rect 17368 58936 17374 58948
rect 18800 58936 18828 58967
rect 18966 58964 18972 58976
rect 19024 58964 19030 59016
rect 22005 59007 22063 59013
rect 22005 58973 22017 59007
rect 22051 59004 22063 59007
rect 22094 59004 22100 59016
rect 22051 58976 22100 59004
rect 22051 58973 22063 58976
rect 22005 58967 22063 58973
rect 22094 58964 22100 58976
rect 22152 58964 22158 59016
rect 23290 59004 23296 59016
rect 23251 58976 23296 59004
rect 23290 58964 23296 58976
rect 23348 58964 23354 59016
rect 17368 58908 18828 58936
rect 17368 58896 17374 58908
rect 19150 58896 19156 58948
rect 19208 58936 19214 58948
rect 20441 58939 20499 58945
rect 20441 58936 20453 58939
rect 19208 58908 20453 58936
rect 19208 58896 19214 58908
rect 20441 58905 20453 58908
rect 20487 58936 20499 58939
rect 20990 58936 20996 58948
rect 20487 58908 20996 58936
rect 20487 58905 20499 58908
rect 20441 58899 20499 58905
rect 20990 58896 20996 58908
rect 21048 58896 21054 58948
rect 14642 58868 14648 58880
rect 14603 58840 14648 58868
rect 14642 58828 14648 58840
rect 14700 58828 14706 58880
rect 18782 58828 18788 58880
rect 18840 58868 18846 58880
rect 19061 58871 19119 58877
rect 19061 58868 19073 58871
rect 18840 58840 19073 58868
rect 18840 58828 18846 58840
rect 19061 58837 19073 58840
rect 19107 58837 19119 58871
rect 19518 58868 19524 58880
rect 19479 58840 19524 58868
rect 19061 58831 19119 58837
rect 19518 58828 19524 58840
rect 19576 58828 19582 58880
rect 24302 58868 24308 58880
rect 24263 58840 24308 58868
rect 24302 58828 24308 58840
rect 24360 58828 24366 58880
rect 1104 58778 28888 58800
rect 1104 58726 5982 58778
rect 6034 58726 6046 58778
rect 6098 58726 6110 58778
rect 6162 58726 6174 58778
rect 6226 58726 15982 58778
rect 16034 58726 16046 58778
rect 16098 58726 16110 58778
rect 16162 58726 16174 58778
rect 16226 58726 25982 58778
rect 26034 58726 26046 58778
rect 26098 58726 26110 58778
rect 26162 58726 26174 58778
rect 26226 58726 28888 58778
rect 1104 58704 28888 58726
rect 2866 58624 2872 58676
rect 2924 58664 2930 58676
rect 2961 58667 3019 58673
rect 2961 58664 2973 58667
rect 2924 58636 2973 58664
rect 2924 58624 2930 58636
rect 2961 58633 2973 58636
rect 3007 58633 3019 58667
rect 14458 58664 14464 58676
rect 14419 58636 14464 58664
rect 2961 58627 3019 58633
rect 2976 58528 3004 58627
rect 14458 58624 14464 58636
rect 14516 58624 14522 58676
rect 15562 58624 15568 58676
rect 15620 58664 15626 58676
rect 16669 58667 16727 58673
rect 16669 58664 16681 58667
rect 15620 58636 16681 58664
rect 15620 58624 15626 58636
rect 16669 58633 16681 58636
rect 16715 58633 16727 58667
rect 16669 58627 16727 58633
rect 19058 58624 19064 58676
rect 19116 58664 19122 58676
rect 20257 58667 20315 58673
rect 20257 58664 20269 58667
rect 19116 58636 20269 58664
rect 19116 58624 19122 58636
rect 20257 58633 20269 58636
rect 20303 58633 20315 58667
rect 21818 58664 21824 58676
rect 21779 58636 21824 58664
rect 20257 58627 20315 58633
rect 3421 58531 3479 58537
rect 3421 58528 3433 58531
rect 2976 58500 3433 58528
rect 3421 58497 3433 58500
rect 3467 58497 3479 58531
rect 3421 58491 3479 58497
rect 16393 58531 16451 58537
rect 16393 58497 16405 58531
rect 16439 58528 16451 58531
rect 16482 58528 16488 58540
rect 16439 58500 16488 58528
rect 16439 58497 16451 58500
rect 16393 58491 16451 58497
rect 16482 58488 16488 58500
rect 16540 58488 16546 58540
rect 18601 58531 18659 58537
rect 18601 58497 18613 58531
rect 18647 58528 18659 58531
rect 18874 58528 18880 58540
rect 18647 58500 18880 58528
rect 18647 58497 18659 58500
rect 18601 58491 18659 58497
rect 18874 58488 18880 58500
rect 18932 58488 18938 58540
rect 18966 58488 18972 58540
rect 19024 58528 19030 58540
rect 19153 58531 19211 58537
rect 19153 58528 19165 58531
rect 19024 58500 19165 58528
rect 19024 58488 19030 58500
rect 19153 58497 19165 58500
rect 19199 58528 19211 58531
rect 19889 58531 19947 58537
rect 19889 58528 19901 58531
rect 19199 58500 19901 58528
rect 19199 58497 19211 58500
rect 19153 58491 19211 58497
rect 19889 58497 19901 58500
rect 19935 58497 19947 58531
rect 20272 58528 20300 58627
rect 21818 58624 21824 58636
rect 21876 58624 21882 58676
rect 22189 58667 22247 58673
rect 22189 58633 22201 58667
rect 22235 58664 22247 58667
rect 22830 58664 22836 58676
rect 22235 58636 22836 58664
rect 22235 58633 22247 58636
rect 22189 58627 22247 58633
rect 22830 58624 22836 58636
rect 22888 58624 22894 58676
rect 23109 58667 23167 58673
rect 23109 58633 23121 58667
rect 23155 58664 23167 58667
rect 23290 58664 23296 58676
rect 23155 58636 23296 58664
rect 23155 58633 23167 58636
rect 23109 58627 23167 58633
rect 23290 58624 23296 58636
rect 23348 58664 23354 58676
rect 23750 58664 23756 58676
rect 23348 58636 23756 58664
rect 23348 58624 23354 58636
rect 23750 58624 23756 58636
rect 23808 58664 23814 58676
rect 23808 58636 24716 58664
rect 23808 58624 23814 58636
rect 22465 58599 22523 58605
rect 22465 58596 22477 58599
rect 21284 58568 22477 58596
rect 21284 58528 21312 58568
rect 22465 58565 22477 58568
rect 22511 58565 22523 58599
rect 22465 58559 22523 58565
rect 23658 58528 23664 58540
rect 20272 58500 21312 58528
rect 23571 58500 23664 58528
rect 19889 58491 19947 58497
rect 3142 58460 3148 58472
rect 3103 58432 3148 58460
rect 3142 58420 3148 58432
rect 3200 58420 3206 58472
rect 14277 58463 14335 58469
rect 14277 58429 14289 58463
rect 14323 58460 14335 58463
rect 15289 58463 15347 58469
rect 14323 58432 14872 58460
rect 14323 58429 14335 58432
rect 14277 58423 14335 58429
rect 4801 58395 4859 58401
rect 4801 58361 4813 58395
rect 4847 58392 4859 58395
rect 5442 58392 5448 58404
rect 4847 58364 5448 58392
rect 4847 58361 4859 58364
rect 4801 58355 4859 58361
rect 5442 58352 5448 58364
rect 5500 58352 5506 58404
rect 14185 58395 14243 58401
rect 14185 58361 14197 58395
rect 14231 58392 14243 58395
rect 14734 58392 14740 58404
rect 14231 58364 14740 58392
rect 14231 58361 14243 58364
rect 14185 58355 14243 58361
rect 14734 58352 14740 58364
rect 14792 58352 14798 58404
rect 14844 58336 14872 58432
rect 15289 58429 15301 58463
rect 15335 58429 15347 58463
rect 15654 58460 15660 58472
rect 15615 58432 15660 58460
rect 15289 58423 15347 58429
rect 14826 58324 14832 58336
rect 14787 58296 14832 58324
rect 14826 58284 14832 58296
rect 14884 58284 14890 58336
rect 15197 58327 15255 58333
rect 15197 58293 15209 58327
rect 15243 58324 15255 58327
rect 15304 58324 15332 58423
rect 15654 58420 15660 58432
rect 15712 58420 15718 58472
rect 16206 58460 16212 58472
rect 16167 58432 16212 58460
rect 16206 58420 16212 58432
rect 16264 58420 16270 58472
rect 19429 58463 19487 58469
rect 19429 58429 19441 58463
rect 19475 58429 19487 58463
rect 19610 58460 19616 58472
rect 19523 58432 19616 58460
rect 19429 58423 19487 58429
rect 16224 58392 16252 58420
rect 16482 58392 16488 58404
rect 16224 58364 16488 58392
rect 16482 58352 16488 58364
rect 16540 58352 16546 58404
rect 17126 58352 17132 58404
rect 17184 58392 17190 58404
rect 17184 58364 17356 58392
rect 17184 58352 17190 58364
rect 15562 58324 15568 58336
rect 15243 58296 15568 58324
rect 15243 58293 15255 58296
rect 15197 58287 15255 58293
rect 15562 58284 15568 58296
rect 15620 58284 15626 58336
rect 17218 58324 17224 58336
rect 17179 58296 17224 58324
rect 17218 58284 17224 58296
rect 17276 58284 17282 58336
rect 17328 58324 17356 58364
rect 17678 58352 17684 58404
rect 17736 58392 17742 58404
rect 18417 58395 18475 58401
rect 18417 58392 18429 58395
rect 17736 58364 18429 58392
rect 17736 58352 17742 58364
rect 18417 58361 18429 58364
rect 18463 58392 18475 58395
rect 19444 58392 19472 58423
rect 19610 58420 19616 58432
rect 19668 58460 19674 58472
rect 20070 58460 20076 58472
rect 19668 58432 20076 58460
rect 19668 58420 19674 58432
rect 20070 58420 20076 58432
rect 20128 58460 20134 58472
rect 20990 58460 20996 58472
rect 20128 58432 20852 58460
rect 20951 58432 20996 58460
rect 20128 58420 20134 58432
rect 19518 58392 19524 58404
rect 18463 58364 19524 58392
rect 18463 58361 18475 58364
rect 18417 58355 18475 58361
rect 19518 58352 19524 58364
rect 19576 58352 19582 58404
rect 17865 58327 17923 58333
rect 17865 58324 17877 58327
rect 17328 58296 17877 58324
rect 17865 58293 17877 58296
rect 17911 58324 17923 58327
rect 19628 58324 19656 58420
rect 19702 58352 19708 58404
rect 19760 58392 19766 58404
rect 20441 58395 20499 58401
rect 20441 58392 20453 58395
rect 19760 58364 20453 58392
rect 19760 58352 19766 58364
rect 20441 58361 20453 58364
rect 20487 58361 20499 58395
rect 20824 58392 20852 58432
rect 20990 58420 20996 58432
rect 21048 58420 21054 58472
rect 21284 58469 21312 58500
rect 23658 58488 23664 58500
rect 23716 58528 23722 58540
rect 24578 58528 24584 58540
rect 23716 58500 24584 58528
rect 23716 58488 23722 58500
rect 24578 58488 24584 58500
rect 24636 58488 24642 58540
rect 24688 58537 24716 58636
rect 24673 58531 24731 58537
rect 24673 58497 24685 58531
rect 24719 58497 24731 58531
rect 24673 58491 24731 58497
rect 21269 58463 21327 58469
rect 21269 58429 21281 58463
rect 21315 58429 21327 58463
rect 21269 58423 21327 58429
rect 21453 58463 21511 58469
rect 21453 58429 21465 58463
rect 21499 58429 21511 58463
rect 21453 58423 21511 58429
rect 22281 58463 22339 58469
rect 22281 58429 22293 58463
rect 22327 58460 22339 58463
rect 22554 58460 22560 58472
rect 22327 58432 22560 58460
rect 22327 58429 22339 58432
rect 22281 58423 22339 58429
rect 21468 58392 21496 58423
rect 22554 58420 22560 58432
rect 22612 58420 22618 58472
rect 23290 58420 23296 58472
rect 23348 58460 23354 58472
rect 24213 58463 24271 58469
rect 24213 58460 24225 58463
rect 23348 58432 24225 58460
rect 23348 58420 23354 58432
rect 24213 58429 24225 58432
rect 24259 58460 24271 58463
rect 24302 58460 24308 58472
rect 24259 58432 24308 58460
rect 24259 58429 24271 58432
rect 24213 58423 24271 58429
rect 24302 58420 24308 58432
rect 24360 58420 24366 58472
rect 24489 58463 24547 58469
rect 24489 58429 24501 58463
rect 24535 58460 24547 58463
rect 24535 58432 24624 58460
rect 24535 58429 24547 58432
rect 24489 58423 24547 58429
rect 20824 58364 21496 58392
rect 20441 58355 20499 58361
rect 17911 58296 19656 58324
rect 17911 58293 17923 58296
rect 17865 58287 17923 58293
rect 21818 58284 21824 58336
rect 21876 58324 21882 58336
rect 23385 58327 23443 58333
rect 23385 58324 23397 58327
rect 21876 58296 23397 58324
rect 21876 58284 21882 58296
rect 23385 58293 23397 58296
rect 23431 58324 23443 58327
rect 23566 58324 23572 58336
rect 23431 58296 23572 58324
rect 23431 58293 23443 58296
rect 23385 58287 23443 58293
rect 23566 58284 23572 58296
rect 23624 58324 23630 58336
rect 24596 58324 24624 58432
rect 23624 58296 24624 58324
rect 23624 58284 23630 58296
rect 1104 58234 28888 58256
rect 1104 58182 10982 58234
rect 11034 58182 11046 58234
rect 11098 58182 11110 58234
rect 11162 58182 11174 58234
rect 11226 58182 20982 58234
rect 21034 58182 21046 58234
rect 21098 58182 21110 58234
rect 21162 58182 21174 58234
rect 21226 58182 28888 58234
rect 1104 58160 28888 58182
rect 11698 58080 11704 58132
rect 11756 58120 11762 58132
rect 11974 58120 11980 58132
rect 11756 58092 11980 58120
rect 11756 58080 11762 58092
rect 11974 58080 11980 58092
rect 12032 58080 12038 58132
rect 14366 58120 14372 58132
rect 14327 58092 14372 58120
rect 14366 58080 14372 58092
rect 14424 58080 14430 58132
rect 15746 58080 15752 58132
rect 15804 58120 15810 58132
rect 15804 58092 16160 58120
rect 15804 58080 15810 58092
rect 15654 58012 15660 58064
rect 15712 58052 15718 58064
rect 15712 58024 15792 58052
rect 15712 58012 15718 58024
rect 12066 57944 12072 57996
rect 12124 57984 12130 57996
rect 12161 57987 12219 57993
rect 12161 57984 12173 57987
rect 12124 57956 12173 57984
rect 12124 57944 12130 57956
rect 12161 57953 12173 57956
rect 12207 57953 12219 57987
rect 14185 57987 14243 57993
rect 14185 57984 14197 57987
rect 12161 57947 12219 57953
rect 13740 57956 14197 57984
rect 3142 57876 3148 57928
rect 3200 57916 3206 57928
rect 3237 57919 3295 57925
rect 3237 57916 3249 57919
rect 3200 57888 3249 57916
rect 3200 57876 3206 57888
rect 3237 57885 3249 57888
rect 3283 57916 3295 57919
rect 3326 57916 3332 57928
rect 3283 57888 3332 57916
rect 3283 57885 3295 57888
rect 3237 57879 3295 57885
rect 3326 57876 3332 57888
rect 3384 57876 3390 57928
rect 13446 57876 13452 57928
rect 13504 57916 13510 57928
rect 13740 57916 13768 57956
rect 14185 57953 14197 57956
rect 14231 57984 14243 57987
rect 15102 57984 15108 57996
rect 14231 57956 15108 57984
rect 14231 57953 14243 57956
rect 14185 57947 14243 57953
rect 15102 57944 15108 57956
rect 15160 57944 15166 57996
rect 15764 57993 15792 58024
rect 16132 57993 16160 58092
rect 20714 58080 20720 58132
rect 20772 58120 20778 58132
rect 20772 58092 21036 58120
rect 20772 58080 20778 58092
rect 21008 58064 21036 58092
rect 23106 58080 23112 58132
rect 23164 58120 23170 58132
rect 23385 58123 23443 58129
rect 23385 58120 23397 58123
rect 23164 58092 23397 58120
rect 23164 58080 23170 58092
rect 23385 58089 23397 58092
rect 23431 58120 23443 58123
rect 23474 58120 23480 58132
rect 23431 58092 23480 58120
rect 23431 58089 23443 58092
rect 23385 58083 23443 58089
rect 23474 58080 23480 58092
rect 23532 58080 23538 58132
rect 17034 58012 17040 58064
rect 17092 58052 17098 58064
rect 17586 58052 17592 58064
rect 17092 58024 17592 58052
rect 17092 58012 17098 58024
rect 17586 58012 17592 58024
rect 17644 58012 17650 58064
rect 20622 58012 20628 58064
rect 20680 58052 20686 58064
rect 20901 58055 20959 58061
rect 20901 58052 20913 58055
rect 20680 58024 20913 58052
rect 20680 58012 20686 58024
rect 20901 58021 20913 58024
rect 20947 58021 20959 58055
rect 20901 58015 20959 58021
rect 20990 58012 20996 58064
rect 21048 58012 21054 58064
rect 15749 57987 15807 57993
rect 15749 57953 15761 57987
rect 15795 57953 15807 57987
rect 15749 57947 15807 57953
rect 16117 57987 16175 57993
rect 16117 57953 16129 57987
rect 16163 57953 16175 57987
rect 16117 57947 16175 57953
rect 16850 57944 16856 57996
rect 16908 57984 16914 57996
rect 17221 57987 17279 57993
rect 17221 57984 17233 57987
rect 16908 57956 17233 57984
rect 16908 57944 16914 57956
rect 17221 57953 17233 57956
rect 17267 57953 17279 57987
rect 18138 57984 18144 57996
rect 17221 57947 17279 57953
rect 17512 57956 18144 57984
rect 13504 57888 13768 57916
rect 13504 57876 13510 57888
rect 14366 57876 14372 57928
rect 14424 57916 14430 57928
rect 15378 57916 15384 57928
rect 14424 57888 15384 57916
rect 14424 57876 14430 57888
rect 15378 57876 15384 57888
rect 15436 57876 15442 57928
rect 16761 57919 16819 57925
rect 16761 57885 16773 57919
rect 16807 57916 16819 57919
rect 17512 57916 17540 57956
rect 18138 57944 18144 57956
rect 18196 57944 18202 57996
rect 19334 57944 19340 57996
rect 19392 57984 19398 57996
rect 19702 57984 19708 57996
rect 19392 57956 19437 57984
rect 19663 57956 19708 57984
rect 19392 57944 19398 57956
rect 19702 57944 19708 57956
rect 19760 57944 19766 57996
rect 21729 57987 21787 57993
rect 21729 57984 21741 57987
rect 20732 57956 21741 57984
rect 20732 57928 20760 57956
rect 21729 57953 21741 57956
rect 21775 57953 21787 57987
rect 23750 57984 23756 57996
rect 23711 57956 23756 57984
rect 21729 57947 21787 57953
rect 23750 57944 23756 57956
rect 23808 57944 23814 57996
rect 23934 57984 23940 57996
rect 23895 57956 23940 57984
rect 23934 57944 23940 57956
rect 23992 57944 23998 57996
rect 24489 57987 24547 57993
rect 24489 57953 24501 57987
rect 24535 57984 24547 57987
rect 24578 57984 24584 57996
rect 24535 57956 24584 57984
rect 24535 57953 24547 57956
rect 24489 57947 24547 57953
rect 24578 57944 24584 57956
rect 24636 57944 24642 57996
rect 16807 57888 17540 57916
rect 16807 57885 16819 57888
rect 16761 57879 16819 57885
rect 17586 57876 17592 57928
rect 17644 57916 17650 57928
rect 17770 57916 17776 57928
rect 17644 57888 17689 57916
rect 17731 57888 17776 57916
rect 17644 57876 17650 57888
rect 17770 57876 17776 57888
rect 17828 57876 17834 57928
rect 18506 57876 18512 57928
rect 18564 57916 18570 57928
rect 18969 57919 19027 57925
rect 18969 57916 18981 57919
rect 18564 57888 18981 57916
rect 18564 57876 18570 57888
rect 18969 57885 18981 57888
rect 19015 57885 19027 57919
rect 18969 57879 19027 57885
rect 20714 57876 20720 57928
rect 20772 57876 20778 57928
rect 21358 57876 21364 57928
rect 21416 57916 21422 57928
rect 21453 57919 21511 57925
rect 21453 57916 21465 57919
rect 21416 57888 21465 57916
rect 21416 57876 21422 57888
rect 21453 57885 21465 57888
rect 21499 57885 21511 57919
rect 21453 57879 21511 57885
rect 21913 57919 21971 57925
rect 21913 57885 21925 57919
rect 21959 57885 21971 57919
rect 21913 57879 21971 57885
rect 2685 57851 2743 57857
rect 2685 57817 2697 57851
rect 2731 57848 2743 57851
rect 3602 57848 3608 57860
rect 2731 57820 3608 57848
rect 2731 57817 2743 57820
rect 2685 57811 2743 57817
rect 3602 57808 3608 57820
rect 3660 57808 3666 57860
rect 13722 57808 13728 57860
rect 13780 57848 13786 57860
rect 14093 57851 14151 57857
rect 14093 57848 14105 57851
rect 13780 57820 14105 57848
rect 13780 57808 13786 57820
rect 14093 57817 14105 57820
rect 14139 57848 14151 57851
rect 15746 57848 15752 57860
rect 14139 57820 15752 57848
rect 14139 57817 14151 57820
rect 14093 57811 14151 57817
rect 15746 57808 15752 57820
rect 15804 57808 15810 57860
rect 16117 57851 16175 57857
rect 16117 57817 16129 57851
rect 16163 57817 16175 57851
rect 16117 57811 16175 57817
rect 17386 57851 17444 57857
rect 17386 57817 17398 57851
rect 17432 57848 17444 57851
rect 17432 57820 17632 57848
rect 17432 57817 17444 57820
rect 17386 57811 17444 57817
rect 13538 57780 13544 57792
rect 13499 57752 13544 57780
rect 13538 57740 13544 57752
rect 13596 57740 13602 57792
rect 14734 57780 14740 57792
rect 14695 57752 14740 57780
rect 14734 57740 14740 57752
rect 14792 57780 14798 57792
rect 15013 57783 15071 57789
rect 15013 57780 15025 57783
rect 14792 57752 15025 57780
rect 14792 57740 14798 57752
rect 15013 57749 15025 57752
rect 15059 57749 15071 57783
rect 15013 57743 15071 57749
rect 15378 57740 15384 57792
rect 15436 57780 15442 57792
rect 16132 57780 16160 57811
rect 17604 57792 17632 57820
rect 19610 57808 19616 57860
rect 19668 57848 19674 57860
rect 19705 57851 19763 57857
rect 19705 57848 19717 57851
rect 19668 57820 19717 57848
rect 19668 57808 19674 57820
rect 19705 57817 19717 57820
rect 19751 57817 19763 57851
rect 19705 57811 19763 57817
rect 20254 57808 20260 57860
rect 20312 57848 20318 57860
rect 21928 57848 21956 57879
rect 22094 57876 22100 57928
rect 22152 57916 22158 57928
rect 22189 57919 22247 57925
rect 22189 57916 22201 57919
rect 22152 57888 22201 57916
rect 22152 57876 22158 57888
rect 22189 57885 22201 57888
rect 22235 57885 22247 57919
rect 22189 57879 22247 57885
rect 22370 57848 22376 57860
rect 20312 57820 22376 57848
rect 20312 57808 20318 57820
rect 22370 57808 22376 57820
rect 22428 57808 22434 57860
rect 24394 57848 24400 57860
rect 24355 57820 24400 57848
rect 24394 57808 24400 57820
rect 24452 57808 24458 57860
rect 17034 57780 17040 57792
rect 15436 57752 16160 57780
rect 16995 57752 17040 57780
rect 15436 57740 15442 57752
rect 17034 57740 17040 57752
rect 17092 57740 17098 57792
rect 17126 57740 17132 57792
rect 17184 57780 17190 57792
rect 17497 57783 17555 57789
rect 17497 57780 17509 57783
rect 17184 57752 17509 57780
rect 17184 57740 17190 57752
rect 17497 57749 17509 57752
rect 17543 57749 17555 57783
rect 17497 57743 17555 57749
rect 17586 57740 17592 57792
rect 17644 57740 17650 57792
rect 18322 57780 18328 57792
rect 18283 57752 18328 57780
rect 18322 57740 18328 57752
rect 18380 57740 18386 57792
rect 18598 57780 18604 57792
rect 18559 57752 18604 57780
rect 18598 57740 18604 57752
rect 18656 57740 18662 57792
rect 20070 57740 20076 57792
rect 20128 57780 20134 57792
rect 20441 57783 20499 57789
rect 20441 57780 20453 57783
rect 20128 57752 20453 57780
rect 20128 57740 20134 57752
rect 20441 57749 20453 57752
rect 20487 57749 20499 57783
rect 22554 57780 22560 57792
rect 22515 57752 22560 57780
rect 20441 57743 20499 57749
rect 22554 57740 22560 57752
rect 22612 57740 22618 57792
rect 23014 57780 23020 57792
rect 22975 57752 23020 57780
rect 23014 57740 23020 57752
rect 23072 57740 23078 57792
rect 1104 57690 28888 57712
rect 1104 57638 5982 57690
rect 6034 57638 6046 57690
rect 6098 57638 6110 57690
rect 6162 57638 6174 57690
rect 6226 57638 15982 57690
rect 16034 57638 16046 57690
rect 16098 57638 16110 57690
rect 16162 57638 16174 57690
rect 16226 57638 25982 57690
rect 26034 57638 26046 57690
rect 26098 57638 26110 57690
rect 26162 57638 26174 57690
rect 26226 57638 28888 57690
rect 1104 57616 28888 57638
rect 5534 57536 5540 57588
rect 5592 57576 5598 57588
rect 6549 57579 6607 57585
rect 6549 57576 6561 57579
rect 5592 57548 6561 57576
rect 5592 57536 5598 57548
rect 6549 57545 6561 57548
rect 6595 57545 6607 57579
rect 13446 57576 13452 57588
rect 13407 57548 13452 57576
rect 6549 57539 6607 57545
rect 2501 57443 2559 57449
rect 2501 57409 2513 57443
rect 2547 57440 2559 57443
rect 2682 57440 2688 57452
rect 2547 57412 2688 57440
rect 2547 57409 2559 57412
rect 2501 57403 2559 57409
rect 2682 57400 2688 57412
rect 2740 57400 2746 57452
rect 2777 57443 2835 57449
rect 2777 57409 2789 57443
rect 2823 57440 2835 57443
rect 2958 57440 2964 57452
rect 2823 57412 2964 57440
rect 2823 57409 2835 57412
rect 2777 57403 2835 57409
rect 2958 57400 2964 57412
rect 3016 57400 3022 57452
rect 6564 57440 6592 57539
rect 13446 57536 13452 57548
rect 13504 57536 13510 57588
rect 17129 57579 17187 57585
rect 17129 57545 17141 57579
rect 17175 57576 17187 57579
rect 17678 57576 17684 57588
rect 17175 57548 17684 57576
rect 17175 57545 17187 57548
rect 17129 57539 17187 57545
rect 17678 57536 17684 57548
rect 17736 57536 17742 57588
rect 18690 57576 18696 57588
rect 18651 57548 18696 57576
rect 18690 57536 18696 57548
rect 18748 57536 18754 57588
rect 19518 57576 19524 57588
rect 19479 57548 19524 57576
rect 19518 57536 19524 57548
rect 19576 57536 19582 57588
rect 20438 57536 20444 57588
rect 20496 57576 20502 57588
rect 20806 57576 20812 57588
rect 20496 57548 20812 57576
rect 20496 57536 20502 57548
rect 20806 57536 20812 57548
rect 20864 57536 20870 57588
rect 22094 57536 22100 57588
rect 22152 57576 22158 57588
rect 22189 57579 22247 57585
rect 22189 57576 22201 57579
rect 22152 57548 22201 57576
rect 22152 57536 22158 57548
rect 22189 57545 22201 57548
rect 22235 57545 22247 57579
rect 22189 57539 22247 57545
rect 22370 57536 22376 57588
rect 22428 57576 22434 57588
rect 22741 57579 22799 57585
rect 22741 57576 22753 57579
rect 22428 57548 22753 57576
rect 22428 57536 22434 57548
rect 22741 57545 22753 57548
rect 22787 57545 22799 57579
rect 22741 57539 22799 57545
rect 23477 57579 23535 57585
rect 23477 57545 23489 57579
rect 23523 57576 23535 57579
rect 23658 57576 23664 57588
rect 23523 57548 23664 57576
rect 23523 57545 23535 57548
rect 23477 57539 23535 57545
rect 23658 57536 23664 57548
rect 23716 57536 23722 57588
rect 23750 57536 23756 57588
rect 23808 57576 23814 57588
rect 24213 57579 24271 57585
rect 24213 57576 24225 57579
rect 23808 57548 24225 57576
rect 23808 57536 23814 57548
rect 24213 57545 24225 57548
rect 24259 57545 24271 57579
rect 24213 57539 24271 57545
rect 18322 57508 18328 57520
rect 18283 57480 18328 57508
rect 18322 57468 18328 57480
rect 18380 57468 18386 57520
rect 7285 57443 7343 57449
rect 7285 57440 7297 57443
rect 6564 57412 7297 57440
rect 7285 57409 7297 57412
rect 7331 57409 7343 57443
rect 7285 57403 7343 57409
rect 13446 57400 13452 57452
rect 13504 57440 13510 57452
rect 14001 57443 14059 57449
rect 14001 57440 14013 57443
rect 13504 57412 14013 57440
rect 13504 57400 13510 57412
rect 14001 57409 14013 57412
rect 14047 57440 14059 57443
rect 14642 57440 14648 57452
rect 14047 57412 14648 57440
rect 14047 57409 14059 57412
rect 14001 57403 14059 57409
rect 14642 57400 14648 57412
rect 14700 57400 14706 57452
rect 17034 57400 17040 57452
rect 17092 57440 17098 57452
rect 18417 57443 18475 57449
rect 18417 57440 18429 57443
rect 17092 57412 18429 57440
rect 17092 57400 17098 57412
rect 18417 57409 18429 57412
rect 18463 57440 18475 57443
rect 18598 57440 18604 57452
rect 18463 57412 18604 57440
rect 18463 57409 18475 57412
rect 18417 57403 18475 57409
rect 18598 57400 18604 57412
rect 18656 57400 18662 57452
rect 19536 57440 19564 57536
rect 21634 57508 21640 57520
rect 20456 57480 21640 57508
rect 19797 57443 19855 57449
rect 19797 57440 19809 57443
rect 19536 57412 19809 57440
rect 19797 57409 19809 57412
rect 19843 57409 19855 57443
rect 19797 57403 19855 57409
rect 3501 57375 3559 57381
rect 3501 57341 3513 57375
rect 3547 57341 3559 57375
rect 3501 57335 3559 57341
rect 3528 57304 3556 57335
rect 3602 57332 3608 57384
rect 3660 57372 3666 57384
rect 7006 57372 7012 57384
rect 3660 57344 3705 57372
rect 6967 57344 7012 57372
rect 3660 57332 3666 57344
rect 7006 57332 7012 57344
rect 7064 57332 7070 57384
rect 13538 57372 13544 57384
rect 13499 57344 13544 57372
rect 13538 57332 13544 57344
rect 13596 57332 13602 57384
rect 14734 57372 14740 57384
rect 14016 57344 14740 57372
rect 2148 57276 3556 57304
rect 8665 57307 8723 57313
rect 2148 57248 2176 57276
rect 8665 57273 8677 57307
rect 8711 57304 8723 57307
rect 9674 57304 9680 57316
rect 8711 57276 9680 57304
rect 8711 57273 8723 57276
rect 8665 57267 8723 57273
rect 9674 57264 9680 57276
rect 9732 57264 9738 57316
rect 14016 57248 14044 57344
rect 14734 57332 14740 57344
rect 14792 57372 14798 57384
rect 14921 57375 14979 57381
rect 14921 57372 14933 57375
rect 14792 57344 14933 57372
rect 14792 57332 14798 57344
rect 14921 57341 14933 57344
rect 14967 57341 14979 57375
rect 14921 57335 14979 57341
rect 15473 57375 15531 57381
rect 15473 57341 15485 57375
rect 15519 57372 15531 57375
rect 15746 57372 15752 57384
rect 15519 57344 15752 57372
rect 15519 57341 15531 57344
rect 15473 57335 15531 57341
rect 15746 57332 15752 57344
rect 15804 57332 15810 57384
rect 16942 57372 16948 57384
rect 16903 57344 16948 57372
rect 16942 57332 16948 57344
rect 17000 57332 17006 57384
rect 18196 57375 18254 57381
rect 18196 57372 18208 57375
rect 17788 57344 18208 57372
rect 15654 57304 15660 57316
rect 15615 57276 15660 57304
rect 15654 57264 15660 57276
rect 15712 57264 15718 57316
rect 17034 57304 17040 57316
rect 16224 57276 17040 57304
rect 16224 57248 16252 57276
rect 17034 57264 17040 57276
rect 17092 57264 17098 57316
rect 2130 57236 2136 57248
rect 2091 57208 2136 57236
rect 2130 57196 2136 57208
rect 2188 57196 2194 57248
rect 12066 57236 12072 57248
rect 12027 57208 12072 57236
rect 12066 57196 12072 57208
rect 12124 57196 12130 57248
rect 13725 57239 13783 57245
rect 13725 57205 13737 57239
rect 13771 57236 13783 57239
rect 13998 57236 14004 57248
rect 13771 57208 14004 57236
rect 13771 57205 13783 57208
rect 13725 57199 13783 57205
rect 13998 57196 14004 57208
rect 14056 57196 14062 57248
rect 14366 57236 14372 57248
rect 14327 57208 14372 57236
rect 14366 57196 14372 57208
rect 14424 57196 14430 57248
rect 16206 57236 16212 57248
rect 16167 57208 16212 57236
rect 16206 57196 16212 57208
rect 16264 57196 16270 57248
rect 16850 57236 16856 57248
rect 16811 57208 16856 57236
rect 16850 57196 16856 57208
rect 16908 57196 16914 57248
rect 17126 57196 17132 57248
rect 17184 57236 17190 57248
rect 17405 57239 17463 57245
rect 17405 57236 17417 57239
rect 17184 57208 17417 57236
rect 17184 57196 17190 57208
rect 17405 57205 17417 57208
rect 17451 57205 17463 57239
rect 17405 57199 17463 57205
rect 17586 57196 17592 57248
rect 17644 57236 17650 57248
rect 17788 57245 17816 57344
rect 18196 57341 18208 57344
rect 18242 57341 18254 57375
rect 18196 57335 18254 57341
rect 19518 57332 19524 57384
rect 19576 57372 19582 57384
rect 20070 57372 20076 57384
rect 19576 57344 20076 57372
rect 19576 57332 19582 57344
rect 20070 57332 20076 57344
rect 20128 57332 20134 57384
rect 20257 57375 20315 57381
rect 20257 57341 20269 57375
rect 20303 57372 20315 57375
rect 20346 57372 20352 57384
rect 20303 57344 20352 57372
rect 20303 57341 20315 57344
rect 20257 57335 20315 57341
rect 20346 57332 20352 57344
rect 20404 57372 20410 57384
rect 20456 57372 20484 57480
rect 21634 57468 21640 57480
rect 21692 57468 21698 57520
rect 23934 57508 23940 57520
rect 23895 57480 23940 57508
rect 23934 57468 23940 57480
rect 23992 57468 23998 57520
rect 20404 57344 20484 57372
rect 20533 57375 20591 57381
rect 20404 57332 20410 57344
rect 20533 57341 20545 57375
rect 20579 57372 20591 57375
rect 20579 57344 20668 57372
rect 20579 57341 20591 57344
rect 20533 57335 20591 57341
rect 18046 57304 18052 57316
rect 18007 57276 18052 57304
rect 18046 57264 18052 57276
rect 18104 57264 18110 57316
rect 20640 57248 20668 57344
rect 20714 57332 20720 57384
rect 20772 57372 20778 57384
rect 21085 57375 21143 57381
rect 21085 57372 21097 57375
rect 20772 57344 21097 57372
rect 20772 57332 20778 57344
rect 21085 57341 21097 57344
rect 21131 57341 21143 57375
rect 21085 57335 21143 57341
rect 21637 57375 21695 57381
rect 21637 57341 21649 57375
rect 21683 57372 21695 57375
rect 22370 57372 22376 57384
rect 21683 57344 22376 57372
rect 21683 57341 21695 57344
rect 21637 57335 21695 57341
rect 22370 57332 22376 57344
rect 22428 57332 22434 57384
rect 20809 57307 20867 57313
rect 20809 57273 20821 57307
rect 20855 57304 20867 57307
rect 21818 57304 21824 57316
rect 20855 57276 21824 57304
rect 20855 57273 20867 57276
rect 20809 57267 20867 57273
rect 21818 57264 21824 57276
rect 21876 57264 21882 57316
rect 17773 57239 17831 57245
rect 17773 57236 17785 57239
rect 17644 57208 17785 57236
rect 17644 57196 17650 57208
rect 17773 57205 17785 57208
rect 17819 57205 17831 57239
rect 19058 57236 19064 57248
rect 19019 57208 19064 57236
rect 17773 57199 17831 57205
rect 19058 57196 19064 57208
rect 19116 57196 19122 57248
rect 20622 57196 20628 57248
rect 20680 57196 20686 57248
rect 1104 57146 28888 57168
rect 1104 57094 10982 57146
rect 11034 57094 11046 57146
rect 11098 57094 11110 57146
rect 11162 57094 11174 57146
rect 11226 57094 20982 57146
rect 21034 57094 21046 57146
rect 21098 57094 21110 57146
rect 21162 57094 21174 57146
rect 21226 57094 28888 57146
rect 1104 57072 28888 57094
rect 2130 56992 2136 57044
rect 2188 57032 2194 57044
rect 2777 57035 2835 57041
rect 2777 57032 2789 57035
rect 2188 57004 2789 57032
rect 2188 56992 2194 57004
rect 2777 57001 2789 57004
rect 2823 57001 2835 57035
rect 7006 57032 7012 57044
rect 6967 57004 7012 57032
rect 2777 56995 2835 57001
rect 7006 56992 7012 57004
rect 7064 56992 7070 57044
rect 13357 57035 13415 57041
rect 13357 57001 13369 57035
rect 13403 57032 13415 57035
rect 13446 57032 13452 57044
rect 13403 57004 13452 57032
rect 13403 57001 13415 57004
rect 13357 56995 13415 57001
rect 13446 56992 13452 57004
rect 13504 56992 13510 57044
rect 13722 57032 13728 57044
rect 13683 57004 13728 57032
rect 13722 56992 13728 57004
rect 13780 56992 13786 57044
rect 14366 57032 14372 57044
rect 14327 57004 14372 57032
rect 14366 56992 14372 57004
rect 14424 56992 14430 57044
rect 16574 56992 16580 57044
rect 16632 57032 16638 57044
rect 17865 57035 17923 57041
rect 17865 57032 17877 57035
rect 16632 57004 17877 57032
rect 16632 56992 16638 57004
rect 17865 57001 17877 57004
rect 17911 57001 17923 57035
rect 20714 57032 20720 57044
rect 20675 57004 20720 57032
rect 17865 56995 17923 57001
rect 20714 56992 20720 57004
rect 20772 56992 20778 57044
rect 21085 57035 21143 57041
rect 21085 57001 21097 57035
rect 21131 57032 21143 57035
rect 21634 57032 21640 57044
rect 21131 57004 21640 57032
rect 21131 57001 21143 57004
rect 21085 56995 21143 57001
rect 21634 56992 21640 57004
rect 21692 57032 21698 57044
rect 21729 57035 21787 57041
rect 21729 57032 21741 57035
rect 21692 57004 21741 57032
rect 21692 56992 21698 57004
rect 21729 57001 21741 57004
rect 21775 57032 21787 57035
rect 22097 57035 22155 57041
rect 22097 57032 22109 57035
rect 21775 57004 22109 57032
rect 21775 57001 21787 57004
rect 21729 56995 21787 57001
rect 22097 57001 22109 57004
rect 22143 57001 22155 57035
rect 22097 56995 22155 57001
rect 23201 57035 23259 57041
rect 23201 57001 23213 57035
rect 23247 57032 23259 57035
rect 23290 57032 23296 57044
rect 23247 57004 23296 57032
rect 23247 57001 23259 57004
rect 23201 56995 23259 57001
rect 23290 56992 23296 57004
rect 23348 56992 23354 57044
rect 14093 56967 14151 56973
rect 14093 56933 14105 56967
rect 14139 56964 14151 56967
rect 17218 56964 17224 56976
rect 14139 56936 16252 56964
rect 17179 56936 17224 56964
rect 14139 56933 14151 56936
rect 14093 56927 14151 56933
rect 1670 56896 1676 56908
rect 1631 56868 1676 56896
rect 1670 56856 1676 56868
rect 1728 56856 1734 56908
rect 13173 56899 13231 56905
rect 13173 56865 13185 56899
rect 13219 56896 13231 56899
rect 13262 56896 13268 56908
rect 13219 56868 13268 56896
rect 13219 56865 13231 56868
rect 13173 56859 13231 56865
rect 13262 56856 13268 56868
rect 13320 56856 13326 56908
rect 14182 56896 14188 56908
rect 14143 56868 14188 56896
rect 14182 56856 14188 56868
rect 14240 56856 14246 56908
rect 14734 56856 14740 56908
rect 14792 56896 14798 56908
rect 16224 56905 16252 56936
rect 17218 56924 17224 56936
rect 17276 56924 17282 56976
rect 19978 56964 19984 56976
rect 18892 56936 19984 56964
rect 15657 56899 15715 56905
rect 15657 56896 15669 56899
rect 14792 56868 15669 56896
rect 14792 56856 14798 56868
rect 15657 56865 15669 56868
rect 15703 56865 15715 56899
rect 15657 56859 15715 56865
rect 16209 56899 16267 56905
rect 16209 56865 16221 56899
rect 16255 56896 16267 56899
rect 16482 56896 16488 56908
rect 16255 56868 16488 56896
rect 16255 56865 16267 56868
rect 16209 56859 16267 56865
rect 16482 56856 16488 56868
rect 16540 56856 16546 56908
rect 16574 56856 16580 56908
rect 16632 56896 16638 56908
rect 17236 56896 17264 56924
rect 16632 56868 17264 56896
rect 16632 56856 16638 56868
rect 18506 56856 18512 56908
rect 18564 56896 18570 56908
rect 18892 56905 18920 56936
rect 19978 56924 19984 56936
rect 20036 56964 20042 56976
rect 20257 56967 20315 56973
rect 20257 56964 20269 56967
rect 20036 56936 20269 56964
rect 20036 56924 20042 56936
rect 20257 56933 20269 56936
rect 20303 56933 20315 56967
rect 21361 56967 21419 56973
rect 21361 56964 21373 56967
rect 20257 56927 20315 56933
rect 20456 56936 21373 56964
rect 20456 56908 20484 56936
rect 21361 56933 21373 56936
rect 21407 56933 21419 56967
rect 21361 56927 21419 56933
rect 18877 56899 18935 56905
rect 18877 56896 18889 56899
rect 18564 56868 18889 56896
rect 18564 56856 18570 56868
rect 18877 56865 18889 56868
rect 18923 56865 18935 56899
rect 19334 56896 19340 56908
rect 19295 56868 19340 56896
rect 18877 56859 18935 56865
rect 19334 56856 19340 56868
rect 19392 56856 19398 56908
rect 19702 56856 19708 56908
rect 19760 56896 19766 56908
rect 19797 56899 19855 56905
rect 19797 56896 19809 56899
rect 19760 56868 19809 56896
rect 19760 56856 19766 56868
rect 19797 56865 19809 56868
rect 19843 56896 19855 56899
rect 20438 56896 20444 56908
rect 19843 56868 20444 56896
rect 19843 56865 19855 56868
rect 19797 56859 19855 56865
rect 20438 56856 20444 56868
rect 20496 56856 20502 56908
rect 20901 56899 20959 56905
rect 20901 56865 20913 56899
rect 20947 56896 20959 56899
rect 20990 56896 20996 56908
rect 20947 56868 20996 56896
rect 20947 56865 20959 56868
rect 20901 56859 20959 56865
rect 20990 56856 20996 56868
rect 21048 56856 21054 56908
rect 22738 56856 22744 56908
rect 22796 56896 22802 56908
rect 22833 56899 22891 56905
rect 22833 56896 22845 56899
rect 22796 56868 22845 56896
rect 22796 56856 22802 56868
rect 22833 56865 22845 56868
rect 22879 56865 22891 56899
rect 22833 56859 22891 56865
rect 1397 56831 1455 56837
rect 1397 56797 1409 56831
rect 1443 56828 1455 56831
rect 1578 56828 1584 56840
rect 1443 56800 1584 56828
rect 1443 56797 1455 56800
rect 1397 56791 1455 56797
rect 1578 56788 1584 56800
rect 1636 56828 1642 56840
rect 2130 56828 2136 56840
rect 1636 56800 2136 56828
rect 1636 56788 1642 56800
rect 2130 56788 2136 56800
rect 2188 56788 2194 56840
rect 14918 56788 14924 56840
rect 14976 56828 14982 56840
rect 15381 56831 15439 56837
rect 15381 56828 15393 56831
rect 14976 56800 15393 56828
rect 14976 56788 14982 56800
rect 15381 56797 15393 56800
rect 15427 56797 15439 56831
rect 15381 56791 15439 56797
rect 17589 56831 17647 56837
rect 17589 56797 17601 56831
rect 17635 56828 17647 56831
rect 17770 56828 17776 56840
rect 17635 56800 17776 56828
rect 17635 56797 17647 56800
rect 17589 56791 17647 56797
rect 17770 56788 17776 56800
rect 17828 56788 17834 56840
rect 19981 56831 20039 56837
rect 19981 56797 19993 56831
rect 20027 56828 20039 56831
rect 20070 56828 20076 56840
rect 20027 56800 20076 56828
rect 20027 56797 20039 56800
rect 19981 56791 20039 56797
rect 20070 56788 20076 56800
rect 20128 56788 20134 56840
rect 21358 56788 21364 56840
rect 21416 56828 21422 56840
rect 21818 56828 21824 56840
rect 21416 56800 21824 56828
rect 21416 56788 21422 56800
rect 21818 56788 21824 56800
rect 21876 56828 21882 56840
rect 22465 56831 22523 56837
rect 22465 56828 22477 56831
rect 21876 56800 22477 56828
rect 21876 56788 21882 56800
rect 22465 56797 22477 56800
rect 22511 56797 22523 56831
rect 22465 56791 22523 56797
rect 15746 56720 15752 56772
rect 15804 56760 15810 56772
rect 16117 56763 16175 56769
rect 16117 56760 16129 56763
rect 15804 56732 16129 56760
rect 15804 56720 15810 56732
rect 16117 56729 16129 56732
rect 16163 56729 16175 56763
rect 16117 56723 16175 56729
rect 16206 56720 16212 56772
rect 16264 56760 16270 56772
rect 16666 56760 16672 56772
rect 16264 56732 16672 56760
rect 16264 56720 16270 56732
rect 16666 56720 16672 56732
rect 16724 56720 16730 56772
rect 16942 56720 16948 56772
rect 17000 56760 17006 56772
rect 17037 56763 17095 56769
rect 17037 56760 17049 56763
rect 17000 56732 17049 56760
rect 17000 56720 17006 56732
rect 17037 56729 17049 56732
rect 17083 56760 17095 56763
rect 17954 56760 17960 56772
rect 17083 56732 17960 56760
rect 17083 56729 17095 56732
rect 17037 56723 17095 56729
rect 17954 56720 17960 56732
rect 18012 56720 18018 56772
rect 18046 56720 18052 56772
rect 18104 56760 18110 56772
rect 18601 56763 18659 56769
rect 18601 56760 18613 56763
rect 18104 56732 18613 56760
rect 18104 56720 18110 56732
rect 18601 56729 18613 56732
rect 18647 56760 18659 56763
rect 19058 56760 19064 56772
rect 18647 56732 19064 56760
rect 18647 56729 18659 56732
rect 18601 56723 18659 56729
rect 19058 56720 19064 56732
rect 19116 56720 19122 56772
rect 19518 56720 19524 56772
rect 19576 56760 19582 56772
rect 19702 56760 19708 56772
rect 19576 56732 19708 56760
rect 19576 56720 19582 56732
rect 19702 56720 19708 56732
rect 19760 56720 19766 56772
rect 14737 56695 14795 56701
rect 14737 56661 14749 56695
rect 14783 56692 14795 56695
rect 15102 56692 15108 56704
rect 14783 56664 15108 56692
rect 14783 56661 14795 56664
rect 14737 56655 14795 56661
rect 15102 56652 15108 56664
rect 15160 56652 15166 56704
rect 17218 56652 17224 56704
rect 17276 56692 17282 56704
rect 17359 56695 17417 56701
rect 17359 56692 17371 56695
rect 17276 56664 17371 56692
rect 17276 56652 17282 56664
rect 17359 56661 17371 56664
rect 17405 56661 17417 56695
rect 17494 56692 17500 56704
rect 17455 56664 17500 56692
rect 17359 56655 17417 56661
rect 17494 56652 17500 56664
rect 17552 56652 17558 56704
rect 17586 56652 17592 56704
rect 17644 56692 17650 56704
rect 18233 56695 18291 56701
rect 18233 56692 18245 56695
rect 17644 56664 18245 56692
rect 17644 56652 17650 56664
rect 18233 56661 18245 56664
rect 18279 56661 18291 56695
rect 18233 56655 18291 56661
rect 23290 56652 23296 56704
rect 23348 56692 23354 56704
rect 23934 56692 23940 56704
rect 23348 56664 23940 56692
rect 23348 56652 23354 56664
rect 23934 56652 23940 56664
rect 23992 56652 23998 56704
rect 1104 56602 28888 56624
rect 1104 56550 5982 56602
rect 6034 56550 6046 56602
rect 6098 56550 6110 56602
rect 6162 56550 6174 56602
rect 6226 56550 15982 56602
rect 16034 56550 16046 56602
rect 16098 56550 16110 56602
rect 16162 56550 16174 56602
rect 16226 56550 25982 56602
rect 26034 56550 26046 56602
rect 26098 56550 26110 56602
rect 26162 56550 26174 56602
rect 26226 56550 28888 56602
rect 1104 56528 28888 56550
rect 1670 56488 1676 56500
rect 1631 56460 1676 56488
rect 1670 56448 1676 56460
rect 1728 56448 1734 56500
rect 2041 56491 2099 56497
rect 2041 56457 2053 56491
rect 2087 56488 2099 56491
rect 2222 56488 2228 56500
rect 2087 56460 2228 56488
rect 2087 56457 2099 56460
rect 2041 56451 2099 56457
rect 2222 56448 2228 56460
rect 2280 56448 2286 56500
rect 15194 56488 15200 56500
rect 15155 56460 15200 56488
rect 15194 56448 15200 56460
rect 15252 56448 15258 56500
rect 17954 56448 17960 56500
rect 18012 56488 18018 56500
rect 18509 56491 18567 56497
rect 18509 56488 18521 56491
rect 18012 56460 18521 56488
rect 18012 56448 18018 56460
rect 18509 56457 18521 56460
rect 18555 56457 18567 56491
rect 18509 56451 18567 56457
rect 19705 56491 19763 56497
rect 19705 56457 19717 56491
rect 19751 56488 19763 56491
rect 20714 56488 20720 56500
rect 19751 56460 20720 56488
rect 19751 56457 19763 56460
rect 19705 56451 19763 56457
rect 20714 56448 20720 56460
rect 20772 56448 20778 56500
rect 20990 56448 20996 56500
rect 21048 56488 21054 56500
rect 21729 56491 21787 56497
rect 21729 56488 21741 56491
rect 21048 56460 21741 56488
rect 21048 56448 21054 56460
rect 21729 56457 21741 56460
rect 21775 56457 21787 56491
rect 21729 56451 21787 56457
rect 23014 56448 23020 56500
rect 23072 56488 23078 56500
rect 23109 56491 23167 56497
rect 23109 56488 23121 56491
rect 23072 56460 23121 56488
rect 23072 56448 23078 56460
rect 23109 56457 23121 56460
rect 23155 56457 23167 56491
rect 23109 56451 23167 56457
rect 25774 56448 25780 56500
rect 25832 56488 25838 56500
rect 26053 56491 26111 56497
rect 26053 56488 26065 56491
rect 25832 56460 26065 56488
rect 25832 56448 25838 56460
rect 26053 56457 26065 56460
rect 26099 56457 26111 56491
rect 26053 56451 26111 56457
rect 13722 56420 13728 56432
rect 13683 56392 13728 56420
rect 13722 56380 13728 56392
rect 13780 56380 13786 56432
rect 14829 56423 14887 56429
rect 14829 56389 14841 56423
rect 14875 56420 14887 56423
rect 15010 56420 15016 56432
rect 14875 56392 15016 56420
rect 14875 56389 14887 56392
rect 14829 56383 14887 56389
rect 15010 56380 15016 56392
rect 15068 56380 15074 56432
rect 15102 56380 15108 56432
rect 15160 56420 15166 56432
rect 15749 56423 15807 56429
rect 15749 56420 15761 56423
rect 15160 56392 15761 56420
rect 15160 56380 15166 56392
rect 15749 56389 15761 56392
rect 15795 56389 15807 56423
rect 15749 56383 15807 56389
rect 16393 56423 16451 56429
rect 16393 56389 16405 56423
rect 16439 56389 16451 56423
rect 16574 56420 16580 56432
rect 16535 56392 16580 56420
rect 16393 56383 16451 56389
rect 14274 56312 14280 56364
rect 14332 56352 14338 56364
rect 14921 56355 14979 56361
rect 14921 56352 14933 56355
rect 14332 56324 14933 56352
rect 14332 56312 14338 56324
rect 14921 56321 14933 56324
rect 14967 56321 14979 56355
rect 14921 56315 14979 56321
rect 15194 56312 15200 56364
rect 15252 56352 15258 56364
rect 15933 56355 15991 56361
rect 15933 56352 15945 56355
rect 15252 56324 15945 56352
rect 15252 56312 15258 56324
rect 15933 56321 15945 56324
rect 15979 56352 15991 56355
rect 16114 56352 16120 56364
rect 15979 56324 16120 56352
rect 15979 56321 15991 56324
rect 15933 56315 15991 56321
rect 16114 56312 16120 56324
rect 16172 56352 16178 56364
rect 16408 56352 16436 56383
rect 16574 56380 16580 56392
rect 16632 56380 16638 56432
rect 17494 56380 17500 56432
rect 17552 56420 17558 56432
rect 18322 56420 18328 56432
rect 17552 56392 18328 56420
rect 17552 56380 17558 56392
rect 18322 56380 18328 56392
rect 18380 56380 18386 56432
rect 19058 56380 19064 56432
rect 19116 56380 19122 56432
rect 19334 56380 19340 56432
rect 19392 56420 19398 56432
rect 21361 56423 21419 56429
rect 21361 56420 21373 56423
rect 19392 56392 21373 56420
rect 19392 56380 19398 56392
rect 21361 56389 21373 56392
rect 21407 56389 21419 56423
rect 21361 56383 21419 56389
rect 16172 56324 16436 56352
rect 16485 56355 16543 56361
rect 16172 56312 16178 56324
rect 16485 56321 16497 56355
rect 16531 56352 16543 56355
rect 16666 56352 16672 56364
rect 16531 56324 16672 56352
rect 16531 56321 16543 56324
rect 16485 56315 16543 56321
rect 14700 56287 14758 56293
rect 14700 56253 14712 56287
rect 14746 56284 14758 56287
rect 16264 56287 16322 56293
rect 16264 56284 16276 56287
rect 14746 56256 16276 56284
rect 14746 56253 14758 56256
rect 14700 56247 14758 56253
rect 14553 56219 14611 56225
rect 14553 56185 14565 56219
rect 14599 56216 14611 56219
rect 15102 56216 15108 56228
rect 14599 56188 15108 56216
rect 14599 56185 14611 56188
rect 14553 56179 14611 56185
rect 15102 56176 15108 56188
rect 15160 56176 15166 56228
rect 15580 56160 15608 56256
rect 16264 56253 16276 56256
rect 16310 56253 16322 56287
rect 16264 56247 16322 56253
rect 15749 56219 15807 56225
rect 15749 56185 15761 56219
rect 15795 56216 15807 56219
rect 16117 56219 16175 56225
rect 16117 56216 16129 56219
rect 15795 56188 16129 56216
rect 15795 56185 15807 56188
rect 15749 56179 15807 56185
rect 16117 56185 16129 56188
rect 16163 56216 16175 56219
rect 16482 56216 16488 56228
rect 16163 56188 16488 56216
rect 16163 56185 16175 56188
rect 16117 56179 16175 56185
rect 16482 56176 16488 56188
rect 16540 56176 16546 56228
rect 13262 56148 13268 56160
rect 13223 56120 13268 56148
rect 13262 56108 13268 56120
rect 13320 56108 13326 56160
rect 14093 56151 14151 56157
rect 14093 56117 14105 56151
rect 14139 56148 14151 56151
rect 14274 56148 14280 56160
rect 14139 56120 14280 56148
rect 14139 56117 14151 56120
rect 14093 56111 14151 56117
rect 14274 56108 14280 56120
rect 14332 56108 14338 56160
rect 14461 56151 14519 56157
rect 14461 56117 14473 56151
rect 14507 56148 14519 56151
rect 15010 56148 15016 56160
rect 14507 56120 15016 56148
rect 14507 56117 14519 56120
rect 14461 56111 14519 56117
rect 15010 56108 15016 56120
rect 15068 56108 15074 56160
rect 15562 56148 15568 56160
rect 15523 56120 15568 56148
rect 15562 56108 15568 56120
rect 15620 56108 15626 56160
rect 16206 56108 16212 56160
rect 16264 56148 16270 56160
rect 16592 56148 16620 56324
rect 16666 56312 16672 56324
rect 16724 56312 16730 56364
rect 17770 56352 17776 56364
rect 17683 56324 17776 56352
rect 17770 56312 17776 56324
rect 17828 56352 17834 56364
rect 18417 56355 18475 56361
rect 18417 56352 18429 56355
rect 17828 56324 18429 56352
rect 17828 56312 17834 56324
rect 18417 56321 18429 56324
rect 18463 56321 18475 56355
rect 19076 56352 19104 56380
rect 19610 56352 19616 56364
rect 19076 56324 19380 56352
rect 19523 56324 19616 56352
rect 18417 56315 18475 56321
rect 16264 56120 16620 56148
rect 16264 56108 16270 56120
rect 16942 56108 16948 56160
rect 17000 56148 17006 56160
rect 17788 56157 17816 56312
rect 18196 56287 18254 56293
rect 18196 56253 18208 56287
rect 18242 56284 18254 56287
rect 19061 56287 19119 56293
rect 19061 56284 19073 56287
rect 18242 56256 19073 56284
rect 18242 56253 18254 56256
rect 18196 56247 18254 56253
rect 18432 56228 18460 56256
rect 19061 56253 19073 56256
rect 19107 56253 19119 56287
rect 19352 56284 19380 56324
rect 19610 56312 19616 56324
rect 19668 56352 19674 56364
rect 20073 56355 20131 56361
rect 20073 56352 20085 56355
rect 19668 56324 20085 56352
rect 19668 56312 19674 56324
rect 20073 56321 20085 56324
rect 20119 56321 20131 56355
rect 23032 56352 23060 56448
rect 20073 56315 20131 56321
rect 20824 56324 23060 56352
rect 19889 56287 19947 56293
rect 19889 56284 19901 56287
rect 19352 56256 19901 56284
rect 19061 56247 19119 56253
rect 19889 56253 19901 56256
rect 19935 56253 19947 56287
rect 20346 56284 20352 56296
rect 20307 56256 20352 56284
rect 19889 56247 19947 56253
rect 18046 56216 18052 56228
rect 18007 56188 18052 56216
rect 18046 56176 18052 56188
rect 18104 56176 18110 56228
rect 18414 56176 18420 56228
rect 18472 56176 18478 56228
rect 17221 56151 17279 56157
rect 17221 56148 17233 56151
rect 17000 56120 17233 56148
rect 17000 56108 17006 56120
rect 17221 56117 17233 56120
rect 17267 56148 17279 56151
rect 17773 56151 17831 56157
rect 17773 56148 17785 56151
rect 17267 56120 17785 56148
rect 17267 56117 17279 56120
rect 17221 56111 17279 56117
rect 17773 56117 17785 56120
rect 17819 56117 17831 56151
rect 19904 56148 19932 56247
rect 20346 56244 20352 56256
rect 20404 56244 20410 56296
rect 20714 56244 20720 56296
rect 20772 56284 20778 56296
rect 20824 56293 20852 56324
rect 25866 56312 25872 56364
rect 25924 56352 25930 56364
rect 26145 56355 26203 56361
rect 26145 56352 26157 56355
rect 25924 56324 26157 56352
rect 25924 56312 25930 56324
rect 26145 56321 26157 56324
rect 26191 56321 26203 56355
rect 26145 56315 26203 56321
rect 20809 56287 20867 56293
rect 20809 56284 20821 56287
rect 20772 56256 20821 56284
rect 20772 56244 20778 56256
rect 20809 56253 20821 56256
rect 20855 56253 20867 56287
rect 20809 56247 20867 56253
rect 21358 56244 21364 56296
rect 21416 56284 21422 56296
rect 21913 56287 21971 56293
rect 21913 56284 21925 56287
rect 21416 56256 21925 56284
rect 21416 56244 21422 56256
rect 21913 56253 21925 56256
rect 21959 56284 21971 56287
rect 22373 56287 22431 56293
rect 22373 56284 22385 56287
rect 21959 56256 22385 56284
rect 21959 56253 21971 56256
rect 21913 56247 21971 56253
rect 22373 56253 22385 56256
rect 22419 56253 22431 56287
rect 22373 56247 22431 56253
rect 25774 56244 25780 56296
rect 25832 56284 25838 56296
rect 26421 56287 26479 56293
rect 26421 56284 26433 56287
rect 25832 56256 26433 56284
rect 25832 56244 25838 56256
rect 26421 56253 26433 56256
rect 26467 56253 26479 56287
rect 26421 56247 26479 56253
rect 21085 56219 21143 56225
rect 21085 56185 21097 56219
rect 21131 56216 21143 56219
rect 21266 56216 21272 56228
rect 21131 56188 21272 56216
rect 21131 56185 21143 56188
rect 21085 56179 21143 56185
rect 21266 56176 21272 56188
rect 21324 56176 21330 56228
rect 22462 56176 22468 56228
rect 22520 56216 22526 56228
rect 22830 56216 22836 56228
rect 22520 56188 22836 56216
rect 22520 56176 22526 56188
rect 22830 56176 22836 56188
rect 22888 56176 22894 56228
rect 21634 56148 21640 56160
rect 19904 56120 21640 56148
rect 17773 56111 17831 56117
rect 21634 56108 21640 56120
rect 21692 56108 21698 56160
rect 22094 56108 22100 56160
rect 22152 56148 22158 56160
rect 22738 56148 22744 56160
rect 22152 56120 22197 56148
rect 22699 56120 22744 56148
rect 22152 56108 22158 56120
rect 22738 56108 22744 56120
rect 22796 56108 22802 56160
rect 24302 56108 24308 56160
rect 24360 56148 24366 56160
rect 24670 56148 24676 56160
rect 24360 56120 24676 56148
rect 24360 56108 24366 56120
rect 24670 56108 24676 56120
rect 24728 56108 24734 56160
rect 27706 56148 27712 56160
rect 27667 56120 27712 56148
rect 27706 56108 27712 56120
rect 27764 56108 27770 56160
rect 1104 56058 28888 56080
rect 1104 56006 10982 56058
rect 11034 56006 11046 56058
rect 11098 56006 11110 56058
rect 11162 56006 11174 56058
rect 11226 56006 20982 56058
rect 21034 56006 21046 56058
rect 21098 56006 21110 56058
rect 21162 56006 21174 56058
rect 21226 56006 28888 56058
rect 1104 55984 28888 56006
rect 13998 55944 14004 55956
rect 13959 55916 14004 55944
rect 13998 55904 14004 55916
rect 14056 55904 14062 55956
rect 14274 55904 14280 55956
rect 14332 55944 14338 55956
rect 14369 55947 14427 55953
rect 14369 55944 14381 55947
rect 14332 55916 14381 55944
rect 14332 55904 14338 55916
rect 14369 55913 14381 55916
rect 14415 55913 14427 55947
rect 14369 55907 14427 55913
rect 16114 55904 16120 55956
rect 16172 55944 16178 55956
rect 17494 55944 17500 55956
rect 16172 55916 17500 55944
rect 16172 55904 16178 55916
rect 17494 55904 17500 55916
rect 17552 55944 17558 55956
rect 17589 55947 17647 55953
rect 17589 55944 17601 55947
rect 17552 55916 17601 55944
rect 17552 55904 17558 55916
rect 17589 55913 17601 55916
rect 17635 55944 17647 55947
rect 18417 55947 18475 55953
rect 18417 55944 18429 55947
rect 17635 55916 18429 55944
rect 17635 55913 17647 55916
rect 17589 55907 17647 55913
rect 18417 55913 18429 55916
rect 18463 55913 18475 55947
rect 18417 55907 18475 55913
rect 19978 55904 19984 55956
rect 20036 55944 20042 55956
rect 20073 55947 20131 55953
rect 20073 55944 20085 55947
rect 20036 55916 20085 55944
rect 20036 55904 20042 55916
rect 20073 55913 20085 55916
rect 20119 55913 20131 55947
rect 20073 55907 20131 55913
rect 20254 55904 20260 55956
rect 20312 55904 20318 55956
rect 20438 55944 20444 55956
rect 20399 55916 20444 55944
rect 20438 55904 20444 55916
rect 20496 55904 20502 55956
rect 21634 55904 21640 55956
rect 21692 55944 21698 55956
rect 22925 55947 22983 55953
rect 22925 55944 22937 55947
rect 21692 55916 22937 55944
rect 21692 55904 21698 55916
rect 22925 55913 22937 55916
rect 22971 55913 22983 55947
rect 22925 55907 22983 55913
rect 25866 55904 25872 55956
rect 25924 55944 25930 55956
rect 26145 55947 26203 55953
rect 26145 55944 26157 55947
rect 25924 55916 26157 55944
rect 25924 55904 25930 55916
rect 26145 55913 26157 55916
rect 26191 55913 26203 55947
rect 26145 55907 26203 55913
rect 14826 55836 14832 55888
rect 14884 55876 14890 55888
rect 16206 55876 16212 55888
rect 14884 55848 16212 55876
rect 14884 55836 14890 55848
rect 16206 55836 16212 55848
rect 16264 55836 16270 55888
rect 17313 55879 17371 55885
rect 17313 55845 17325 55879
rect 17359 55876 17371 55879
rect 17770 55876 17776 55888
rect 17359 55848 17776 55876
rect 17359 55845 17371 55848
rect 17313 55839 17371 55845
rect 17770 55836 17776 55848
rect 17828 55836 17834 55888
rect 18782 55876 18788 55888
rect 18743 55848 18788 55876
rect 18782 55836 18788 55848
rect 18840 55836 18846 55888
rect 19334 55836 19340 55888
rect 19392 55836 19398 55888
rect 9674 55768 9680 55820
rect 9732 55808 9738 55820
rect 10594 55808 10600 55820
rect 9732 55780 10600 55808
rect 9732 55768 9738 55780
rect 10594 55768 10600 55780
rect 10652 55808 10658 55820
rect 10781 55811 10839 55817
rect 10781 55808 10793 55811
rect 10652 55780 10793 55808
rect 10652 55768 10658 55780
rect 10781 55777 10793 55780
rect 10827 55777 10839 55811
rect 13170 55808 13176 55820
rect 13131 55780 13176 55808
rect 10781 55771 10839 55777
rect 13170 55768 13176 55780
rect 13228 55768 13234 55820
rect 13998 55768 14004 55820
rect 14056 55808 14062 55820
rect 14185 55811 14243 55817
rect 14185 55808 14197 55811
rect 14056 55780 14197 55808
rect 14056 55768 14062 55780
rect 14185 55777 14197 55780
rect 14231 55777 14243 55811
rect 15565 55811 15623 55817
rect 15565 55808 15577 55811
rect 14185 55771 14243 55777
rect 14660 55780 15577 55808
rect 10505 55743 10563 55749
rect 10505 55709 10517 55743
rect 10551 55740 10563 55743
rect 10870 55740 10876 55752
rect 10551 55712 10876 55740
rect 10551 55709 10563 55712
rect 10505 55703 10563 55709
rect 10870 55700 10876 55712
rect 10928 55700 10934 55752
rect 13357 55675 13415 55681
rect 13357 55641 13369 55675
rect 13403 55672 13415 55675
rect 14366 55672 14372 55684
rect 13403 55644 14372 55672
rect 13403 55641 13415 55644
rect 13357 55635 13415 55641
rect 14366 55632 14372 55644
rect 14424 55632 14430 55684
rect 12066 55604 12072 55616
rect 12027 55576 12072 55604
rect 12066 55564 12072 55576
rect 12124 55564 12130 55616
rect 13078 55564 13084 55616
rect 13136 55604 13142 55616
rect 13633 55607 13691 55613
rect 13633 55604 13645 55607
rect 13136 55576 13645 55604
rect 13136 55564 13142 55576
rect 13633 55573 13645 55576
rect 13679 55604 13691 55607
rect 14660 55604 14688 55780
rect 15565 55777 15577 55780
rect 15611 55777 15623 55811
rect 15565 55771 15623 55777
rect 16577 55811 16635 55817
rect 16577 55777 16589 55811
rect 16623 55808 16635 55811
rect 16850 55808 16856 55820
rect 16623 55780 16856 55808
rect 16623 55777 16635 55780
rect 16577 55771 16635 55777
rect 16850 55768 16856 55780
rect 16908 55768 16914 55820
rect 19352 55808 19380 55836
rect 19613 55811 19671 55817
rect 19613 55808 19625 55811
rect 19352 55780 19625 55808
rect 19613 55777 19625 55780
rect 19659 55777 19671 55811
rect 19613 55771 19671 55777
rect 16942 55740 16948 55752
rect 16903 55712 16948 55740
rect 16942 55700 16948 55712
rect 17000 55740 17006 55752
rect 18049 55743 18107 55749
rect 18049 55740 18061 55743
rect 17000 55712 18061 55740
rect 17000 55700 17006 55712
rect 18049 55709 18061 55712
rect 18095 55709 18107 55743
rect 18049 55703 18107 55709
rect 19058 55700 19064 55752
rect 19116 55740 19122 55752
rect 19337 55743 19395 55749
rect 19337 55740 19349 55743
rect 19116 55712 19349 55740
rect 19116 55700 19122 55712
rect 19337 55709 19349 55712
rect 19383 55709 19395 55743
rect 19337 55703 19395 55709
rect 19797 55743 19855 55749
rect 19797 55709 19809 55743
rect 19843 55740 19855 55743
rect 20272 55740 20300 55904
rect 22738 55876 22744 55888
rect 21928 55848 22744 55876
rect 20898 55808 20904 55820
rect 20859 55780 20904 55808
rect 20898 55768 20904 55780
rect 20956 55808 20962 55820
rect 21361 55811 21419 55817
rect 21361 55808 21373 55811
rect 20956 55780 21373 55808
rect 20956 55768 20962 55780
rect 21361 55777 21373 55780
rect 21407 55777 21419 55811
rect 21361 55771 21419 55777
rect 21634 55768 21640 55820
rect 21692 55808 21698 55820
rect 21928 55817 21956 55848
rect 22738 55836 22744 55848
rect 22796 55836 22802 55888
rect 21913 55811 21971 55817
rect 21913 55808 21925 55811
rect 21692 55780 21925 55808
rect 21692 55768 21698 55780
rect 21913 55777 21925 55780
rect 21959 55777 21971 55811
rect 22370 55808 22376 55820
rect 22331 55780 22376 55808
rect 21913 55771 21971 55777
rect 22370 55768 22376 55780
rect 22428 55768 22434 55820
rect 23753 55811 23811 55817
rect 23753 55777 23765 55811
rect 23799 55808 23811 55811
rect 23842 55808 23848 55820
rect 23799 55780 23848 55808
rect 23799 55777 23811 55780
rect 23753 55771 23811 55777
rect 23842 55768 23848 55780
rect 23900 55768 23906 55820
rect 20346 55740 20352 55752
rect 19843 55712 20352 55740
rect 19843 55709 19855 55712
rect 19797 55703 19855 55709
rect 14737 55675 14795 55681
rect 14737 55641 14749 55675
rect 14783 55672 14795 55675
rect 16853 55675 16911 55681
rect 14783 55644 15608 55672
rect 14783 55641 14795 55644
rect 14737 55635 14795 55641
rect 15580 55616 15608 55644
rect 16853 55641 16865 55675
rect 16899 55672 16911 55675
rect 17034 55672 17040 55684
rect 16899 55644 17040 55672
rect 16899 55641 16911 55644
rect 16853 55635 16911 55641
rect 17034 55632 17040 55644
rect 17092 55632 17098 55684
rect 19352 55672 19380 55703
rect 20346 55700 20352 55712
rect 20404 55700 20410 55752
rect 22649 55743 22707 55749
rect 22649 55709 22661 55743
rect 22695 55740 22707 55743
rect 22738 55740 22744 55752
rect 22695 55712 22744 55740
rect 22695 55709 22707 55712
rect 22649 55703 22707 55709
rect 22738 55700 22744 55712
rect 22796 55700 22802 55752
rect 23385 55743 23443 55749
rect 23385 55709 23397 55743
rect 23431 55740 23443 55743
rect 23477 55743 23535 55749
rect 23477 55740 23489 55743
rect 23431 55712 23489 55740
rect 23431 55709 23443 55712
rect 23385 55703 23443 55709
rect 23477 55709 23489 55712
rect 23523 55740 23535 55743
rect 26326 55740 26332 55752
rect 23523 55712 26332 55740
rect 23523 55709 23535 55712
rect 23477 55703 23535 55709
rect 26326 55700 26332 55712
rect 26384 55700 26390 55752
rect 20162 55672 20168 55684
rect 19352 55644 20168 55672
rect 20162 55632 20168 55644
rect 20220 55632 20226 55684
rect 13679 55576 14688 55604
rect 13679 55573 13691 55576
rect 13633 55567 13691 55573
rect 14918 55564 14924 55616
rect 14976 55604 14982 55616
rect 15102 55604 15108 55616
rect 14976 55576 15108 55604
rect 14976 55564 14982 55576
rect 15102 55564 15108 55576
rect 15160 55564 15166 55616
rect 15562 55564 15568 55616
rect 15620 55604 15626 55616
rect 15749 55607 15807 55613
rect 15749 55604 15761 55607
rect 15620 55576 15761 55604
rect 15620 55564 15626 55576
rect 15749 55573 15761 55576
rect 15795 55604 15807 55607
rect 16117 55607 16175 55613
rect 16117 55604 16129 55607
rect 15795 55576 16129 55604
rect 15795 55573 15807 55576
rect 15749 55567 15807 55573
rect 16117 55573 16129 55576
rect 16163 55604 16175 55607
rect 16482 55604 16488 55616
rect 16163 55576 16488 55604
rect 16163 55573 16175 55576
rect 16117 55567 16175 55573
rect 16482 55564 16488 55576
rect 16540 55564 16546 55616
rect 16742 55607 16800 55613
rect 16742 55573 16754 55607
rect 16788 55604 16800 55607
rect 17126 55604 17132 55616
rect 16788 55576 17132 55604
rect 16788 55573 16800 55576
rect 16742 55567 16800 55573
rect 17126 55564 17132 55576
rect 17184 55564 17190 55616
rect 21082 55604 21088 55616
rect 21043 55576 21088 55604
rect 21082 55564 21088 55576
rect 21140 55564 21146 55616
rect 21821 55607 21879 55613
rect 21821 55573 21833 55607
rect 21867 55604 21879 55607
rect 22646 55604 22652 55616
rect 21867 55576 22652 55604
rect 21867 55573 21879 55576
rect 21821 55567 21879 55573
rect 22646 55564 22652 55576
rect 22704 55564 22710 55616
rect 24854 55604 24860 55616
rect 24815 55576 24860 55604
rect 24854 55564 24860 55576
rect 24912 55564 24918 55616
rect 1104 55514 28888 55536
rect 1104 55462 5982 55514
rect 6034 55462 6046 55514
rect 6098 55462 6110 55514
rect 6162 55462 6174 55514
rect 6226 55462 15982 55514
rect 16034 55462 16046 55514
rect 16098 55462 16110 55514
rect 16162 55462 16174 55514
rect 16226 55462 25982 55514
rect 26034 55462 26046 55514
rect 26098 55462 26110 55514
rect 26162 55462 26174 55514
rect 26226 55462 28888 55514
rect 1104 55440 28888 55462
rect 10594 55400 10600 55412
rect 10555 55372 10600 55400
rect 10594 55360 10600 55372
rect 10652 55360 10658 55412
rect 10870 55400 10876 55412
rect 10831 55372 10876 55400
rect 10870 55360 10876 55372
rect 10928 55360 10934 55412
rect 12989 55403 13047 55409
rect 12989 55369 13001 55403
rect 13035 55400 13047 55403
rect 13170 55400 13176 55412
rect 13035 55372 13176 55400
rect 13035 55369 13047 55372
rect 12989 55363 13047 55369
rect 13170 55360 13176 55372
rect 13228 55400 13234 55412
rect 14921 55403 14979 55409
rect 14921 55400 14933 55403
rect 13228 55372 14933 55400
rect 13228 55360 13234 55372
rect 14921 55369 14933 55372
rect 14967 55369 14979 55403
rect 14921 55363 14979 55369
rect 15010 55360 15016 55412
rect 15068 55400 15074 55412
rect 16190 55403 16248 55409
rect 15068 55372 15976 55400
rect 15068 55360 15074 55372
rect 15948 55344 15976 55372
rect 16190 55369 16202 55403
rect 16236 55400 16248 55403
rect 16482 55400 16488 55412
rect 16236 55372 16488 55400
rect 16236 55369 16248 55372
rect 16190 55363 16248 55369
rect 16482 55360 16488 55372
rect 16540 55360 16546 55412
rect 16666 55400 16672 55412
rect 16627 55372 16672 55400
rect 16666 55360 16672 55372
rect 16724 55360 16730 55412
rect 16942 55360 16948 55412
rect 17000 55400 17006 55412
rect 17405 55403 17463 55409
rect 17405 55400 17417 55403
rect 17000 55372 17417 55400
rect 17000 55360 17006 55372
rect 17405 55369 17417 55372
rect 17451 55369 17463 55403
rect 17405 55363 17463 55369
rect 14734 55332 14740 55344
rect 14695 55304 14740 55332
rect 14734 55292 14740 55304
rect 14792 55332 14798 55344
rect 15194 55332 15200 55344
rect 14792 55304 15200 55332
rect 14792 55292 14798 55304
rect 15194 55292 15200 55304
rect 15252 55292 15258 55344
rect 15930 55292 15936 55344
rect 15988 55332 15994 55344
rect 16301 55335 16359 55341
rect 16301 55332 16313 55335
rect 15988 55304 16313 55332
rect 15988 55292 15994 55304
rect 16301 55301 16313 55304
rect 16347 55301 16359 55335
rect 17034 55332 17040 55344
rect 16995 55304 17040 55332
rect 16301 55295 16359 55301
rect 17034 55292 17040 55304
rect 17092 55292 17098 55344
rect 14642 55273 14648 55276
rect 14608 55267 14648 55273
rect 14608 55233 14620 55267
rect 14608 55227 14648 55233
rect 14642 55224 14648 55227
rect 14700 55224 14706 55276
rect 14826 55224 14832 55276
rect 14884 55264 14890 55276
rect 15289 55267 15347 55273
rect 15289 55264 15301 55267
rect 14884 55236 15301 55264
rect 14884 55224 14890 55236
rect 15289 55233 15301 55236
rect 15335 55264 15347 55267
rect 16393 55267 16451 55273
rect 16393 55264 16405 55267
rect 15335 55236 16405 55264
rect 15335 55233 15347 55236
rect 15289 55227 15347 55233
rect 16393 55233 16405 55236
rect 16439 55233 16451 55267
rect 17420 55264 17448 55363
rect 17954 55360 17960 55412
rect 18012 55400 18018 55412
rect 18214 55403 18272 55409
rect 18214 55400 18226 55403
rect 18012 55372 18226 55400
rect 18012 55360 18018 55372
rect 18214 55369 18226 55372
rect 18260 55400 18272 55403
rect 19429 55403 19487 55409
rect 19429 55400 19441 55403
rect 18260 55372 19441 55400
rect 18260 55369 18272 55372
rect 18214 55363 18272 55369
rect 19429 55369 19441 55372
rect 19475 55369 19487 55403
rect 23106 55400 23112 55412
rect 23067 55372 23112 55400
rect 19429 55363 19487 55369
rect 23106 55360 23112 55372
rect 23164 55360 23170 55412
rect 23842 55400 23848 55412
rect 23803 55372 23848 55400
rect 23842 55360 23848 55372
rect 23900 55360 23906 55412
rect 17681 55335 17739 55341
rect 17681 55301 17693 55335
rect 17727 55332 17739 55335
rect 18325 55335 18383 55341
rect 18325 55332 18337 55335
rect 17727 55304 18337 55332
rect 17727 55301 17739 55304
rect 17681 55295 17739 55301
rect 18325 55301 18337 55304
rect 18371 55301 18383 55335
rect 18325 55295 18383 55301
rect 22005 55335 22063 55341
rect 22005 55301 22017 55335
rect 22051 55332 22063 55335
rect 22370 55332 22376 55344
rect 22051 55304 22376 55332
rect 22051 55301 22063 55304
rect 22005 55295 22063 55301
rect 22370 55292 22376 55304
rect 22428 55292 22434 55344
rect 18417 55267 18475 55273
rect 18417 55264 18429 55267
rect 17420 55236 18429 55264
rect 16393 55227 16451 55233
rect 18417 55233 18429 55236
rect 18463 55233 18475 55267
rect 22646 55264 22652 55276
rect 22607 55236 22652 55264
rect 18417 55227 18475 55233
rect 22646 55224 22652 55236
rect 22704 55224 22710 55276
rect 24026 55224 24032 55276
rect 24084 55264 24090 55276
rect 25225 55267 25283 55273
rect 25225 55264 25237 55267
rect 24084 55236 25237 55264
rect 24084 55224 24090 55236
rect 25225 55233 25237 55236
rect 25271 55233 25283 55267
rect 25225 55227 25283 55233
rect 26053 55267 26111 55273
rect 26053 55233 26065 55267
rect 26099 55264 26111 55267
rect 26421 55267 26479 55273
rect 26421 55264 26433 55267
rect 26099 55236 26433 55264
rect 26099 55233 26111 55236
rect 26053 55227 26111 55233
rect 26421 55233 26433 55236
rect 26467 55264 26479 55267
rect 27522 55264 27528 55276
rect 26467 55236 27528 55264
rect 26467 55233 26479 55236
rect 26421 55227 26479 55233
rect 27522 55224 27528 55236
rect 27580 55224 27586 55276
rect 13449 55199 13507 55205
rect 13449 55196 13461 55199
rect 13280 55168 13461 55196
rect 13280 55072 13308 55168
rect 13449 55165 13461 55168
rect 13495 55165 13507 55199
rect 14458 55196 14464 55208
rect 14371 55168 14464 55196
rect 13449 55159 13507 55165
rect 14458 55156 14464 55168
rect 14516 55196 14522 55208
rect 16025 55199 16083 55205
rect 16025 55196 16037 55199
rect 14516 55168 16037 55196
rect 14516 55156 14522 55168
rect 16025 55165 16037 55168
rect 16071 55196 16083 55199
rect 16574 55196 16580 55208
rect 16071 55168 16580 55196
rect 16071 55165 16083 55168
rect 16025 55159 16083 55165
rect 16574 55156 16580 55168
rect 16632 55156 16638 55208
rect 16850 55156 16856 55208
rect 16908 55196 16914 55208
rect 18046 55196 18052 55208
rect 16908 55168 18052 55196
rect 16908 55156 16914 55168
rect 18046 55156 18052 55168
rect 18104 55196 18110 55208
rect 19061 55199 19119 55205
rect 19061 55196 19073 55199
rect 18104 55168 19073 55196
rect 18104 55156 18110 55168
rect 19061 55165 19073 55168
rect 19107 55165 19119 55199
rect 19061 55159 19119 55165
rect 19981 55199 20039 55205
rect 19981 55165 19993 55199
rect 20027 55196 20039 55199
rect 20622 55196 20628 55208
rect 20027 55168 20628 55196
rect 20027 55165 20039 55168
rect 19981 55159 20039 55165
rect 20622 55156 20628 55168
rect 20680 55156 20686 55208
rect 21269 55199 21327 55205
rect 21269 55165 21281 55199
rect 21315 55196 21327 55199
rect 22002 55196 22008 55208
rect 21315 55168 22008 55196
rect 21315 55165 21327 55168
rect 21269 55159 21327 55165
rect 22002 55156 22008 55168
rect 22060 55156 22066 55208
rect 22189 55199 22247 55205
rect 22189 55165 22201 55199
rect 22235 55165 22247 55199
rect 22189 55159 22247 55165
rect 22557 55199 22615 55205
rect 22557 55165 22569 55199
rect 22603 55196 22615 55199
rect 23106 55196 23112 55208
rect 22603 55168 23112 55196
rect 22603 55165 22615 55168
rect 22557 55159 22615 55165
rect 14476 55128 14504 55156
rect 13648 55100 14504 55128
rect 13262 55060 13268 55072
rect 13223 55032 13268 55060
rect 13262 55020 13268 55032
rect 13320 55020 13326 55072
rect 13648 55069 13676 55100
rect 17034 55088 17040 55140
rect 17092 55128 17098 55140
rect 17494 55128 17500 55140
rect 17092 55100 17500 55128
rect 17092 55088 17098 55100
rect 17494 55088 17500 55100
rect 17552 55128 17558 55140
rect 17681 55131 17739 55137
rect 17681 55128 17693 55131
rect 17552 55100 17693 55128
rect 17552 55088 17558 55100
rect 17681 55097 17693 55100
rect 17727 55128 17739 55131
rect 17773 55131 17831 55137
rect 17773 55128 17785 55131
rect 17727 55100 17785 55128
rect 17727 55097 17739 55100
rect 17681 55091 17739 55097
rect 17773 55097 17785 55100
rect 17819 55097 17831 55131
rect 18782 55128 18788 55140
rect 18743 55100 18788 55128
rect 17773 55091 17831 55097
rect 18782 55088 18788 55100
rect 18840 55088 18846 55140
rect 20073 55131 20131 55137
rect 20073 55097 20085 55131
rect 20119 55097 20131 55131
rect 22020 55128 22048 55156
rect 22204 55128 22232 55159
rect 23106 55156 23112 55168
rect 23164 55156 23170 55208
rect 24118 55156 24124 55208
rect 24176 55196 24182 55208
rect 24305 55199 24363 55205
rect 24305 55196 24317 55199
rect 24176 55168 24317 55196
rect 24176 55156 24182 55168
rect 24305 55165 24317 55168
rect 24351 55165 24363 55199
rect 24305 55159 24363 55165
rect 24397 55199 24455 55205
rect 24397 55165 24409 55199
rect 24443 55196 24455 55199
rect 24486 55196 24492 55208
rect 24443 55168 24492 55196
rect 24443 55165 24455 55168
rect 24397 55159 24455 55165
rect 24486 55156 24492 55168
rect 24544 55156 24550 55208
rect 25133 55199 25191 55205
rect 25133 55165 25145 55199
rect 25179 55165 25191 55199
rect 25133 55159 25191 55165
rect 26145 55199 26203 55205
rect 26145 55165 26157 55199
rect 26191 55196 26203 55199
rect 26234 55196 26240 55208
rect 26191 55168 26240 55196
rect 26191 55165 26203 55168
rect 26145 55159 26203 55165
rect 22020 55100 22232 55128
rect 20073 55091 20131 55097
rect 13633 55063 13691 55069
rect 13633 55029 13645 55063
rect 13679 55029 13691 55063
rect 13633 55023 13691 55029
rect 13998 55020 14004 55072
rect 14056 55060 14062 55072
rect 14185 55063 14243 55069
rect 14185 55060 14197 55063
rect 14056 55032 14197 55060
rect 14056 55020 14062 55032
rect 14185 55029 14197 55032
rect 14231 55029 14243 55063
rect 14185 55023 14243 55029
rect 15102 55020 15108 55072
rect 15160 55060 15166 55072
rect 15289 55063 15347 55069
rect 15289 55060 15301 55063
rect 15160 55032 15301 55060
rect 15160 55020 15166 55032
rect 15289 55029 15301 55032
rect 15335 55060 15347 55063
rect 15473 55063 15531 55069
rect 15473 55060 15485 55063
rect 15335 55032 15485 55060
rect 15335 55029 15347 55032
rect 15289 55023 15347 55029
rect 15473 55029 15485 55032
rect 15519 55029 15531 55063
rect 15930 55060 15936 55072
rect 15891 55032 15936 55060
rect 15473 55023 15531 55029
rect 15930 55020 15936 55032
rect 15988 55020 15994 55072
rect 18046 55020 18052 55072
rect 18104 55060 18110 55072
rect 19150 55060 19156 55072
rect 18104 55032 19156 55060
rect 18104 55020 18110 55032
rect 19150 55020 19156 55032
rect 19208 55020 19214 55072
rect 19978 55020 19984 55072
rect 20036 55060 20042 55072
rect 20088 55060 20116 55091
rect 24670 55088 24676 55140
rect 24728 55128 24734 55140
rect 25148 55128 25176 55159
rect 26234 55156 26240 55168
rect 26292 55156 26298 55208
rect 24728 55100 26096 55128
rect 24728 55088 24734 55100
rect 21634 55060 21640 55072
rect 20036 55032 20116 55060
rect 21595 55032 21640 55060
rect 20036 55020 20042 55032
rect 21634 55020 21640 55032
rect 21692 55020 21698 55072
rect 21910 55020 21916 55072
rect 21968 55060 21974 55072
rect 23477 55063 23535 55069
rect 23477 55060 23489 55063
rect 21968 55032 23489 55060
rect 21968 55020 21974 55032
rect 23477 55029 23489 55032
rect 23523 55060 23535 55063
rect 24026 55060 24032 55072
rect 23523 55032 24032 55060
rect 23523 55029 23535 55032
rect 23477 55023 23535 55029
rect 24026 55020 24032 55032
rect 24084 55020 24090 55072
rect 26068 55060 26096 55100
rect 27709 55063 27767 55069
rect 27709 55060 27721 55063
rect 26068 55032 27721 55060
rect 27709 55029 27721 55032
rect 27755 55029 27767 55063
rect 27709 55023 27767 55029
rect 1104 54970 28888 54992
rect 1104 54918 10982 54970
rect 11034 54918 11046 54970
rect 11098 54918 11110 54970
rect 11162 54918 11174 54970
rect 11226 54918 20982 54970
rect 21034 54918 21046 54970
rect 21098 54918 21110 54970
rect 21162 54918 21174 54970
rect 21226 54918 28888 54970
rect 1104 54896 28888 54918
rect 14093 54859 14151 54865
rect 14093 54825 14105 54859
rect 14139 54856 14151 54859
rect 14458 54856 14464 54868
rect 14139 54828 14464 54856
rect 14139 54825 14151 54828
rect 14093 54819 14151 54825
rect 14458 54816 14464 54828
rect 14516 54816 14522 54868
rect 15286 54816 15292 54868
rect 15344 54856 15350 54868
rect 15562 54856 15568 54868
rect 15344 54828 15568 54856
rect 15344 54816 15350 54828
rect 15562 54816 15568 54828
rect 15620 54816 15626 54868
rect 17126 54856 17132 54868
rect 15672 54828 17132 54856
rect 12066 54788 12072 54800
rect 11979 54760 12072 54788
rect 12066 54748 12072 54760
rect 12124 54788 12130 54800
rect 12713 54791 12771 54797
rect 12713 54788 12725 54791
rect 12124 54760 12725 54788
rect 12124 54748 12130 54760
rect 12713 54757 12725 54760
rect 12759 54788 12771 54791
rect 12759 54760 14228 54788
rect 12759 54757 12771 54760
rect 12713 54751 12771 54757
rect 12161 54723 12219 54729
rect 12161 54689 12173 54723
rect 12207 54720 12219 54723
rect 12250 54720 12256 54732
rect 12207 54692 12256 54720
rect 12207 54689 12219 54692
rect 12161 54683 12219 54689
rect 12250 54680 12256 54692
rect 12308 54680 12314 54732
rect 13173 54723 13231 54729
rect 13173 54689 13185 54723
rect 13219 54720 13231 54723
rect 13814 54720 13820 54732
rect 13219 54692 13820 54720
rect 13219 54689 13231 54692
rect 13173 54683 13231 54689
rect 13814 54680 13820 54692
rect 13872 54680 13878 54732
rect 14200 54729 14228 54760
rect 14642 54748 14648 54800
rect 14700 54788 14706 54800
rect 15010 54788 15016 54800
rect 14700 54760 15016 54788
rect 14700 54748 14706 54760
rect 15010 54748 15016 54760
rect 15068 54788 15074 54800
rect 15105 54791 15163 54797
rect 15105 54788 15117 54791
rect 15068 54760 15117 54788
rect 15068 54748 15074 54760
rect 15105 54757 15117 54760
rect 15151 54788 15163 54791
rect 15381 54791 15439 54797
rect 15381 54788 15393 54791
rect 15151 54760 15393 54788
rect 15151 54757 15163 54760
rect 15105 54751 15163 54757
rect 15381 54757 15393 54760
rect 15427 54788 15439 54791
rect 15672 54788 15700 54828
rect 17126 54816 17132 54828
rect 17184 54816 17190 54868
rect 17586 54816 17592 54868
rect 17644 54856 17650 54868
rect 18141 54859 18199 54865
rect 18141 54856 18153 54859
rect 17644 54828 18153 54856
rect 17644 54816 17650 54828
rect 18141 54825 18153 54828
rect 18187 54825 18199 54859
rect 19334 54856 19340 54868
rect 19295 54828 19340 54856
rect 18141 54819 18199 54825
rect 19334 54816 19340 54828
rect 19392 54816 19398 54868
rect 19610 54856 19616 54868
rect 19571 54828 19616 54856
rect 19610 54816 19616 54828
rect 19668 54816 19674 54868
rect 20162 54816 20168 54868
rect 20220 54856 20226 54868
rect 20717 54859 20775 54865
rect 20717 54856 20729 54859
rect 20220 54828 20729 54856
rect 20220 54816 20226 54828
rect 20717 54825 20729 54828
rect 20763 54856 20775 54859
rect 21818 54856 21824 54868
rect 20763 54828 21824 54856
rect 20763 54825 20775 54828
rect 20717 54819 20775 54825
rect 21818 54816 21824 54828
rect 21876 54816 21882 54868
rect 22370 54856 22376 54868
rect 22331 54828 22376 54856
rect 22370 54816 22376 54828
rect 22428 54816 22434 54868
rect 24118 54816 24124 54868
rect 24176 54856 24182 54868
rect 24213 54859 24271 54865
rect 24213 54856 24225 54859
rect 24176 54828 24225 54856
rect 24176 54816 24182 54828
rect 24213 54825 24225 54828
rect 24259 54825 24271 54859
rect 24670 54856 24676 54868
rect 24631 54828 24676 54856
rect 24213 54819 24271 54825
rect 24670 54816 24676 54828
rect 24728 54816 24734 54868
rect 16666 54788 16672 54800
rect 15427 54760 15700 54788
rect 16627 54760 16672 54788
rect 15427 54757 15439 54760
rect 15381 54751 15439 54757
rect 16666 54748 16672 54760
rect 16724 54788 16730 54800
rect 16850 54788 16856 54800
rect 16724 54760 16856 54788
rect 16724 54748 16730 54760
rect 16850 54748 16856 54760
rect 16908 54748 16914 54800
rect 17678 54748 17684 54800
rect 17736 54788 17742 54800
rect 18233 54791 18291 54797
rect 18233 54788 18245 54791
rect 17736 54760 18245 54788
rect 17736 54748 17742 54760
rect 18233 54757 18245 54760
rect 18279 54757 18291 54791
rect 18233 54751 18291 54757
rect 23017 54791 23075 54797
rect 23017 54757 23029 54791
rect 23063 54788 23075 54791
rect 23198 54788 23204 54800
rect 23063 54760 23204 54788
rect 23063 54757 23075 54760
rect 23017 54751 23075 54757
rect 23198 54748 23204 54760
rect 23256 54748 23262 54800
rect 24762 54788 24768 54800
rect 23768 54760 24768 54788
rect 14185 54723 14243 54729
rect 14185 54689 14197 54723
rect 14231 54720 14243 54723
rect 14826 54720 14832 54732
rect 14231 54692 14832 54720
rect 14231 54689 14243 54692
rect 14185 54683 14243 54689
rect 14826 54680 14832 54692
rect 14884 54680 14890 54732
rect 15286 54680 15292 54732
rect 15344 54720 15350 54732
rect 15657 54723 15715 54729
rect 15657 54720 15669 54723
rect 15344 54692 15669 54720
rect 15344 54680 15350 54692
rect 15657 54689 15669 54692
rect 15703 54689 15715 54723
rect 18049 54723 18107 54729
rect 18049 54720 18061 54723
rect 15657 54683 15715 54689
rect 17696 54692 18061 54720
rect 14645 54655 14703 54661
rect 14645 54652 14657 54655
rect 13372 54624 14657 54652
rect 11974 54544 11980 54596
rect 12032 54584 12038 54596
rect 12989 54587 13047 54593
rect 12989 54584 13001 54587
rect 12032 54556 13001 54584
rect 12032 54544 12038 54556
rect 12989 54553 13001 54556
rect 13035 54584 13047 54587
rect 13078 54584 13084 54596
rect 13035 54556 13084 54584
rect 13035 54553 13047 54556
rect 12989 54547 13047 54553
rect 13078 54544 13084 54556
rect 13136 54544 13142 54596
rect 13372 54593 13400 54624
rect 14645 54621 14657 54624
rect 14691 54652 14703 54655
rect 14734 54652 14740 54664
rect 14691 54624 14740 54652
rect 14691 54621 14703 54624
rect 14645 54615 14703 54621
rect 14734 54612 14740 54624
rect 14792 54612 14798 54664
rect 15194 54612 15200 54664
rect 15252 54652 15258 54664
rect 16025 54655 16083 54661
rect 16025 54652 16037 54655
rect 15252 54624 16037 54652
rect 15252 54612 15258 54624
rect 16025 54621 16037 54624
rect 16071 54621 16083 54655
rect 16025 54615 16083 54621
rect 16298 54612 16304 54664
rect 16356 54652 16362 54664
rect 16482 54652 16488 54664
rect 16356 54624 16488 54652
rect 16356 54612 16362 54624
rect 16482 54612 16488 54624
rect 16540 54612 16546 54664
rect 17494 54612 17500 54664
rect 17552 54652 17558 54664
rect 17696 54661 17724 54692
rect 18049 54689 18061 54692
rect 18095 54689 18107 54723
rect 18049 54683 18107 54689
rect 17681 54655 17739 54661
rect 17681 54652 17693 54655
rect 17552 54624 17693 54652
rect 17552 54612 17558 54624
rect 17681 54621 17693 54624
rect 17727 54621 17739 54655
rect 17681 54615 17739 54621
rect 17865 54655 17923 54661
rect 17865 54621 17877 54655
rect 17911 54652 17923 54655
rect 17954 54652 17960 54664
rect 17911 54624 17960 54652
rect 17911 54621 17923 54624
rect 17865 54615 17923 54621
rect 17954 54612 17960 54624
rect 18012 54612 18018 54664
rect 18064 54652 18092 54683
rect 18782 54680 18788 54732
rect 18840 54720 18846 54732
rect 19429 54723 19487 54729
rect 19429 54720 19441 54723
rect 18840 54692 19441 54720
rect 18840 54680 18846 54692
rect 19429 54689 19441 54692
rect 19475 54720 19487 54723
rect 19889 54723 19947 54729
rect 19889 54720 19901 54723
rect 19475 54692 19901 54720
rect 19475 54689 19487 54692
rect 19429 54683 19487 54689
rect 19889 54689 19901 54692
rect 19935 54689 19947 54723
rect 21082 54720 21088 54732
rect 21043 54692 21088 54720
rect 19889 54683 19947 54689
rect 21082 54680 21088 54692
rect 21140 54680 21146 54732
rect 21818 54720 21824 54732
rect 21779 54692 21824 54720
rect 21818 54680 21824 54692
rect 21876 54680 21882 54732
rect 21910 54680 21916 54732
rect 21968 54720 21974 54732
rect 23768 54729 23796 54760
rect 24762 54748 24768 54760
rect 24820 54748 24826 54800
rect 22741 54723 22799 54729
rect 21968 54692 22013 54720
rect 21968 54680 21974 54692
rect 22741 54689 22753 54723
rect 22787 54720 22799 54723
rect 23753 54723 23811 54729
rect 23753 54720 23765 54723
rect 22787 54692 23765 54720
rect 22787 54689 22799 54692
rect 22741 54683 22799 54689
rect 23753 54689 23765 54692
rect 23799 54689 23811 54723
rect 23753 54683 23811 54689
rect 24210 54680 24216 54732
rect 24268 54720 24274 54732
rect 24670 54720 24676 54732
rect 24268 54692 24676 54720
rect 24268 54680 24274 54692
rect 24670 54680 24676 54692
rect 24728 54680 24734 54732
rect 27433 54723 27491 54729
rect 27433 54689 27445 54723
rect 27479 54720 27491 54723
rect 27706 54720 27712 54732
rect 27479 54692 27712 54720
rect 27479 54689 27491 54692
rect 27433 54683 27491 54689
rect 27706 54680 27712 54692
rect 27764 54680 27770 54732
rect 18230 54652 18236 54664
rect 18064 54624 18236 54652
rect 18230 54612 18236 54624
rect 18288 54612 18294 54664
rect 18601 54655 18659 54661
rect 18601 54621 18613 54655
rect 18647 54652 18659 54655
rect 19150 54652 19156 54664
rect 18647 54624 19156 54652
rect 18647 54621 18659 54624
rect 18601 54615 18659 54621
rect 19150 54612 19156 54624
rect 19208 54612 19214 54664
rect 20714 54612 20720 54664
rect 20772 54652 20778 54664
rect 20993 54655 21051 54661
rect 20993 54652 21005 54655
rect 20772 54624 21005 54652
rect 20772 54612 20778 54624
rect 20993 54621 21005 54624
rect 21039 54652 21051 54655
rect 21358 54652 21364 54664
rect 21039 54624 21364 54652
rect 21039 54621 21051 54624
rect 20993 54615 21051 54621
rect 21358 54612 21364 54624
rect 21416 54612 21422 54664
rect 22925 54655 22983 54661
rect 22925 54621 22937 54655
rect 22971 54652 22983 54655
rect 23106 54652 23112 54664
rect 22971 54624 23112 54652
rect 22971 54621 22983 54624
rect 22925 54615 22983 54621
rect 23106 54612 23112 54624
rect 23164 54612 23170 54664
rect 23566 54612 23572 54664
rect 23624 54652 23630 54664
rect 23845 54655 23903 54661
rect 23845 54652 23857 54655
rect 23624 54624 23857 54652
rect 23624 54612 23630 54624
rect 23845 54621 23857 54624
rect 23891 54621 23903 54655
rect 26602 54652 26608 54664
rect 26563 54624 26608 54652
rect 23845 54615 23903 54621
rect 26602 54612 26608 54624
rect 26660 54612 26666 54664
rect 26697 54655 26755 54661
rect 26697 54621 26709 54655
rect 26743 54652 26755 54655
rect 26970 54652 26976 54664
rect 26743 54624 26976 54652
rect 26743 54621 26755 54624
rect 26697 54615 26755 54621
rect 26970 54612 26976 54624
rect 27028 54612 27034 54664
rect 27522 54652 27528 54664
rect 27483 54624 27528 54652
rect 27522 54612 27528 54624
rect 27580 54612 27586 54664
rect 13357 54587 13415 54593
rect 13357 54553 13369 54587
rect 13403 54553 13415 54587
rect 13357 54547 13415 54553
rect 14369 54587 14427 54593
rect 14369 54553 14381 54587
rect 14415 54584 14427 54587
rect 14918 54584 14924 54596
rect 14415 54556 14924 54584
rect 14415 54553 14427 54556
rect 14369 54547 14427 54553
rect 14918 54544 14924 54556
rect 14976 54544 14982 54596
rect 15381 54587 15439 54593
rect 15381 54553 15393 54587
rect 15427 54584 15439 54587
rect 15930 54584 15936 54596
rect 15427 54556 15608 54584
rect 15843 54556 15936 54584
rect 15427 54553 15439 54556
rect 15381 54547 15439 54553
rect 12342 54516 12348 54528
rect 12303 54488 12348 54516
rect 12342 54476 12348 54488
rect 12400 54476 12406 54528
rect 13725 54519 13783 54525
rect 13725 54485 13737 54519
rect 13771 54516 13783 54519
rect 13906 54516 13912 54528
rect 13771 54488 13912 54516
rect 13771 54485 13783 54488
rect 13725 54479 13783 54485
rect 13906 54476 13912 54488
rect 13964 54476 13970 54528
rect 15102 54476 15108 54528
rect 15160 54516 15166 54528
rect 15473 54519 15531 54525
rect 15473 54516 15485 54519
rect 15160 54488 15485 54516
rect 15160 54476 15166 54488
rect 15473 54485 15485 54488
rect 15519 54485 15531 54519
rect 15580 54516 15608 54556
rect 15930 54544 15936 54556
rect 15988 54584 15994 54596
rect 16666 54584 16672 54596
rect 15988 54556 16672 54584
rect 15988 54544 15994 54556
rect 16666 54544 16672 54556
rect 16724 54544 16730 54596
rect 18248 54584 18276 54612
rect 18877 54587 18935 54593
rect 18877 54584 18889 54587
rect 18248 54556 18889 54584
rect 18877 54553 18889 54556
rect 18923 54553 18935 54587
rect 18877 54547 18935 54553
rect 15795 54519 15853 54525
rect 15795 54516 15807 54519
rect 15580 54488 15807 54516
rect 15473 54479 15531 54485
rect 15795 54485 15807 54488
rect 15841 54485 15853 54519
rect 16298 54516 16304 54528
rect 16259 54488 16304 54516
rect 15795 54479 15853 54485
rect 16298 54476 16304 54488
rect 16356 54476 16362 54528
rect 20346 54516 20352 54528
rect 20307 54488 20352 54516
rect 20346 54476 20352 54488
rect 20404 54476 20410 54528
rect 26237 54519 26295 54525
rect 26237 54485 26249 54519
rect 26283 54516 26295 54519
rect 26326 54516 26332 54528
rect 26283 54488 26332 54516
rect 26283 54485 26295 54488
rect 26237 54479 26295 54485
rect 26326 54476 26332 54488
rect 26384 54476 26390 54528
rect 1104 54426 28888 54448
rect 1104 54374 5982 54426
rect 6034 54374 6046 54426
rect 6098 54374 6110 54426
rect 6162 54374 6174 54426
rect 6226 54374 15982 54426
rect 16034 54374 16046 54426
rect 16098 54374 16110 54426
rect 16162 54374 16174 54426
rect 16226 54374 25982 54426
rect 26034 54374 26046 54426
rect 26098 54374 26110 54426
rect 26162 54374 26174 54426
rect 26226 54374 28888 54426
rect 1104 54352 28888 54374
rect 12250 54312 12256 54324
rect 12211 54284 12256 54312
rect 12250 54272 12256 54284
rect 12308 54272 12314 54324
rect 13814 54272 13820 54324
rect 13872 54312 13878 54324
rect 15841 54315 15899 54321
rect 15841 54312 15853 54315
rect 13872 54284 15853 54312
rect 13872 54272 13878 54284
rect 15841 54281 15853 54284
rect 15887 54281 15899 54315
rect 16574 54312 16580 54324
rect 16535 54284 16580 54312
rect 15841 54275 15899 54281
rect 16574 54272 16580 54284
rect 16632 54272 16638 54324
rect 18506 54312 18512 54324
rect 18467 54284 18512 54312
rect 18506 54272 18512 54284
rect 18564 54272 18570 54324
rect 19334 54272 19340 54324
rect 19392 54312 19398 54324
rect 19521 54315 19579 54321
rect 19521 54312 19533 54315
rect 19392 54284 19533 54312
rect 19392 54272 19398 54284
rect 19521 54281 19533 54284
rect 19567 54281 19579 54315
rect 19521 54275 19579 54281
rect 20901 54315 20959 54321
rect 20901 54281 20913 54315
rect 20947 54312 20959 54315
rect 21910 54312 21916 54324
rect 20947 54284 21916 54312
rect 20947 54281 20959 54284
rect 20901 54275 20959 54281
rect 11882 54176 11888 54188
rect 11348 54148 11888 54176
rect 11348 54117 11376 54148
rect 11882 54136 11888 54148
rect 11940 54136 11946 54188
rect 12268 54176 12296 54272
rect 13173 54247 13231 54253
rect 13173 54213 13185 54247
rect 13219 54244 13231 54247
rect 15102 54244 15108 54256
rect 13219 54216 15108 54244
rect 13219 54213 13231 54216
rect 13173 54207 13231 54213
rect 15102 54204 15108 54216
rect 15160 54204 15166 54256
rect 16022 54244 16028 54256
rect 15983 54216 16028 54244
rect 16022 54204 16028 54216
rect 16080 54204 16086 54256
rect 12897 54179 12955 54185
rect 12897 54176 12909 54179
rect 12268 54148 12909 54176
rect 12897 54145 12909 54148
rect 12943 54176 12955 54179
rect 15933 54179 15991 54185
rect 15933 54176 15945 54179
rect 12943 54148 13952 54176
rect 12943 54145 12955 54148
rect 12897 54139 12955 54145
rect 13924 54120 13952 54148
rect 14660 54148 15945 54176
rect 11333 54111 11391 54117
rect 11333 54077 11345 54111
rect 11379 54077 11391 54111
rect 11333 54071 11391 54077
rect 12342 54068 12348 54120
rect 12400 54108 12406 54120
rect 12989 54111 13047 54117
rect 12989 54108 13001 54111
rect 12400 54080 13001 54108
rect 12400 54068 12406 54080
rect 12989 54077 13001 54080
rect 13035 54108 13047 54111
rect 13446 54108 13452 54120
rect 13035 54080 13452 54108
rect 13035 54077 13047 54080
rect 12989 54071 13047 54077
rect 13446 54068 13452 54080
rect 13504 54068 13510 54120
rect 13906 54068 13912 54120
rect 13964 54108 13970 54120
rect 14660 54117 14688 54148
rect 15933 54145 15945 54148
rect 15979 54145 15991 54179
rect 15933 54139 15991 54145
rect 17129 54179 17187 54185
rect 17129 54145 17141 54179
rect 17175 54176 17187 54179
rect 17954 54176 17960 54188
rect 17175 54148 17960 54176
rect 17175 54145 17187 54148
rect 17129 54139 17187 54145
rect 17954 54136 17960 54148
rect 18012 54176 18018 54188
rect 18049 54179 18107 54185
rect 18049 54176 18061 54179
rect 18012 54148 18061 54176
rect 18012 54136 18018 54148
rect 18049 54145 18061 54148
rect 18095 54176 18107 54179
rect 18782 54176 18788 54188
rect 18095 54148 18788 54176
rect 18095 54145 18107 54148
rect 18049 54139 18107 54145
rect 18782 54136 18788 54148
rect 18840 54136 18846 54188
rect 14645 54111 14703 54117
rect 14645 54108 14657 54111
rect 13964 54080 14657 54108
rect 13964 54068 13970 54080
rect 14645 54077 14657 54080
rect 14691 54077 14703 54111
rect 14645 54071 14703 54077
rect 14826 54068 14832 54120
rect 14884 54108 14890 54120
rect 15712 54111 15770 54117
rect 14884 54080 15608 54108
rect 14884 54068 14890 54080
rect 13998 54040 14004 54052
rect 13959 54012 14004 54040
rect 13998 54000 14004 54012
rect 14056 54000 14062 54052
rect 15010 54040 15016 54052
rect 14971 54012 15016 54040
rect 15010 54000 15016 54012
rect 15068 54000 15074 54052
rect 15194 54000 15200 54052
rect 15252 54040 15258 54052
rect 15580 54049 15608 54080
rect 15712 54077 15724 54111
rect 15758 54108 15770 54111
rect 16114 54108 16120 54120
rect 15758 54080 16120 54108
rect 15758 54077 15770 54080
rect 15712 54071 15770 54077
rect 16114 54068 16120 54080
rect 16172 54068 16178 54120
rect 18325 54111 18383 54117
rect 18325 54108 18337 54111
rect 17420 54080 18337 54108
rect 15381 54043 15439 54049
rect 15381 54040 15393 54043
rect 15252 54012 15393 54040
rect 15252 54000 15258 54012
rect 15381 54009 15393 54012
rect 15427 54009 15439 54043
rect 15381 54003 15439 54009
rect 15565 54043 15623 54049
rect 15565 54009 15577 54043
rect 15611 54040 15623 54043
rect 16206 54040 16212 54052
rect 15611 54012 16212 54040
rect 15611 54009 15623 54012
rect 15565 54003 15623 54009
rect 16206 54000 16212 54012
rect 16264 54000 16270 54052
rect 11514 53972 11520 53984
rect 11475 53944 11520 53972
rect 11514 53932 11520 53944
rect 11572 53932 11578 53984
rect 13814 53972 13820 53984
rect 13775 53944 13820 53972
rect 13814 53932 13820 53944
rect 13872 53932 13878 53984
rect 16850 53932 16856 53984
rect 16908 53972 16914 53984
rect 17420 53981 17448 54080
rect 18325 54077 18337 54080
rect 18371 54077 18383 54111
rect 19536 54108 19564 54275
rect 21910 54272 21916 54284
rect 21968 54272 21974 54324
rect 27706 54272 27712 54324
rect 27764 54312 27770 54324
rect 27893 54315 27951 54321
rect 27893 54312 27905 54315
rect 27764 54284 27905 54312
rect 27764 54272 27770 54284
rect 27893 54281 27905 54284
rect 27939 54281 27951 54315
rect 27893 54275 27951 54281
rect 22005 54247 22063 54253
rect 22005 54213 22017 54247
rect 22051 54213 22063 54247
rect 22005 54207 22063 54213
rect 22020 54176 22048 54207
rect 25866 54176 25872 54188
rect 22020 54148 24164 54176
rect 25827 54148 25872 54176
rect 19797 54111 19855 54117
rect 19797 54108 19809 54111
rect 19536 54080 19809 54108
rect 18325 54071 18383 54077
rect 19797 54077 19809 54080
rect 19843 54077 19855 54111
rect 19797 54071 19855 54077
rect 21269 54111 21327 54117
rect 21269 54077 21281 54111
rect 21315 54108 21327 54111
rect 22186 54108 22192 54120
rect 21315 54080 22192 54108
rect 21315 54077 21327 54080
rect 21269 54071 21327 54077
rect 22186 54068 22192 54080
rect 22244 54068 22250 54120
rect 22370 54068 22376 54120
rect 22428 54108 22434 54120
rect 22511 54111 22569 54117
rect 22511 54108 22523 54111
rect 22428 54080 22523 54108
rect 22428 54068 22434 54080
rect 22511 54077 22523 54080
rect 22557 54077 22569 54111
rect 22646 54108 22652 54120
rect 22607 54080 22652 54108
rect 22511 54071 22569 54077
rect 22646 54068 22652 54080
rect 22704 54068 22710 54120
rect 23017 54111 23075 54117
rect 23017 54077 23029 54111
rect 23063 54108 23075 54111
rect 23566 54108 23572 54120
rect 23063 54080 23572 54108
rect 23063 54077 23075 54080
rect 23017 54071 23075 54077
rect 23566 54068 23572 54080
rect 23624 54068 23630 54120
rect 23658 54068 23664 54120
rect 23716 54108 23722 54120
rect 24136 54117 24164 54148
rect 25866 54136 25872 54148
rect 25924 54176 25930 54188
rect 26237 54179 26295 54185
rect 26237 54176 26249 54179
rect 25924 54148 26249 54176
rect 25924 54136 25930 54148
rect 26237 54145 26249 54148
rect 26283 54145 26295 54179
rect 26237 54139 26295 54145
rect 24121 54111 24179 54117
rect 23716 54080 23761 54108
rect 23716 54068 23722 54080
rect 24121 54077 24133 54111
rect 24167 54108 24179 54111
rect 24673 54111 24731 54117
rect 24673 54108 24685 54111
rect 24167 54080 24685 54108
rect 24167 54077 24179 54080
rect 24121 54071 24179 54077
rect 24673 54077 24685 54080
rect 24719 54077 24731 54111
rect 25958 54108 25964 54120
rect 25919 54080 25964 54108
rect 24673 54071 24731 54077
rect 25958 54068 25964 54080
rect 26016 54108 26022 54120
rect 26326 54108 26332 54120
rect 26016 54080 26332 54108
rect 26016 54068 26022 54080
rect 26326 54068 26332 54080
rect 26384 54068 26390 54120
rect 18230 54000 18236 54052
rect 18288 54040 18294 54052
rect 18288 54012 18333 54040
rect 18288 54000 18294 54012
rect 19334 54000 19340 54052
rect 19392 54040 19398 54052
rect 19702 54040 19708 54052
rect 19392 54012 19708 54040
rect 19392 54000 19398 54012
rect 19702 54000 19708 54012
rect 19760 54000 19766 54052
rect 20441 54043 20499 54049
rect 20441 54009 20453 54043
rect 20487 54040 20499 54043
rect 20622 54040 20628 54052
rect 20487 54012 20628 54040
rect 20487 54009 20499 54012
rect 20441 54003 20499 54009
rect 20622 54000 20628 54012
rect 20680 54000 20686 54052
rect 21637 54043 21695 54049
rect 21637 54009 21649 54043
rect 21683 54040 21695 54043
rect 22664 54040 22692 54068
rect 21683 54012 22692 54040
rect 21683 54009 21695 54012
rect 21637 54003 21695 54009
rect 23106 54000 23112 54052
rect 23164 54040 23170 54052
rect 23164 54012 23796 54040
rect 23164 54000 23170 54012
rect 17405 53975 17463 53981
rect 17405 53972 17417 53975
rect 16908 53944 17417 53972
rect 16908 53932 16914 53944
rect 17405 53941 17417 53944
rect 17451 53941 17463 53975
rect 17405 53935 17463 53941
rect 17678 53932 17684 53984
rect 17736 53972 17742 53984
rect 17773 53975 17831 53981
rect 17773 53972 17785 53975
rect 17736 53944 17785 53972
rect 17736 53932 17742 53944
rect 17773 53941 17785 53944
rect 17819 53941 17831 53975
rect 17773 53935 17831 53941
rect 18782 53932 18788 53984
rect 18840 53972 18846 53984
rect 19061 53975 19119 53981
rect 19061 53972 19073 53975
rect 18840 53944 19073 53972
rect 18840 53932 18846 53944
rect 19061 53941 19073 53944
rect 19107 53941 19119 53975
rect 19061 53935 19119 53941
rect 22462 53932 22468 53984
rect 22520 53972 22526 53984
rect 23014 53972 23020 53984
rect 22520 53944 23020 53972
rect 22520 53932 22526 53944
rect 23014 53932 23020 53944
rect 23072 53972 23078 53984
rect 23477 53975 23535 53981
rect 23477 53972 23489 53975
rect 23072 53944 23489 53972
rect 23072 53932 23078 53944
rect 23477 53941 23489 53944
rect 23523 53972 23535 53975
rect 23658 53972 23664 53984
rect 23523 53944 23664 53972
rect 23523 53941 23535 53944
rect 23477 53935 23535 53941
rect 23658 53932 23664 53944
rect 23716 53932 23722 53984
rect 23768 53981 23796 54012
rect 23753 53975 23811 53981
rect 23753 53941 23765 53975
rect 23799 53941 23811 53975
rect 27338 53972 27344 53984
rect 27299 53944 27344 53972
rect 23753 53935 23811 53941
rect 27338 53932 27344 53944
rect 27396 53932 27402 53984
rect 1104 53882 28888 53904
rect 1104 53830 10982 53882
rect 11034 53830 11046 53882
rect 11098 53830 11110 53882
rect 11162 53830 11174 53882
rect 11226 53830 20982 53882
rect 21034 53830 21046 53882
rect 21098 53830 21110 53882
rect 21162 53830 21174 53882
rect 21226 53830 28888 53882
rect 1104 53808 28888 53830
rect 11793 53771 11851 53777
rect 11793 53737 11805 53771
rect 11839 53768 11851 53771
rect 12066 53768 12072 53780
rect 11839 53740 12072 53768
rect 11839 53737 11851 53740
rect 11793 53731 11851 53737
rect 12066 53728 12072 53740
rect 12124 53728 12130 53780
rect 18049 53771 18107 53777
rect 18049 53737 18061 53771
rect 18095 53768 18107 53771
rect 18138 53768 18144 53780
rect 18095 53740 18144 53768
rect 18095 53737 18107 53740
rect 18049 53731 18107 53737
rect 18138 53728 18144 53740
rect 18196 53728 18202 53780
rect 18690 53768 18696 53780
rect 18432 53740 18696 53768
rect 13906 53700 13912 53712
rect 13867 53672 13912 53700
rect 13906 53660 13912 53672
rect 13964 53660 13970 53712
rect 16945 53703 17003 53709
rect 16945 53669 16957 53703
rect 16991 53700 17003 53703
rect 17770 53700 17776 53712
rect 16991 53672 17776 53700
rect 16991 53669 17003 53672
rect 16945 53663 17003 53669
rect 17770 53660 17776 53672
rect 17828 53660 17834 53712
rect 11238 53632 11244 53644
rect 11199 53604 11244 53632
rect 11238 53592 11244 53604
rect 11296 53592 11302 53644
rect 12066 53592 12072 53644
rect 12124 53632 12130 53644
rect 12529 53635 12587 53641
rect 12529 53632 12541 53635
rect 12124 53604 12541 53632
rect 12124 53592 12130 53604
rect 12529 53601 12541 53604
rect 12575 53601 12587 53635
rect 16206 53632 16212 53644
rect 16119 53604 16212 53632
rect 12529 53595 12587 53601
rect 16206 53592 16212 53604
rect 16264 53632 16270 53644
rect 18046 53632 18052 53644
rect 16264 53604 16988 53632
rect 18007 53604 18052 53632
rect 16264 53592 16270 53604
rect 16960 53576 16988 53604
rect 18046 53592 18052 53604
rect 18104 53592 18110 53644
rect 18230 53632 18236 53644
rect 18191 53604 18236 53632
rect 18230 53592 18236 53604
rect 18288 53592 18294 53644
rect 12253 53567 12311 53573
rect 12253 53533 12265 53567
rect 12299 53564 12311 53567
rect 12434 53564 12440 53576
rect 12299 53536 12440 53564
rect 12299 53533 12311 53536
rect 12253 53527 12311 53533
rect 12434 53524 12440 53536
rect 12492 53524 12498 53576
rect 15194 53524 15200 53576
rect 15252 53564 15258 53576
rect 16577 53567 16635 53573
rect 16577 53564 16589 53567
rect 15252 53536 16589 53564
rect 15252 53524 15258 53536
rect 16577 53533 16589 53536
rect 16623 53533 16635 53567
rect 16577 53527 16635 53533
rect 16942 53524 16948 53576
rect 17000 53524 17006 53576
rect 17310 53524 17316 53576
rect 17368 53564 17374 53576
rect 17586 53564 17592 53576
rect 17368 53536 17592 53564
rect 17368 53524 17374 53536
rect 17586 53524 17592 53536
rect 17644 53524 17650 53576
rect 18138 53524 18144 53576
rect 18196 53564 18202 53576
rect 18432 53564 18460 53740
rect 18690 53728 18696 53740
rect 18748 53728 18754 53780
rect 19150 53728 19156 53780
rect 19208 53768 19214 53780
rect 20257 53771 20315 53777
rect 20257 53768 20269 53771
rect 19208 53740 20269 53768
rect 19208 53728 19214 53740
rect 20257 53737 20269 53740
rect 20303 53737 20315 53771
rect 20714 53768 20720 53780
rect 20675 53740 20720 53768
rect 20257 53731 20315 53737
rect 19245 53703 19303 53709
rect 19245 53669 19257 53703
rect 19291 53700 19303 53703
rect 19610 53700 19616 53712
rect 19291 53672 19616 53700
rect 19291 53669 19303 53672
rect 19245 53663 19303 53669
rect 19610 53660 19616 53672
rect 19668 53660 19674 53712
rect 20272 53700 20300 53731
rect 20714 53728 20720 53740
rect 20772 53728 20778 53780
rect 21818 53728 21824 53780
rect 21876 53768 21882 53780
rect 21913 53771 21971 53777
rect 21913 53768 21925 53771
rect 21876 53740 21925 53768
rect 21876 53728 21882 53740
rect 21913 53737 21925 53740
rect 21959 53737 21971 53771
rect 22370 53768 22376 53780
rect 22331 53740 22376 53768
rect 21913 53731 21971 53737
rect 22370 53728 22376 53740
rect 22428 53728 22434 53780
rect 23934 53728 23940 53780
rect 23992 53728 23998 53780
rect 26602 53728 26608 53780
rect 26660 53768 26666 53780
rect 26697 53771 26755 53777
rect 26697 53768 26709 53771
rect 26660 53740 26709 53768
rect 26660 53728 26666 53740
rect 26697 53737 26709 53740
rect 26743 53737 26755 53771
rect 26697 53731 26755 53737
rect 23952 53700 23980 53728
rect 27065 53703 27123 53709
rect 27065 53700 27077 53703
rect 20272 53672 21036 53700
rect 23952 53672 27077 53700
rect 18601 53635 18659 53641
rect 18601 53601 18613 53635
rect 18647 53632 18659 53635
rect 18690 53632 18696 53644
rect 18647 53604 18696 53632
rect 18647 53601 18659 53604
rect 18601 53595 18659 53601
rect 18690 53592 18696 53604
rect 18748 53592 18754 53644
rect 19426 53592 19432 53644
rect 19484 53632 19490 53644
rect 19521 53635 19579 53641
rect 19521 53632 19533 53635
rect 19484 53604 19533 53632
rect 19484 53592 19490 53604
rect 19521 53601 19533 53604
rect 19567 53601 19579 53635
rect 19702 53632 19708 53644
rect 19663 53604 19708 53632
rect 19521 53595 19579 53601
rect 19702 53592 19708 53604
rect 19760 53592 19766 53644
rect 20162 53592 20168 53644
rect 20220 53632 20226 53644
rect 21008 53641 21036 53672
rect 20901 53635 20959 53641
rect 20901 53632 20913 53635
rect 20220 53604 20913 53632
rect 20220 53592 20226 53604
rect 20901 53601 20913 53604
rect 20947 53601 20959 53635
rect 20901 53595 20959 53601
rect 20993 53635 21051 53641
rect 20993 53601 21005 53635
rect 21039 53601 21051 53635
rect 20993 53595 21051 53601
rect 21082 53592 21088 53644
rect 21140 53632 21146 53644
rect 21177 53635 21235 53641
rect 21177 53632 21189 53635
rect 21140 53604 21189 53632
rect 21140 53592 21146 53604
rect 21177 53601 21189 53604
rect 21223 53601 21235 53635
rect 21177 53595 21235 53601
rect 22925 53635 22983 53641
rect 22925 53601 22937 53635
rect 22971 53632 22983 53635
rect 23106 53632 23112 53644
rect 22971 53604 23112 53632
rect 22971 53601 22983 53604
rect 22925 53595 22983 53601
rect 23106 53592 23112 53604
rect 23164 53592 23170 53644
rect 23934 53632 23940 53644
rect 23895 53604 23940 53632
rect 23934 53592 23940 53604
rect 23992 53592 23998 53644
rect 24044 53641 24072 53672
rect 27065 53669 27077 53672
rect 27111 53700 27123 53703
rect 27522 53700 27528 53712
rect 27111 53672 27528 53700
rect 27111 53669 27123 53672
rect 27065 53663 27123 53669
rect 27522 53660 27528 53672
rect 27580 53660 27586 53712
rect 24029 53635 24087 53641
rect 24029 53601 24041 53635
rect 24075 53601 24087 53635
rect 24029 53595 24087 53601
rect 21358 53564 21364 53576
rect 18196 53536 18460 53564
rect 21319 53536 21364 53564
rect 18196 53524 18202 53536
rect 21358 53524 21364 53536
rect 21416 53524 21422 53576
rect 22370 53524 22376 53576
rect 22428 53564 22434 53576
rect 23201 53567 23259 53573
rect 23201 53564 23213 53567
rect 22428 53536 23213 53564
rect 22428 53524 22434 53536
rect 23201 53533 23213 53536
rect 23247 53533 23259 53567
rect 25958 53564 25964 53576
rect 23201 53527 23259 53533
rect 24780 53536 25964 53564
rect 15286 53456 15292 53508
rect 15344 53496 15350 53508
rect 16025 53499 16083 53505
rect 16025 53496 16037 53499
rect 15344 53468 16037 53496
rect 15344 53456 15350 53468
rect 16025 53465 16037 53468
rect 16071 53465 16083 53499
rect 16025 53459 16083 53465
rect 16114 53456 16120 53508
rect 16172 53496 16178 53508
rect 16347 53499 16405 53505
rect 16347 53496 16359 53499
rect 16172 53468 16359 53496
rect 16172 53456 16178 53468
rect 16347 53465 16359 53468
rect 16393 53496 16405 53499
rect 16666 53496 16672 53508
rect 16393 53468 16672 53496
rect 16393 53465 16405 53468
rect 16347 53459 16405 53465
rect 16666 53456 16672 53468
rect 16724 53456 16730 53508
rect 19889 53499 19947 53505
rect 19889 53465 19901 53499
rect 19935 53496 19947 53499
rect 20346 53496 20352 53508
rect 19935 53468 20352 53496
rect 19935 53465 19947 53468
rect 19889 53459 19947 53465
rect 20346 53456 20352 53468
rect 20404 53456 20410 53508
rect 24780 53440 24808 53536
rect 25958 53524 25964 53536
rect 26016 53524 26022 53576
rect 11422 53428 11428 53440
rect 11383 53400 11428 53428
rect 11422 53388 11428 53400
rect 11480 53388 11486 53440
rect 11974 53388 11980 53440
rect 12032 53428 12038 53440
rect 12069 53431 12127 53437
rect 12069 53428 12081 53431
rect 12032 53400 12081 53428
rect 12032 53388 12038 53400
rect 12069 53397 12081 53400
rect 12115 53397 12127 53431
rect 12069 53391 12127 53397
rect 13998 53388 14004 53440
rect 14056 53428 14062 53440
rect 14277 53431 14335 53437
rect 14277 53428 14289 53431
rect 14056 53400 14289 53428
rect 14056 53388 14062 53400
rect 14277 53397 14289 53400
rect 14323 53428 14335 53431
rect 14645 53431 14703 53437
rect 14645 53428 14657 53431
rect 14323 53400 14657 53428
rect 14323 53397 14335 53400
rect 14277 53391 14335 53397
rect 14645 53397 14657 53400
rect 14691 53397 14703 53431
rect 14645 53391 14703 53397
rect 14734 53388 14740 53440
rect 14792 53428 14798 53440
rect 15013 53431 15071 53437
rect 15013 53428 15025 53431
rect 14792 53400 15025 53428
rect 14792 53388 14798 53400
rect 15013 53397 15025 53400
rect 15059 53397 15071 53431
rect 15013 53391 15071 53397
rect 15102 53388 15108 53440
rect 15160 53428 15166 53440
rect 15657 53431 15715 53437
rect 15657 53428 15669 53431
rect 15160 53400 15669 53428
rect 15160 53388 15166 53400
rect 15657 53397 15669 53400
rect 15703 53428 15715 53431
rect 16485 53431 16543 53437
rect 16485 53428 16497 53431
rect 15703 53400 16497 53428
rect 15703 53397 15715 53400
rect 15657 53391 15715 53397
rect 16485 53397 16497 53400
rect 16531 53428 16543 53431
rect 16574 53428 16580 53440
rect 16531 53400 16580 53428
rect 16531 53397 16543 53400
rect 16485 53391 16543 53397
rect 16574 53388 16580 53400
rect 16632 53428 16638 53440
rect 17034 53428 17040 53440
rect 16632 53400 17040 53428
rect 16632 53388 16638 53400
rect 17034 53388 17040 53400
rect 17092 53388 17098 53440
rect 17313 53431 17371 53437
rect 17313 53397 17325 53431
rect 17359 53428 17371 53431
rect 17770 53428 17776 53440
rect 17359 53400 17776 53428
rect 17359 53397 17371 53400
rect 17313 53391 17371 53397
rect 17770 53388 17776 53400
rect 17828 53388 17834 53440
rect 21818 53388 21824 53440
rect 21876 53428 21882 53440
rect 22094 53428 22100 53440
rect 21876 53400 22100 53428
rect 21876 53388 21882 53400
rect 22094 53388 22100 53400
rect 22152 53388 22158 53440
rect 24489 53431 24547 53437
rect 24489 53397 24501 53431
rect 24535 53428 24547 53431
rect 24762 53428 24768 53440
rect 24535 53400 24768 53428
rect 24535 53397 24547 53400
rect 24489 53391 24547 53397
rect 24762 53388 24768 53400
rect 24820 53388 24826 53440
rect 1104 53338 28888 53360
rect 1104 53286 5982 53338
rect 6034 53286 6046 53338
rect 6098 53286 6110 53338
rect 6162 53286 6174 53338
rect 6226 53286 15982 53338
rect 16034 53286 16046 53338
rect 16098 53286 16110 53338
rect 16162 53286 16174 53338
rect 16226 53286 25982 53338
rect 26034 53286 26046 53338
rect 26098 53286 26110 53338
rect 26162 53286 26174 53338
rect 26226 53286 28888 53338
rect 1104 53264 28888 53286
rect 10410 53184 10416 53236
rect 10468 53224 10474 53236
rect 10505 53227 10563 53233
rect 10505 53224 10517 53227
rect 10468 53196 10517 53224
rect 10468 53184 10474 53196
rect 10505 53193 10517 53196
rect 10551 53224 10563 53227
rect 10870 53224 10876 53236
rect 10551 53196 10876 53224
rect 10551 53193 10563 53196
rect 10505 53187 10563 53193
rect 10870 53184 10876 53196
rect 10928 53184 10934 53236
rect 11882 53224 11888 53236
rect 11843 53196 11888 53224
rect 11882 53184 11888 53196
rect 11940 53184 11946 53236
rect 14458 53224 14464 53236
rect 14419 53196 14464 53224
rect 14458 53184 14464 53196
rect 14516 53184 14522 53236
rect 15194 53184 15200 53236
rect 15252 53224 15258 53236
rect 16209 53227 16267 53233
rect 16209 53224 16221 53227
rect 15252 53196 16221 53224
rect 15252 53184 15258 53196
rect 16209 53193 16221 53196
rect 16255 53193 16267 53227
rect 16209 53187 16267 53193
rect 16482 53184 16488 53236
rect 16540 53224 16546 53236
rect 16669 53227 16727 53233
rect 16669 53224 16681 53227
rect 16540 53196 16681 53224
rect 16540 53184 16546 53196
rect 16669 53193 16681 53196
rect 16715 53193 16727 53227
rect 17034 53224 17040 53236
rect 16995 53196 17040 53224
rect 16669 53187 16727 53193
rect 17034 53184 17040 53196
rect 17092 53184 17098 53236
rect 17770 53184 17776 53236
rect 17828 53224 17834 53236
rect 17828 53196 18920 53224
rect 17828 53184 17834 53196
rect 16942 53116 16948 53168
rect 17000 53156 17006 53168
rect 17865 53159 17923 53165
rect 17865 53156 17877 53159
rect 17000 53128 17877 53156
rect 17000 53116 17006 53128
rect 17865 53125 17877 53128
rect 17911 53156 17923 53159
rect 18782 53156 18788 53168
rect 17911 53128 18788 53156
rect 17911 53125 17923 53128
rect 17865 53119 17923 53125
rect 12434 53048 12440 53100
rect 12492 53088 12498 53100
rect 12802 53088 12808 53100
rect 12492 53060 12808 53088
rect 12492 53048 12498 53060
rect 12802 53048 12808 53060
rect 12860 53048 12866 53100
rect 18064 53097 18092 53128
rect 18782 53116 18788 53128
rect 18840 53116 18846 53168
rect 18049 53091 18107 53097
rect 18049 53057 18061 53091
rect 18095 53057 18107 53091
rect 18414 53088 18420 53100
rect 18049 53051 18107 53057
rect 18340 53060 18420 53088
rect 11333 53023 11391 53029
rect 11333 52989 11345 53023
rect 11379 53020 11391 53023
rect 11882 53020 11888 53032
rect 11379 52992 11888 53020
rect 11379 52989 11391 52992
rect 11333 52983 11391 52989
rect 11882 52980 11888 52992
rect 11940 52980 11946 53032
rect 12158 52980 12164 53032
rect 12216 52980 12222 53032
rect 12526 52980 12532 53032
rect 12584 53020 12590 53032
rect 12713 53023 12771 53029
rect 12713 53020 12725 53023
rect 12584 52992 12725 53020
rect 12584 52980 12590 52992
rect 12713 52989 12725 52992
rect 12759 52989 12771 53023
rect 12713 52983 12771 52989
rect 13998 52980 14004 53032
rect 14056 53020 14062 53032
rect 15013 53023 15071 53029
rect 15013 53020 15025 53023
rect 14056 52992 15025 53020
rect 14056 52980 14062 52992
rect 15013 52989 15025 52992
rect 15059 52989 15071 53023
rect 15013 52983 15071 52989
rect 16298 52980 16304 53032
rect 16356 53020 16362 53032
rect 18340 53029 18368 53060
rect 18414 53048 18420 53060
rect 18472 53048 18478 53100
rect 16485 53023 16543 53029
rect 16485 53020 16497 53023
rect 16356 52992 16497 53020
rect 16356 52980 16362 52992
rect 16485 52989 16497 52992
rect 16531 52989 16543 53023
rect 16485 52983 16543 52989
rect 18325 53023 18383 53029
rect 18325 52989 18337 53023
rect 18371 52989 18383 53023
rect 18325 52983 18383 52989
rect 18785 53023 18843 53029
rect 18785 52989 18797 53023
rect 18831 53020 18843 53023
rect 18892 53020 18920 53196
rect 20714 53184 20720 53236
rect 20772 53224 20778 53236
rect 21453 53227 21511 53233
rect 21453 53224 21465 53227
rect 20772 53196 21465 53224
rect 20772 53184 20778 53196
rect 21453 53193 21465 53196
rect 21499 53193 21511 53227
rect 23106 53224 23112 53236
rect 23067 53196 23112 53224
rect 21453 53187 21511 53193
rect 19058 53048 19064 53100
rect 19116 53088 19122 53100
rect 19610 53088 19616 53100
rect 19116 53060 19616 53088
rect 19116 53048 19122 53060
rect 19610 53048 19616 53060
rect 19668 53088 19674 53100
rect 20622 53088 20628 53100
rect 19668 53060 20116 53088
rect 20583 53060 20628 53088
rect 19668 53048 19674 53060
rect 20088 53029 20116 53060
rect 20622 53048 20628 53060
rect 20680 53048 20686 53100
rect 21468 53088 21496 53187
rect 23106 53184 23112 53196
rect 23164 53184 23170 53236
rect 23477 53227 23535 53233
rect 23477 53193 23489 53227
rect 23523 53224 23535 53227
rect 23842 53224 23848 53236
rect 23523 53196 23848 53224
rect 23523 53193 23535 53196
rect 23477 53187 23535 53193
rect 22738 53116 22744 53168
rect 22796 53156 22802 53168
rect 23492 53156 23520 53187
rect 23842 53184 23848 53196
rect 23900 53184 23906 53236
rect 22796 53128 23520 53156
rect 22796 53116 22802 53128
rect 24121 53091 24179 53097
rect 21468 53060 21772 53088
rect 21744 53029 21772 53060
rect 24121 53057 24133 53091
rect 24167 53088 24179 53091
rect 24486 53088 24492 53100
rect 24167 53060 24492 53088
rect 24167 53057 24179 53060
rect 24121 53051 24179 53057
rect 24486 53048 24492 53060
rect 24544 53048 24550 53100
rect 19705 53023 19763 53029
rect 19705 53020 19717 53023
rect 18831 52992 18920 53020
rect 19168 52992 19717 53020
rect 18831 52989 18843 52992
rect 18785 52983 18843 52989
rect 11238 52952 11244 52964
rect 11151 52924 11244 52952
rect 11238 52912 11244 52924
rect 11296 52952 11302 52964
rect 11422 52952 11428 52964
rect 11296 52924 11428 52952
rect 11296 52912 11302 52924
rect 11422 52912 11428 52924
rect 11480 52912 11486 52964
rect 12176 52952 12204 52980
rect 17586 52952 17592 52964
rect 11900 52924 12204 52952
rect 17420 52924 17592 52952
rect 11900 52896 11928 52924
rect 11514 52884 11520 52896
rect 11475 52856 11520 52884
rect 11514 52844 11520 52856
rect 11572 52844 11578 52896
rect 11882 52844 11888 52896
rect 11940 52844 11946 52896
rect 12066 52844 12072 52896
rect 12124 52884 12130 52896
rect 12161 52887 12219 52893
rect 12161 52884 12173 52887
rect 12124 52856 12173 52884
rect 12124 52844 12130 52856
rect 12161 52853 12173 52856
rect 12207 52853 12219 52887
rect 13998 52884 14004 52896
rect 13959 52856 14004 52884
rect 12161 52847 12219 52853
rect 13998 52844 14004 52856
rect 14056 52844 14062 52896
rect 14829 52887 14887 52893
rect 14829 52853 14841 52887
rect 14875 52884 14887 52887
rect 15010 52884 15016 52896
rect 14875 52856 15016 52884
rect 14875 52853 14887 52856
rect 14829 52847 14887 52853
rect 15010 52844 15016 52856
rect 15068 52844 15074 52896
rect 15194 52884 15200 52896
rect 15155 52856 15200 52884
rect 15194 52844 15200 52856
rect 15252 52844 15258 52896
rect 17218 52844 17224 52896
rect 17276 52884 17282 52896
rect 17420 52893 17448 52924
rect 17586 52912 17592 52924
rect 17644 52952 17650 52964
rect 18417 52955 18475 52961
rect 18417 52952 18429 52955
rect 17644 52924 18429 52952
rect 17644 52912 17650 52924
rect 18417 52921 18429 52924
rect 18463 52921 18475 52955
rect 18417 52915 18475 52921
rect 17405 52887 17463 52893
rect 17405 52884 17417 52887
rect 17276 52856 17417 52884
rect 17276 52844 17282 52856
rect 17405 52853 17417 52856
rect 17451 52853 17463 52887
rect 17405 52847 17463 52853
rect 18230 52844 18236 52896
rect 18288 52884 18294 52896
rect 18288 52856 18333 52884
rect 18288 52844 18294 52856
rect 18874 52844 18880 52896
rect 18932 52884 18938 52896
rect 19168 52893 19196 52992
rect 19705 52989 19717 52992
rect 19751 52989 19763 53023
rect 19705 52983 19763 52989
rect 20073 53023 20131 53029
rect 20073 52989 20085 53023
rect 20119 52989 20131 53023
rect 20073 52983 20131 52989
rect 20533 53023 20591 53029
rect 20533 52989 20545 53023
rect 20579 52989 20591 53023
rect 20533 52983 20591 52989
rect 21637 53023 21695 53029
rect 21637 52989 21649 53023
rect 21683 52989 21695 53023
rect 21637 52983 21695 52989
rect 21729 53023 21787 53029
rect 21729 52989 21741 53023
rect 21775 53020 21787 53023
rect 21910 53020 21916 53032
rect 21775 52992 21916 53020
rect 21775 52989 21787 52992
rect 21729 52983 21787 52989
rect 19426 52912 19432 52964
rect 19484 52952 19490 52964
rect 20548 52952 20576 52983
rect 20714 52952 20720 52964
rect 19484 52924 20720 52952
rect 19484 52912 19490 52924
rect 20714 52912 20720 52924
rect 20772 52912 20778 52964
rect 21082 52952 21088 52964
rect 21043 52924 21088 52952
rect 21082 52912 21088 52924
rect 21140 52912 21146 52964
rect 19153 52887 19211 52893
rect 19153 52884 19165 52887
rect 18932 52856 19165 52884
rect 18932 52844 18938 52856
rect 19153 52853 19165 52856
rect 19199 52853 19211 52887
rect 19153 52847 19211 52853
rect 19613 52887 19671 52893
rect 19613 52853 19625 52887
rect 19659 52884 19671 52887
rect 19702 52884 19708 52896
rect 19659 52856 19708 52884
rect 19659 52853 19671 52856
rect 19613 52847 19671 52853
rect 19702 52844 19708 52856
rect 19760 52884 19766 52896
rect 20070 52884 20076 52896
rect 19760 52856 20076 52884
rect 19760 52844 19766 52856
rect 20070 52844 20076 52856
rect 20128 52844 20134 52896
rect 21652 52884 21680 52983
rect 21910 52980 21916 52992
rect 21968 52980 21974 53032
rect 24213 53023 24271 53029
rect 24213 52989 24225 53023
rect 24259 53020 24271 53023
rect 24762 53020 24768 53032
rect 24259 52992 24768 53020
rect 24259 52989 24271 52992
rect 24213 52983 24271 52989
rect 24762 52980 24768 52992
rect 24820 52980 24826 53032
rect 22186 52952 22192 52964
rect 22147 52924 22192 52952
rect 22186 52912 22192 52924
rect 22244 52912 22250 52964
rect 22465 52887 22523 52893
rect 22465 52884 22477 52887
rect 21652 52856 22477 52884
rect 22465 52853 22477 52856
rect 22511 52884 22523 52887
rect 22554 52884 22560 52896
rect 22511 52856 22560 52884
rect 22511 52853 22523 52856
rect 22465 52847 22523 52853
rect 22554 52844 22560 52856
rect 22612 52844 22618 52896
rect 23934 52844 23940 52896
rect 23992 52884 23998 52896
rect 25593 52887 25651 52893
rect 25593 52884 25605 52887
rect 23992 52856 25605 52884
rect 23992 52844 23998 52856
rect 25593 52853 25605 52856
rect 25639 52853 25651 52887
rect 25593 52847 25651 52853
rect 1104 52794 28888 52816
rect 1104 52742 10982 52794
rect 11034 52742 11046 52794
rect 11098 52742 11110 52794
rect 11162 52742 11174 52794
rect 11226 52742 20982 52794
rect 21034 52742 21046 52794
rect 21098 52742 21110 52794
rect 21162 52742 21174 52794
rect 21226 52742 28888 52794
rect 1104 52720 28888 52742
rect 10781 52683 10839 52689
rect 10781 52649 10793 52683
rect 10827 52680 10839 52683
rect 10870 52680 10876 52692
rect 10827 52652 10876 52680
rect 10827 52649 10839 52652
rect 10781 52643 10839 52649
rect 10870 52640 10876 52652
rect 10928 52640 10934 52692
rect 11790 52680 11796 52692
rect 11751 52652 11796 52680
rect 11790 52640 11796 52652
rect 11848 52640 11854 52692
rect 13814 52680 13820 52692
rect 13727 52652 13820 52680
rect 13814 52640 13820 52652
rect 13872 52680 13878 52692
rect 15102 52680 15108 52692
rect 13872 52652 15108 52680
rect 13872 52640 13878 52652
rect 15102 52640 15108 52652
rect 15160 52640 15166 52692
rect 16298 52640 16304 52692
rect 16356 52680 16362 52692
rect 16485 52683 16543 52689
rect 16485 52680 16497 52683
rect 16356 52652 16497 52680
rect 16356 52640 16362 52652
rect 16485 52649 16497 52652
rect 16531 52649 16543 52683
rect 16485 52643 16543 52649
rect 18141 52683 18199 52689
rect 18141 52649 18153 52683
rect 18187 52680 18199 52683
rect 18414 52680 18420 52692
rect 18187 52652 18420 52680
rect 18187 52649 18199 52652
rect 18141 52643 18199 52649
rect 18414 52640 18420 52652
rect 18472 52640 18478 52692
rect 19150 52680 19156 52692
rect 19111 52652 19156 52680
rect 19150 52640 19156 52652
rect 19208 52640 19214 52692
rect 19705 52683 19763 52689
rect 19705 52649 19717 52683
rect 19751 52680 19763 52683
rect 19978 52680 19984 52692
rect 19751 52652 19984 52680
rect 19751 52649 19763 52652
rect 19705 52643 19763 52649
rect 19978 52640 19984 52652
rect 20036 52640 20042 52692
rect 20073 52683 20131 52689
rect 20073 52649 20085 52683
rect 20119 52680 20131 52683
rect 20162 52680 20168 52692
rect 20119 52652 20168 52680
rect 20119 52649 20131 52652
rect 20073 52643 20131 52649
rect 20162 52640 20168 52652
rect 20220 52640 20226 52692
rect 20714 52640 20720 52692
rect 20772 52680 20778 52692
rect 20993 52683 21051 52689
rect 20993 52680 21005 52683
rect 20772 52652 21005 52680
rect 20772 52640 20778 52652
rect 20993 52649 21005 52652
rect 21039 52649 21051 52683
rect 20993 52643 21051 52649
rect 22833 52683 22891 52689
rect 22833 52649 22845 52683
rect 22879 52680 22891 52683
rect 23934 52680 23940 52692
rect 22879 52652 23940 52680
rect 22879 52649 22891 52652
rect 22833 52643 22891 52649
rect 23934 52640 23940 52652
rect 23992 52640 23998 52692
rect 11517 52615 11575 52621
rect 11517 52581 11529 52615
rect 11563 52612 11575 52615
rect 11882 52612 11888 52624
rect 11563 52584 11888 52612
rect 11563 52581 11575 52584
rect 11517 52575 11575 52581
rect 11882 52572 11888 52584
rect 11940 52572 11946 52624
rect 13173 52615 13231 52621
rect 13173 52581 13185 52615
rect 13219 52612 13231 52615
rect 14001 52615 14059 52621
rect 14001 52612 14013 52615
rect 13219 52584 14013 52612
rect 13219 52581 13231 52584
rect 13173 52575 13231 52581
rect 14001 52581 14013 52584
rect 14047 52612 14059 52615
rect 14274 52612 14280 52624
rect 14047 52584 14280 52612
rect 14047 52581 14059 52584
rect 14001 52575 14059 52581
rect 14274 52572 14280 52584
rect 14332 52572 14338 52624
rect 14369 52615 14427 52621
rect 14369 52581 14381 52615
rect 14415 52612 14427 52615
rect 14458 52612 14464 52624
rect 14415 52584 14464 52612
rect 14415 52581 14427 52584
rect 14369 52575 14427 52581
rect 14458 52572 14464 52584
rect 14516 52572 14522 52624
rect 14734 52612 14740 52624
rect 14695 52584 14740 52612
rect 14734 52572 14740 52584
rect 14792 52572 14798 52624
rect 15010 52612 15016 52624
rect 14971 52584 15016 52612
rect 15010 52572 15016 52584
rect 15068 52572 15074 52624
rect 18046 52572 18052 52624
rect 18104 52612 18110 52624
rect 19996 52612 20024 52640
rect 21726 52612 21732 52624
rect 18104 52584 18736 52612
rect 19996 52584 21732 52612
rect 18104 52572 18110 52584
rect 1670 52544 1676 52556
rect 1631 52516 1676 52544
rect 1670 52504 1676 52516
rect 1728 52504 1734 52556
rect 3053 52547 3111 52553
rect 3053 52513 3065 52547
rect 3099 52544 3111 52547
rect 4062 52544 4068 52556
rect 3099 52516 4068 52544
rect 3099 52513 3111 52516
rect 3053 52507 3111 52513
rect 4062 52504 4068 52516
rect 4120 52504 4126 52556
rect 10597 52547 10655 52553
rect 10597 52513 10609 52547
rect 10643 52513 10655 52547
rect 10597 52507 10655 52513
rect 1397 52479 1455 52485
rect 1397 52445 1409 52479
rect 1443 52476 1455 52479
rect 1578 52476 1584 52488
rect 1443 52448 1584 52476
rect 1443 52445 1455 52448
rect 1397 52439 1455 52445
rect 1578 52436 1584 52448
rect 1636 52436 1642 52488
rect 10612 52476 10640 52507
rect 11422 52504 11428 52556
rect 11480 52544 11486 52556
rect 11609 52547 11667 52553
rect 11609 52544 11621 52547
rect 11480 52516 11621 52544
rect 11480 52504 11486 52516
rect 11609 52513 11621 52516
rect 11655 52544 11667 52547
rect 12250 52544 12256 52556
rect 11655 52516 12256 52544
rect 11655 52513 11667 52516
rect 11609 52507 11667 52513
rect 12250 52504 12256 52516
rect 12308 52504 12314 52556
rect 12618 52544 12624 52556
rect 12579 52516 12624 52544
rect 12618 52504 12624 52516
rect 12676 52504 12682 52556
rect 13541 52547 13599 52553
rect 13541 52513 13553 52547
rect 13587 52544 13599 52547
rect 13906 52544 13912 52556
rect 13587 52516 13912 52544
rect 13587 52513 13599 52516
rect 13541 52507 13599 52513
rect 13906 52504 13912 52516
rect 13964 52504 13970 52556
rect 15933 52547 15991 52553
rect 15933 52513 15945 52547
rect 15979 52513 15991 52547
rect 15933 52507 15991 52513
rect 10612 52448 11100 52476
rect 11072 52408 11100 52448
rect 12434 52436 12440 52488
rect 12492 52476 12498 52488
rect 13633 52479 13691 52485
rect 12492 52448 12537 52476
rect 12492 52436 12498 52448
rect 13633 52445 13645 52479
rect 13679 52445 13691 52479
rect 13633 52439 13691 52445
rect 11330 52408 11336 52420
rect 11072 52380 11336 52408
rect 11330 52368 11336 52380
rect 11388 52368 11394 52420
rect 11974 52300 11980 52352
rect 12032 52340 12038 52352
rect 12069 52343 12127 52349
rect 12069 52340 12081 52343
rect 12032 52312 12081 52340
rect 12032 52300 12038 52312
rect 12069 52309 12081 52312
rect 12115 52309 12127 52343
rect 12069 52303 12127 52309
rect 12805 52343 12863 52349
rect 12805 52309 12817 52343
rect 12851 52340 12863 52343
rect 12986 52340 12992 52352
rect 12851 52312 12992 52340
rect 12851 52309 12863 52312
rect 12805 52303 12863 52309
rect 12986 52300 12992 52312
rect 13044 52300 13050 52352
rect 13648 52340 13676 52439
rect 14366 52436 14372 52488
rect 14424 52476 14430 52488
rect 14734 52476 14740 52488
rect 14424 52448 14740 52476
rect 14424 52436 14430 52448
rect 14734 52436 14740 52448
rect 14792 52436 14798 52488
rect 15194 52436 15200 52488
rect 15252 52476 15258 52488
rect 15289 52479 15347 52485
rect 15289 52476 15301 52479
rect 15252 52448 15301 52476
rect 15252 52436 15258 52448
rect 15289 52445 15301 52448
rect 15335 52445 15347 52479
rect 15948 52476 15976 52507
rect 16298 52504 16304 52556
rect 16356 52544 16362 52556
rect 16853 52547 16911 52553
rect 16853 52544 16865 52547
rect 16356 52516 16865 52544
rect 16356 52504 16362 52516
rect 16853 52513 16865 52516
rect 16899 52513 16911 52547
rect 17034 52544 17040 52556
rect 16995 52516 17040 52544
rect 16853 52507 16911 52513
rect 17034 52504 17040 52516
rect 17092 52504 17098 52556
rect 17770 52504 17776 52556
rect 17828 52544 17834 52556
rect 18708 52553 18736 52584
rect 21726 52572 21732 52584
rect 21784 52612 21790 52624
rect 22281 52615 22339 52621
rect 22281 52612 22293 52615
rect 21784 52584 22293 52612
rect 21784 52572 21790 52584
rect 22281 52581 22293 52584
rect 22327 52581 22339 52615
rect 22281 52575 22339 52581
rect 18233 52547 18291 52553
rect 18233 52544 18245 52547
rect 17828 52516 18245 52544
rect 17828 52504 17834 52516
rect 18233 52513 18245 52516
rect 18279 52513 18291 52547
rect 18233 52507 18291 52513
rect 18693 52547 18751 52553
rect 18693 52513 18705 52547
rect 18739 52513 18751 52547
rect 18693 52507 18751 52513
rect 18782 52504 18788 52556
rect 18840 52544 18846 52556
rect 19061 52547 19119 52553
rect 19061 52544 19073 52547
rect 18840 52516 19073 52544
rect 18840 52504 18846 52516
rect 19061 52513 19073 52516
rect 19107 52513 19119 52547
rect 19061 52507 19119 52513
rect 21085 52547 21143 52553
rect 21085 52513 21097 52547
rect 21131 52544 21143 52547
rect 21358 52544 21364 52556
rect 21131 52516 21364 52544
rect 21131 52513 21143 52516
rect 21085 52507 21143 52513
rect 21358 52504 21364 52516
rect 21416 52504 21422 52556
rect 21453 52547 21511 52553
rect 21453 52513 21465 52547
rect 21499 52544 21511 52547
rect 22554 52544 22560 52556
rect 21499 52516 22560 52544
rect 21499 52513 21511 52516
rect 21453 52507 21511 52513
rect 16482 52476 16488 52488
rect 15948 52448 16488 52476
rect 15289 52439 15347 52445
rect 16482 52436 16488 52448
rect 16540 52436 16546 52488
rect 17218 52436 17224 52488
rect 17276 52476 17282 52488
rect 17313 52479 17371 52485
rect 17313 52476 17325 52479
rect 17276 52448 17325 52476
rect 17276 52436 17282 52448
rect 17313 52445 17325 52448
rect 17359 52445 17371 52479
rect 17313 52439 17371 52445
rect 19334 52436 19340 52488
rect 19392 52476 19398 52488
rect 20162 52476 20168 52488
rect 19392 52448 20168 52476
rect 19392 52436 19398 52448
rect 20162 52436 20168 52448
rect 20220 52436 20226 52488
rect 20714 52436 20720 52488
rect 20772 52476 20778 52488
rect 21468 52476 21496 52507
rect 22554 52504 22560 52516
rect 22612 52504 22618 52556
rect 23290 52544 23296 52556
rect 23251 52516 23296 52544
rect 23290 52504 23296 52516
rect 23348 52504 23354 52556
rect 23845 52547 23903 52553
rect 23845 52513 23857 52547
rect 23891 52544 23903 52547
rect 24118 52544 24124 52556
rect 23891 52516 24124 52544
rect 23891 52513 23903 52516
rect 23845 52507 23903 52513
rect 21726 52476 21732 52488
rect 20772 52448 21496 52476
rect 21687 52448 21732 52476
rect 20772 52436 20778 52448
rect 21726 52436 21732 52448
rect 21784 52436 21790 52488
rect 23106 52476 23112 52488
rect 23067 52448 23112 52476
rect 23106 52436 23112 52448
rect 23164 52436 23170 52488
rect 23860 52476 23888 52507
rect 24118 52504 24124 52516
rect 24176 52504 24182 52556
rect 23400 52448 23888 52476
rect 13722 52368 13728 52420
rect 13780 52408 13786 52420
rect 15562 52408 15568 52420
rect 13780 52380 15568 52408
rect 13780 52368 13786 52380
rect 15562 52368 15568 52380
rect 15620 52368 15626 52420
rect 19426 52368 19432 52420
rect 19484 52408 19490 52420
rect 19978 52408 19984 52420
rect 19484 52380 19984 52408
rect 19484 52368 19490 52380
rect 19978 52368 19984 52380
rect 20036 52368 20042 52420
rect 23198 52368 23204 52420
rect 23256 52408 23262 52420
rect 23400 52408 23428 52448
rect 23750 52408 23756 52420
rect 23256 52380 23428 52408
rect 23711 52380 23756 52408
rect 23256 52368 23262 52380
rect 23750 52368 23756 52380
rect 23808 52368 23814 52420
rect 14826 52340 14832 52352
rect 13648 52312 14832 52340
rect 14826 52300 14832 52312
rect 14884 52300 14890 52352
rect 16574 52300 16580 52352
rect 16632 52340 16638 52352
rect 17681 52343 17739 52349
rect 17681 52340 17693 52343
rect 16632 52312 17693 52340
rect 16632 52300 16638 52312
rect 17681 52309 17693 52312
rect 17727 52340 17739 52343
rect 18230 52340 18236 52352
rect 17727 52312 18236 52340
rect 17727 52309 17739 52312
rect 17681 52303 17739 52309
rect 18230 52300 18236 52312
rect 18288 52300 18294 52352
rect 20346 52340 20352 52352
rect 20307 52312 20352 52340
rect 20346 52300 20352 52312
rect 20404 52340 20410 52352
rect 22186 52340 22192 52352
rect 20404 52312 22192 52340
rect 20404 52300 20410 52312
rect 22186 52300 22192 52312
rect 22244 52300 22250 52352
rect 23842 52300 23848 52352
rect 23900 52340 23906 52352
rect 24305 52343 24363 52349
rect 24305 52340 24317 52343
rect 23900 52312 24317 52340
rect 23900 52300 23906 52312
rect 24305 52309 24317 52312
rect 24351 52309 24363 52343
rect 24305 52303 24363 52309
rect 1104 52250 28888 52272
rect 1104 52198 5982 52250
rect 6034 52198 6046 52250
rect 6098 52198 6110 52250
rect 6162 52198 6174 52250
rect 6226 52198 15982 52250
rect 16034 52198 16046 52250
rect 16098 52198 16110 52250
rect 16162 52198 16174 52250
rect 16226 52198 25982 52250
rect 26034 52198 26046 52250
rect 26098 52198 26110 52250
rect 26162 52198 26174 52250
rect 26226 52198 28888 52250
rect 1104 52176 28888 52198
rect 1670 52136 1676 52148
rect 1631 52108 1676 52136
rect 1670 52096 1676 52108
rect 1728 52096 1734 52148
rect 8386 52136 8392 52148
rect 8347 52108 8392 52136
rect 8386 52096 8392 52108
rect 8444 52096 8450 52148
rect 10873 52139 10931 52145
rect 10873 52105 10885 52139
rect 10919 52136 10931 52139
rect 10962 52136 10968 52148
rect 10919 52108 10968 52136
rect 10919 52105 10931 52108
rect 10873 52099 10931 52105
rect 8021 51935 8079 51941
rect 8021 51901 8033 51935
rect 8067 51932 8079 51935
rect 8386 51932 8392 51944
rect 8067 51904 8392 51932
rect 8067 51901 8079 51904
rect 8021 51895 8079 51901
rect 8386 51892 8392 51904
rect 8444 51892 8450 51944
rect 10321 51935 10379 51941
rect 10321 51901 10333 51935
rect 10367 51932 10379 51935
rect 10888 51932 10916 52099
rect 10962 52096 10968 52108
rect 11020 52096 11026 52148
rect 11241 52139 11299 52145
rect 11241 52105 11253 52139
rect 11287 52136 11299 52139
rect 11330 52136 11336 52148
rect 11287 52108 11336 52136
rect 11287 52105 11299 52108
rect 11241 52099 11299 52105
rect 11330 52096 11336 52108
rect 11388 52096 11394 52148
rect 11885 52139 11943 52145
rect 11885 52136 11897 52139
rect 11440 52108 11897 52136
rect 10367 51904 10916 51932
rect 11333 51935 11391 51941
rect 10367 51901 10379 51904
rect 10321 51895 10379 51901
rect 11333 51901 11345 51935
rect 11379 51932 11391 51935
rect 11440 51932 11468 52108
rect 11885 52105 11897 52108
rect 11931 52136 11943 52139
rect 12250 52136 12256 52148
rect 11931 52108 12256 52136
rect 11931 52105 11943 52108
rect 11885 52099 11943 52105
rect 12250 52096 12256 52108
rect 12308 52096 12314 52148
rect 14826 52136 14832 52148
rect 14787 52108 14832 52136
rect 14826 52096 14832 52108
rect 14884 52096 14890 52148
rect 15102 52096 15108 52148
rect 15160 52136 15166 52148
rect 15197 52139 15255 52145
rect 15197 52136 15209 52139
rect 15160 52108 15209 52136
rect 15160 52096 15166 52108
rect 15197 52105 15209 52108
rect 15243 52136 15255 52139
rect 15562 52136 15568 52148
rect 15243 52108 15568 52136
rect 15243 52105 15255 52108
rect 15197 52099 15255 52105
rect 15562 52096 15568 52108
rect 15620 52096 15626 52148
rect 18325 52139 18383 52145
rect 18325 52105 18337 52139
rect 18371 52136 18383 52139
rect 18506 52136 18512 52148
rect 18371 52108 18512 52136
rect 18371 52105 18383 52108
rect 18325 52099 18383 52105
rect 18506 52096 18512 52108
rect 18564 52096 18570 52148
rect 18598 52096 18604 52148
rect 18656 52136 18662 52148
rect 18782 52136 18788 52148
rect 18656 52108 18788 52136
rect 18656 52096 18662 52108
rect 18782 52096 18788 52108
rect 18840 52096 18846 52148
rect 20257 52139 20315 52145
rect 20257 52105 20269 52139
rect 20303 52136 20315 52139
rect 20714 52136 20720 52148
rect 20303 52108 20720 52136
rect 20303 52105 20315 52108
rect 20257 52099 20315 52105
rect 20714 52096 20720 52108
rect 20772 52096 20778 52148
rect 21358 52096 21364 52148
rect 21416 52136 21422 52148
rect 21542 52136 21548 52148
rect 21416 52108 21548 52136
rect 21416 52096 21422 52108
rect 21542 52096 21548 52108
rect 21600 52136 21606 52148
rect 21821 52139 21879 52145
rect 21821 52136 21833 52139
rect 21600 52108 21833 52136
rect 21600 52096 21606 52108
rect 21821 52105 21833 52108
rect 21867 52105 21879 52139
rect 21821 52099 21879 52105
rect 22462 52096 22468 52148
rect 22520 52136 22526 52148
rect 22557 52139 22615 52145
rect 22557 52136 22569 52139
rect 22520 52108 22569 52136
rect 22520 52096 22526 52108
rect 22557 52105 22569 52108
rect 22603 52105 22615 52139
rect 22557 52099 22615 52105
rect 23106 52096 23112 52148
rect 23164 52136 23170 52148
rect 23293 52139 23351 52145
rect 23293 52136 23305 52139
rect 23164 52108 23305 52136
rect 23164 52096 23170 52108
rect 23293 52105 23305 52108
rect 23339 52105 23351 52139
rect 23293 52099 23351 52105
rect 13906 52028 13912 52080
rect 13964 52068 13970 52080
rect 17037 52071 17095 52077
rect 17037 52068 17049 52071
rect 13964 52040 17049 52068
rect 13964 52028 13970 52040
rect 17037 52037 17049 52040
rect 17083 52068 17095 52071
rect 18414 52068 18420 52080
rect 17083 52040 18420 52068
rect 17083 52037 17095 52040
rect 17037 52031 17095 52037
rect 18414 52028 18420 52040
rect 18472 52028 18478 52080
rect 18966 52028 18972 52080
rect 19024 52068 19030 52080
rect 19245 52071 19303 52077
rect 19245 52068 19257 52071
rect 19024 52040 19257 52068
rect 19024 52028 19030 52040
rect 19245 52037 19257 52040
rect 19291 52037 19303 52071
rect 19245 52031 19303 52037
rect 11974 51960 11980 52012
rect 12032 52000 12038 52012
rect 14185 52003 14243 52009
rect 14185 52000 14197 52003
rect 12032 51972 14197 52000
rect 12032 51960 12038 51972
rect 14185 51969 14197 51972
rect 14231 51969 14243 52003
rect 15286 52000 15292 52012
rect 15247 51972 15292 52000
rect 14185 51963 14243 51969
rect 12802 51932 12808 51944
rect 11379 51904 11468 51932
rect 12763 51904 12808 51932
rect 11379 51901 11391 51904
rect 11333 51895 11391 51901
rect 12802 51892 12808 51904
rect 12860 51892 12866 51944
rect 13081 51935 13139 51941
rect 13081 51932 13093 51935
rect 12912 51904 13093 51932
rect 1578 51756 1584 51808
rect 1636 51796 1642 51808
rect 1949 51799 2007 51805
rect 1949 51796 1961 51799
rect 1636 51768 1961 51796
rect 1636 51756 1642 51768
rect 1949 51765 1961 51768
rect 1995 51765 2007 51799
rect 7834 51796 7840 51808
rect 7795 51768 7840 51796
rect 1949 51759 2007 51765
rect 7834 51756 7840 51768
rect 7892 51756 7898 51808
rect 10502 51796 10508 51808
rect 10463 51768 10508 51796
rect 10502 51756 10508 51768
rect 10560 51756 10566 51808
rect 11517 51799 11575 51805
rect 11517 51765 11529 51799
rect 11563 51796 11575 51799
rect 12342 51796 12348 51808
rect 11563 51768 12348 51796
rect 11563 51765 11575 51768
rect 11517 51759 11575 51765
rect 12342 51756 12348 51768
rect 12400 51756 12406 51808
rect 12618 51796 12624 51808
rect 12579 51768 12624 51796
rect 12618 51756 12624 51768
rect 12676 51796 12682 51808
rect 12912 51796 12940 51904
rect 13081 51901 13093 51904
rect 13127 51901 13139 51935
rect 14200 51932 14228 51963
rect 15286 51960 15292 51972
rect 15344 52000 15350 52012
rect 16114 52000 16120 52012
rect 15344 51972 16120 52000
rect 15344 51960 15350 51972
rect 16114 51960 16120 51972
rect 16172 51960 16178 52012
rect 17497 52003 17555 52009
rect 17497 51969 17509 52003
rect 17543 52000 17555 52003
rect 19150 52000 19156 52012
rect 17543 51972 19156 52000
rect 17543 51969 17555 51972
rect 17497 51963 17555 51969
rect 19150 51960 19156 51972
rect 19208 51960 19214 52012
rect 19889 52003 19947 52009
rect 19889 51969 19901 52003
rect 19935 52000 19947 52003
rect 21376 52000 21404 52096
rect 23308 52068 23336 52099
rect 24854 52096 24860 52148
rect 24912 52136 24918 52148
rect 25041 52139 25099 52145
rect 25041 52136 25053 52139
rect 24912 52108 25053 52136
rect 24912 52096 24918 52108
rect 25041 52105 25053 52108
rect 25087 52105 25099 52139
rect 25041 52099 25099 52105
rect 23750 52068 23756 52080
rect 23308 52040 23756 52068
rect 23750 52028 23756 52040
rect 23808 52028 23814 52080
rect 23934 52028 23940 52080
rect 23992 52068 23998 52080
rect 24118 52068 24124 52080
rect 23992 52040 24124 52068
rect 23992 52028 23998 52040
rect 24118 52028 24124 52040
rect 24176 52028 24182 52080
rect 19935 51972 21404 52000
rect 23017 52003 23075 52009
rect 19935 51969 19947 51972
rect 19889 51963 19947 51969
rect 15381 51935 15439 51941
rect 15381 51932 15393 51935
rect 14200 51904 15393 51932
rect 13081 51895 13139 51901
rect 15381 51901 15393 51904
rect 15427 51932 15439 51935
rect 16666 51932 16672 51944
rect 15427 51904 16672 51932
rect 15427 51901 15439 51904
rect 15381 51895 15439 51901
rect 16666 51892 16672 51904
rect 16724 51932 16730 51944
rect 16853 51935 16911 51941
rect 16853 51932 16865 51935
rect 16724 51904 16865 51932
rect 16724 51892 16730 51904
rect 16853 51901 16865 51904
rect 16899 51901 16911 51935
rect 16853 51895 16911 51901
rect 17034 51892 17040 51944
rect 17092 51892 17098 51944
rect 17865 51935 17923 51941
rect 17865 51901 17877 51935
rect 17911 51932 17923 51935
rect 18506 51932 18512 51944
rect 17911 51904 18368 51932
rect 18467 51904 18512 51932
rect 17911 51901 17923 51904
rect 17865 51895 17923 51901
rect 16022 51824 16028 51876
rect 16080 51864 16086 51876
rect 16482 51864 16488 51876
rect 16080 51836 16488 51864
rect 16080 51824 16086 51836
rect 16482 51824 16488 51836
rect 16540 51824 16546 51876
rect 16761 51867 16819 51873
rect 16761 51833 16773 51867
rect 16807 51864 16819 51867
rect 17052 51864 17080 51892
rect 18046 51864 18052 51876
rect 16807 51836 18052 51864
rect 16807 51833 16819 51836
rect 16761 51827 16819 51833
rect 18046 51824 18052 51836
rect 18104 51824 18110 51876
rect 18340 51864 18368 51904
rect 18506 51892 18512 51904
rect 18564 51892 18570 51944
rect 18598 51892 18604 51944
rect 18656 51932 18662 51944
rect 19245 51935 19303 51941
rect 19245 51932 19257 51935
rect 18656 51904 19257 51932
rect 18656 51892 18662 51904
rect 19245 51901 19257 51904
rect 19291 51932 19303 51935
rect 19334 51932 19340 51944
rect 19291 51904 19340 51932
rect 19291 51901 19303 51904
rect 19245 51895 19303 51901
rect 19334 51892 19340 51904
rect 19392 51892 19398 51944
rect 20162 51892 20168 51944
rect 20220 51932 20226 51944
rect 21008 51941 21036 51972
rect 23017 51969 23029 52003
rect 23063 52000 23075 52003
rect 23290 52000 23296 52012
rect 23063 51972 23296 52000
rect 23063 51969 23075 51972
rect 23017 51963 23075 51969
rect 23290 51960 23296 51972
rect 23348 51960 23354 52012
rect 23474 51960 23480 52012
rect 23532 52000 23538 52012
rect 24397 52003 24455 52009
rect 24397 52000 24409 52003
rect 23532 51972 24409 52000
rect 23532 51960 23538 51972
rect 24397 51969 24409 51972
rect 24443 51969 24455 52003
rect 24397 51963 24455 51969
rect 20349 51935 20407 51941
rect 20349 51932 20361 51935
rect 20220 51904 20361 51932
rect 20220 51892 20226 51904
rect 20349 51901 20361 51904
rect 20395 51901 20407 51935
rect 20349 51895 20407 51901
rect 20993 51935 21051 51941
rect 20993 51901 21005 51935
rect 21039 51901 21051 51935
rect 20993 51895 21051 51901
rect 21085 51935 21143 51941
rect 21085 51901 21097 51935
rect 21131 51901 21143 51935
rect 21358 51932 21364 51944
rect 21319 51904 21364 51932
rect 21085 51895 21143 51901
rect 18616 51864 18644 51892
rect 18340 51836 18644 51864
rect 12676 51768 12940 51796
rect 12676 51756 12682 51768
rect 15286 51756 15292 51808
rect 15344 51796 15350 51808
rect 16298 51796 16304 51808
rect 15344 51768 16304 51796
rect 15344 51756 15350 51768
rect 16298 51756 16304 51768
rect 16356 51756 16362 51808
rect 18506 51756 18512 51808
rect 18564 51796 18570 51808
rect 18966 51796 18972 51808
rect 18564 51768 18972 51796
rect 18564 51756 18570 51768
rect 18966 51756 18972 51768
rect 19024 51756 19030 51808
rect 20346 51756 20352 51808
rect 20404 51796 20410 51808
rect 21100 51796 21128 51895
rect 21358 51892 21364 51904
rect 21416 51892 21422 51944
rect 21545 51935 21603 51941
rect 21545 51901 21557 51935
rect 21591 51932 21603 51935
rect 21726 51932 21732 51944
rect 21591 51904 21732 51932
rect 21591 51901 21603 51904
rect 21545 51895 21603 51901
rect 21726 51892 21732 51904
rect 21784 51892 21790 51944
rect 22373 51935 22431 51941
rect 22373 51932 22385 51935
rect 22204 51904 22385 51932
rect 20404 51768 21128 51796
rect 20404 51756 20410 51768
rect 21726 51756 21732 51808
rect 21784 51796 21790 51808
rect 22204 51805 22232 51904
rect 22373 51901 22385 51904
rect 22419 51901 22431 51935
rect 24673 51935 24731 51941
rect 24673 51932 24685 51935
rect 22373 51895 22431 51901
rect 23676 51904 24685 51932
rect 23676 51876 23704 51904
rect 24673 51901 24685 51904
rect 24719 51901 24731 51935
rect 24673 51895 24731 51901
rect 23658 51864 23664 51876
rect 23619 51836 23664 51864
rect 23658 51824 23664 51836
rect 23716 51824 23722 51876
rect 23842 51864 23848 51876
rect 23803 51836 23848 51864
rect 23842 51824 23848 51836
rect 23900 51824 23906 51876
rect 24029 51867 24087 51873
rect 24029 51833 24041 51867
rect 24075 51864 24087 51867
rect 24854 51864 24860 51876
rect 24075 51836 24860 51864
rect 24075 51833 24087 51836
rect 24029 51827 24087 51833
rect 24854 51824 24860 51836
rect 24912 51824 24918 51876
rect 22189 51799 22247 51805
rect 22189 51796 22201 51799
rect 21784 51768 22201 51796
rect 21784 51756 21790 51768
rect 22189 51765 22201 51768
rect 22235 51765 22247 51799
rect 23934 51796 23940 51808
rect 23895 51768 23940 51796
rect 22189 51759 22247 51765
rect 23934 51756 23940 51768
rect 23992 51756 23998 51808
rect 1104 51706 28888 51728
rect 1104 51654 10982 51706
rect 11034 51654 11046 51706
rect 11098 51654 11110 51706
rect 11162 51654 11174 51706
rect 11226 51654 20982 51706
rect 21034 51654 21046 51706
rect 21098 51654 21110 51706
rect 21162 51654 21174 51706
rect 21226 51654 28888 51706
rect 1104 51632 28888 51654
rect 10410 51592 10416 51604
rect 10371 51564 10416 51592
rect 10410 51552 10416 51564
rect 10468 51592 10474 51604
rect 10778 51592 10784 51604
rect 10468 51564 10784 51592
rect 10468 51552 10474 51564
rect 10778 51552 10784 51564
rect 10836 51592 10842 51604
rect 11057 51595 11115 51601
rect 11057 51592 11069 51595
rect 10836 51564 11069 51592
rect 10836 51552 10842 51564
rect 11057 51561 11069 51564
rect 11103 51561 11115 51595
rect 11057 51555 11115 51561
rect 11517 51595 11575 51601
rect 11517 51561 11529 51595
rect 11563 51592 11575 51595
rect 11974 51592 11980 51604
rect 11563 51564 11980 51592
rect 11563 51561 11575 51564
rect 11517 51555 11575 51561
rect 11974 51552 11980 51564
rect 12032 51552 12038 51604
rect 12710 51552 12716 51604
rect 12768 51592 12774 51604
rect 13081 51595 13139 51601
rect 13081 51592 13093 51595
rect 12768 51564 13093 51592
rect 12768 51552 12774 51564
rect 13081 51561 13093 51564
rect 13127 51592 13139 51595
rect 13538 51592 13544 51604
rect 13127 51564 13544 51592
rect 13127 51561 13139 51564
rect 13081 51555 13139 51561
rect 13538 51552 13544 51564
rect 13596 51552 13602 51604
rect 14826 51592 14832 51604
rect 14787 51564 14832 51592
rect 14826 51552 14832 51564
rect 14884 51552 14890 51604
rect 16666 51592 16672 51604
rect 16627 51564 16672 51592
rect 16666 51552 16672 51564
rect 16724 51552 16730 51604
rect 17865 51595 17923 51601
rect 17865 51561 17877 51595
rect 17911 51592 17923 51595
rect 17954 51592 17960 51604
rect 17911 51564 17960 51592
rect 17911 51561 17923 51564
rect 17865 51555 17923 51561
rect 17954 51552 17960 51564
rect 18012 51552 18018 51604
rect 19058 51592 19064 51604
rect 19019 51564 19064 51592
rect 19058 51552 19064 51564
rect 19116 51592 19122 51604
rect 19518 51592 19524 51604
rect 19116 51564 19524 51592
rect 19116 51552 19122 51564
rect 19518 51552 19524 51564
rect 19576 51552 19582 51604
rect 20441 51595 20499 51601
rect 20441 51561 20453 51595
rect 20487 51592 20499 51595
rect 21358 51592 21364 51604
rect 20487 51564 21364 51592
rect 20487 51561 20499 51564
rect 20441 51555 20499 51561
rect 21358 51552 21364 51564
rect 21416 51592 21422 51604
rect 23842 51592 23848 51604
rect 21416 51564 22048 51592
rect 21416 51552 21422 51564
rect 12161 51527 12219 51533
rect 12161 51493 12173 51527
rect 12207 51524 12219 51527
rect 13262 51524 13268 51536
rect 12207 51496 13268 51524
rect 12207 51493 12219 51496
rect 12161 51487 12219 51493
rect 13262 51484 13268 51496
rect 13320 51524 13326 51536
rect 13633 51527 13691 51533
rect 13633 51524 13645 51527
rect 13320 51496 13645 51524
rect 13320 51484 13326 51496
rect 13633 51493 13645 51496
rect 13679 51524 13691 51527
rect 13906 51524 13912 51536
rect 13679 51496 13912 51524
rect 13679 51493 13691 51496
rect 13633 51487 13691 51493
rect 13906 51484 13912 51496
rect 13964 51484 13970 51536
rect 14844 51524 14872 51552
rect 14918 51524 14924 51536
rect 14844 51496 14924 51524
rect 6089 51459 6147 51465
rect 6089 51425 6101 51459
rect 6135 51456 6147 51459
rect 6270 51456 6276 51468
rect 6135 51428 6276 51456
rect 6135 51425 6147 51428
rect 6089 51419 6147 51425
rect 6270 51416 6276 51428
rect 6328 51416 6334 51468
rect 10410 51416 10416 51468
rect 10468 51456 10474 51468
rect 10597 51459 10655 51465
rect 10597 51456 10609 51459
rect 10468 51428 10609 51456
rect 10468 51416 10474 51428
rect 10597 51425 10609 51428
rect 10643 51425 10655 51459
rect 10597 51419 10655 51425
rect 11609 51459 11667 51465
rect 11609 51425 11621 51459
rect 11655 51456 11667 51459
rect 12250 51456 12256 51468
rect 11655 51428 12256 51456
rect 11655 51425 11667 51428
rect 11609 51419 11667 51425
rect 12250 51416 12256 51428
rect 12308 51416 12314 51468
rect 12621 51459 12679 51465
rect 12621 51425 12633 51459
rect 12667 51456 12679 51459
rect 12710 51456 12716 51468
rect 12667 51428 12716 51456
rect 12667 51425 12679 51428
rect 12621 51419 12679 51425
rect 12710 51416 12716 51428
rect 12768 51416 12774 51468
rect 12986 51416 12992 51468
rect 13044 51456 13050 51468
rect 13780 51459 13838 51465
rect 13780 51456 13792 51459
rect 13044 51428 13792 51456
rect 13044 51416 13050 51428
rect 13780 51425 13792 51428
rect 13826 51456 13838 51459
rect 14844 51456 14872 51496
rect 14918 51484 14924 51496
rect 14976 51484 14982 51536
rect 15933 51527 15991 51533
rect 15933 51493 15945 51527
rect 15979 51524 15991 51527
rect 17034 51524 17040 51536
rect 15979 51496 17040 51524
rect 15979 51493 15991 51496
rect 15933 51487 15991 51493
rect 17034 51484 17040 51496
rect 17092 51484 17098 51536
rect 19426 51484 19432 51536
rect 19484 51524 19490 51536
rect 21726 51524 21732 51536
rect 19484 51496 21732 51524
rect 19484 51484 19490 51496
rect 21726 51484 21732 51496
rect 21784 51484 21790 51536
rect 13826 51428 14872 51456
rect 15105 51459 15163 51465
rect 13826 51425 13838 51428
rect 13780 51419 13838 51425
rect 15105 51425 15117 51459
rect 15151 51456 15163 51459
rect 16022 51456 16028 51468
rect 15151 51428 16028 51456
rect 15151 51425 15163 51428
rect 15105 51419 15163 51425
rect 16022 51416 16028 51428
rect 16080 51416 16086 51468
rect 16114 51416 16120 51468
rect 16172 51465 16178 51468
rect 16172 51459 16230 51465
rect 16172 51425 16184 51459
rect 16218 51456 16230 51459
rect 17497 51459 17555 51465
rect 16218 51428 16528 51456
rect 16218 51425 16230 51428
rect 16172 51419 16230 51425
rect 16172 51416 16178 51419
rect 12529 51391 12587 51397
rect 12529 51357 12541 51391
rect 12575 51388 12587 51391
rect 13004 51388 13032 51416
rect 13998 51388 14004 51400
rect 12575 51360 13032 51388
rect 13372 51360 14004 51388
rect 12575 51357 12587 51360
rect 12529 51351 12587 51357
rect 11514 51280 11520 51332
rect 11572 51320 11578 51332
rect 13372 51320 13400 51360
rect 13998 51348 14004 51360
rect 14056 51348 14062 51400
rect 14182 51348 14188 51400
rect 14240 51388 14246 51400
rect 15470 51388 15476 51400
rect 14240 51360 15476 51388
rect 14240 51348 14246 51360
rect 15470 51348 15476 51360
rect 15528 51348 15534 51400
rect 16298 51348 16304 51400
rect 16356 51388 16362 51400
rect 16393 51391 16451 51397
rect 16393 51388 16405 51391
rect 16356 51360 16405 51388
rect 16356 51348 16362 51360
rect 16393 51357 16405 51360
rect 16439 51357 16451 51391
rect 16500 51388 16528 51428
rect 17497 51425 17509 51459
rect 17543 51456 17555 51459
rect 17770 51456 17776 51468
rect 17543 51428 17776 51456
rect 17543 51425 17555 51428
rect 17497 51419 17555 51425
rect 17770 51416 17776 51428
rect 17828 51416 17834 51468
rect 18046 51456 18052 51468
rect 18007 51428 18052 51456
rect 18046 51416 18052 51428
rect 18104 51416 18110 51468
rect 18417 51459 18475 51465
rect 18417 51425 18429 51459
rect 18463 51456 18475 51459
rect 18598 51456 18604 51468
rect 18463 51428 18604 51456
rect 18463 51425 18475 51428
rect 18417 51419 18475 51425
rect 18598 51416 18604 51428
rect 18656 51416 18662 51468
rect 19334 51416 19340 51468
rect 19392 51456 19398 51468
rect 19521 51459 19579 51465
rect 19521 51456 19533 51459
rect 19392 51428 19533 51456
rect 19392 51416 19398 51428
rect 19521 51425 19533 51428
rect 19567 51425 19579 51459
rect 19521 51419 19579 51425
rect 20073 51459 20131 51465
rect 20073 51425 20085 51459
rect 20119 51456 20131 51459
rect 21542 51456 21548 51468
rect 20119 51428 21548 51456
rect 20119 51425 20131 51428
rect 20073 51419 20131 51425
rect 21542 51416 21548 51428
rect 21600 51416 21606 51468
rect 21910 51456 21916 51468
rect 21871 51428 21916 51456
rect 21910 51416 21916 51428
rect 21968 51416 21974 51468
rect 22020 51465 22048 51564
rect 23492 51564 23848 51592
rect 22094 51484 22100 51536
rect 22152 51484 22158 51536
rect 22005 51459 22063 51465
rect 22005 51425 22017 51459
rect 22051 51425 22063 51459
rect 22112 51456 22140 51484
rect 22373 51459 22431 51465
rect 22373 51456 22385 51459
rect 22112 51428 22385 51456
rect 22005 51419 22063 51425
rect 16666 51388 16672 51400
rect 16500 51360 16672 51388
rect 16393 51351 16451 51357
rect 16666 51348 16672 51360
rect 16724 51348 16730 51400
rect 18138 51348 18144 51400
rect 18196 51388 18202 51400
rect 18966 51388 18972 51400
rect 18196 51360 18972 51388
rect 18196 51348 18202 51360
rect 18966 51348 18972 51360
rect 19024 51348 19030 51400
rect 20346 51348 20352 51400
rect 20404 51388 20410 51400
rect 21453 51391 21511 51397
rect 21453 51388 21465 51391
rect 20404 51360 21465 51388
rect 20404 51348 20410 51360
rect 21453 51357 21465 51360
rect 21499 51357 21511 51391
rect 21928 51388 21956 51416
rect 22094 51388 22100 51400
rect 21928 51360 22100 51388
rect 21453 51351 21511 51357
rect 22094 51348 22100 51360
rect 22152 51348 22158 51400
rect 11572 51292 13400 51320
rect 11572 51280 11578 51292
rect 13446 51280 13452 51332
rect 13504 51320 13510 51332
rect 13541 51323 13599 51329
rect 13541 51320 13553 51323
rect 13504 51292 13553 51320
rect 13504 51280 13510 51292
rect 13541 51289 13553 51292
rect 13587 51320 13599 51323
rect 13909 51323 13967 51329
rect 13909 51320 13921 51323
rect 13587 51292 13921 51320
rect 13587 51289 13599 51292
rect 13541 51283 13599 51289
rect 13909 51289 13921 51292
rect 13955 51320 13967 51323
rect 16574 51320 16580 51332
rect 13955 51292 16580 51320
rect 13955 51289 13967 51292
rect 13909 51283 13967 51289
rect 5810 51212 5816 51264
rect 5868 51252 5874 51264
rect 5905 51255 5963 51261
rect 5905 51252 5917 51255
rect 5868 51224 5917 51252
rect 5868 51212 5874 51224
rect 5905 51221 5917 51224
rect 5951 51221 5963 51255
rect 5905 51215 5963 51221
rect 11793 51255 11851 51261
rect 11793 51221 11805 51255
rect 11839 51252 11851 51255
rect 11974 51252 11980 51264
rect 11839 51224 11980 51252
rect 11839 51221 11851 51224
rect 11793 51215 11851 51221
rect 11974 51212 11980 51224
rect 12032 51212 12038 51264
rect 12805 51255 12863 51261
rect 12805 51221 12817 51255
rect 12851 51252 12863 51255
rect 13078 51252 13084 51264
rect 12851 51224 13084 51252
rect 12851 51221 12863 51224
rect 12805 51215 12863 51221
rect 13078 51212 13084 51224
rect 13136 51212 13142 51264
rect 14274 51252 14280 51264
rect 14235 51224 14280 51252
rect 14274 51212 14280 51224
rect 14332 51212 14338 51264
rect 14826 51212 14832 51264
rect 14884 51252 14890 51264
rect 15105 51255 15163 51261
rect 15105 51252 15117 51255
rect 14884 51224 15117 51252
rect 14884 51212 14890 51224
rect 15105 51221 15117 51224
rect 15151 51221 15163 51255
rect 15105 51215 15163 51221
rect 15194 51212 15200 51264
rect 15252 51252 15258 51264
rect 16316 51261 16344 51292
rect 16574 51280 16580 51292
rect 16632 51280 16638 51332
rect 17034 51280 17040 51332
rect 17092 51320 17098 51332
rect 17586 51320 17592 51332
rect 17092 51292 17592 51320
rect 17092 51280 17098 51292
rect 17586 51280 17592 51292
rect 17644 51280 17650 51332
rect 19705 51323 19763 51329
rect 19705 51320 19717 51323
rect 19352 51292 19717 51320
rect 15473 51255 15531 51261
rect 15473 51252 15485 51255
rect 15252 51224 15485 51252
rect 15252 51212 15258 51224
rect 15473 51221 15485 51224
rect 15519 51221 15531 51255
rect 15473 51215 15531 51221
rect 16301 51255 16359 51261
rect 16301 51221 16313 51255
rect 16347 51221 16359 51255
rect 16301 51215 16359 51221
rect 16482 51212 16488 51264
rect 16540 51252 16546 51264
rect 17129 51255 17187 51261
rect 17129 51252 17141 51255
rect 16540 51224 17141 51252
rect 16540 51212 16546 51224
rect 17129 51221 17141 51224
rect 17175 51221 17187 51255
rect 17129 51215 17187 51221
rect 19150 51212 19156 51264
rect 19208 51252 19214 51264
rect 19352 51252 19380 51292
rect 19705 51289 19717 51292
rect 19751 51289 19763 51323
rect 19705 51283 19763 51289
rect 21542 51280 21548 51332
rect 21600 51320 21606 51332
rect 22204 51320 22232 51428
rect 22373 51425 22385 51428
rect 22419 51425 22431 51459
rect 22373 51419 22431 51425
rect 23017 51459 23075 51465
rect 23017 51425 23029 51459
rect 23063 51456 23075 51459
rect 23198 51456 23204 51468
rect 23063 51428 23204 51456
rect 23063 51425 23075 51428
rect 23017 51419 23075 51425
rect 23198 51416 23204 51428
rect 23256 51416 23262 51468
rect 23492 51456 23520 51564
rect 23842 51552 23848 51564
rect 23900 51552 23906 51604
rect 23934 51552 23940 51604
rect 23992 51592 23998 51604
rect 24489 51595 24547 51601
rect 24489 51592 24501 51595
rect 23992 51564 24501 51592
rect 23992 51552 23998 51564
rect 24489 51561 24501 51564
rect 24535 51561 24547 51595
rect 24489 51555 24547 51561
rect 25498 51552 25504 51604
rect 25556 51592 25562 51604
rect 25682 51592 25688 51604
rect 25556 51564 25688 51592
rect 25556 51552 25562 51564
rect 25682 51552 25688 51564
rect 25740 51552 25746 51604
rect 23750 51484 23756 51536
rect 23808 51524 23814 51536
rect 23808 51496 24256 51524
rect 23808 51484 23814 51496
rect 23400 51428 23520 51456
rect 24029 51459 24087 51465
rect 23106 51348 23112 51400
rect 23164 51388 23170 51400
rect 23290 51388 23296 51400
rect 23164 51360 23296 51388
rect 23164 51348 23170 51360
rect 23290 51348 23296 51360
rect 23348 51348 23354 51400
rect 21600 51292 22232 51320
rect 21600 51280 21606 51292
rect 19208 51224 19380 51252
rect 19429 51255 19487 51261
rect 19208 51212 19214 51224
rect 19429 51221 19441 51255
rect 19475 51252 19487 51255
rect 19978 51252 19984 51264
rect 19475 51224 19984 51252
rect 19475 51221 19487 51224
rect 19429 51215 19487 51221
rect 19978 51212 19984 51224
rect 20036 51212 20042 51264
rect 20993 51255 21051 51261
rect 20993 51221 21005 51255
rect 21039 51252 21051 51255
rect 21726 51252 21732 51264
rect 21039 51224 21732 51252
rect 21039 51221 21051 51224
rect 20993 51215 21051 51221
rect 21726 51212 21732 51224
rect 21784 51212 21790 51264
rect 23290 51212 23296 51264
rect 23348 51252 23354 51264
rect 23400 51252 23428 51428
rect 24029 51425 24041 51459
rect 24075 51456 24087 51459
rect 24118 51456 24124 51468
rect 24075 51428 24124 51456
rect 24075 51425 24087 51428
rect 24029 51419 24087 51425
rect 24118 51416 24124 51428
rect 24176 51416 24182 51468
rect 24228 51465 24256 51496
rect 24213 51459 24271 51465
rect 24213 51425 24225 51459
rect 24259 51425 24271 51459
rect 24213 51419 24271 51425
rect 23474 51348 23480 51400
rect 23532 51388 23538 51400
rect 23753 51391 23811 51397
rect 23753 51388 23765 51391
rect 23532 51360 23765 51388
rect 23532 51348 23538 51360
rect 23753 51357 23765 51360
rect 23799 51357 23811 51391
rect 23753 51351 23811 51357
rect 23842 51280 23848 51332
rect 23900 51320 23906 51332
rect 24026 51320 24032 51332
rect 23900 51292 24032 51320
rect 23900 51280 23906 51292
rect 24026 51280 24032 51292
rect 24084 51280 24090 51332
rect 23348 51224 23428 51252
rect 23348 51212 23354 51224
rect 24762 51212 24768 51264
rect 24820 51252 24826 51264
rect 24949 51255 25007 51261
rect 24949 51252 24961 51255
rect 24820 51224 24961 51252
rect 24820 51212 24826 51224
rect 24949 51221 24961 51224
rect 24995 51252 25007 51255
rect 25774 51252 25780 51264
rect 24995 51224 25780 51252
rect 24995 51221 25007 51224
rect 24949 51215 25007 51221
rect 25774 51212 25780 51224
rect 25832 51212 25838 51264
rect 1104 51162 28888 51184
rect 1104 51110 5982 51162
rect 6034 51110 6046 51162
rect 6098 51110 6110 51162
rect 6162 51110 6174 51162
rect 6226 51110 15982 51162
rect 16034 51110 16046 51162
rect 16098 51110 16110 51162
rect 16162 51110 16174 51162
rect 16226 51110 25982 51162
rect 26034 51110 26046 51162
rect 26098 51110 26110 51162
rect 26162 51110 26174 51162
rect 26226 51110 28888 51162
rect 1104 51088 28888 51110
rect 5997 51051 6055 51057
rect 5997 51017 6009 51051
rect 6043 51048 6055 51051
rect 6270 51048 6276 51060
rect 6043 51020 6276 51048
rect 6043 51017 6055 51020
rect 5997 51011 6055 51017
rect 6270 51008 6276 51020
rect 6328 51008 6334 51060
rect 10410 51048 10416 51060
rect 10371 51020 10416 51048
rect 10410 51008 10416 51020
rect 10468 51008 10474 51060
rect 11241 51051 11299 51057
rect 11241 51017 11253 51051
rect 11287 51048 11299 51051
rect 11882 51048 11888 51060
rect 11287 51020 11888 51048
rect 11287 51017 11299 51020
rect 11241 51011 11299 51017
rect 11882 51008 11888 51020
rect 11940 51008 11946 51060
rect 12250 51048 12256 51060
rect 12163 51020 12256 51048
rect 12250 51008 12256 51020
rect 12308 51048 12314 51060
rect 12986 51048 12992 51060
rect 12308 51020 12992 51048
rect 12308 51008 12314 51020
rect 12986 51008 12992 51020
rect 13044 51048 13050 51060
rect 13044 51020 13308 51048
rect 13044 51008 13050 51020
rect 11514 50980 11520 50992
rect 11475 50952 11520 50980
rect 11514 50940 11520 50952
rect 11572 50940 11578 50992
rect 13280 50921 13308 51020
rect 13998 51008 14004 51060
rect 14056 51048 14062 51060
rect 14277 51051 14335 51057
rect 14277 51048 14289 51051
rect 14056 51020 14289 51048
rect 14056 51008 14062 51020
rect 14277 51017 14289 51020
rect 14323 51048 14335 51051
rect 14737 51051 14795 51057
rect 14737 51048 14749 51051
rect 14323 51020 14749 51048
rect 14323 51017 14335 51020
rect 14277 51011 14335 51017
rect 13265 50915 13323 50921
rect 13265 50881 13277 50915
rect 13311 50881 13323 50915
rect 13446 50912 13452 50924
rect 13265 50875 13323 50881
rect 13372 50884 13452 50912
rect 11054 50804 11060 50856
rect 11112 50844 11118 50856
rect 11333 50847 11391 50853
rect 11333 50844 11345 50847
rect 11112 50816 11345 50844
rect 11112 50804 11118 50816
rect 11333 50813 11345 50816
rect 11379 50844 11391 50847
rect 11793 50847 11851 50853
rect 11793 50844 11805 50847
rect 11379 50816 11805 50844
rect 11379 50813 11391 50816
rect 11333 50807 11391 50813
rect 11793 50813 11805 50816
rect 11839 50844 11851 50847
rect 12805 50847 12863 50853
rect 12805 50844 12817 50847
rect 11839 50816 12817 50844
rect 11839 50813 11851 50816
rect 11793 50807 11851 50813
rect 12805 50813 12817 50816
rect 12851 50844 12863 50847
rect 13372 50844 13400 50884
rect 13446 50872 13452 50884
rect 13504 50872 13510 50924
rect 14568 50912 14596 51020
rect 14737 51017 14749 51020
rect 14783 51017 14795 51051
rect 14737 51011 14795 51017
rect 14918 51008 14924 51060
rect 14976 51057 14982 51060
rect 14976 51051 15025 51057
rect 14976 51017 14979 51051
rect 15013 51017 15025 51051
rect 14976 51011 15025 51017
rect 14976 51008 14982 51011
rect 17586 51008 17592 51060
rect 17644 51048 17650 51060
rect 18325 51051 18383 51057
rect 18325 51048 18337 51051
rect 17644 51020 18337 51048
rect 17644 51008 17650 51020
rect 18325 51017 18337 51020
rect 18371 51048 18383 51051
rect 18598 51048 18604 51060
rect 18371 51020 18604 51048
rect 18371 51017 18383 51020
rect 18325 51011 18383 51017
rect 18598 51008 18604 51020
rect 18656 51008 18662 51060
rect 19518 51008 19524 51060
rect 19576 51048 19582 51060
rect 19576 51020 19748 51048
rect 19576 51008 19582 51020
rect 14642 50940 14648 50992
rect 14700 50980 14706 50992
rect 15105 50983 15163 50989
rect 15105 50980 15117 50983
rect 14700 50952 15117 50980
rect 14700 50940 14706 50952
rect 15105 50949 15117 50952
rect 15151 50949 15163 50983
rect 16298 50980 16304 50992
rect 15105 50943 15163 50949
rect 15856 50952 16304 50980
rect 15856 50921 15884 50952
rect 16298 50940 16304 50952
rect 16356 50980 16362 50992
rect 16393 50983 16451 50989
rect 16393 50980 16405 50983
rect 16356 50952 16405 50980
rect 16356 50940 16362 50952
rect 16393 50949 16405 50952
rect 16439 50980 16451 50983
rect 19426 50980 19432 50992
rect 16439 50952 19432 50980
rect 16439 50949 16451 50952
rect 16393 50943 16451 50949
rect 19426 50940 19432 50952
rect 19484 50940 19490 50992
rect 15197 50915 15255 50921
rect 15197 50912 15209 50915
rect 14568 50884 15209 50912
rect 15197 50881 15209 50884
rect 15243 50912 15255 50915
rect 15841 50915 15899 50921
rect 15841 50912 15853 50915
rect 15243 50884 15853 50912
rect 15243 50881 15255 50884
rect 15197 50875 15255 50881
rect 15841 50881 15853 50884
rect 15887 50881 15899 50915
rect 15841 50875 15899 50881
rect 16209 50915 16267 50921
rect 16209 50881 16221 50915
rect 16255 50912 16267 50915
rect 17126 50912 17132 50924
rect 16255 50884 16712 50912
rect 17087 50884 17132 50912
rect 16255 50881 16267 50884
rect 16209 50875 16267 50881
rect 13538 50844 13544 50856
rect 12851 50816 13400 50844
rect 13499 50816 13544 50844
rect 12851 50813 12863 50816
rect 12805 50807 12863 50813
rect 13372 50776 13400 50816
rect 13538 50804 13544 50816
rect 13596 50804 13602 50856
rect 13906 50804 13912 50856
rect 13964 50844 13970 50856
rect 14829 50847 14887 50853
rect 14829 50844 14841 50847
rect 13964 50816 14841 50844
rect 13964 50804 13970 50816
rect 14829 50813 14841 50816
rect 14875 50844 14887 50847
rect 15102 50844 15108 50856
rect 14875 50816 15108 50844
rect 14875 50813 14887 50816
rect 14829 50807 14887 50813
rect 15102 50804 15108 50816
rect 15160 50804 15166 50856
rect 16574 50844 16580 50856
rect 16535 50816 16580 50844
rect 16574 50804 16580 50816
rect 16632 50804 16638 50856
rect 16684 50853 16712 50884
rect 17126 50872 17132 50884
rect 17184 50872 17190 50924
rect 19058 50872 19064 50924
rect 19116 50912 19122 50924
rect 19334 50912 19340 50924
rect 19116 50884 19340 50912
rect 19116 50872 19122 50884
rect 19334 50872 19340 50884
rect 19392 50872 19398 50924
rect 16669 50847 16727 50853
rect 16669 50813 16681 50847
rect 16715 50844 16727 50847
rect 16942 50844 16948 50856
rect 16715 50816 16948 50844
rect 16715 50813 16727 50816
rect 16669 50807 16727 50813
rect 16942 50804 16948 50816
rect 17000 50804 17006 50856
rect 18506 50804 18512 50856
rect 18564 50844 18570 50856
rect 19720 50853 19748 51020
rect 22094 51008 22100 51060
rect 22152 51048 22158 51060
rect 22189 51051 22247 51057
rect 22189 51048 22201 51051
rect 22152 51020 22201 51048
rect 22152 51008 22158 51020
rect 22189 51017 22201 51020
rect 22235 51017 22247 51051
rect 22189 51011 22247 51017
rect 22925 51051 22983 51057
rect 22925 51017 22937 51051
rect 22971 51048 22983 51051
rect 23474 51048 23480 51060
rect 22971 51020 23480 51048
rect 22971 51017 22983 51020
rect 22925 51011 22983 51017
rect 23474 51008 23480 51020
rect 23532 51008 23538 51060
rect 24302 51048 24308 51060
rect 24263 51020 24308 51048
rect 24302 51008 24308 51020
rect 24360 51008 24366 51060
rect 20806 50940 20812 50992
rect 20864 50980 20870 50992
rect 21450 50980 21456 50992
rect 20864 50952 21456 50980
rect 20864 50940 20870 50952
rect 21450 50940 21456 50952
rect 21508 50940 21514 50992
rect 23293 50983 23351 50989
rect 23293 50949 23305 50983
rect 23339 50980 23351 50983
rect 24118 50980 24124 50992
rect 23339 50952 24124 50980
rect 23339 50949 23351 50952
rect 23293 50943 23351 50949
rect 24118 50940 24124 50952
rect 24176 50940 24182 50992
rect 20349 50915 20407 50921
rect 20349 50881 20361 50915
rect 20395 50912 20407 50915
rect 20901 50915 20959 50921
rect 20901 50912 20913 50915
rect 20395 50884 20913 50912
rect 20395 50881 20407 50884
rect 20349 50875 20407 50881
rect 20901 50881 20913 50884
rect 20947 50881 20959 50915
rect 20901 50875 20959 50881
rect 21913 50915 21971 50921
rect 21913 50881 21925 50915
rect 21959 50912 21971 50915
rect 22002 50912 22008 50924
rect 21959 50884 22008 50912
rect 21959 50881 21971 50884
rect 21913 50875 21971 50881
rect 22002 50872 22008 50884
rect 22060 50872 22066 50924
rect 22554 50872 22560 50924
rect 22612 50912 22618 50924
rect 24397 50915 24455 50921
rect 22612 50884 23520 50912
rect 22612 50872 22618 50884
rect 19429 50847 19487 50853
rect 19429 50844 19441 50847
rect 18564 50816 19441 50844
rect 18564 50804 18570 50816
rect 19429 50813 19441 50816
rect 19475 50813 19487 50847
rect 19429 50807 19487 50813
rect 19705 50847 19763 50853
rect 19705 50813 19717 50847
rect 19751 50813 19763 50847
rect 19705 50807 19763 50813
rect 19889 50847 19947 50853
rect 19889 50813 19901 50847
rect 19935 50844 19947 50847
rect 19978 50844 19984 50856
rect 19935 50816 19984 50844
rect 19935 50813 19947 50816
rect 19889 50807 19947 50813
rect 13449 50779 13507 50785
rect 13449 50776 13461 50779
rect 13372 50748 13461 50776
rect 13449 50745 13461 50748
rect 13495 50745 13507 50779
rect 13449 50739 13507 50745
rect 13633 50779 13691 50785
rect 13633 50745 13645 50779
rect 13679 50745 13691 50779
rect 13633 50739 13691 50745
rect 14001 50779 14059 50785
rect 14001 50745 14013 50779
rect 14047 50776 14059 50779
rect 15286 50776 15292 50788
rect 14047 50748 15292 50776
rect 14047 50745 14059 50748
rect 14001 50739 14059 50745
rect 13173 50711 13231 50717
rect 13173 50677 13185 50711
rect 13219 50708 13231 50711
rect 13648 50708 13676 50739
rect 15286 50736 15292 50748
rect 15344 50736 15350 50788
rect 16592 50776 16620 50804
rect 17405 50779 17463 50785
rect 17405 50776 17417 50779
rect 16592 50748 17417 50776
rect 17405 50745 17417 50748
rect 17451 50776 17463 50779
rect 17773 50779 17831 50785
rect 17773 50776 17785 50779
rect 17451 50748 17785 50776
rect 17451 50745 17463 50748
rect 17405 50739 17463 50745
rect 17773 50745 17785 50748
rect 17819 50745 17831 50779
rect 17773 50739 17831 50745
rect 18877 50779 18935 50785
rect 18877 50745 18889 50779
rect 18923 50776 18935 50779
rect 19334 50776 19340 50788
rect 18923 50748 19340 50776
rect 18923 50745 18935 50748
rect 18877 50739 18935 50745
rect 19334 50736 19340 50748
rect 19392 50736 19398 50788
rect 14458 50708 14464 50720
rect 13219 50680 14464 50708
rect 13219 50677 13231 50680
rect 13173 50671 13231 50677
rect 14458 50668 14464 50680
rect 14516 50668 14522 50720
rect 15470 50708 15476 50720
rect 15431 50680 15476 50708
rect 15470 50668 15476 50680
rect 15528 50668 15534 50720
rect 18785 50711 18843 50717
rect 18785 50677 18797 50711
rect 18831 50708 18843 50711
rect 19058 50708 19064 50720
rect 18831 50680 19064 50708
rect 18831 50677 18843 50680
rect 18785 50671 18843 50677
rect 19058 50668 19064 50680
rect 19116 50668 19122 50720
rect 19426 50668 19432 50720
rect 19484 50708 19490 50720
rect 19904 50708 19932 50807
rect 19978 50804 19984 50816
rect 20036 50804 20042 50856
rect 21361 50847 21419 50853
rect 21361 50844 21373 50847
rect 20640 50816 21373 50844
rect 19484 50680 19932 50708
rect 19484 50668 19490 50680
rect 20438 50668 20444 50720
rect 20496 50708 20502 50720
rect 20640 50717 20668 50816
rect 21361 50813 21373 50816
rect 21407 50844 21419 50847
rect 21407 50816 22048 50844
rect 21407 50813 21419 50816
rect 21361 50807 21419 50813
rect 22020 50788 22048 50816
rect 23014 50804 23020 50856
rect 23072 50844 23078 50856
rect 23072 50816 23336 50844
rect 23072 50804 23078 50816
rect 20806 50736 20812 50788
rect 20864 50776 20870 50788
rect 20993 50779 21051 50785
rect 20993 50776 21005 50779
rect 20864 50748 21005 50776
rect 20864 50736 20870 50748
rect 20993 50745 21005 50748
rect 21039 50776 21051 50779
rect 21174 50776 21180 50788
rect 21039 50748 21180 50776
rect 21039 50745 21051 50748
rect 20993 50739 21051 50745
rect 21174 50736 21180 50748
rect 21232 50736 21238 50788
rect 21542 50776 21548 50788
rect 21503 50748 21548 50776
rect 21542 50736 21548 50748
rect 21600 50736 21606 50788
rect 22002 50736 22008 50788
rect 22060 50736 22066 50788
rect 23308 50720 23336 50816
rect 23492 50776 23520 50884
rect 24397 50881 24409 50915
rect 24443 50912 24455 50915
rect 24762 50912 24768 50924
rect 24443 50884 24768 50912
rect 24443 50881 24455 50884
rect 24397 50875 24455 50881
rect 24762 50872 24768 50884
rect 24820 50872 24826 50924
rect 23750 50844 23756 50856
rect 23711 50816 23756 50844
rect 23750 50804 23756 50816
rect 23808 50804 23814 50856
rect 24302 50804 24308 50856
rect 24360 50844 24366 50856
rect 24673 50847 24731 50853
rect 24673 50844 24685 50847
rect 24360 50816 24685 50844
rect 24360 50804 24366 50816
rect 24673 50813 24685 50816
rect 24719 50813 24731 50847
rect 24673 50807 24731 50813
rect 24486 50776 24492 50788
rect 23492 50748 24492 50776
rect 24486 50736 24492 50748
rect 24544 50736 24550 50788
rect 20625 50711 20683 50717
rect 20625 50708 20637 50711
rect 20496 50680 20637 50708
rect 20496 50668 20502 50680
rect 20625 50677 20637 50680
rect 20671 50677 20683 50711
rect 20625 50671 20683 50677
rect 20714 50668 20720 50720
rect 20772 50708 20778 50720
rect 20901 50711 20959 50717
rect 20901 50708 20913 50711
rect 20772 50680 20913 50708
rect 20772 50668 20778 50680
rect 20901 50677 20913 50680
rect 20947 50708 20959 50711
rect 21453 50711 21511 50717
rect 21453 50708 21465 50711
rect 20947 50680 21465 50708
rect 20947 50677 20959 50680
rect 20901 50671 20959 50677
rect 21453 50677 21465 50680
rect 21499 50677 21511 50711
rect 21453 50671 21511 50677
rect 22738 50668 22744 50720
rect 22796 50708 22802 50720
rect 23014 50708 23020 50720
rect 22796 50680 23020 50708
rect 22796 50668 22802 50680
rect 23014 50668 23020 50680
rect 23072 50668 23078 50720
rect 23290 50668 23296 50720
rect 23348 50668 23354 50720
rect 23753 50711 23811 50717
rect 23753 50677 23765 50711
rect 23799 50708 23811 50711
rect 23937 50711 23995 50717
rect 23937 50708 23949 50711
rect 23799 50680 23949 50708
rect 23799 50677 23811 50680
rect 23753 50671 23811 50677
rect 23937 50677 23949 50680
rect 23983 50708 23995 50711
rect 24302 50708 24308 50720
rect 23983 50680 24308 50708
rect 23983 50677 23995 50680
rect 23937 50671 23995 50677
rect 24302 50668 24308 50680
rect 24360 50668 24366 50720
rect 25130 50668 25136 50720
rect 25188 50708 25194 50720
rect 25777 50711 25835 50717
rect 25777 50708 25789 50711
rect 25188 50680 25789 50708
rect 25188 50668 25194 50680
rect 25777 50677 25789 50680
rect 25823 50677 25835 50711
rect 25777 50671 25835 50677
rect 1104 50618 28888 50640
rect 1104 50566 10982 50618
rect 11034 50566 11046 50618
rect 11098 50566 11110 50618
rect 11162 50566 11174 50618
rect 11226 50566 20982 50618
rect 21034 50566 21046 50618
rect 21098 50566 21110 50618
rect 21162 50566 21174 50618
rect 21226 50566 28888 50618
rect 1104 50544 28888 50566
rect 12621 50507 12679 50513
rect 12621 50473 12633 50507
rect 12667 50504 12679 50507
rect 12710 50504 12716 50516
rect 12667 50476 12716 50504
rect 12667 50473 12679 50476
rect 12621 50467 12679 50473
rect 12710 50464 12716 50476
rect 12768 50464 12774 50516
rect 12986 50504 12992 50516
rect 12947 50476 12992 50504
rect 12986 50464 12992 50476
rect 13044 50464 13050 50516
rect 13357 50507 13415 50513
rect 13357 50473 13369 50507
rect 13403 50504 13415 50507
rect 13538 50504 13544 50516
rect 13403 50476 13544 50504
rect 13403 50473 13415 50476
rect 13357 50467 13415 50473
rect 13538 50464 13544 50476
rect 13596 50464 13602 50516
rect 14642 50464 14648 50516
rect 14700 50504 14706 50516
rect 14829 50507 14887 50513
rect 14829 50504 14841 50507
rect 14700 50476 14841 50504
rect 14700 50464 14706 50476
rect 14829 50473 14841 50476
rect 14875 50473 14887 50507
rect 14829 50467 14887 50473
rect 15286 50464 15292 50516
rect 15344 50504 15350 50516
rect 15746 50504 15752 50516
rect 15344 50476 15752 50504
rect 15344 50464 15350 50476
rect 15746 50464 15752 50476
rect 15804 50464 15810 50516
rect 16298 50464 16304 50516
rect 16356 50504 16362 50516
rect 16485 50507 16543 50513
rect 16485 50504 16497 50507
rect 16356 50476 16497 50504
rect 16356 50464 16362 50476
rect 16485 50473 16497 50476
rect 16531 50473 16543 50507
rect 16485 50467 16543 50473
rect 16666 50464 16672 50516
rect 16724 50504 16730 50516
rect 16853 50507 16911 50513
rect 16853 50504 16865 50507
rect 16724 50476 16865 50504
rect 16724 50464 16730 50476
rect 16853 50473 16865 50476
rect 16899 50473 16911 50507
rect 18506 50504 18512 50516
rect 18467 50476 18512 50504
rect 16853 50467 16911 50473
rect 18506 50464 18512 50476
rect 18564 50464 18570 50516
rect 20346 50504 20352 50516
rect 20307 50476 20352 50504
rect 20346 50464 20352 50476
rect 20404 50464 20410 50516
rect 20717 50507 20775 50513
rect 20717 50473 20729 50507
rect 20763 50504 20775 50507
rect 21177 50507 21235 50513
rect 21177 50504 21189 50507
rect 20763 50476 21189 50504
rect 20763 50473 20775 50476
rect 20717 50467 20775 50473
rect 21177 50473 21189 50476
rect 21223 50504 21235 50507
rect 21266 50504 21272 50516
rect 21223 50476 21272 50504
rect 21223 50473 21235 50476
rect 21177 50467 21235 50473
rect 21266 50464 21272 50476
rect 21324 50464 21330 50516
rect 21450 50464 21456 50516
rect 21508 50504 21514 50516
rect 23477 50507 23535 50513
rect 23477 50504 23489 50507
rect 21508 50476 23489 50504
rect 21508 50464 21514 50476
rect 23477 50473 23489 50476
rect 23523 50473 23535 50507
rect 24302 50504 24308 50516
rect 24263 50476 24308 50504
rect 23477 50467 23535 50473
rect 24302 50464 24308 50476
rect 24360 50464 24366 50516
rect 12342 50396 12348 50448
rect 12400 50436 12406 50448
rect 14918 50436 14924 50448
rect 12400 50408 14924 50436
rect 12400 50396 12406 50408
rect 14918 50396 14924 50408
rect 14976 50436 14982 50448
rect 14976 50408 15148 50436
rect 14976 50396 14982 50408
rect 10413 50371 10471 50377
rect 10413 50337 10425 50371
rect 10459 50368 10471 50371
rect 10778 50368 10784 50380
rect 10459 50340 10784 50368
rect 10459 50337 10471 50340
rect 10413 50331 10471 50337
rect 10778 50328 10784 50340
rect 10836 50368 10842 50380
rect 11422 50368 11428 50380
rect 10836 50340 11428 50368
rect 10836 50328 10842 50340
rect 11422 50328 11428 50340
rect 11480 50328 11486 50380
rect 13909 50371 13967 50377
rect 13909 50337 13921 50371
rect 13955 50368 13967 50371
rect 13998 50368 14004 50380
rect 13955 50340 14004 50368
rect 13955 50337 13967 50340
rect 13909 50331 13967 50337
rect 13998 50328 14004 50340
rect 14056 50328 14062 50380
rect 14182 50368 14188 50380
rect 14143 50340 14188 50368
rect 14182 50328 14188 50340
rect 14240 50328 14246 50380
rect 15120 50368 15148 50408
rect 15194 50396 15200 50448
rect 15252 50436 15258 50448
rect 16209 50439 16267 50445
rect 16209 50436 16221 50439
rect 15252 50408 16221 50436
rect 15252 50396 15258 50408
rect 16209 50405 16221 50408
rect 16255 50405 16267 50439
rect 16209 50399 16267 50405
rect 17405 50439 17463 50445
rect 17405 50405 17417 50439
rect 17451 50436 17463 50439
rect 17494 50436 17500 50448
rect 17451 50408 17500 50436
rect 17451 50405 17463 50408
rect 17405 50399 17463 50405
rect 17494 50396 17500 50408
rect 17552 50396 17558 50448
rect 17770 50436 17776 50448
rect 17731 50408 17776 50436
rect 17770 50396 17776 50408
rect 17828 50396 17834 50448
rect 22002 50396 22008 50448
rect 22060 50436 22066 50448
rect 22462 50436 22468 50448
rect 22060 50408 22140 50436
rect 22423 50408 22468 50436
rect 22060 50396 22066 50408
rect 15657 50371 15715 50377
rect 15657 50368 15669 50371
rect 15120 50340 15669 50368
rect 15657 50337 15669 50340
rect 15703 50337 15715 50371
rect 15657 50331 15715 50337
rect 10689 50303 10747 50309
rect 10689 50269 10701 50303
rect 10735 50300 10747 50303
rect 10870 50300 10876 50312
rect 10735 50272 10876 50300
rect 10735 50269 10747 50272
rect 10689 50263 10747 50269
rect 10870 50260 10876 50272
rect 10928 50260 10934 50312
rect 14369 50303 14427 50309
rect 14369 50269 14381 50303
rect 14415 50300 14427 50303
rect 15102 50300 15108 50312
rect 14415 50272 15108 50300
rect 14415 50269 14427 50272
rect 14369 50263 14427 50269
rect 15102 50260 15108 50272
rect 15160 50260 15166 50312
rect 15672 50300 15700 50331
rect 15746 50328 15752 50380
rect 15804 50368 15810 50380
rect 17221 50371 17279 50377
rect 17221 50368 17233 50371
rect 15804 50340 15849 50368
rect 16960 50340 17233 50368
rect 15804 50328 15810 50340
rect 16482 50300 16488 50312
rect 15672 50272 16488 50300
rect 16482 50260 16488 50272
rect 16540 50300 16546 50312
rect 16666 50300 16672 50312
rect 16540 50272 16672 50300
rect 16540 50260 16546 50272
rect 16666 50260 16672 50272
rect 16724 50300 16730 50312
rect 16960 50300 16988 50340
rect 17221 50337 17233 50340
rect 17267 50337 17279 50371
rect 17221 50331 17279 50337
rect 17310 50328 17316 50380
rect 17368 50368 17374 50380
rect 17368 50340 17413 50368
rect 17368 50328 17374 50340
rect 17954 50328 17960 50380
rect 18012 50368 18018 50380
rect 18969 50371 19027 50377
rect 18969 50368 18981 50371
rect 18012 50340 18981 50368
rect 18012 50328 18018 50340
rect 18969 50337 18981 50340
rect 19015 50337 19027 50371
rect 18969 50331 19027 50337
rect 19334 50328 19340 50380
rect 19392 50368 19398 50380
rect 19429 50371 19487 50377
rect 19429 50368 19441 50371
rect 19392 50340 19441 50368
rect 19392 50328 19398 50340
rect 19429 50337 19441 50340
rect 19475 50337 19487 50371
rect 19429 50331 19487 50337
rect 21545 50371 21603 50377
rect 21545 50337 21557 50371
rect 21591 50337 21603 50371
rect 21545 50331 21603 50337
rect 16724 50272 16988 50300
rect 17037 50303 17095 50309
rect 16724 50260 16730 50272
rect 17037 50269 17049 50303
rect 17083 50269 17095 50303
rect 17037 50263 17095 50269
rect 11790 50164 11796 50176
rect 11751 50136 11796 50164
rect 11790 50124 11796 50136
rect 11848 50124 11854 50176
rect 15473 50167 15531 50173
rect 15473 50133 15485 50167
rect 15519 50164 15531 50167
rect 15746 50164 15752 50176
rect 15519 50136 15752 50164
rect 15519 50133 15531 50136
rect 15473 50127 15531 50133
rect 15746 50124 15752 50136
rect 15804 50164 15810 50176
rect 17052 50164 17080 50263
rect 18414 50260 18420 50312
rect 18472 50300 18478 50312
rect 18785 50303 18843 50309
rect 18785 50300 18797 50303
rect 18472 50272 18797 50300
rect 18472 50260 18478 50272
rect 18785 50269 18797 50272
rect 18831 50300 18843 50303
rect 19150 50300 19156 50312
rect 18831 50272 19156 50300
rect 18831 50269 18843 50272
rect 18785 50263 18843 50269
rect 19150 50260 19156 50272
rect 19208 50260 19214 50312
rect 19702 50300 19708 50312
rect 19663 50272 19708 50300
rect 19702 50260 19708 50272
rect 19760 50260 19766 50312
rect 20346 50260 20352 50312
rect 20404 50300 20410 50312
rect 21560 50300 21588 50331
rect 22002 50300 22008 50312
rect 20404 50272 22008 50300
rect 20404 50260 20410 50272
rect 22002 50260 22008 50272
rect 22060 50260 22066 50312
rect 22112 50300 22140 50408
rect 22462 50396 22468 50408
rect 22520 50396 22526 50448
rect 22830 50436 22836 50448
rect 22791 50408 22836 50436
rect 22830 50396 22836 50408
rect 22888 50396 22894 50448
rect 23198 50436 23204 50448
rect 23159 50408 23204 50436
rect 23198 50396 23204 50408
rect 23256 50396 23262 50448
rect 22186 50328 22192 50380
rect 22244 50368 22250 50380
rect 22649 50371 22707 50377
rect 22649 50368 22661 50371
rect 22244 50340 22661 50368
rect 22244 50328 22250 50340
rect 22649 50337 22661 50340
rect 22695 50337 22707 50371
rect 22649 50331 22707 50337
rect 22738 50328 22744 50380
rect 22796 50368 22802 50380
rect 24302 50368 24308 50380
rect 22796 50340 22841 50368
rect 24263 50340 24308 50368
rect 22796 50328 22802 50340
rect 24302 50328 24308 50340
rect 24360 50328 24366 50380
rect 22756 50300 22784 50328
rect 22112 50272 22784 50300
rect 18138 50164 18144 50176
rect 15804 50136 17080 50164
rect 18099 50136 18144 50164
rect 15804 50124 15810 50136
rect 18138 50124 18144 50136
rect 18196 50124 18202 50176
rect 21542 50124 21548 50176
rect 21600 50164 21606 50176
rect 21913 50167 21971 50173
rect 21913 50164 21925 50167
rect 21600 50136 21925 50164
rect 21600 50124 21606 50136
rect 21913 50133 21925 50136
rect 21959 50133 21971 50167
rect 22278 50164 22284 50176
rect 22239 50136 22284 50164
rect 21913 50127 21971 50133
rect 22278 50124 22284 50136
rect 22336 50124 22342 50176
rect 1104 50074 28888 50096
rect 1104 50022 5982 50074
rect 6034 50022 6046 50074
rect 6098 50022 6110 50074
rect 6162 50022 6174 50074
rect 6226 50022 15982 50074
rect 16034 50022 16046 50074
rect 16098 50022 16110 50074
rect 16162 50022 16174 50074
rect 16226 50022 25982 50074
rect 26034 50022 26046 50074
rect 26098 50022 26110 50074
rect 26162 50022 26174 50074
rect 26226 50022 28888 50074
rect 1104 50000 28888 50022
rect 8938 49960 8944 49972
rect 8899 49932 8944 49960
rect 8938 49920 8944 49932
rect 8996 49920 9002 49972
rect 9861 49963 9919 49969
rect 9861 49929 9873 49963
rect 9907 49960 9919 49963
rect 10870 49960 10876 49972
rect 9907 49932 10876 49960
rect 9907 49929 9919 49932
rect 9861 49923 9919 49929
rect 10870 49920 10876 49932
rect 10928 49960 10934 49972
rect 12250 49960 12256 49972
rect 10928 49932 11284 49960
rect 12211 49932 12256 49960
rect 10928 49920 10934 49932
rect 10229 49895 10287 49901
rect 10229 49861 10241 49895
rect 10275 49892 10287 49895
rect 10275 49864 11192 49892
rect 10275 49861 10287 49864
rect 10229 49855 10287 49861
rect 7374 49824 7380 49836
rect 7335 49796 7380 49824
rect 7374 49784 7380 49796
rect 7432 49784 7438 49836
rect 10318 49824 10324 49836
rect 10279 49796 10324 49824
rect 10318 49784 10324 49796
rect 10376 49784 10382 49836
rect 7653 49759 7711 49765
rect 7653 49756 7665 49759
rect 7208 49728 7665 49756
rect 7208 49632 7236 49728
rect 7653 49725 7665 49728
rect 7699 49725 7711 49759
rect 10778 49756 10784 49768
rect 10739 49728 10784 49756
rect 7653 49719 7711 49725
rect 10778 49716 10784 49728
rect 10836 49716 10842 49768
rect 11164 49765 11192 49864
rect 11256 49833 11284 49932
rect 12250 49920 12256 49932
rect 12308 49920 12314 49972
rect 12897 49963 12955 49969
rect 12897 49929 12909 49963
rect 12943 49960 12955 49963
rect 13446 49960 13452 49972
rect 12943 49932 13452 49960
rect 12943 49929 12955 49932
rect 12897 49923 12955 49929
rect 13446 49920 13452 49932
rect 13504 49960 13510 49972
rect 13998 49960 14004 49972
rect 13504 49932 14004 49960
rect 13504 49920 13510 49932
rect 13998 49920 14004 49932
rect 14056 49920 14062 49972
rect 15286 49920 15292 49972
rect 15344 49960 15350 49972
rect 15381 49963 15439 49969
rect 15381 49960 15393 49963
rect 15344 49932 15393 49960
rect 15344 49920 15350 49932
rect 15381 49929 15393 49932
rect 15427 49960 15439 49963
rect 17494 49960 17500 49972
rect 15427 49932 16528 49960
rect 17455 49932 17500 49960
rect 15427 49929 15439 49932
rect 15381 49923 15439 49929
rect 15562 49852 15568 49904
rect 15620 49892 15626 49904
rect 16393 49895 16451 49901
rect 16393 49892 16405 49895
rect 15620 49864 16405 49892
rect 15620 49852 15626 49864
rect 16393 49861 16405 49864
rect 16439 49861 16451 49895
rect 16393 49855 16451 49861
rect 11241 49827 11299 49833
rect 11241 49793 11253 49827
rect 11287 49824 11299 49827
rect 12158 49824 12164 49836
rect 11287 49796 12164 49824
rect 11287 49793 11299 49796
rect 11241 49787 11299 49793
rect 12158 49784 12164 49796
rect 12216 49784 12222 49836
rect 12802 49784 12808 49836
rect 12860 49824 12866 49836
rect 12989 49827 13047 49833
rect 12989 49824 13001 49827
rect 12860 49796 13001 49824
rect 12860 49784 12866 49796
rect 12989 49793 13001 49796
rect 13035 49793 13047 49827
rect 13262 49824 13268 49836
rect 13175 49796 13268 49824
rect 12989 49787 13047 49793
rect 13262 49784 13268 49796
rect 13320 49824 13326 49836
rect 13722 49824 13728 49836
rect 13320 49796 13728 49824
rect 13320 49784 13326 49796
rect 13722 49784 13728 49796
rect 13780 49784 13786 49836
rect 13906 49784 13912 49836
rect 13964 49824 13970 49836
rect 14369 49827 14427 49833
rect 14369 49824 14381 49827
rect 13964 49796 14381 49824
rect 13964 49784 13970 49796
rect 14369 49793 14381 49796
rect 14415 49793 14427 49827
rect 16500 49824 16528 49932
rect 17494 49920 17500 49932
rect 17552 49920 17558 49972
rect 17865 49963 17923 49969
rect 17865 49929 17877 49963
rect 17911 49960 17923 49963
rect 17954 49960 17960 49972
rect 17911 49932 17960 49960
rect 17911 49929 17923 49932
rect 17865 49923 17923 49929
rect 17954 49920 17960 49932
rect 18012 49920 18018 49972
rect 18414 49960 18420 49972
rect 18375 49932 18420 49960
rect 18414 49920 18420 49932
rect 18472 49920 18478 49972
rect 20257 49963 20315 49969
rect 20257 49929 20269 49963
rect 20303 49960 20315 49963
rect 20346 49960 20352 49972
rect 20303 49932 20352 49960
rect 20303 49929 20315 49932
rect 20257 49923 20315 49929
rect 20346 49920 20352 49932
rect 20404 49920 20410 49972
rect 22186 49960 22192 49972
rect 22147 49932 22192 49960
rect 22186 49920 22192 49932
rect 22244 49920 22250 49972
rect 22462 49960 22468 49972
rect 22423 49932 22468 49960
rect 22462 49920 22468 49932
rect 22520 49920 22526 49972
rect 22738 49920 22744 49972
rect 22796 49960 22802 49972
rect 22833 49963 22891 49969
rect 22833 49960 22845 49963
rect 22796 49932 22845 49960
rect 22796 49920 22802 49932
rect 22833 49929 22845 49932
rect 22879 49929 22891 49963
rect 22833 49923 22891 49929
rect 23477 49963 23535 49969
rect 23477 49929 23489 49963
rect 23523 49960 23535 49963
rect 23566 49960 23572 49972
rect 23523 49932 23572 49960
rect 23523 49929 23535 49932
rect 23477 49923 23535 49929
rect 23566 49920 23572 49932
rect 23624 49920 23630 49972
rect 16850 49852 16856 49904
rect 16908 49892 16914 49904
rect 17037 49895 17095 49901
rect 17037 49892 17049 49895
rect 16908 49864 17049 49892
rect 16908 49852 16914 49864
rect 17037 49861 17049 49864
rect 17083 49892 17095 49895
rect 17310 49892 17316 49904
rect 17083 49864 17316 49892
rect 17083 49861 17095 49864
rect 17037 49855 17095 49861
rect 17310 49852 17316 49864
rect 17368 49852 17374 49904
rect 18874 49852 18880 49904
rect 18932 49892 18938 49904
rect 20898 49892 20904 49904
rect 18932 49864 20904 49892
rect 18932 49852 18938 49864
rect 20898 49852 20904 49864
rect 20956 49852 20962 49904
rect 22002 49852 22008 49904
rect 22060 49892 22066 49904
rect 25409 49895 25467 49901
rect 25409 49892 25421 49895
rect 22060 49864 25421 49892
rect 22060 49852 22066 49864
rect 25409 49861 25421 49864
rect 25455 49861 25467 49895
rect 25409 49855 25467 49861
rect 16500 49796 16620 49824
rect 14369 49787 14427 49793
rect 11149 49759 11207 49765
rect 11149 49725 11161 49759
rect 11195 49756 11207 49759
rect 11698 49756 11704 49768
rect 11195 49728 11704 49756
rect 11195 49725 11207 49728
rect 11149 49719 11207 49725
rect 11698 49716 11704 49728
rect 11756 49716 11762 49768
rect 14642 49716 14648 49768
rect 14700 49756 14706 49768
rect 14921 49759 14979 49765
rect 14921 49756 14933 49759
rect 14700 49728 14933 49756
rect 14700 49716 14706 49728
rect 14921 49725 14933 49728
rect 14967 49756 14979 49759
rect 15286 49756 15292 49768
rect 14967 49728 15292 49756
rect 14967 49725 14979 49728
rect 14921 49719 14979 49725
rect 15286 49716 15292 49728
rect 15344 49756 15350 49768
rect 15473 49759 15531 49765
rect 15473 49756 15485 49759
rect 15344 49728 15485 49756
rect 15344 49716 15350 49728
rect 15473 49725 15485 49728
rect 15519 49725 15531 49759
rect 16022 49756 16028 49768
rect 15983 49728 16028 49756
rect 15473 49719 15531 49725
rect 16022 49716 16028 49728
rect 16080 49716 16086 49768
rect 16393 49759 16451 49765
rect 16393 49725 16405 49759
rect 16439 49756 16451 49759
rect 16482 49756 16488 49768
rect 16439 49728 16488 49756
rect 16439 49725 16451 49728
rect 16393 49719 16451 49725
rect 16482 49716 16488 49728
rect 16540 49716 16546 49768
rect 15010 49648 15016 49700
rect 15068 49688 15074 49700
rect 16040 49688 16068 49716
rect 15068 49660 16068 49688
rect 16592 49688 16620 49796
rect 18138 49784 18144 49836
rect 18196 49824 18202 49836
rect 19334 49824 19340 49836
rect 18196 49796 19340 49824
rect 18196 49784 18202 49796
rect 19334 49784 19340 49796
rect 19392 49824 19398 49836
rect 19392 49796 19472 49824
rect 19392 49784 19398 49796
rect 17770 49716 17776 49768
rect 17828 49756 17834 49768
rect 18690 49756 18696 49768
rect 17828 49728 18696 49756
rect 17828 49716 17834 49728
rect 18690 49716 18696 49728
rect 18748 49716 18754 49768
rect 18966 49756 18972 49768
rect 18927 49728 18972 49756
rect 18966 49716 18972 49728
rect 19024 49716 19030 49768
rect 19444 49765 19472 49796
rect 22554 49784 22560 49836
rect 22612 49824 22618 49836
rect 22738 49824 22744 49836
rect 22612 49796 22744 49824
rect 22612 49784 22618 49796
rect 22738 49784 22744 49796
rect 22796 49784 22802 49836
rect 23198 49784 23204 49836
rect 23256 49824 23262 49836
rect 24397 49827 24455 49833
rect 24397 49824 24409 49827
rect 23256 49796 24409 49824
rect 23256 49784 23262 49796
rect 24397 49793 24409 49796
rect 24443 49824 24455 49827
rect 24486 49824 24492 49836
rect 24443 49796 24492 49824
rect 24443 49793 24455 49796
rect 24397 49787 24455 49793
rect 24486 49784 24492 49796
rect 24544 49784 24550 49836
rect 19429 49759 19487 49765
rect 19429 49725 19441 49759
rect 19475 49725 19487 49759
rect 19429 49719 19487 49725
rect 20438 49716 20444 49768
rect 20496 49756 20502 49768
rect 20533 49759 20591 49765
rect 20533 49756 20545 49759
rect 20496 49728 20545 49756
rect 20496 49716 20502 49728
rect 20533 49725 20545 49728
rect 20579 49756 20591 49759
rect 21269 49759 21327 49765
rect 21269 49756 21281 49759
rect 20579 49728 21281 49756
rect 20579 49725 20591 49728
rect 20533 49719 20591 49725
rect 21269 49725 21281 49728
rect 21315 49725 21327 49759
rect 21269 49719 21327 49725
rect 23566 49716 23572 49768
rect 23624 49756 23630 49768
rect 23753 49759 23811 49765
rect 23753 49756 23765 49759
rect 23624 49728 23765 49756
rect 23624 49716 23630 49728
rect 23753 49725 23765 49728
rect 23799 49725 23811 49759
rect 23753 49719 23811 49725
rect 24302 49716 24308 49768
rect 24360 49756 24366 49768
rect 24673 49759 24731 49765
rect 24673 49756 24685 49759
rect 24360 49728 24685 49756
rect 24360 49716 24366 49728
rect 24673 49725 24685 49728
rect 24719 49725 24731 49759
rect 24673 49719 24731 49725
rect 25225 49759 25283 49765
rect 25225 49725 25237 49759
rect 25271 49725 25283 49759
rect 25225 49719 25283 49725
rect 17310 49688 17316 49700
rect 16592 49660 17316 49688
rect 15068 49648 15074 49660
rect 17310 49648 17316 49660
rect 17368 49648 17374 49700
rect 19518 49648 19524 49700
rect 19576 49688 19582 49700
rect 19613 49691 19671 49697
rect 19613 49688 19625 49691
rect 19576 49660 19625 49688
rect 19576 49648 19582 49660
rect 19613 49657 19625 49660
rect 19659 49657 19671 49691
rect 19613 49651 19671 49657
rect 20806 49648 20812 49700
rect 20864 49688 20870 49700
rect 20901 49691 20959 49697
rect 20901 49688 20913 49691
rect 20864 49660 20913 49688
rect 20864 49648 20870 49660
rect 20901 49657 20913 49660
rect 20947 49688 20959 49691
rect 21085 49691 21143 49697
rect 21085 49688 21097 49691
rect 20947 49660 21097 49688
rect 20947 49657 20959 49660
rect 20901 49651 20959 49657
rect 21085 49657 21097 49660
rect 21131 49657 21143 49691
rect 21450 49688 21456 49700
rect 21411 49660 21456 49688
rect 21085 49651 21143 49657
rect 21450 49648 21456 49660
rect 21508 49648 21514 49700
rect 21821 49691 21879 49697
rect 21821 49657 21833 49691
rect 21867 49657 21879 49691
rect 21821 49651 21879 49657
rect 7190 49620 7196 49632
rect 7151 49592 7196 49620
rect 7190 49580 7196 49592
rect 7248 49580 7254 49632
rect 11422 49580 11428 49632
rect 11480 49620 11486 49632
rect 11793 49623 11851 49629
rect 11793 49620 11805 49623
rect 11480 49592 11805 49620
rect 11480 49580 11486 49592
rect 11793 49589 11805 49592
rect 11839 49589 11851 49623
rect 11793 49583 11851 49589
rect 20714 49580 20720 49632
rect 20772 49620 20778 49632
rect 21266 49620 21272 49632
rect 20772 49592 21272 49620
rect 20772 49580 20778 49592
rect 21266 49580 21272 49592
rect 21324 49620 21330 49632
rect 21361 49623 21419 49629
rect 21361 49620 21373 49623
rect 21324 49592 21373 49620
rect 21324 49580 21330 49592
rect 21361 49589 21373 49592
rect 21407 49589 21419 49623
rect 21836 49620 21864 49651
rect 25240 49632 25268 49719
rect 22370 49620 22376 49632
rect 21836 49592 22376 49620
rect 21361 49583 21419 49589
rect 22370 49580 22376 49592
rect 22428 49580 22434 49632
rect 25222 49580 25228 49632
rect 25280 49620 25286 49632
rect 25685 49623 25743 49629
rect 25685 49620 25697 49623
rect 25280 49592 25697 49620
rect 25280 49580 25286 49592
rect 25685 49589 25697 49592
rect 25731 49589 25743 49623
rect 25685 49583 25743 49589
rect 1104 49530 28888 49552
rect 1104 49478 10982 49530
rect 11034 49478 11046 49530
rect 11098 49478 11110 49530
rect 11162 49478 11174 49530
rect 11226 49478 20982 49530
rect 21034 49478 21046 49530
rect 21098 49478 21110 49530
rect 21162 49478 21174 49530
rect 21226 49478 28888 49530
rect 1104 49456 28888 49478
rect 7374 49416 7380 49428
rect 7335 49388 7380 49416
rect 7374 49376 7380 49388
rect 7432 49376 7438 49428
rect 10781 49419 10839 49425
rect 10781 49385 10793 49419
rect 10827 49416 10839 49419
rect 10870 49416 10876 49428
rect 10827 49388 10876 49416
rect 10827 49385 10839 49388
rect 10781 49379 10839 49385
rect 10870 49376 10876 49388
rect 10928 49376 10934 49428
rect 12621 49419 12679 49425
rect 12621 49385 12633 49419
rect 12667 49416 12679 49419
rect 13262 49416 13268 49428
rect 12667 49388 13268 49416
rect 12667 49385 12679 49388
rect 12621 49379 12679 49385
rect 13262 49376 13268 49388
rect 13320 49376 13326 49428
rect 14737 49419 14795 49425
rect 14737 49385 14749 49419
rect 14783 49416 14795 49419
rect 16482 49416 16488 49428
rect 14783 49388 16488 49416
rect 14783 49385 14795 49388
rect 14737 49379 14795 49385
rect 16482 49376 16488 49388
rect 16540 49376 16546 49428
rect 17770 49416 17776 49428
rect 17731 49388 17776 49416
rect 17770 49376 17776 49388
rect 17828 49376 17834 49428
rect 18138 49416 18144 49428
rect 18099 49388 18144 49416
rect 18138 49376 18144 49388
rect 18196 49376 18202 49428
rect 18506 49376 18512 49428
rect 18564 49416 18570 49428
rect 19794 49416 19800 49428
rect 18564 49388 19800 49416
rect 18564 49376 18570 49388
rect 19794 49376 19800 49388
rect 19852 49416 19858 49428
rect 19981 49419 20039 49425
rect 19981 49416 19993 49419
rect 19852 49388 19993 49416
rect 19852 49376 19858 49388
rect 19981 49385 19993 49388
rect 20027 49385 20039 49419
rect 21266 49416 21272 49428
rect 19981 49379 20039 49385
rect 20916 49388 21272 49416
rect 14918 49308 14924 49360
rect 14976 49348 14982 49360
rect 15013 49351 15071 49357
rect 15013 49348 15025 49351
rect 14976 49320 15025 49348
rect 14976 49308 14982 49320
rect 15013 49317 15025 49320
rect 15059 49317 15071 49351
rect 15013 49311 15071 49317
rect 15746 49308 15752 49360
rect 15804 49348 15810 49360
rect 15841 49351 15899 49357
rect 15841 49348 15853 49351
rect 15804 49320 15853 49348
rect 15804 49308 15810 49320
rect 15841 49317 15853 49320
rect 15887 49348 15899 49351
rect 16209 49351 16267 49357
rect 16209 49348 16221 49351
rect 15887 49320 16221 49348
rect 15887 49317 15899 49320
rect 15841 49311 15899 49317
rect 16209 49317 16221 49320
rect 16255 49348 16267 49351
rect 16298 49348 16304 49360
rect 16255 49320 16304 49348
rect 16255 49317 16267 49320
rect 16209 49311 16267 49317
rect 16298 49308 16304 49320
rect 16356 49308 16362 49360
rect 17586 49348 17592 49360
rect 16684 49320 17592 49348
rect 11425 49283 11483 49289
rect 11425 49249 11437 49283
rect 11471 49280 11483 49283
rect 11790 49280 11796 49292
rect 11471 49252 11796 49280
rect 11471 49249 11483 49252
rect 11425 49243 11483 49249
rect 11790 49240 11796 49252
rect 11848 49240 11854 49292
rect 12250 49240 12256 49292
rect 12308 49280 12314 49292
rect 12989 49283 13047 49289
rect 12989 49280 13001 49283
rect 12308 49252 13001 49280
rect 12308 49240 12314 49252
rect 12989 49249 13001 49252
rect 13035 49280 13047 49283
rect 13722 49280 13728 49292
rect 13035 49252 13728 49280
rect 13035 49249 13047 49252
rect 12989 49243 13047 49249
rect 13722 49240 13728 49252
rect 13780 49240 13786 49292
rect 15286 49240 15292 49292
rect 15344 49280 15350 49292
rect 15381 49283 15439 49289
rect 15381 49280 15393 49283
rect 15344 49252 15393 49280
rect 15344 49240 15350 49252
rect 15381 49249 15393 49252
rect 15427 49249 15439 49283
rect 15381 49243 15439 49249
rect 16574 49240 16580 49292
rect 16632 49280 16638 49292
rect 16684 49289 16712 49320
rect 17586 49308 17592 49320
rect 17644 49308 17650 49360
rect 16669 49283 16727 49289
rect 16669 49280 16681 49283
rect 16632 49252 16681 49280
rect 16632 49240 16638 49252
rect 16669 49249 16681 49252
rect 16715 49249 16727 49283
rect 16850 49280 16856 49292
rect 16811 49252 16856 49280
rect 16669 49243 16727 49249
rect 16850 49240 16856 49252
rect 16908 49240 16914 49292
rect 17218 49280 17224 49292
rect 17179 49252 17224 49280
rect 17218 49240 17224 49252
rect 17276 49240 17282 49292
rect 17954 49240 17960 49292
rect 18012 49280 18018 49292
rect 18877 49283 18935 49289
rect 18877 49280 18889 49283
rect 18012 49252 18889 49280
rect 18012 49240 18018 49252
rect 18877 49249 18889 49252
rect 18923 49249 18935 49283
rect 18877 49243 18935 49249
rect 18966 49240 18972 49292
rect 19024 49280 19030 49292
rect 19153 49283 19211 49289
rect 19153 49280 19165 49283
rect 19024 49252 19165 49280
rect 19024 49240 19030 49252
rect 19153 49249 19165 49252
rect 19199 49280 19211 49283
rect 19426 49280 19432 49292
rect 19199 49252 19432 49280
rect 19199 49249 19211 49252
rect 19153 49243 19211 49249
rect 19426 49240 19432 49252
rect 19484 49280 19490 49292
rect 19613 49283 19671 49289
rect 19613 49280 19625 49283
rect 19484 49252 19625 49280
rect 19484 49240 19490 49252
rect 19613 49249 19625 49252
rect 19659 49249 19671 49283
rect 19613 49243 19671 49249
rect 20346 49240 20352 49292
rect 20404 49280 20410 49292
rect 20916 49289 20944 49388
rect 21266 49376 21272 49388
rect 21324 49416 21330 49428
rect 21361 49419 21419 49425
rect 21361 49416 21373 49419
rect 21324 49388 21373 49416
rect 21324 49376 21330 49388
rect 21361 49385 21373 49388
rect 21407 49385 21419 49419
rect 21361 49379 21419 49385
rect 21545 49351 21603 49357
rect 21545 49317 21557 49351
rect 21591 49348 21603 49351
rect 21910 49348 21916 49360
rect 21591 49320 21916 49348
rect 21591 49317 21603 49320
rect 21545 49311 21603 49317
rect 21910 49308 21916 49320
rect 21968 49348 21974 49360
rect 23934 49348 23940 49360
rect 21968 49320 23940 49348
rect 21968 49308 21974 49320
rect 23934 49308 23940 49320
rect 23992 49308 23998 49360
rect 20901 49283 20959 49289
rect 20901 49280 20913 49283
rect 20404 49252 20913 49280
rect 20404 49240 20410 49252
rect 20901 49249 20913 49252
rect 20947 49249 20959 49283
rect 22370 49280 22376 49292
rect 22331 49252 22376 49280
rect 20901 49243 20959 49249
rect 22370 49240 22376 49252
rect 22428 49240 22434 49292
rect 22554 49280 22560 49292
rect 22515 49252 22560 49280
rect 22554 49240 22560 49252
rect 22612 49240 22618 49292
rect 22741 49283 22799 49289
rect 22741 49249 22753 49283
rect 22787 49280 22799 49283
rect 23661 49283 23719 49289
rect 23661 49280 23673 49283
rect 22787 49252 23673 49280
rect 22787 49249 22799 49252
rect 22741 49243 22799 49249
rect 23661 49249 23673 49252
rect 23707 49280 23719 49283
rect 24762 49280 24768 49292
rect 23707 49252 24768 49280
rect 23707 49249 23719 49252
rect 23661 49243 23719 49249
rect 24762 49240 24768 49252
rect 24820 49280 24826 49292
rect 25130 49280 25136 49292
rect 24820 49252 25136 49280
rect 24820 49240 24826 49252
rect 25130 49240 25136 49252
rect 25188 49240 25194 49292
rect 11330 49212 11336 49224
rect 11291 49184 11336 49212
rect 11330 49172 11336 49184
rect 11388 49172 11394 49224
rect 11514 49172 11520 49224
rect 11572 49212 11578 49224
rect 12710 49212 12716 49224
rect 11572 49184 12716 49212
rect 11572 49172 11578 49184
rect 12710 49172 12716 49184
rect 12768 49172 12774 49224
rect 18138 49172 18144 49224
rect 18196 49212 18202 49224
rect 18325 49215 18383 49221
rect 18325 49212 18337 49215
rect 18196 49184 18337 49212
rect 18196 49172 18202 49184
rect 18325 49181 18337 49184
rect 18371 49181 18383 49215
rect 18325 49175 18383 49181
rect 18414 49172 18420 49224
rect 18472 49212 18478 49224
rect 19334 49212 19340 49224
rect 18472 49184 19340 49212
rect 18472 49172 18478 49184
rect 19334 49172 19340 49184
rect 19392 49172 19398 49224
rect 23934 49172 23940 49224
rect 23992 49212 23998 49224
rect 24394 49212 24400 49224
rect 23992 49184 24400 49212
rect 23992 49172 23998 49184
rect 24394 49172 24400 49184
rect 24452 49172 24458 49224
rect 10413 49147 10471 49153
rect 10413 49113 10425 49147
rect 10459 49144 10471 49147
rect 10778 49144 10784 49156
rect 10459 49116 10784 49144
rect 10459 49113 10471 49116
rect 10413 49107 10471 49113
rect 10778 49104 10784 49116
rect 10836 49144 10842 49156
rect 21085 49147 21143 49153
rect 10836 49116 11652 49144
rect 10836 49104 10842 49116
rect 11149 49079 11207 49085
rect 11149 49045 11161 49079
rect 11195 49076 11207 49079
rect 11422 49076 11428 49088
rect 11195 49048 11428 49076
rect 11195 49045 11207 49048
rect 11149 49039 11207 49045
rect 11422 49036 11428 49048
rect 11480 49036 11486 49088
rect 11624 49085 11652 49116
rect 21085 49113 21097 49147
rect 21131 49144 21143 49147
rect 21545 49147 21603 49153
rect 21545 49144 21557 49147
rect 21131 49116 21557 49144
rect 21131 49113 21143 49116
rect 21085 49107 21143 49113
rect 21545 49113 21557 49116
rect 21591 49113 21603 49147
rect 21545 49107 21603 49113
rect 21634 49104 21640 49156
rect 21692 49144 21698 49156
rect 21729 49147 21787 49153
rect 21729 49144 21741 49147
rect 21692 49116 21741 49144
rect 21692 49104 21698 49116
rect 21729 49113 21741 49116
rect 21775 49113 21787 49147
rect 21729 49107 21787 49113
rect 11609 49079 11667 49085
rect 11609 49045 11621 49079
rect 11655 49045 11667 49079
rect 11609 49039 11667 49045
rect 13906 49036 13912 49088
rect 13964 49076 13970 49088
rect 14093 49079 14151 49085
rect 14093 49076 14105 49079
rect 13964 49048 14105 49076
rect 13964 49036 13970 49048
rect 14093 49045 14105 49048
rect 14139 49045 14151 49079
rect 14093 49039 14151 49045
rect 14826 49036 14832 49088
rect 14884 49076 14890 49088
rect 15286 49076 15292 49088
rect 14884 49048 15292 49076
rect 14884 49036 14890 49048
rect 15286 49036 15292 49048
rect 15344 49036 15350 49088
rect 15565 49079 15623 49085
rect 15565 49045 15577 49079
rect 15611 49076 15623 49079
rect 15654 49076 15660 49088
rect 15611 49048 15660 49076
rect 15611 49045 15623 49048
rect 15565 49039 15623 49045
rect 15654 49036 15660 49048
rect 15712 49036 15718 49088
rect 19058 49036 19064 49088
rect 19116 49076 19122 49088
rect 19334 49076 19340 49088
rect 19116 49048 19340 49076
rect 19116 49036 19122 49048
rect 19334 49036 19340 49048
rect 19392 49036 19398 49088
rect 19978 49036 19984 49088
rect 20036 49076 20042 49088
rect 20625 49079 20683 49085
rect 20625 49076 20637 49079
rect 20036 49048 20637 49076
rect 20036 49036 20042 49048
rect 20625 49045 20637 49048
rect 20671 49045 20683 49079
rect 21744 49076 21772 49107
rect 22094 49104 22100 49156
rect 22152 49144 22158 49156
rect 22189 49147 22247 49153
rect 22189 49144 22201 49147
rect 22152 49116 22201 49144
rect 22152 49104 22158 49116
rect 22189 49113 22201 49116
rect 22235 49113 22247 49147
rect 22189 49107 22247 49113
rect 22830 49076 22836 49088
rect 21744 49048 22836 49076
rect 20625 49039 20683 49045
rect 22830 49036 22836 49048
rect 22888 49076 22894 49088
rect 23201 49079 23259 49085
rect 23201 49076 23213 49079
rect 22888 49048 23213 49076
rect 22888 49036 22894 49048
rect 23201 49045 23213 49048
rect 23247 49045 23259 49079
rect 23201 49039 23259 49045
rect 23474 49036 23480 49088
rect 23532 49076 23538 49088
rect 23937 49079 23995 49085
rect 23937 49076 23949 49079
rect 23532 49048 23949 49076
rect 23532 49036 23538 49048
rect 23937 49045 23949 49048
rect 23983 49045 23995 49079
rect 24394 49076 24400 49088
rect 24355 49048 24400 49076
rect 23937 49039 23995 49045
rect 24394 49036 24400 49048
rect 24452 49036 24458 49088
rect 1104 48986 28888 49008
rect 1104 48934 5982 48986
rect 6034 48934 6046 48986
rect 6098 48934 6110 48986
rect 6162 48934 6174 48986
rect 6226 48934 15982 48986
rect 16034 48934 16046 48986
rect 16098 48934 16110 48986
rect 16162 48934 16174 48986
rect 16226 48934 25982 48986
rect 26034 48934 26046 48986
rect 26098 48934 26110 48986
rect 26162 48934 26174 48986
rect 26226 48934 28888 48986
rect 1104 48912 28888 48934
rect 11790 48872 11796 48884
rect 11751 48844 11796 48872
rect 11790 48832 11796 48844
rect 11848 48832 11854 48884
rect 12250 48872 12256 48884
rect 12211 48844 12256 48872
rect 12250 48832 12256 48844
rect 12308 48832 12314 48884
rect 12894 48832 12900 48884
rect 12952 48872 12958 48884
rect 13081 48875 13139 48881
rect 13081 48872 13093 48875
rect 12952 48844 13093 48872
rect 12952 48832 12958 48844
rect 13081 48841 13093 48844
rect 13127 48841 13139 48875
rect 13538 48872 13544 48884
rect 13499 48844 13544 48872
rect 13081 48835 13139 48841
rect 13538 48832 13544 48844
rect 13596 48832 13602 48884
rect 15194 48832 15200 48884
rect 15252 48872 15258 48884
rect 16025 48875 16083 48881
rect 16025 48872 16037 48875
rect 15252 48844 16037 48872
rect 15252 48832 15258 48844
rect 16025 48841 16037 48844
rect 16071 48872 16083 48875
rect 16850 48872 16856 48884
rect 16071 48844 16856 48872
rect 16071 48841 16083 48844
rect 16025 48835 16083 48841
rect 16850 48832 16856 48844
rect 16908 48832 16914 48884
rect 17865 48875 17923 48881
rect 17865 48841 17877 48875
rect 17911 48872 17923 48875
rect 18414 48872 18420 48884
rect 17911 48844 18420 48872
rect 17911 48841 17923 48844
rect 17865 48835 17923 48841
rect 18414 48832 18420 48844
rect 18472 48832 18478 48884
rect 19426 48872 19432 48884
rect 19387 48844 19432 48872
rect 19426 48832 19432 48844
rect 19484 48832 19490 48884
rect 21085 48875 21143 48881
rect 19628 48844 20576 48872
rect 15470 48804 15476 48816
rect 15431 48776 15476 48804
rect 15470 48764 15476 48776
rect 15528 48764 15534 48816
rect 16485 48807 16543 48813
rect 16485 48773 16497 48807
rect 16531 48804 16543 48807
rect 16574 48804 16580 48816
rect 16531 48776 16580 48804
rect 16531 48773 16543 48776
rect 16485 48767 16543 48773
rect 16574 48764 16580 48776
rect 16632 48764 16638 48816
rect 14185 48739 14243 48745
rect 14185 48705 14197 48739
rect 14231 48736 14243 48739
rect 14231 48708 15608 48736
rect 14231 48705 14243 48708
rect 14185 48699 14243 48705
rect 12621 48671 12679 48677
rect 12621 48637 12633 48671
rect 12667 48668 12679 48671
rect 12894 48668 12900 48680
rect 12667 48640 12900 48668
rect 12667 48637 12679 48640
rect 12621 48631 12679 48637
rect 12894 48628 12900 48640
rect 12952 48628 12958 48680
rect 13630 48668 13636 48680
rect 13591 48640 13636 48668
rect 13630 48628 13636 48640
rect 13688 48628 13694 48680
rect 14553 48671 14611 48677
rect 14553 48637 14565 48671
rect 14599 48668 14611 48671
rect 14642 48668 14648 48680
rect 14599 48640 14648 48668
rect 14599 48637 14611 48640
rect 14553 48631 14611 48637
rect 14642 48628 14648 48640
rect 14700 48628 14706 48680
rect 14734 48628 14740 48680
rect 14792 48668 14798 48680
rect 15580 48677 15608 48708
rect 16298 48696 16304 48748
rect 16356 48736 16362 48748
rect 16761 48739 16819 48745
rect 16761 48736 16773 48739
rect 16356 48708 16773 48736
rect 16356 48696 16362 48708
rect 16761 48705 16773 48708
rect 16807 48736 16819 48739
rect 17126 48736 17132 48748
rect 16807 48708 17132 48736
rect 16807 48705 16819 48708
rect 16761 48699 16819 48705
rect 17126 48696 17132 48708
rect 17184 48696 17190 48748
rect 19628 48736 19656 48844
rect 20548 48804 20576 48844
rect 21085 48841 21097 48875
rect 21131 48872 21143 48875
rect 21266 48872 21272 48884
rect 21131 48844 21272 48872
rect 21131 48841 21143 48844
rect 21085 48835 21143 48841
rect 21266 48832 21272 48844
rect 21324 48832 21330 48884
rect 22370 48832 22376 48884
rect 22428 48872 22434 48884
rect 22925 48875 22983 48881
rect 22925 48872 22937 48875
rect 22428 48844 22937 48872
rect 22428 48832 22434 48844
rect 22925 48841 22937 48844
rect 22971 48841 22983 48875
rect 24762 48872 24768 48884
rect 24723 48844 24768 48872
rect 22925 48835 22983 48841
rect 24762 48832 24768 48844
rect 24820 48832 24826 48884
rect 25406 48872 25412 48884
rect 25367 48844 25412 48872
rect 25406 48832 25412 48844
rect 25464 48832 25470 48884
rect 21453 48807 21511 48813
rect 20548 48776 20760 48804
rect 18064 48708 19656 48736
rect 18064 48680 18092 48708
rect 19978 48696 19984 48748
rect 20036 48736 20042 48748
rect 20732 48745 20760 48776
rect 21453 48773 21465 48807
rect 21499 48804 21511 48807
rect 21499 48776 22140 48804
rect 21499 48773 21511 48776
rect 21453 48767 21511 48773
rect 20717 48739 20775 48745
rect 20036 48708 20081 48736
rect 20036 48696 20042 48708
rect 20717 48705 20729 48739
rect 20763 48705 20775 48739
rect 22112 48736 22140 48776
rect 22649 48739 22707 48745
rect 22112 48708 22508 48736
rect 20717 48699 20775 48705
rect 22480 48680 22508 48708
rect 22649 48705 22661 48739
rect 22695 48736 22707 48739
rect 22922 48736 22928 48748
rect 22695 48708 22928 48736
rect 22695 48705 22707 48708
rect 22649 48699 22707 48705
rect 22922 48696 22928 48708
rect 22980 48696 22986 48748
rect 23658 48736 23664 48748
rect 23619 48708 23664 48736
rect 23658 48696 23664 48708
rect 23716 48696 23722 48748
rect 15013 48671 15071 48677
rect 15013 48668 15025 48671
rect 14792 48640 15025 48668
rect 14792 48628 14798 48640
rect 15013 48637 15025 48640
rect 15059 48637 15071 48671
rect 15013 48631 15071 48637
rect 15565 48671 15623 48677
rect 15565 48637 15577 48671
rect 15611 48668 15623 48671
rect 16482 48668 16488 48680
rect 15611 48640 16488 48668
rect 15611 48637 15623 48640
rect 15565 48631 15623 48637
rect 16482 48628 16488 48640
rect 16540 48628 16546 48680
rect 16942 48668 16948 48680
rect 16855 48640 16948 48668
rect 16942 48628 16948 48640
rect 17000 48668 17006 48680
rect 18046 48668 18052 48680
rect 17000 48640 17540 48668
rect 18007 48640 18052 48668
rect 17000 48628 17006 48640
rect 14660 48600 14688 48628
rect 15102 48600 15108 48612
rect 14660 48572 15108 48600
rect 15102 48560 15108 48572
rect 15160 48560 15166 48612
rect 11330 48492 11336 48544
rect 11388 48532 11394 48544
rect 11425 48535 11483 48541
rect 11425 48532 11437 48535
rect 11388 48504 11437 48532
rect 11388 48492 11394 48504
rect 11425 48501 11437 48504
rect 11471 48532 11483 48535
rect 12802 48532 12808 48544
rect 11471 48504 12808 48532
rect 11471 48501 11483 48504
rect 11425 48495 11483 48501
rect 12802 48492 12808 48504
rect 12860 48492 12866 48544
rect 13814 48532 13820 48544
rect 13775 48504 13820 48532
rect 13814 48492 13820 48504
rect 13872 48492 13878 48544
rect 17129 48535 17187 48541
rect 17129 48501 17141 48535
rect 17175 48532 17187 48535
rect 17310 48532 17316 48544
rect 17175 48504 17316 48532
rect 17175 48501 17187 48504
rect 17129 48495 17187 48501
rect 17310 48492 17316 48504
rect 17368 48492 17374 48544
rect 17512 48541 17540 48640
rect 18046 48628 18052 48640
rect 18104 48628 18110 48680
rect 18230 48628 18236 48680
rect 18288 48668 18294 48680
rect 18598 48668 18604 48680
rect 18288 48640 18604 48668
rect 18288 48628 18294 48640
rect 18598 48628 18604 48640
rect 18656 48668 18662 48680
rect 18877 48671 18935 48677
rect 18877 48668 18889 48671
rect 18656 48640 18889 48668
rect 18656 48628 18662 48640
rect 18877 48637 18889 48640
rect 18923 48637 18935 48671
rect 19058 48668 19064 48680
rect 19019 48640 19064 48668
rect 18877 48631 18935 48637
rect 19058 48628 19064 48640
rect 19116 48628 19122 48680
rect 19794 48628 19800 48680
rect 19852 48668 19858 48680
rect 20257 48671 20315 48677
rect 20257 48668 20269 48671
rect 19852 48640 20269 48668
rect 19852 48628 19858 48640
rect 20257 48637 20269 48640
rect 20303 48637 20315 48671
rect 20257 48631 20315 48637
rect 21450 48628 21456 48680
rect 21508 48668 21514 48680
rect 22002 48668 22008 48680
rect 21508 48640 22008 48668
rect 21508 48628 21514 48640
rect 22002 48628 22008 48640
rect 22060 48628 22066 48680
rect 22189 48671 22247 48677
rect 22189 48637 22201 48671
rect 22235 48637 22247 48671
rect 22189 48631 22247 48637
rect 17678 48560 17684 48612
rect 17736 48600 17742 48612
rect 17736 48572 19104 48600
rect 17736 48560 17742 48572
rect 17497 48535 17555 48541
rect 17497 48501 17509 48535
rect 17543 48532 17555 48535
rect 17770 48532 17776 48544
rect 17543 48504 17776 48532
rect 17543 48501 17555 48504
rect 17497 48495 17555 48501
rect 17770 48492 17776 48504
rect 17828 48492 17834 48544
rect 18322 48532 18328 48544
rect 18283 48504 18328 48532
rect 18322 48492 18328 48504
rect 18380 48492 18386 48544
rect 19076 48532 19104 48572
rect 19150 48560 19156 48612
rect 19208 48600 19214 48612
rect 20165 48603 20223 48609
rect 20165 48600 20177 48603
rect 19208 48572 20177 48600
rect 19208 48560 19214 48572
rect 20165 48569 20177 48572
rect 20211 48569 20223 48603
rect 20165 48563 20223 48569
rect 20349 48603 20407 48609
rect 20349 48569 20361 48603
rect 20395 48569 20407 48603
rect 21821 48603 21879 48609
rect 21821 48600 21833 48603
rect 20349 48563 20407 48569
rect 21468 48572 21833 48600
rect 19797 48535 19855 48541
rect 19797 48532 19809 48535
rect 19076 48504 19809 48532
rect 19797 48501 19809 48504
rect 19843 48532 19855 48535
rect 20364 48532 20392 48563
rect 21468 48544 21496 48572
rect 21821 48569 21833 48572
rect 21867 48600 21879 48603
rect 22204 48600 22232 48631
rect 22462 48628 22468 48680
rect 22520 48668 22526 48680
rect 23477 48671 23535 48677
rect 22520 48640 22613 48668
rect 22520 48628 22526 48640
rect 23477 48637 23489 48671
rect 23523 48668 23535 48671
rect 23753 48671 23811 48677
rect 23753 48668 23765 48671
rect 23523 48640 23765 48668
rect 23523 48637 23535 48640
rect 23477 48631 23535 48637
rect 23753 48637 23765 48640
rect 23799 48637 23811 48671
rect 25222 48668 25228 48680
rect 25183 48640 25228 48668
rect 23753 48631 23811 48637
rect 23492 48600 23520 48631
rect 25222 48628 25228 48640
rect 25280 48668 25286 48680
rect 25685 48671 25743 48677
rect 25685 48668 25697 48671
rect 25280 48640 25697 48668
rect 25280 48628 25286 48640
rect 25685 48637 25697 48640
rect 25731 48637 25743 48671
rect 25685 48631 25743 48637
rect 21867 48572 23520 48600
rect 21867 48569 21879 48572
rect 21821 48563 21879 48569
rect 19843 48504 20392 48532
rect 19843 48501 19855 48504
rect 19797 48495 19855 48501
rect 21450 48492 21456 48544
rect 21508 48492 21514 48544
rect 1104 48442 28888 48464
rect 1104 48390 10982 48442
rect 11034 48390 11046 48442
rect 11098 48390 11110 48442
rect 11162 48390 11174 48442
rect 11226 48390 20982 48442
rect 21034 48390 21046 48442
rect 21098 48390 21110 48442
rect 21162 48390 21174 48442
rect 21226 48390 28888 48442
rect 1104 48368 28888 48390
rect 11422 48288 11428 48340
rect 11480 48328 11486 48340
rect 12437 48331 12495 48337
rect 12437 48328 12449 48331
rect 11480 48300 12449 48328
rect 11480 48288 11486 48300
rect 12437 48297 12449 48300
rect 12483 48297 12495 48331
rect 12437 48291 12495 48297
rect 13265 48331 13323 48337
rect 13265 48297 13277 48331
rect 13311 48328 13323 48331
rect 13630 48328 13636 48340
rect 13311 48300 13636 48328
rect 13311 48297 13323 48300
rect 13265 48291 13323 48297
rect 13630 48288 13636 48300
rect 13688 48288 13694 48340
rect 14734 48328 14740 48340
rect 14695 48300 14740 48328
rect 14734 48288 14740 48300
rect 14792 48288 14798 48340
rect 15654 48328 15660 48340
rect 14844 48300 15660 48328
rect 12897 48263 12955 48269
rect 12897 48229 12909 48263
rect 12943 48260 12955 48263
rect 13170 48260 13176 48272
rect 12943 48232 13176 48260
rect 12943 48229 12955 48232
rect 12897 48223 12955 48229
rect 13170 48220 13176 48232
rect 13228 48220 13234 48272
rect 13354 48260 13360 48272
rect 13315 48232 13360 48260
rect 13354 48220 13360 48232
rect 13412 48220 13418 48272
rect 14844 48260 14872 48300
rect 15654 48288 15660 48300
rect 15712 48288 15718 48340
rect 17497 48331 17555 48337
rect 17497 48328 17509 48331
rect 16500 48300 17509 48328
rect 15746 48260 15752 48272
rect 14200 48232 14872 48260
rect 15120 48232 15752 48260
rect 14200 48204 14228 48232
rect 14182 48192 14188 48204
rect 14095 48164 14188 48192
rect 14182 48152 14188 48164
rect 14240 48152 14246 48204
rect 14292 48164 14596 48192
rect 13722 48084 13728 48136
rect 13780 48124 13786 48136
rect 13909 48127 13967 48133
rect 13909 48124 13921 48127
rect 13780 48096 13921 48124
rect 13780 48084 13786 48096
rect 13909 48093 13921 48096
rect 13955 48124 13967 48127
rect 14292 48124 14320 48164
rect 13955 48096 14320 48124
rect 14369 48127 14427 48133
rect 13955 48093 13967 48096
rect 13909 48087 13967 48093
rect 14369 48093 14381 48127
rect 14415 48093 14427 48127
rect 14568 48124 14596 48164
rect 14826 48152 14832 48204
rect 14884 48192 14890 48204
rect 15120 48192 15148 48232
rect 15746 48220 15752 48232
rect 15804 48220 15810 48272
rect 16500 48260 16528 48300
rect 17497 48297 17509 48300
rect 17543 48297 17555 48331
rect 19058 48328 19064 48340
rect 17497 48291 17555 48297
rect 17880 48300 19064 48328
rect 16132 48232 16528 48260
rect 16945 48263 17003 48269
rect 16132 48201 16160 48232
rect 16945 48229 16957 48263
rect 16991 48260 17003 48263
rect 17218 48260 17224 48272
rect 16991 48232 17224 48260
rect 16991 48229 17003 48232
rect 16945 48223 17003 48229
rect 17218 48220 17224 48232
rect 17276 48220 17282 48272
rect 16117 48195 16175 48201
rect 16117 48192 16129 48195
rect 14884 48164 15148 48192
rect 15304 48164 16129 48192
rect 14884 48152 14890 48164
rect 15304 48124 15332 48164
rect 16117 48161 16129 48164
rect 16163 48161 16175 48195
rect 16117 48155 16175 48161
rect 16393 48195 16451 48201
rect 16393 48161 16405 48195
rect 16439 48161 16451 48195
rect 17678 48192 17684 48204
rect 17591 48164 17684 48192
rect 16393 48155 16451 48161
rect 14568 48096 15332 48124
rect 15565 48127 15623 48133
rect 14369 48087 14427 48093
rect 15565 48093 15577 48127
rect 15611 48124 15623 48127
rect 15746 48124 15752 48136
rect 15611 48096 15752 48124
rect 15611 48093 15623 48096
rect 15565 48087 15623 48093
rect 13446 48016 13452 48068
rect 13504 48056 13510 48068
rect 14384 48056 14412 48087
rect 15746 48084 15752 48096
rect 15804 48084 15810 48136
rect 14642 48056 14648 48068
rect 13504 48028 14648 48056
rect 13504 48016 13510 48028
rect 14642 48016 14648 48028
rect 14700 48016 14706 48068
rect 15010 48056 15016 48068
rect 14971 48028 15016 48056
rect 15010 48016 15016 48028
rect 15068 48016 15074 48068
rect 15102 48016 15108 48068
rect 15160 48056 15166 48068
rect 15286 48056 15292 48068
rect 15160 48028 15292 48056
rect 15160 48016 15166 48028
rect 15286 48016 15292 48028
rect 15344 48016 15350 48068
rect 15470 48016 15476 48068
rect 15528 48056 15534 48068
rect 16408 48056 16436 48155
rect 17678 48152 17684 48164
rect 17736 48192 17742 48204
rect 17880 48192 17908 48300
rect 19058 48288 19064 48300
rect 19116 48288 19122 48340
rect 19794 48288 19800 48340
rect 19852 48328 19858 48340
rect 20257 48331 20315 48337
rect 20257 48328 20269 48331
rect 19852 48300 20269 48328
rect 19852 48288 19858 48300
rect 20257 48297 20269 48300
rect 20303 48297 20315 48331
rect 21177 48331 21235 48337
rect 21177 48328 21189 48331
rect 20257 48291 20315 48297
rect 20916 48300 21189 48328
rect 18874 48260 18880 48272
rect 18835 48232 18880 48260
rect 18874 48220 18880 48232
rect 18932 48220 18938 48272
rect 18966 48220 18972 48272
rect 19024 48260 19030 48272
rect 20165 48263 20223 48269
rect 20165 48260 20177 48263
rect 19024 48232 20177 48260
rect 19024 48220 19030 48232
rect 20165 48229 20177 48232
rect 20211 48229 20223 48263
rect 20272 48260 20300 48291
rect 20916 48260 20944 48300
rect 21177 48297 21189 48300
rect 21223 48297 21235 48331
rect 22554 48328 22560 48340
rect 21177 48291 21235 48297
rect 22112 48300 22560 48328
rect 21542 48260 21548 48272
rect 20272 48232 20944 48260
rect 21376 48232 21548 48260
rect 20165 48223 20223 48229
rect 18046 48192 18052 48204
rect 17736 48164 17908 48192
rect 18007 48164 18052 48192
rect 17736 48152 17742 48164
rect 18046 48152 18052 48164
rect 18104 48152 18110 48204
rect 18230 48192 18236 48204
rect 18191 48164 18236 48192
rect 18230 48152 18236 48164
rect 18288 48152 18294 48204
rect 19521 48195 19579 48201
rect 19521 48161 19533 48195
rect 19567 48192 19579 48195
rect 19886 48192 19892 48204
rect 19567 48164 19892 48192
rect 19567 48161 19579 48164
rect 19521 48155 19579 48161
rect 19886 48152 19892 48164
rect 19944 48152 19950 48204
rect 20070 48152 20076 48204
rect 20128 48192 20134 48204
rect 20901 48195 20959 48201
rect 20901 48192 20913 48195
rect 20128 48164 20913 48192
rect 20128 48152 20134 48164
rect 20901 48161 20913 48164
rect 20947 48161 20959 48195
rect 20901 48155 20959 48161
rect 21085 48195 21143 48201
rect 21085 48161 21097 48195
rect 21131 48161 21143 48195
rect 21253 48195 21311 48201
rect 21253 48192 21265 48195
rect 21085 48155 21143 48161
rect 21192 48164 21265 48192
rect 16577 48127 16635 48133
rect 16577 48124 16589 48127
rect 15528 48028 16436 48056
rect 16500 48096 16589 48124
rect 15528 48016 15534 48028
rect 14660 47988 14688 48016
rect 16500 47988 16528 48096
rect 16577 48093 16589 48096
rect 16623 48093 16635 48127
rect 16577 48087 16635 48093
rect 16666 48084 16672 48136
rect 16724 48124 16730 48136
rect 17221 48127 17279 48133
rect 17221 48124 17233 48127
rect 16724 48096 17233 48124
rect 16724 48084 16730 48096
rect 17221 48093 17233 48096
rect 17267 48124 17279 48127
rect 19150 48124 19156 48136
rect 17267 48096 19156 48124
rect 17267 48093 17279 48096
rect 17221 48087 17279 48093
rect 19150 48084 19156 48096
rect 19208 48084 19214 48136
rect 19429 48127 19487 48133
rect 19429 48093 19441 48127
rect 19475 48124 19487 48127
rect 19794 48124 19800 48136
rect 19475 48096 19800 48124
rect 19475 48093 19487 48096
rect 19429 48087 19487 48093
rect 19794 48084 19800 48096
rect 19852 48084 19858 48136
rect 19978 48124 19984 48136
rect 19939 48096 19984 48124
rect 19978 48084 19984 48096
rect 20036 48084 20042 48136
rect 21100 48124 21128 48155
rect 20732 48096 21128 48124
rect 18874 48016 18880 48068
rect 18932 48056 18938 48068
rect 20732 48065 20760 48096
rect 20717 48059 20775 48065
rect 20717 48056 20729 48059
rect 18932 48028 20729 48056
rect 18932 48016 18938 48028
rect 20717 48025 20729 48028
rect 20763 48025 20775 48059
rect 20717 48019 20775 48025
rect 16850 47988 16856 48000
rect 14660 47960 16856 47988
rect 16850 47948 16856 47960
rect 16908 47948 16914 48000
rect 19150 47988 19156 48000
rect 19111 47960 19156 47988
rect 19150 47948 19156 47960
rect 19208 47948 19214 48000
rect 20165 47991 20223 47997
rect 20165 47957 20177 47991
rect 20211 47988 20223 47991
rect 21192 47988 21220 48164
rect 21253 48161 21265 48164
rect 21299 48192 21311 48195
rect 21376 48192 21404 48232
rect 21542 48220 21548 48232
rect 21600 48220 21606 48272
rect 22112 48192 22140 48300
rect 22554 48288 22560 48300
rect 22612 48328 22618 48340
rect 22612 48300 23428 48328
rect 22612 48288 22618 48300
rect 22373 48263 22431 48269
rect 22373 48229 22385 48263
rect 22419 48260 22431 48263
rect 22922 48260 22928 48272
rect 22419 48232 22928 48260
rect 22419 48229 22431 48232
rect 22373 48223 22431 48229
rect 22646 48192 22652 48204
rect 21299 48164 21404 48192
rect 21928 48164 22140 48192
rect 22607 48164 22652 48192
rect 21299 48161 21311 48164
rect 21253 48155 21311 48161
rect 21542 48084 21548 48136
rect 21600 48124 21606 48136
rect 21637 48127 21695 48133
rect 21637 48124 21649 48127
rect 21600 48096 21649 48124
rect 21600 48084 21606 48096
rect 21637 48093 21649 48096
rect 21683 48093 21695 48127
rect 21637 48087 21695 48093
rect 20211 47960 21220 47988
rect 20211 47957 20223 47960
rect 20165 47951 20223 47957
rect 21542 47948 21548 48000
rect 21600 47988 21606 48000
rect 21928 47997 21956 48164
rect 22646 48152 22652 48164
rect 22704 48152 22710 48204
rect 22848 48201 22876 48232
rect 22922 48220 22928 48232
rect 22980 48220 22986 48272
rect 23400 48260 23428 48300
rect 25130 48260 25136 48272
rect 23400 48232 24716 48260
rect 25091 48232 25136 48260
rect 24688 48204 24716 48232
rect 25130 48220 25136 48232
rect 25188 48220 25194 48272
rect 22833 48195 22891 48201
rect 22833 48161 22845 48195
rect 22879 48161 22891 48195
rect 22833 48155 22891 48161
rect 23566 48152 23572 48204
rect 23624 48192 23630 48204
rect 23661 48195 23719 48201
rect 23661 48192 23673 48195
rect 23624 48164 23673 48192
rect 23624 48152 23630 48164
rect 23661 48161 23673 48164
rect 23707 48192 23719 48195
rect 24121 48195 24179 48201
rect 24121 48192 24133 48195
rect 23707 48164 24133 48192
rect 23707 48161 23719 48164
rect 23661 48155 23719 48161
rect 24121 48161 24133 48164
rect 24167 48192 24179 48195
rect 24489 48195 24547 48201
rect 24489 48192 24501 48195
rect 24167 48164 24501 48192
rect 24167 48161 24179 48164
rect 24121 48155 24179 48161
rect 24489 48161 24501 48164
rect 24535 48161 24547 48195
rect 24670 48192 24676 48204
rect 24583 48164 24676 48192
rect 24489 48155 24547 48161
rect 24670 48152 24676 48164
rect 24728 48152 24734 48204
rect 22925 48127 22983 48133
rect 22925 48093 22937 48127
rect 22971 48093 22983 48127
rect 23750 48124 23756 48136
rect 23711 48096 23756 48124
rect 22925 48087 22983 48093
rect 22830 48016 22836 48068
rect 22888 48056 22894 48068
rect 22940 48056 22968 48087
rect 23750 48084 23756 48096
rect 23808 48084 23814 48136
rect 22888 48028 22968 48056
rect 22888 48016 22894 48028
rect 21913 47991 21971 47997
rect 21913 47988 21925 47991
rect 21600 47960 21925 47988
rect 21600 47948 21606 47960
rect 21913 47957 21925 47960
rect 21959 47957 21971 47991
rect 21913 47951 21971 47957
rect 22465 47991 22523 47997
rect 22465 47957 22477 47991
rect 22511 47988 22523 47991
rect 23474 47988 23480 48000
rect 22511 47960 23480 47988
rect 22511 47957 22523 47960
rect 22465 47951 22523 47957
rect 23474 47948 23480 47960
rect 23532 47948 23538 48000
rect 24854 47988 24860 48000
rect 24815 47960 24860 47988
rect 24854 47948 24860 47960
rect 24912 47948 24918 48000
rect 26237 47991 26295 47997
rect 26237 47957 26249 47991
rect 26283 47988 26295 47991
rect 26326 47988 26332 48000
rect 26283 47960 26332 47988
rect 26283 47957 26295 47960
rect 26237 47951 26295 47957
rect 26326 47948 26332 47960
rect 26384 47948 26390 48000
rect 1104 47898 28888 47920
rect 1104 47846 5982 47898
rect 6034 47846 6046 47898
rect 6098 47846 6110 47898
rect 6162 47846 6174 47898
rect 6226 47846 15982 47898
rect 16034 47846 16046 47898
rect 16098 47846 16110 47898
rect 16162 47846 16174 47898
rect 16226 47846 25982 47898
rect 26034 47846 26046 47898
rect 26098 47846 26110 47898
rect 26162 47846 26174 47898
rect 26226 47846 28888 47898
rect 1104 47824 28888 47846
rect 7834 47744 7840 47796
rect 7892 47784 7898 47796
rect 8021 47787 8079 47793
rect 8021 47784 8033 47787
rect 7892 47756 8033 47784
rect 7892 47744 7898 47756
rect 8021 47753 8033 47756
rect 8067 47753 8079 47787
rect 13078 47784 13084 47796
rect 13039 47756 13084 47784
rect 8021 47747 8079 47753
rect 8036 47648 8064 47747
rect 13078 47744 13084 47756
rect 13136 47744 13142 47796
rect 13446 47784 13452 47796
rect 13407 47756 13452 47784
rect 13446 47744 13452 47756
rect 13504 47744 13510 47796
rect 13814 47744 13820 47796
rect 13872 47784 13878 47796
rect 14277 47787 14335 47793
rect 14277 47784 14289 47787
rect 13872 47756 14289 47784
rect 13872 47744 13878 47756
rect 14277 47753 14289 47756
rect 14323 47784 14335 47787
rect 14458 47784 14464 47796
rect 14323 47756 14464 47784
rect 14323 47753 14335 47756
rect 14277 47747 14335 47753
rect 14458 47744 14464 47756
rect 14516 47744 14522 47796
rect 14642 47784 14648 47796
rect 14603 47756 14648 47784
rect 14642 47744 14648 47756
rect 14700 47744 14706 47796
rect 15194 47744 15200 47796
rect 15252 47784 15258 47796
rect 15289 47787 15347 47793
rect 15289 47784 15301 47787
rect 15252 47756 15301 47784
rect 15252 47744 15258 47756
rect 15289 47753 15301 47756
rect 15335 47784 15347 47787
rect 16850 47784 16856 47796
rect 15335 47756 15608 47784
rect 16811 47756 16856 47784
rect 15335 47753 15347 47756
rect 15289 47747 15347 47753
rect 12713 47719 12771 47725
rect 12713 47685 12725 47719
rect 12759 47716 12771 47719
rect 13722 47716 13728 47728
rect 12759 47688 13728 47716
rect 12759 47685 12771 47688
rect 12713 47679 12771 47685
rect 13722 47676 13728 47688
rect 13780 47676 13786 47728
rect 8481 47651 8539 47657
rect 8481 47648 8493 47651
rect 8036 47620 8493 47648
rect 8481 47617 8493 47620
rect 8527 47617 8539 47651
rect 8481 47611 8539 47617
rect 13817 47651 13875 47657
rect 13817 47617 13829 47651
rect 13863 47648 13875 47651
rect 14182 47648 14188 47660
rect 13863 47620 14188 47648
rect 13863 47617 13875 47620
rect 13817 47611 13875 47617
rect 14182 47608 14188 47620
rect 14240 47608 14246 47660
rect 15580 47657 15608 47756
rect 16850 47744 16856 47756
rect 16908 47744 16914 47796
rect 17034 47744 17040 47796
rect 17092 47784 17098 47796
rect 17405 47787 17463 47793
rect 17405 47784 17417 47787
rect 17092 47756 17417 47784
rect 17092 47744 17098 47756
rect 17405 47753 17417 47756
rect 17451 47753 17463 47787
rect 19794 47784 19800 47796
rect 19755 47756 19800 47784
rect 17405 47747 17463 47753
rect 19794 47744 19800 47756
rect 19852 47744 19858 47796
rect 19886 47744 19892 47796
rect 19944 47784 19950 47796
rect 20165 47787 20223 47793
rect 20165 47784 20177 47787
rect 19944 47756 20177 47784
rect 19944 47744 19950 47756
rect 20165 47753 20177 47756
rect 20211 47753 20223 47787
rect 23106 47784 23112 47796
rect 23067 47756 23112 47784
rect 20165 47747 20223 47753
rect 23106 47744 23112 47756
rect 23164 47784 23170 47796
rect 24486 47784 24492 47796
rect 23164 47756 24492 47784
rect 23164 47744 23170 47756
rect 24486 47744 24492 47756
rect 24544 47744 24550 47796
rect 24670 47744 24676 47796
rect 24728 47784 24734 47796
rect 24949 47787 25007 47793
rect 24949 47784 24961 47787
rect 24728 47756 24961 47784
rect 24728 47744 24734 47756
rect 24949 47753 24961 47756
rect 24995 47753 25007 47787
rect 27706 47784 27712 47796
rect 27667 47756 27712 47784
rect 24949 47747 25007 47753
rect 27706 47744 27712 47756
rect 27764 47744 27770 47796
rect 17310 47676 17316 47728
rect 17368 47716 17374 47728
rect 17586 47716 17592 47728
rect 17368 47688 17592 47716
rect 17368 47676 17374 47688
rect 17586 47676 17592 47688
rect 17644 47676 17650 47728
rect 19904 47716 19932 47744
rect 19076 47688 19932 47716
rect 15565 47651 15623 47657
rect 15565 47617 15577 47651
rect 15611 47617 15623 47651
rect 16482 47648 16488 47660
rect 16443 47620 16488 47648
rect 15565 47611 15623 47617
rect 16482 47608 16488 47620
rect 16540 47608 16546 47660
rect 18046 47608 18052 47660
rect 18104 47648 18110 47660
rect 18325 47651 18383 47657
rect 18325 47648 18337 47651
rect 18104 47620 18337 47648
rect 18104 47608 18110 47620
rect 18325 47617 18337 47620
rect 18371 47648 18383 47651
rect 19076 47648 19104 47688
rect 19978 47676 19984 47728
rect 20036 47716 20042 47728
rect 20346 47716 20352 47728
rect 20036 47688 20352 47716
rect 20036 47676 20042 47688
rect 20346 47676 20352 47688
rect 20404 47676 20410 47728
rect 22646 47676 22652 47728
rect 22704 47716 22710 47728
rect 23566 47716 23572 47728
rect 22704 47688 23572 47716
rect 22704 47676 22710 47688
rect 23566 47676 23572 47688
rect 23624 47716 23630 47728
rect 23750 47716 23756 47728
rect 23624 47688 23756 47716
rect 23624 47676 23630 47688
rect 23750 47676 23756 47688
rect 23808 47676 23814 47728
rect 18371 47620 19104 47648
rect 18371 47617 18383 47620
rect 18325 47611 18383 47617
rect 8202 47580 8208 47592
rect 8163 47552 8208 47580
rect 8202 47540 8208 47552
rect 8260 47540 8266 47592
rect 14461 47583 14519 47589
rect 14461 47549 14473 47583
rect 14507 47580 14519 47583
rect 14507 47552 15056 47580
rect 14507 47549 14519 47552
rect 14461 47543 14519 47549
rect 15028 47456 15056 47552
rect 15654 47540 15660 47592
rect 15712 47580 15718 47592
rect 16025 47583 16083 47589
rect 16025 47580 16037 47583
rect 15712 47552 16037 47580
rect 15712 47540 15718 47552
rect 16025 47549 16037 47552
rect 16071 47549 16083 47583
rect 16298 47580 16304 47592
rect 16259 47552 16304 47580
rect 16025 47543 16083 47549
rect 16040 47512 16068 47543
rect 16298 47540 16304 47552
rect 16356 47540 16362 47592
rect 17586 47580 17592 47592
rect 17547 47552 17592 47580
rect 17586 47540 17592 47552
rect 17644 47540 17650 47592
rect 18601 47583 18659 47589
rect 18601 47549 18613 47583
rect 18647 47580 18659 47583
rect 18782 47580 18788 47592
rect 18647 47552 18788 47580
rect 18647 47549 18659 47552
rect 18601 47543 18659 47549
rect 18782 47540 18788 47552
rect 18840 47540 18846 47592
rect 18966 47580 18972 47592
rect 18879 47552 18972 47580
rect 18966 47540 18972 47552
rect 19024 47580 19030 47592
rect 19076 47580 19104 47620
rect 19521 47651 19579 47657
rect 19521 47617 19533 47651
rect 19567 47648 19579 47651
rect 19610 47648 19616 47660
rect 19567 47620 19616 47648
rect 19567 47617 19579 47620
rect 19521 47611 19579 47617
rect 19610 47608 19616 47620
rect 19668 47608 19674 47660
rect 22833 47651 22891 47657
rect 22833 47617 22845 47651
rect 22879 47648 22891 47651
rect 24394 47648 24400 47660
rect 22879 47620 24400 47648
rect 22879 47617 22891 47620
rect 22833 47611 22891 47617
rect 24394 47608 24400 47620
rect 24452 47648 24458 47660
rect 24673 47651 24731 47657
rect 24673 47648 24685 47651
rect 24452 47620 24685 47648
rect 24452 47608 24458 47620
rect 24673 47617 24685 47620
rect 24719 47617 24731 47651
rect 25774 47648 25780 47660
rect 24673 47611 24731 47617
rect 25332 47620 25780 47648
rect 19024 47552 19104 47580
rect 19024 47540 19030 47552
rect 19150 47540 19156 47592
rect 19208 47580 19214 47592
rect 19245 47583 19303 47589
rect 19245 47580 19257 47583
rect 19208 47552 19257 47580
rect 19208 47540 19214 47552
rect 19245 47549 19257 47552
rect 19291 47549 19303 47583
rect 19245 47543 19303 47549
rect 20441 47583 20499 47589
rect 20441 47549 20453 47583
rect 20487 47580 20499 47583
rect 20714 47580 20720 47592
rect 20487 47552 20720 47580
rect 20487 47549 20499 47552
rect 20441 47543 20499 47549
rect 20714 47540 20720 47552
rect 20772 47580 20778 47592
rect 20901 47583 20959 47589
rect 20901 47580 20913 47583
rect 20772 47552 20913 47580
rect 20772 47540 20778 47552
rect 20901 47549 20913 47552
rect 20947 47549 20959 47583
rect 20901 47543 20959 47549
rect 21266 47540 21272 47592
rect 21324 47580 21330 47592
rect 21361 47583 21419 47589
rect 21361 47580 21373 47583
rect 21324 47552 21373 47580
rect 21324 47540 21330 47552
rect 21361 47549 21373 47552
rect 21407 47580 21419 47583
rect 21450 47580 21456 47592
rect 21407 47552 21456 47580
rect 21407 47549 21419 47552
rect 21361 47543 21419 47549
rect 21450 47540 21456 47552
rect 21508 47540 21514 47592
rect 21634 47540 21640 47592
rect 21692 47580 21698 47592
rect 21913 47583 21971 47589
rect 21913 47580 21925 47583
rect 21692 47552 21925 47580
rect 21692 47540 21698 47552
rect 21913 47549 21925 47552
rect 21959 47549 21971 47583
rect 23474 47580 23480 47592
rect 23435 47552 23480 47580
rect 21913 47543 21971 47549
rect 23474 47540 23480 47552
rect 23532 47540 23538 47592
rect 23750 47540 23756 47592
rect 23808 47580 23814 47592
rect 24213 47583 24271 47589
rect 24213 47580 24225 47583
rect 23808 47552 24225 47580
rect 23808 47540 23814 47552
rect 24213 47549 24225 47552
rect 24259 47549 24271 47583
rect 24486 47580 24492 47592
rect 24447 47552 24492 47580
rect 24213 47543 24271 47549
rect 24486 47540 24492 47552
rect 24544 47540 24550 47592
rect 16206 47512 16212 47524
rect 16040 47484 16212 47512
rect 16206 47472 16212 47484
rect 16264 47512 16270 47524
rect 17221 47515 17279 47521
rect 17221 47512 17233 47515
rect 16264 47484 17233 47512
rect 16264 47472 16270 47484
rect 17221 47481 17233 47484
rect 17267 47481 17279 47515
rect 17221 47475 17279 47481
rect 22554 47472 22560 47524
rect 22612 47512 22618 47524
rect 23198 47512 23204 47524
rect 22612 47484 23204 47512
rect 22612 47472 22618 47484
rect 23198 47472 23204 47484
rect 23256 47472 23262 47524
rect 23661 47515 23719 47521
rect 23661 47481 23673 47515
rect 23707 47512 23719 47515
rect 24118 47512 24124 47524
rect 23707 47484 24124 47512
rect 23707 47481 23719 47484
rect 23661 47475 23719 47481
rect 24118 47472 24124 47484
rect 24176 47472 24182 47524
rect 9766 47444 9772 47456
rect 9727 47416 9772 47444
rect 9766 47404 9772 47416
rect 9824 47404 9830 47456
rect 11974 47404 11980 47456
rect 12032 47444 12038 47456
rect 12161 47447 12219 47453
rect 12161 47444 12173 47447
rect 12032 47416 12173 47444
rect 12032 47404 12038 47416
rect 12161 47413 12173 47416
rect 12207 47413 12219 47447
rect 15010 47444 15016 47456
rect 14971 47416 15016 47444
rect 12161 47407 12219 47413
rect 15010 47404 15016 47416
rect 15068 47404 15074 47456
rect 20438 47404 20444 47456
rect 20496 47444 20502 47456
rect 20625 47447 20683 47453
rect 20625 47444 20637 47447
rect 20496 47416 20637 47444
rect 20496 47404 20502 47416
rect 20625 47413 20637 47416
rect 20671 47413 20683 47447
rect 21542 47444 21548 47456
rect 21503 47416 21548 47444
rect 20625 47407 20683 47413
rect 21542 47404 21548 47416
rect 21600 47404 21606 47456
rect 23293 47447 23351 47453
rect 23293 47413 23305 47447
rect 23339 47444 23351 47447
rect 25332 47444 25360 47620
rect 25774 47608 25780 47620
rect 25832 47648 25838 47660
rect 26145 47651 26203 47657
rect 26145 47648 26157 47651
rect 25832 47620 26157 47648
rect 25832 47608 25838 47620
rect 26145 47617 26157 47620
rect 26191 47648 26203 47651
rect 26326 47648 26332 47660
rect 26191 47620 26332 47648
rect 26191 47617 26203 47620
rect 26145 47611 26203 47617
rect 26326 47608 26332 47620
rect 26384 47648 26390 47660
rect 26878 47648 26884 47660
rect 26384 47620 26884 47648
rect 26384 47608 26390 47620
rect 26878 47608 26884 47620
rect 26936 47608 26942 47660
rect 25409 47583 25467 47589
rect 25409 47549 25421 47583
rect 25455 47580 25467 47583
rect 25866 47580 25872 47592
rect 25455 47552 25872 47580
rect 25455 47549 25467 47552
rect 25409 47543 25467 47549
rect 25866 47540 25872 47552
rect 25924 47540 25930 47592
rect 26421 47583 26479 47589
rect 26421 47580 26433 47583
rect 25976 47552 26433 47580
rect 23339 47416 25360 47444
rect 23339 47413 23351 47416
rect 23293 47407 23351 47413
rect 25406 47404 25412 47456
rect 25464 47444 25470 47456
rect 25976 47453 26004 47552
rect 26421 47549 26433 47552
rect 26467 47549 26479 47583
rect 26421 47543 26479 47549
rect 25961 47447 26019 47453
rect 25961 47444 25973 47447
rect 25464 47416 25973 47444
rect 25464 47404 25470 47416
rect 25961 47413 25973 47416
rect 26007 47413 26019 47447
rect 25961 47407 26019 47413
rect 1104 47354 28888 47376
rect 1104 47302 10982 47354
rect 11034 47302 11046 47354
rect 11098 47302 11110 47354
rect 11162 47302 11174 47354
rect 11226 47302 20982 47354
rect 21034 47302 21046 47354
rect 21098 47302 21110 47354
rect 21162 47302 21174 47354
rect 21226 47302 28888 47354
rect 1104 47280 28888 47302
rect 8202 47240 8208 47252
rect 8163 47212 8208 47240
rect 8202 47200 8208 47212
rect 8260 47200 8266 47252
rect 13722 47240 13728 47252
rect 13683 47212 13728 47240
rect 13722 47200 13728 47212
rect 13780 47200 13786 47252
rect 13998 47240 14004 47252
rect 13959 47212 14004 47240
rect 13998 47200 14004 47212
rect 14056 47200 14062 47252
rect 14090 47200 14096 47252
rect 14148 47240 14154 47252
rect 14369 47243 14427 47249
rect 14369 47240 14381 47243
rect 14148 47212 14381 47240
rect 14148 47200 14154 47212
rect 14369 47209 14381 47212
rect 14415 47209 14427 47243
rect 14734 47240 14740 47252
rect 14695 47212 14740 47240
rect 14369 47203 14427 47209
rect 14734 47200 14740 47212
rect 14792 47200 14798 47252
rect 16945 47243 17003 47249
rect 16945 47209 16957 47243
rect 16991 47240 17003 47243
rect 17494 47240 17500 47252
rect 16991 47212 17500 47240
rect 16991 47209 17003 47212
rect 16945 47203 17003 47209
rect 17494 47200 17500 47212
rect 17552 47240 17558 47252
rect 17954 47240 17960 47252
rect 17552 47212 17960 47240
rect 17552 47200 17558 47212
rect 17954 47200 17960 47212
rect 18012 47200 18018 47252
rect 20717 47243 20775 47249
rect 20717 47209 20729 47243
rect 20763 47240 20775 47243
rect 21634 47240 21640 47252
rect 20763 47212 21640 47240
rect 20763 47209 20775 47212
rect 20717 47203 20775 47209
rect 21634 47200 21640 47212
rect 21692 47200 21698 47252
rect 22373 47243 22431 47249
rect 22373 47209 22385 47243
rect 22419 47240 22431 47243
rect 22646 47240 22652 47252
rect 22419 47212 22652 47240
rect 22419 47209 22431 47212
rect 22373 47203 22431 47209
rect 22646 47200 22652 47212
rect 22704 47200 22710 47252
rect 22738 47200 22744 47252
rect 22796 47200 22802 47252
rect 23658 47200 23664 47252
rect 23716 47240 23722 47252
rect 23753 47243 23811 47249
rect 23753 47240 23765 47243
rect 23716 47212 23765 47240
rect 23716 47200 23722 47212
rect 23753 47209 23765 47212
rect 23799 47209 23811 47243
rect 24118 47240 24124 47252
rect 24079 47212 24124 47240
rect 23753 47203 23811 47209
rect 24118 47200 24124 47212
rect 24176 47240 24182 47252
rect 26694 47240 26700 47252
rect 24176 47212 24532 47240
rect 26655 47212 26700 47240
rect 24176 47200 24182 47212
rect 14918 47132 14924 47184
rect 14976 47172 14982 47184
rect 15105 47175 15163 47181
rect 15105 47172 15117 47175
rect 14976 47144 15117 47172
rect 14976 47132 14982 47144
rect 15105 47141 15117 47144
rect 15151 47172 15163 47175
rect 15151 47144 16252 47172
rect 15151 47141 15163 47144
rect 15105 47135 15163 47141
rect 12526 47104 12532 47116
rect 12439 47076 12532 47104
rect 12526 47064 12532 47076
rect 12584 47104 12590 47116
rect 13265 47107 13323 47113
rect 13265 47104 13277 47107
rect 12584 47076 13277 47104
rect 12584 47064 12590 47076
rect 13265 47073 13277 47076
rect 13311 47104 13323 47107
rect 13722 47104 13728 47116
rect 13311 47076 13728 47104
rect 13311 47073 13323 47076
rect 13265 47067 13323 47073
rect 13722 47064 13728 47076
rect 13780 47064 13786 47116
rect 14182 47104 14188 47116
rect 14143 47076 14188 47104
rect 14182 47064 14188 47076
rect 14240 47064 14246 47116
rect 14458 47064 14464 47116
rect 14516 47104 14522 47116
rect 15470 47104 15476 47116
rect 14516 47076 15476 47104
rect 14516 47064 14522 47076
rect 15470 47064 15476 47076
rect 15528 47104 15534 47116
rect 16224 47113 16252 47144
rect 17126 47132 17132 47184
rect 17184 47172 17190 47184
rect 17221 47175 17279 47181
rect 17221 47172 17233 47175
rect 17184 47144 17233 47172
rect 17184 47132 17190 47144
rect 17221 47141 17233 47144
rect 17267 47172 17279 47175
rect 17267 47144 17724 47172
rect 17267 47141 17279 47144
rect 17221 47135 17279 47141
rect 15657 47107 15715 47113
rect 15657 47104 15669 47107
rect 15528 47076 15669 47104
rect 15528 47064 15534 47076
rect 15657 47073 15669 47076
rect 15703 47073 15715 47107
rect 15657 47067 15715 47073
rect 16209 47107 16267 47113
rect 16209 47073 16221 47107
rect 16255 47104 16267 47107
rect 16298 47104 16304 47116
rect 16255 47076 16304 47104
rect 16255 47073 16267 47076
rect 16209 47067 16267 47073
rect 16298 47064 16304 47076
rect 16356 47064 16362 47116
rect 17310 47064 17316 47116
rect 17368 47104 17374 47116
rect 17405 47107 17463 47113
rect 17405 47104 17417 47107
rect 17368 47076 17417 47104
rect 17368 47064 17374 47076
rect 17405 47073 17417 47076
rect 17451 47073 17463 47107
rect 17696 47104 17724 47144
rect 17770 47132 17776 47184
rect 17828 47172 17834 47184
rect 18141 47175 18199 47181
rect 18141 47172 18153 47175
rect 17828 47144 18153 47172
rect 17828 47132 17834 47144
rect 18141 47141 18153 47144
rect 18187 47172 18199 47175
rect 18322 47172 18328 47184
rect 18187 47144 18328 47172
rect 18187 47141 18199 47144
rect 18141 47135 18199 47141
rect 18322 47132 18328 47144
rect 18380 47172 18386 47184
rect 20901 47175 20959 47181
rect 20901 47172 20913 47175
rect 18380 47144 20913 47172
rect 18380 47132 18386 47144
rect 20901 47141 20913 47144
rect 20947 47141 20959 47175
rect 22462 47172 22468 47184
rect 22423 47144 22468 47172
rect 20901 47135 20959 47141
rect 22462 47132 22468 47144
rect 22520 47132 22526 47184
rect 22756 47172 22784 47200
rect 23198 47172 23204 47184
rect 22756 47144 23204 47172
rect 17954 47104 17960 47116
rect 17696 47076 17960 47104
rect 17405 47067 17463 47073
rect 17954 47064 17960 47076
rect 18012 47064 18018 47116
rect 18966 47104 18972 47116
rect 18927 47076 18972 47104
rect 18966 47064 18972 47076
rect 19024 47064 19030 47116
rect 19150 47064 19156 47116
rect 19208 47104 19214 47116
rect 19245 47107 19303 47113
rect 19245 47104 19257 47107
rect 19208 47076 19257 47104
rect 19208 47064 19214 47076
rect 19245 47073 19257 47076
rect 19291 47104 19303 47107
rect 19702 47104 19708 47116
rect 19291 47076 19708 47104
rect 19291 47073 19303 47076
rect 19245 47067 19303 47073
rect 19702 47064 19708 47076
rect 19760 47104 19766 47116
rect 20165 47107 20223 47113
rect 20165 47104 20177 47107
rect 19760 47076 20177 47104
rect 19760 47064 19766 47076
rect 20165 47073 20177 47076
rect 20211 47073 20223 47107
rect 20990 47104 20996 47116
rect 20951 47076 20996 47104
rect 20165 47067 20223 47073
rect 20990 47064 20996 47076
rect 21048 47064 21054 47116
rect 21634 47064 21640 47116
rect 21692 47104 21698 47116
rect 22002 47104 22008 47116
rect 21692 47076 22008 47104
rect 21692 47064 21698 47076
rect 22002 47064 22008 47076
rect 22060 47064 22066 47116
rect 22738 47064 22744 47116
rect 22796 47104 22802 47116
rect 23124 47113 23152 47144
rect 23198 47132 23204 47144
rect 23256 47132 23262 47184
rect 22925 47107 22983 47113
rect 22925 47104 22937 47107
rect 22796 47076 22937 47104
rect 22796 47064 22802 47076
rect 22925 47073 22937 47076
rect 22971 47073 22983 47107
rect 22925 47067 22983 47073
rect 23109 47107 23167 47113
rect 23109 47073 23121 47107
rect 23155 47073 23167 47107
rect 23290 47104 23296 47116
rect 23251 47076 23296 47104
rect 23109 47067 23167 47073
rect 23290 47064 23296 47076
rect 23348 47064 23354 47116
rect 24504 47113 24532 47212
rect 26694 47200 26700 47212
rect 26752 47200 26758 47252
rect 24489 47107 24547 47113
rect 24489 47073 24501 47107
rect 24535 47104 24547 47107
rect 24762 47104 24768 47116
rect 24535 47076 24768 47104
rect 24535 47073 24547 47076
rect 24489 47067 24547 47073
rect 24762 47064 24768 47076
rect 24820 47064 24826 47116
rect 25314 47104 25320 47116
rect 25275 47076 25320 47104
rect 25314 47064 25320 47076
rect 25372 47064 25378 47116
rect 25682 47064 25688 47116
rect 25740 47064 25746 47116
rect 26510 47104 26516 47116
rect 26471 47076 26516 47104
rect 26510 47064 26516 47076
rect 26568 47064 26574 47116
rect 12618 47036 12624 47048
rect 12579 47008 12624 47036
rect 12618 46996 12624 47008
rect 12676 46996 12682 47048
rect 15194 46996 15200 47048
rect 15252 47036 15258 47048
rect 15381 47039 15439 47045
rect 15381 47036 15393 47039
rect 15252 47008 15393 47036
rect 15252 46996 15258 47008
rect 15381 47005 15393 47008
rect 15427 47005 15439 47039
rect 15381 46999 15439 47005
rect 16666 46996 16672 47048
rect 16724 47036 16730 47048
rect 18509 47039 18567 47045
rect 18509 47036 18521 47039
rect 16724 47008 18521 47036
rect 16724 46996 16730 47008
rect 18509 47005 18521 47008
rect 18555 47005 18567 47039
rect 18509 46999 18567 47005
rect 24302 46996 24308 47048
rect 24360 47036 24366 47048
rect 24581 47039 24639 47045
rect 24581 47036 24593 47039
rect 24360 47008 24593 47036
rect 24360 46996 24366 47008
rect 24581 47005 24593 47008
rect 24627 47005 24639 47039
rect 24581 46999 24639 47005
rect 25409 47039 25467 47045
rect 25409 47005 25421 47039
rect 25455 47005 25467 47039
rect 25409 46999 25467 47005
rect 16114 46968 16120 46980
rect 16075 46940 16120 46968
rect 16114 46928 16120 46940
rect 16172 46928 16178 46980
rect 17586 46968 17592 46980
rect 17547 46940 17592 46968
rect 17586 46928 17592 46940
rect 17644 46928 17650 46980
rect 18230 46928 18236 46980
rect 18288 46968 18294 46980
rect 19245 46971 19303 46977
rect 19245 46968 19257 46971
rect 18288 46940 19257 46968
rect 18288 46928 18294 46940
rect 19245 46937 19257 46940
rect 19291 46937 19303 46971
rect 19245 46931 19303 46937
rect 24486 46928 24492 46980
rect 24544 46968 24550 46980
rect 25424 46968 25452 46999
rect 25700 46968 25728 47064
rect 25777 46971 25835 46977
rect 25777 46968 25789 46971
rect 24544 46940 25789 46968
rect 24544 46928 24550 46940
rect 25777 46937 25789 46940
rect 25823 46937 25835 46971
rect 25777 46931 25835 46937
rect 19886 46900 19892 46912
rect 19847 46872 19892 46900
rect 19886 46860 19892 46872
rect 19944 46860 19950 46912
rect 21450 46860 21456 46912
rect 21508 46900 21514 46912
rect 21726 46900 21732 46912
rect 21508 46872 21732 46900
rect 21508 46860 21514 46872
rect 21726 46860 21732 46872
rect 21784 46860 21790 46912
rect 22002 46900 22008 46912
rect 21963 46872 22008 46900
rect 22002 46860 22008 46872
rect 22060 46860 22066 46912
rect 25866 46860 25872 46912
rect 25924 46900 25930 46912
rect 26145 46903 26203 46909
rect 26145 46900 26157 46903
rect 25924 46872 26157 46900
rect 25924 46860 25930 46872
rect 26145 46869 26157 46872
rect 26191 46869 26203 46903
rect 26145 46863 26203 46869
rect 1104 46810 28888 46832
rect 1104 46758 5982 46810
rect 6034 46758 6046 46810
rect 6098 46758 6110 46810
rect 6162 46758 6174 46810
rect 6226 46758 15982 46810
rect 16034 46758 16046 46810
rect 16098 46758 16110 46810
rect 16162 46758 16174 46810
rect 16226 46758 25982 46810
rect 26034 46758 26046 46810
rect 26098 46758 26110 46810
rect 26162 46758 26174 46810
rect 26226 46758 28888 46810
rect 1104 46736 28888 46758
rect 13541 46699 13599 46705
rect 13541 46665 13553 46699
rect 13587 46696 13599 46699
rect 13722 46696 13728 46708
rect 13587 46668 13728 46696
rect 13587 46665 13599 46668
rect 13541 46659 13599 46665
rect 13722 46656 13728 46668
rect 13780 46656 13786 46708
rect 14458 46696 14464 46708
rect 14419 46668 14464 46696
rect 14458 46656 14464 46668
rect 14516 46656 14522 46708
rect 14918 46696 14924 46708
rect 14879 46668 14924 46696
rect 14918 46656 14924 46668
rect 14976 46656 14982 46708
rect 15010 46656 15016 46708
rect 15068 46696 15074 46708
rect 15197 46699 15255 46705
rect 15197 46696 15209 46699
rect 15068 46668 15209 46696
rect 15068 46656 15074 46668
rect 15197 46665 15209 46668
rect 15243 46665 15255 46699
rect 15197 46659 15255 46665
rect 17310 46656 17316 46708
rect 17368 46696 17374 46708
rect 17405 46699 17463 46705
rect 17405 46696 17417 46699
rect 17368 46668 17417 46696
rect 17368 46656 17374 46668
rect 17405 46665 17417 46668
rect 17451 46696 17463 46699
rect 17678 46696 17684 46708
rect 17451 46668 17684 46696
rect 17451 46665 17463 46668
rect 17405 46659 17463 46665
rect 17678 46656 17684 46668
rect 17736 46656 17742 46708
rect 17865 46699 17923 46705
rect 17865 46665 17877 46699
rect 17911 46696 17923 46699
rect 18046 46696 18052 46708
rect 17911 46668 18052 46696
rect 17911 46665 17923 46668
rect 17865 46659 17923 46665
rect 18046 46656 18052 46668
rect 18104 46656 18110 46708
rect 23566 46696 23572 46708
rect 20548 46668 23572 46696
rect 12526 46628 12532 46640
rect 12487 46600 12532 46628
rect 12526 46588 12532 46600
rect 12584 46588 12590 46640
rect 19613 46631 19671 46637
rect 19613 46597 19625 46631
rect 19659 46628 19671 46631
rect 19659 46600 20300 46628
rect 19659 46597 19671 46600
rect 19613 46591 19671 46597
rect 15194 46520 15200 46572
rect 15252 46560 15258 46572
rect 15841 46563 15899 46569
rect 15841 46560 15853 46563
rect 15252 46532 15853 46560
rect 15252 46520 15258 46532
rect 15841 46529 15853 46532
rect 15887 46529 15899 46563
rect 15841 46523 15899 46529
rect 16114 46520 16120 46572
rect 16172 46560 16178 46572
rect 16172 46532 16436 46560
rect 16172 46520 16178 46532
rect 12253 46495 12311 46501
rect 12253 46461 12265 46495
rect 12299 46492 12311 46495
rect 12434 46492 12440 46504
rect 12299 46464 12440 46492
rect 12299 46461 12311 46464
rect 12253 46455 12311 46461
rect 12434 46452 12440 46464
rect 12492 46492 12498 46504
rect 12710 46492 12716 46504
rect 12492 46464 12585 46492
rect 12671 46464 12716 46492
rect 12492 46452 12498 46464
rect 12710 46452 12716 46464
rect 12768 46452 12774 46504
rect 15013 46495 15071 46501
rect 15013 46461 15025 46495
rect 15059 46492 15071 46495
rect 16206 46492 16212 46504
rect 15059 46464 15608 46492
rect 16167 46464 16212 46492
rect 15059 46461 15071 46464
rect 15013 46455 15071 46461
rect 15580 46368 15608 46464
rect 16206 46452 16212 46464
rect 16264 46452 16270 46504
rect 16408 46501 16436 46532
rect 17954 46520 17960 46572
rect 18012 46560 18018 46572
rect 18049 46563 18107 46569
rect 18049 46560 18061 46563
rect 18012 46532 18061 46560
rect 18012 46520 18018 46532
rect 18049 46529 18061 46532
rect 18095 46529 18107 46563
rect 18049 46523 18107 46529
rect 18785 46563 18843 46569
rect 18785 46529 18797 46563
rect 18831 46560 18843 46563
rect 19058 46560 19064 46572
rect 18831 46532 19064 46560
rect 18831 46529 18843 46532
rect 18785 46523 18843 46529
rect 19058 46520 19064 46532
rect 19116 46520 19122 46572
rect 19702 46560 19708 46572
rect 19663 46532 19708 46560
rect 19702 46520 19708 46532
rect 19760 46520 19766 46572
rect 20272 46569 20300 46600
rect 20257 46563 20315 46569
rect 20257 46529 20269 46563
rect 20303 46560 20315 46563
rect 20548 46560 20576 46668
rect 23566 46656 23572 46668
rect 23624 46656 23630 46708
rect 23676 46668 24532 46696
rect 21545 46631 21603 46637
rect 21545 46597 21557 46631
rect 21591 46597 21603 46631
rect 21545 46591 21603 46597
rect 20714 46560 20720 46572
rect 20303 46532 20576 46560
rect 20675 46532 20720 46560
rect 20303 46529 20315 46532
rect 20257 46523 20315 46529
rect 20714 46520 20720 46532
rect 20772 46520 20778 46572
rect 21560 46560 21588 46591
rect 21726 46588 21732 46640
rect 21784 46628 21790 46640
rect 21821 46631 21879 46637
rect 21821 46628 21833 46631
rect 21784 46600 21833 46628
rect 21784 46588 21790 46600
rect 21821 46597 21833 46600
rect 21867 46597 21879 46631
rect 21821 46591 21879 46597
rect 22094 46588 22100 46640
rect 22152 46628 22158 46640
rect 22462 46628 22468 46640
rect 22152 46600 22468 46628
rect 22152 46588 22158 46600
rect 22462 46588 22468 46600
rect 22520 46588 22526 46640
rect 23198 46588 23204 46640
rect 23256 46628 23262 46640
rect 23385 46631 23443 46637
rect 23385 46628 23397 46631
rect 23256 46600 23397 46628
rect 23256 46588 23262 46600
rect 23385 46597 23397 46600
rect 23431 46597 23443 46631
rect 23385 46591 23443 46597
rect 23474 46588 23480 46640
rect 23532 46628 23538 46640
rect 23676 46628 23704 46668
rect 24394 46628 24400 46640
rect 23532 46600 23704 46628
rect 24228 46600 24400 46628
rect 23532 46588 23538 46600
rect 22370 46560 22376 46572
rect 21560 46532 22376 46560
rect 22370 46520 22376 46532
rect 22428 46520 22434 46572
rect 24228 46569 24256 46600
rect 24394 46588 24400 46600
rect 24452 46588 24458 46640
rect 24504 46628 24532 46668
rect 26510 46656 26516 46708
rect 26568 46696 26574 46708
rect 26789 46699 26847 46705
rect 26789 46696 26801 46699
rect 26568 46668 26801 46696
rect 26568 46656 26574 46668
rect 26789 46665 26801 46668
rect 26835 46665 26847 46699
rect 26789 46659 26847 46665
rect 27157 46631 27215 46637
rect 27157 46628 27169 46631
rect 24504 46600 27169 46628
rect 27157 46597 27169 46600
rect 27203 46597 27215 46631
rect 27157 46591 27215 46597
rect 24213 46563 24271 46569
rect 24213 46529 24225 46563
rect 24259 46529 24271 46563
rect 24213 46523 24271 46529
rect 16393 46495 16451 46501
rect 16393 46461 16405 46495
rect 16439 46461 16451 46495
rect 16393 46455 16451 46461
rect 16853 46495 16911 46501
rect 16853 46461 16865 46495
rect 16899 46461 16911 46495
rect 18322 46492 18328 46504
rect 18283 46464 18328 46492
rect 16853 46455 16911 46461
rect 15746 46384 15752 46436
rect 15804 46424 15810 46436
rect 16868 46424 16896 46455
rect 18322 46452 18328 46464
rect 18380 46452 18386 46504
rect 19886 46452 19892 46504
rect 19944 46492 19950 46504
rect 20533 46495 20591 46501
rect 20533 46492 20545 46495
rect 19944 46464 20545 46492
rect 19944 46452 19950 46464
rect 20533 46461 20545 46464
rect 20579 46461 20591 46495
rect 20533 46455 20591 46461
rect 21729 46495 21787 46501
rect 21729 46461 21741 46495
rect 21775 46492 21787 46495
rect 21821 46495 21879 46501
rect 21821 46492 21833 46495
rect 21775 46464 21833 46492
rect 21775 46461 21787 46464
rect 21729 46455 21787 46461
rect 21821 46461 21833 46464
rect 21867 46461 21879 46495
rect 22189 46495 22247 46501
rect 22189 46492 22201 46495
rect 21821 46455 21879 46461
rect 21928 46464 22201 46492
rect 17126 46424 17132 46436
rect 15804 46396 16896 46424
rect 17087 46396 17132 46424
rect 15804 46384 15810 46396
rect 17126 46384 17132 46396
rect 17184 46384 17190 46436
rect 18233 46427 18291 46433
rect 18233 46393 18245 46427
rect 18279 46424 18291 46427
rect 18782 46424 18788 46436
rect 18279 46396 18788 46424
rect 18279 46393 18291 46396
rect 18233 46387 18291 46393
rect 18782 46384 18788 46396
rect 18840 46384 18846 46436
rect 19334 46384 19340 46436
rect 19392 46424 19398 46436
rect 19702 46424 19708 46436
rect 19392 46396 19708 46424
rect 19392 46384 19398 46396
rect 19702 46384 19708 46396
rect 19760 46384 19766 46436
rect 19794 46384 19800 46436
rect 19852 46424 19858 46436
rect 20990 46424 20996 46436
rect 19852 46396 20996 46424
rect 19852 46384 19858 46396
rect 20990 46384 20996 46396
rect 21048 46384 21054 46436
rect 21928 46424 21956 46464
rect 22189 46461 22201 46464
rect 22235 46492 22247 46495
rect 23474 46492 23480 46504
rect 22235 46464 23480 46492
rect 22235 46461 22247 46464
rect 22189 46455 22247 46461
rect 23474 46452 23480 46464
rect 23532 46452 23538 46504
rect 23753 46495 23811 46501
rect 23753 46461 23765 46495
rect 23799 46492 23811 46495
rect 24397 46495 24455 46501
rect 24397 46492 24409 46495
rect 23799 46464 24409 46492
rect 23799 46461 23811 46464
rect 23753 46455 23811 46461
rect 24397 46461 24409 46464
rect 24443 46461 24455 46495
rect 24854 46492 24860 46504
rect 24815 46464 24860 46492
rect 24397 46455 24455 46461
rect 24854 46452 24860 46464
rect 24912 46492 24918 46504
rect 25409 46495 25467 46501
rect 25409 46492 25421 46495
rect 24912 46464 25421 46492
rect 24912 46452 24918 46464
rect 25409 46461 25421 46464
rect 25455 46461 25467 46495
rect 25958 46492 25964 46504
rect 25919 46464 25964 46492
rect 25409 46455 25467 46461
rect 25958 46452 25964 46464
rect 26016 46452 26022 46504
rect 26053 46495 26111 46501
rect 26053 46461 26065 46495
rect 26099 46461 26111 46495
rect 26053 46455 26111 46461
rect 21376 46396 21956 46424
rect 22005 46427 22063 46433
rect 11882 46356 11888 46368
rect 11843 46328 11888 46356
rect 11882 46316 11888 46328
rect 11940 46316 11946 46368
rect 12342 46316 12348 46368
rect 12400 46356 12406 46368
rect 12897 46359 12955 46365
rect 12897 46356 12909 46359
rect 12400 46328 12909 46356
rect 12400 46316 12406 46328
rect 12897 46325 12909 46328
rect 12943 46325 12955 46359
rect 14182 46356 14188 46368
rect 14143 46328 14188 46356
rect 12897 46319 12955 46325
rect 14182 46316 14188 46328
rect 14240 46316 14246 46368
rect 15562 46356 15568 46368
rect 15523 46328 15568 46356
rect 15562 46316 15568 46328
rect 15620 46316 15626 46368
rect 19150 46356 19156 46368
rect 19111 46328 19156 46356
rect 19150 46316 19156 46328
rect 19208 46316 19214 46368
rect 20346 46316 20352 46368
rect 20404 46356 20410 46368
rect 21376 46365 21404 46396
rect 22005 46393 22017 46427
rect 22051 46393 22063 46427
rect 22373 46427 22431 46433
rect 22373 46424 22385 46427
rect 22005 46387 22063 46393
rect 22204 46396 22385 46424
rect 21361 46359 21419 46365
rect 21361 46356 21373 46359
rect 20404 46328 21373 46356
rect 20404 46316 20410 46328
rect 21361 46325 21373 46328
rect 21407 46325 21419 46359
rect 22020 46356 22048 46387
rect 22204 46368 22232 46396
rect 22373 46393 22385 46396
rect 22419 46393 22431 46427
rect 22738 46424 22744 46436
rect 22699 46396 22744 46424
rect 22373 46387 22431 46393
rect 22738 46384 22744 46396
rect 22796 46384 22802 46436
rect 25130 46424 25136 46436
rect 23032 46396 24992 46424
rect 25091 46396 25136 46424
rect 22094 46356 22100 46368
rect 22020 46328 22100 46356
rect 21361 46319 21419 46325
rect 22094 46316 22100 46328
rect 22152 46316 22158 46368
rect 22186 46316 22192 46368
rect 22244 46316 22250 46368
rect 22281 46359 22339 46365
rect 22281 46325 22293 46359
rect 22327 46356 22339 46359
rect 22462 46356 22468 46368
rect 22327 46328 22468 46356
rect 22327 46325 22339 46328
rect 22281 46319 22339 46325
rect 22462 46316 22468 46328
rect 22520 46356 22526 46368
rect 23032 46365 23060 46396
rect 23017 46359 23075 46365
rect 23017 46356 23029 46359
rect 22520 46328 23029 46356
rect 22520 46316 22526 46328
rect 23017 46325 23029 46328
rect 23063 46325 23075 46359
rect 23017 46319 23075 46325
rect 23566 46316 23572 46368
rect 23624 46356 23630 46368
rect 23753 46359 23811 46365
rect 23753 46356 23765 46359
rect 23624 46328 23765 46356
rect 23624 46316 23630 46328
rect 23753 46325 23765 46328
rect 23799 46356 23811 46359
rect 23845 46359 23903 46365
rect 23845 46356 23857 46359
rect 23799 46328 23857 46356
rect 23799 46325 23811 46328
rect 23753 46319 23811 46325
rect 23845 46325 23857 46328
rect 23891 46325 23903 46359
rect 23845 46319 23903 46325
rect 23934 46316 23940 46368
rect 23992 46356 23998 46368
rect 24762 46356 24768 46368
rect 23992 46328 24768 46356
rect 23992 46316 23998 46328
rect 24762 46316 24768 46328
rect 24820 46316 24826 46368
rect 24964 46356 24992 46396
rect 25130 46384 25136 46396
rect 25188 46384 25194 46436
rect 25038 46356 25044 46368
rect 24964 46328 25044 46356
rect 25038 46316 25044 46328
rect 25096 46316 25102 46368
rect 25869 46359 25927 46365
rect 25869 46325 25881 46359
rect 25915 46356 25927 46359
rect 26068 46356 26096 46455
rect 26510 46424 26516 46436
rect 26471 46396 26516 46424
rect 26510 46384 26516 46396
rect 26568 46384 26574 46436
rect 26326 46356 26332 46368
rect 25915 46328 26332 46356
rect 25915 46325 25927 46328
rect 25869 46319 25927 46325
rect 26326 46316 26332 46328
rect 26384 46316 26390 46368
rect 1104 46266 28888 46288
rect 1104 46214 10982 46266
rect 11034 46214 11046 46266
rect 11098 46214 11110 46266
rect 11162 46214 11174 46266
rect 11226 46214 20982 46266
rect 21034 46214 21046 46266
rect 21098 46214 21110 46266
rect 21162 46214 21174 46266
rect 21226 46214 28888 46266
rect 1104 46192 28888 46214
rect 11882 46152 11888 46164
rect 11843 46124 11888 46152
rect 11882 46112 11888 46124
rect 11940 46152 11946 46164
rect 12253 46155 12311 46161
rect 12253 46152 12265 46155
rect 11940 46124 12265 46152
rect 11940 46112 11946 46124
rect 12253 46121 12265 46124
rect 12299 46121 12311 46155
rect 12253 46115 12311 46121
rect 12268 45948 12296 46115
rect 14090 46112 14096 46164
rect 14148 46152 14154 46164
rect 15013 46155 15071 46161
rect 15013 46152 15025 46155
rect 14148 46124 15025 46152
rect 14148 46112 14154 46124
rect 15013 46121 15025 46124
rect 15059 46152 15071 46155
rect 16114 46152 16120 46164
rect 15059 46124 16120 46152
rect 15059 46121 15071 46124
rect 15013 46115 15071 46121
rect 16114 46112 16120 46124
rect 16172 46112 16178 46164
rect 16206 46112 16212 46164
rect 16264 46152 16270 46164
rect 16669 46155 16727 46161
rect 16669 46152 16681 46155
rect 16264 46124 16681 46152
rect 16264 46112 16270 46124
rect 16669 46121 16681 46124
rect 16715 46121 16727 46155
rect 16669 46115 16727 46121
rect 17218 46112 17224 46164
rect 17276 46112 17282 46164
rect 17494 46152 17500 46164
rect 17455 46124 17500 46152
rect 17494 46112 17500 46124
rect 17552 46112 17558 46164
rect 18693 46155 18751 46161
rect 18693 46121 18705 46155
rect 18739 46152 18751 46155
rect 18782 46152 18788 46164
rect 18739 46124 18788 46152
rect 18739 46121 18751 46124
rect 18693 46115 18751 46121
rect 18782 46112 18788 46124
rect 18840 46112 18846 46164
rect 19705 46155 19763 46161
rect 19705 46121 19717 46155
rect 19751 46152 19763 46155
rect 19794 46152 19800 46164
rect 19751 46124 19800 46152
rect 19751 46121 19763 46124
rect 19705 46115 19763 46121
rect 19794 46112 19800 46124
rect 19852 46112 19858 46164
rect 23198 46112 23204 46164
rect 23256 46152 23262 46164
rect 23256 46124 23428 46152
rect 23256 46112 23262 46124
rect 13262 46044 13268 46096
rect 13320 46084 13326 46096
rect 15562 46084 15568 46096
rect 13320 46056 15568 46084
rect 13320 46044 13326 46056
rect 15562 46044 15568 46056
rect 15620 46044 15626 46096
rect 17236 46084 17264 46112
rect 20625 46087 20683 46093
rect 17236 46056 17724 46084
rect 12434 45976 12440 46028
rect 12492 46016 12498 46028
rect 12492 45988 12537 46016
rect 12492 45976 12498 45988
rect 12710 45976 12716 46028
rect 12768 46016 12774 46028
rect 13446 46016 13452 46028
rect 12768 45988 13452 46016
rect 12768 45976 12774 45988
rect 13446 45976 13452 45988
rect 13504 45976 13510 46028
rect 15470 46016 15476 46028
rect 15431 45988 15476 46016
rect 15470 45976 15476 45988
rect 15528 45976 15534 46028
rect 15657 46019 15715 46025
rect 15657 45985 15669 46019
rect 15703 45985 15715 46019
rect 15657 45979 15715 45985
rect 12728 45948 12756 45976
rect 12268 45920 12756 45948
rect 13173 45951 13231 45957
rect 13173 45917 13185 45951
rect 13219 45948 13231 45951
rect 13814 45948 13820 45960
rect 13219 45920 13820 45948
rect 13219 45917 13231 45920
rect 13173 45911 13231 45917
rect 13814 45908 13820 45920
rect 13872 45908 13878 45960
rect 14182 45908 14188 45960
rect 14240 45948 14246 45960
rect 15672 45948 15700 45979
rect 15746 45976 15752 46028
rect 15804 46016 15810 46028
rect 16117 46019 16175 46025
rect 16117 46016 16129 46019
rect 15804 45988 16129 46016
rect 15804 45976 15810 45988
rect 16117 45985 16129 45988
rect 16163 45985 16175 46019
rect 16117 45979 16175 45985
rect 16574 45976 16580 46028
rect 16632 46016 16638 46028
rect 17034 46016 17040 46028
rect 16632 45988 17040 46016
rect 16632 45976 16638 45988
rect 17034 45976 17040 45988
rect 17092 46016 17098 46028
rect 17696 46025 17724 46056
rect 20625 46053 20637 46087
rect 20671 46084 20683 46087
rect 22738 46084 22744 46096
rect 20671 46056 22744 46084
rect 20671 46053 20683 46056
rect 20625 46047 20683 46053
rect 22738 46044 22744 46056
rect 22796 46044 22802 46096
rect 17221 46019 17279 46025
rect 17221 46016 17233 46019
rect 17092 45988 17233 46016
rect 17092 45976 17098 45988
rect 17221 45985 17233 45988
rect 17267 45985 17279 46019
rect 17221 45979 17279 45985
rect 17681 46019 17739 46025
rect 17681 45985 17693 46019
rect 17727 45985 17739 46019
rect 17681 45979 17739 45985
rect 19058 45976 19064 46028
rect 19116 46016 19122 46028
rect 19245 46019 19303 46025
rect 19245 46016 19257 46019
rect 19116 45988 19257 46016
rect 19116 45976 19122 45988
rect 19245 45985 19257 45988
rect 19291 45985 19303 46019
rect 19245 45979 19303 45985
rect 19426 45976 19432 46028
rect 19484 46016 19490 46028
rect 19521 46019 19579 46025
rect 19521 46016 19533 46019
rect 19484 45988 19533 46016
rect 19484 45976 19490 45988
rect 19521 45985 19533 45988
rect 19567 45985 19579 46019
rect 19521 45979 19579 45985
rect 20714 45976 20720 46028
rect 20772 46016 20778 46028
rect 20901 46019 20959 46025
rect 20901 46016 20913 46019
rect 20772 45988 20913 46016
rect 20772 45976 20778 45988
rect 20901 45985 20913 45988
rect 20947 45985 20959 46019
rect 21082 46016 21088 46028
rect 21043 45988 21088 46016
rect 20901 45979 20959 45985
rect 21082 45976 21088 45988
rect 21140 45976 21146 46028
rect 22925 46019 22983 46025
rect 22925 45985 22937 46019
rect 22971 46016 22983 46019
rect 23198 46016 23204 46028
rect 22971 45988 23204 46016
rect 22971 45985 22983 45988
rect 22925 45979 22983 45985
rect 23198 45976 23204 45988
rect 23256 45976 23262 46028
rect 23400 46025 23428 46124
rect 23474 46112 23480 46164
rect 23532 46112 23538 46164
rect 24121 46155 24179 46161
rect 24121 46121 24133 46155
rect 24167 46152 24179 46155
rect 24394 46152 24400 46164
rect 24167 46124 24400 46152
rect 24167 46121 24179 46124
rect 24121 46115 24179 46121
rect 24394 46112 24400 46124
rect 24452 46112 24458 46164
rect 24581 46155 24639 46161
rect 24581 46121 24593 46155
rect 24627 46152 24639 46155
rect 24670 46152 24676 46164
rect 24627 46124 24676 46152
rect 24627 46121 24639 46124
rect 24581 46115 24639 46121
rect 24670 46112 24676 46124
rect 24728 46112 24734 46164
rect 25314 46112 25320 46164
rect 25372 46152 25378 46164
rect 25961 46155 26019 46161
rect 25961 46152 25973 46155
rect 25372 46124 25973 46152
rect 25372 46112 25378 46124
rect 25961 46121 25973 46124
rect 26007 46121 26019 46155
rect 25961 46115 26019 46121
rect 23492 46084 23520 46112
rect 25593 46087 25651 46093
rect 25593 46084 25605 46087
rect 23492 46056 25605 46084
rect 25593 46053 25605 46056
rect 25639 46084 25651 46087
rect 25774 46084 25780 46096
rect 25639 46056 25780 46084
rect 25639 46053 25651 46056
rect 25593 46047 25651 46053
rect 25774 46044 25780 46056
rect 25832 46044 25838 46096
rect 23293 46019 23351 46025
rect 23293 45985 23305 46019
rect 23339 45985 23351 46019
rect 23293 45979 23351 45985
rect 23385 46019 23443 46025
rect 23385 45985 23397 46019
rect 23431 46016 23443 46019
rect 23474 46016 23480 46028
rect 23431 45988 23480 46016
rect 23431 45985 23443 45988
rect 23385 45979 23443 45985
rect 16482 45948 16488 45960
rect 14240 45920 16488 45948
rect 14240 45908 14246 45920
rect 16482 45908 16488 45920
rect 16540 45908 16546 45960
rect 19150 45948 19156 45960
rect 19063 45920 19156 45948
rect 19150 45908 19156 45920
rect 19208 45948 19214 45960
rect 19337 45951 19395 45957
rect 19337 45948 19349 45951
rect 19208 45920 19349 45948
rect 19208 45908 19214 45920
rect 19337 45917 19349 45920
rect 19383 45948 19395 45951
rect 20732 45948 20760 45976
rect 19383 45920 20760 45948
rect 19383 45917 19395 45920
rect 19337 45911 19395 45917
rect 22554 45908 22560 45960
rect 22612 45948 22618 45960
rect 23308 45948 23336 45979
rect 23474 45976 23480 45988
rect 23532 45976 23538 46028
rect 24118 45976 24124 46028
rect 24176 46016 24182 46028
rect 24305 46019 24363 46025
rect 24305 46016 24317 46019
rect 24176 45988 24317 46016
rect 24176 45976 24182 45988
rect 24305 45985 24317 45988
rect 24351 45985 24363 46019
rect 24305 45979 24363 45985
rect 24857 46019 24915 46025
rect 24857 45985 24869 46019
rect 24903 45985 24915 46019
rect 25958 46016 25964 46028
rect 24857 45979 24915 45985
rect 25884 45988 25964 46016
rect 22612 45920 23336 45948
rect 24320 45948 24348 45979
rect 24486 45948 24492 45960
rect 24320 45920 24492 45948
rect 22612 45908 22618 45920
rect 24486 45908 24492 45920
rect 24544 45908 24550 45960
rect 24872 45892 24900 45979
rect 12529 45883 12587 45889
rect 12529 45849 12541 45883
rect 12575 45880 12587 45883
rect 12618 45880 12624 45892
rect 12575 45852 12624 45880
rect 12575 45849 12587 45852
rect 12529 45843 12587 45849
rect 12618 45840 12624 45852
rect 12676 45840 12682 45892
rect 16114 45880 16120 45892
rect 16075 45852 16120 45880
rect 16114 45840 16120 45852
rect 16172 45840 16178 45892
rect 16666 45840 16672 45892
rect 16724 45880 16730 45892
rect 17037 45883 17095 45889
rect 17037 45880 17049 45883
rect 16724 45852 17049 45880
rect 16724 45840 16730 45852
rect 17037 45849 17049 45852
rect 17083 45849 17095 45883
rect 17037 45843 17095 45849
rect 22741 45883 22799 45889
rect 22741 45849 22753 45883
rect 22787 45880 22799 45883
rect 24854 45880 24860 45892
rect 22787 45852 24860 45880
rect 22787 45849 22799 45852
rect 22741 45843 22799 45849
rect 24854 45840 24860 45852
rect 24912 45840 24918 45892
rect 25884 45824 25912 45988
rect 25958 45976 25964 45988
rect 26016 45976 26022 46028
rect 1578 45812 1584 45824
rect 1539 45784 1584 45812
rect 1578 45772 1584 45784
rect 1636 45772 1642 45824
rect 14458 45812 14464 45824
rect 14419 45784 14464 45812
rect 14458 45772 14464 45784
rect 14516 45772 14522 45824
rect 18322 45812 18328 45824
rect 18283 45784 18328 45812
rect 18322 45772 18328 45784
rect 18380 45772 18386 45824
rect 20070 45772 20076 45824
rect 20128 45812 20134 45824
rect 20257 45815 20315 45821
rect 20257 45812 20269 45815
rect 20128 45784 20269 45812
rect 20128 45772 20134 45784
rect 20257 45781 20269 45784
rect 20303 45812 20315 45815
rect 20898 45812 20904 45824
rect 20303 45784 20904 45812
rect 20303 45781 20315 45784
rect 20257 45775 20315 45781
rect 20898 45772 20904 45784
rect 20956 45812 20962 45824
rect 22005 45815 22063 45821
rect 22005 45812 22017 45815
rect 20956 45784 22017 45812
rect 20956 45772 20962 45784
rect 22005 45781 22017 45784
rect 22051 45812 22063 45815
rect 22094 45812 22100 45824
rect 22051 45784 22100 45812
rect 22051 45781 22063 45784
rect 22005 45775 22063 45781
rect 22094 45772 22100 45784
rect 22152 45812 22158 45824
rect 23290 45812 23296 45824
rect 22152 45784 23296 45812
rect 22152 45772 22158 45784
rect 23290 45772 23296 45784
rect 23348 45772 23354 45824
rect 23934 45772 23940 45824
rect 23992 45812 23998 45824
rect 24394 45812 24400 45824
rect 23992 45784 24400 45812
rect 23992 45772 23998 45784
rect 24394 45772 24400 45784
rect 24452 45772 24458 45824
rect 25866 45772 25872 45824
rect 25924 45772 25930 45824
rect 1104 45722 28888 45744
rect 1104 45670 5982 45722
rect 6034 45670 6046 45722
rect 6098 45670 6110 45722
rect 6162 45670 6174 45722
rect 6226 45670 15982 45722
rect 16034 45670 16046 45722
rect 16098 45670 16110 45722
rect 16162 45670 16174 45722
rect 16226 45670 25982 45722
rect 26034 45670 26046 45722
rect 26098 45670 26110 45722
rect 26162 45670 26174 45722
rect 26226 45670 28888 45722
rect 1104 45648 28888 45670
rect 12250 45568 12256 45620
rect 12308 45608 12314 45620
rect 12529 45611 12587 45617
rect 12529 45608 12541 45611
rect 12308 45580 12541 45608
rect 12308 45568 12314 45580
rect 12529 45577 12541 45580
rect 12575 45577 12587 45611
rect 12529 45571 12587 45577
rect 14921 45611 14979 45617
rect 14921 45577 14933 45611
rect 14967 45577 14979 45611
rect 15470 45608 15476 45620
rect 15431 45580 15476 45608
rect 14921 45571 14979 45577
rect 11241 45543 11299 45549
rect 11241 45509 11253 45543
rect 11287 45540 11299 45543
rect 12342 45540 12348 45552
rect 11287 45512 12348 45540
rect 11287 45509 11299 45512
rect 11241 45503 11299 45509
rect 1397 45475 1455 45481
rect 1397 45441 1409 45475
rect 1443 45472 1455 45475
rect 1578 45472 1584 45484
rect 1443 45444 1584 45472
rect 1443 45441 1455 45444
rect 1397 45435 1455 45441
rect 1578 45432 1584 45444
rect 1636 45432 1642 45484
rect 1673 45475 1731 45481
rect 1673 45441 1685 45475
rect 1719 45472 1731 45475
rect 1762 45472 1768 45484
rect 1719 45444 1768 45472
rect 1719 45441 1731 45444
rect 1673 45435 1731 45441
rect 1762 45432 1768 45444
rect 1820 45432 1826 45484
rect 11348 45413 11376 45512
rect 12342 45500 12348 45512
rect 12400 45500 12406 45552
rect 13906 45500 13912 45552
rect 13964 45540 13970 45552
rect 14936 45540 14964 45571
rect 15470 45568 15476 45580
rect 15528 45568 15534 45620
rect 17218 45608 17224 45620
rect 16500 45580 17224 45608
rect 16500 45549 16528 45580
rect 17218 45568 17224 45580
rect 17276 45568 17282 45620
rect 17678 45568 17684 45620
rect 17736 45608 17742 45620
rect 18690 45608 18696 45620
rect 17736 45580 18696 45608
rect 17736 45568 17742 45580
rect 18690 45568 18696 45580
rect 18748 45568 18754 45620
rect 18874 45568 18880 45620
rect 18932 45608 18938 45620
rect 19705 45611 19763 45617
rect 19705 45608 19717 45611
rect 18932 45580 19717 45608
rect 18932 45568 18938 45580
rect 19705 45577 19717 45580
rect 19751 45577 19763 45611
rect 19705 45571 19763 45577
rect 20714 45568 20720 45620
rect 20772 45608 20778 45620
rect 21082 45608 21088 45620
rect 20772 45580 21088 45608
rect 20772 45568 20778 45580
rect 21082 45568 21088 45580
rect 21140 45608 21146 45620
rect 21361 45611 21419 45617
rect 21361 45608 21373 45611
rect 21140 45580 21373 45608
rect 21140 45568 21146 45580
rect 21361 45577 21373 45580
rect 21407 45577 21419 45611
rect 21361 45571 21419 45577
rect 22738 45568 22744 45620
rect 22796 45608 22802 45620
rect 23017 45611 23075 45617
rect 23017 45608 23029 45611
rect 22796 45580 23029 45608
rect 22796 45568 22802 45580
rect 23017 45577 23029 45580
rect 23063 45608 23075 45611
rect 23474 45608 23480 45620
rect 23063 45580 23480 45608
rect 23063 45577 23075 45580
rect 23017 45571 23075 45577
rect 23474 45568 23480 45580
rect 23532 45568 23538 45620
rect 23658 45568 23664 45620
rect 23716 45568 23722 45620
rect 24486 45568 24492 45620
rect 24544 45608 24550 45620
rect 25041 45611 25099 45617
rect 25041 45608 25053 45611
rect 24544 45580 25053 45608
rect 24544 45568 24550 45580
rect 25041 45577 25053 45580
rect 25087 45577 25099 45611
rect 25041 45571 25099 45577
rect 13964 45512 14964 45540
rect 16485 45543 16543 45549
rect 13964 45500 13970 45512
rect 16485 45509 16497 45543
rect 16531 45509 16543 45543
rect 16485 45503 16543 45509
rect 17129 45543 17187 45549
rect 17129 45509 17141 45543
rect 17175 45540 17187 45543
rect 17770 45540 17776 45552
rect 17175 45512 17776 45540
rect 17175 45509 17187 45512
rect 17129 45503 17187 45509
rect 17770 45500 17776 45512
rect 17828 45500 17834 45552
rect 17865 45543 17923 45549
rect 17865 45509 17877 45543
rect 17911 45540 17923 45543
rect 18141 45543 18199 45549
rect 18141 45540 18153 45543
rect 17911 45512 18153 45540
rect 17911 45509 17923 45512
rect 17865 45503 17923 45509
rect 18141 45509 18153 45512
rect 18187 45540 18199 45543
rect 19794 45540 19800 45552
rect 18187 45512 19800 45540
rect 18187 45509 18199 45512
rect 18141 45503 18199 45509
rect 13630 45472 13636 45484
rect 12544 45444 13636 45472
rect 11333 45407 11391 45413
rect 11333 45373 11345 45407
rect 11379 45373 11391 45407
rect 11333 45367 11391 45373
rect 11885 45407 11943 45413
rect 11885 45373 11897 45407
rect 11931 45404 11943 45407
rect 12434 45404 12440 45416
rect 11931 45376 12440 45404
rect 11931 45373 11943 45376
rect 11885 45367 11943 45373
rect 12434 45364 12440 45376
rect 12492 45404 12498 45416
rect 12544 45413 12572 45444
rect 13630 45432 13636 45444
rect 13688 45472 13694 45484
rect 14001 45475 14059 45481
rect 14001 45472 14013 45475
rect 13688 45444 14013 45472
rect 13688 45432 13694 45444
rect 14001 45441 14013 45444
rect 14047 45472 14059 45475
rect 14369 45475 14427 45481
rect 14369 45472 14381 45475
rect 14047 45444 14381 45472
rect 14047 45441 14059 45444
rect 14001 45435 14059 45441
rect 14369 45441 14381 45444
rect 14415 45472 14427 45475
rect 14415 45444 14780 45472
rect 14415 45441 14427 45444
rect 14369 45435 14427 45441
rect 12529 45407 12587 45413
rect 12529 45404 12541 45407
rect 12492 45376 12541 45404
rect 12492 45364 12498 45376
rect 12529 45373 12541 45376
rect 12575 45373 12587 45407
rect 12529 45367 12587 45373
rect 12618 45364 12624 45416
rect 12676 45404 12682 45416
rect 12805 45407 12863 45413
rect 12805 45404 12817 45407
rect 12676 45376 12817 45404
rect 12676 45364 12682 45376
rect 12805 45373 12817 45376
rect 12851 45373 12863 45407
rect 13446 45404 13452 45416
rect 13359 45376 13452 45404
rect 12805 45367 12863 45373
rect 13446 45364 13452 45376
rect 13504 45404 13510 45416
rect 14090 45404 14096 45416
rect 13504 45376 14096 45404
rect 13504 45364 13510 45376
rect 14090 45364 14096 45376
rect 14148 45404 14154 45416
rect 14458 45404 14464 45416
rect 14148 45376 14464 45404
rect 14148 45364 14154 45376
rect 14458 45364 14464 45376
rect 14516 45364 14522 45416
rect 14752 45413 14780 45444
rect 17402 45432 17408 45484
rect 17460 45472 17466 45484
rect 17880 45472 17908 45503
rect 19794 45500 19800 45512
rect 19852 45500 19858 45552
rect 23676 45540 23704 45568
rect 24670 45540 24676 45552
rect 23492 45512 23704 45540
rect 23768 45512 24676 45540
rect 17460 45444 17908 45472
rect 18785 45475 18843 45481
rect 17460 45432 17466 45444
rect 18785 45441 18797 45475
rect 18831 45472 18843 45475
rect 18966 45472 18972 45484
rect 18831 45444 18972 45472
rect 18831 45441 18843 45444
rect 18785 45435 18843 45441
rect 18966 45432 18972 45444
rect 19024 45432 19030 45484
rect 23492 45481 23520 45512
rect 23477 45475 23535 45481
rect 23477 45441 23489 45475
rect 23523 45441 23535 45475
rect 23477 45435 23535 45441
rect 14737 45407 14795 45413
rect 14737 45373 14749 45407
rect 14783 45373 14795 45407
rect 14737 45367 14795 45373
rect 15933 45407 15991 45413
rect 15933 45373 15945 45407
rect 15979 45404 15991 45407
rect 16482 45404 16488 45416
rect 15979 45376 16488 45404
rect 15979 45373 15991 45376
rect 15933 45367 15991 45373
rect 16482 45364 16488 45376
rect 16540 45364 16546 45416
rect 16853 45407 16911 45413
rect 16853 45373 16865 45407
rect 16899 45404 16911 45407
rect 16945 45407 17003 45413
rect 16945 45404 16957 45407
rect 16899 45376 16957 45404
rect 16899 45373 16911 45376
rect 16853 45367 16911 45373
rect 16945 45373 16957 45376
rect 16991 45404 17003 45407
rect 17218 45404 17224 45416
rect 16991 45376 17224 45404
rect 16991 45373 17003 45376
rect 16945 45367 17003 45373
rect 17218 45364 17224 45376
rect 17276 45364 17282 45416
rect 18049 45407 18107 45413
rect 18049 45373 18061 45407
rect 18095 45373 18107 45407
rect 18322 45404 18328 45416
rect 18283 45376 18328 45404
rect 18049 45367 18107 45373
rect 3053 45339 3111 45345
rect 3053 45305 3065 45339
rect 3099 45336 3111 45339
rect 4062 45336 4068 45348
rect 3099 45308 4068 45336
rect 3099 45305 3111 45308
rect 3053 45299 3111 45305
rect 4062 45296 4068 45308
rect 4120 45296 4126 45348
rect 12253 45339 12311 45345
rect 12253 45305 12265 45339
rect 12299 45336 12311 45339
rect 12636 45336 12664 45364
rect 12299 45308 12664 45336
rect 12299 45305 12311 45308
rect 12253 45299 12311 45305
rect 13998 45296 14004 45348
rect 14056 45336 14062 45348
rect 14550 45336 14556 45348
rect 14056 45308 14556 45336
rect 14056 45296 14062 45308
rect 14550 45296 14556 45308
rect 14608 45336 14614 45348
rect 14645 45339 14703 45345
rect 14645 45336 14657 45339
rect 14608 45308 14657 45336
rect 14608 45296 14614 45308
rect 14645 45305 14657 45308
rect 14691 45305 14703 45339
rect 14645 45299 14703 45305
rect 17497 45339 17555 45345
rect 17497 45305 17509 45339
rect 17543 45336 17555 45339
rect 17586 45336 17592 45348
rect 17543 45308 17592 45336
rect 17543 45305 17555 45308
rect 17497 45299 17555 45305
rect 17586 45296 17592 45308
rect 17644 45336 17650 45348
rect 18064 45336 18092 45367
rect 18322 45364 18328 45376
rect 18380 45364 18386 45416
rect 19426 45364 19432 45416
rect 19484 45404 19490 45416
rect 19613 45407 19671 45413
rect 19613 45404 19625 45407
rect 19484 45376 19625 45404
rect 19484 45364 19490 45376
rect 19613 45373 19625 45376
rect 19659 45373 19671 45407
rect 19978 45404 19984 45416
rect 19939 45376 19984 45404
rect 19613 45367 19671 45373
rect 19978 45364 19984 45376
rect 20036 45364 20042 45416
rect 20346 45404 20352 45416
rect 20307 45376 20352 45404
rect 20346 45364 20352 45376
rect 20404 45364 20410 45416
rect 20898 45404 20904 45416
rect 20859 45376 20904 45404
rect 20898 45364 20904 45376
rect 20956 45364 20962 45416
rect 21913 45407 21971 45413
rect 21913 45404 21925 45407
rect 21744 45376 21925 45404
rect 19058 45336 19064 45348
rect 17644 45308 19064 45336
rect 17644 45296 17650 45308
rect 19058 45296 19064 45308
rect 19116 45296 19122 45348
rect 21744 45280 21772 45376
rect 21913 45373 21925 45376
rect 21959 45373 21971 45407
rect 21913 45367 21971 45373
rect 22002 45364 22008 45416
rect 22060 45404 22066 45416
rect 22370 45404 22376 45416
rect 22060 45376 22376 45404
rect 22060 45364 22066 45376
rect 22370 45364 22376 45376
rect 22428 45364 22434 45416
rect 22646 45336 22652 45348
rect 22607 45308 22652 45336
rect 22646 45296 22652 45308
rect 22704 45296 22710 45348
rect 11514 45268 11520 45280
rect 11475 45240 11520 45268
rect 11514 45228 11520 45240
rect 11572 45228 11578 45280
rect 19334 45268 19340 45280
rect 19295 45240 19340 45268
rect 19334 45228 19340 45240
rect 19392 45228 19398 45280
rect 21726 45268 21732 45280
rect 21687 45240 21732 45268
rect 21726 45228 21732 45240
rect 21784 45228 21790 45280
rect 23492 45268 23520 45435
rect 23658 45432 23664 45484
rect 23716 45472 23722 45484
rect 23768 45481 23796 45512
rect 24670 45500 24676 45512
rect 24728 45500 24734 45552
rect 23753 45475 23811 45481
rect 23753 45472 23765 45475
rect 23716 45444 23765 45472
rect 23716 45432 23722 45444
rect 23753 45441 23765 45444
rect 23799 45441 23811 45475
rect 23753 45435 23811 45441
rect 24596 45444 26004 45472
rect 24486 45364 24492 45416
rect 24544 45404 24550 45416
rect 24596 45413 24624 45444
rect 24581 45407 24639 45413
rect 24581 45404 24593 45407
rect 24544 45376 24593 45404
rect 24544 45364 24550 45376
rect 24581 45373 24593 45376
rect 24627 45373 24639 45407
rect 24581 45367 24639 45373
rect 24673 45407 24731 45413
rect 24673 45373 24685 45407
rect 24719 45373 24731 45407
rect 24673 45367 24731 45373
rect 23842 45336 23848 45348
rect 23803 45308 23848 45336
rect 23842 45296 23848 45308
rect 23900 45296 23906 45348
rect 24688 45280 24716 45367
rect 25038 45364 25044 45416
rect 25096 45404 25102 45416
rect 25869 45407 25927 45413
rect 25869 45404 25881 45407
rect 25096 45376 25881 45404
rect 25096 45364 25102 45376
rect 25869 45373 25881 45376
rect 25915 45373 25927 45407
rect 25869 45367 25927 45373
rect 25976 45404 26004 45444
rect 26973 45407 27031 45413
rect 26973 45404 26985 45407
rect 25976 45376 26985 45404
rect 25130 45296 25136 45348
rect 25188 45336 25194 45348
rect 25409 45339 25467 45345
rect 25409 45336 25421 45339
rect 25188 45308 25421 45336
rect 25188 45296 25194 45308
rect 25409 45305 25421 45308
rect 25455 45336 25467 45339
rect 25593 45339 25651 45345
rect 25593 45336 25605 45339
rect 25455 45308 25605 45336
rect 25455 45305 25467 45308
rect 25409 45299 25467 45305
rect 25593 45305 25605 45308
rect 25639 45305 25651 45339
rect 25593 45299 25651 45305
rect 24670 45268 24676 45280
rect 23492 45240 24676 45268
rect 24670 45228 24676 45240
rect 24728 45228 24734 45280
rect 25038 45228 25044 45280
rect 25096 45268 25102 45280
rect 25222 45268 25228 45280
rect 25096 45240 25228 45268
rect 25096 45228 25102 45240
rect 25222 45228 25228 45240
rect 25280 45228 25286 45280
rect 25774 45268 25780 45280
rect 25735 45240 25780 45268
rect 25774 45228 25780 45240
rect 25832 45228 25838 45280
rect 25884 45268 25912 45367
rect 25976 45345 26004 45376
rect 26973 45373 26985 45376
rect 27019 45404 27031 45407
rect 27341 45407 27399 45413
rect 27341 45404 27353 45407
rect 27019 45376 27353 45404
rect 27019 45373 27031 45376
rect 26973 45367 27031 45373
rect 27341 45373 27353 45376
rect 27387 45373 27399 45407
rect 27341 45367 27399 45373
rect 25961 45339 26019 45345
rect 25961 45305 25973 45339
rect 26007 45305 26019 45339
rect 26326 45336 26332 45348
rect 26287 45308 26332 45336
rect 25961 45299 26019 45305
rect 26326 45296 26332 45308
rect 26384 45296 26390 45348
rect 26050 45268 26056 45280
rect 25884 45240 26056 45268
rect 26050 45228 26056 45240
rect 26108 45228 26114 45280
rect 26602 45268 26608 45280
rect 26563 45240 26608 45268
rect 26602 45228 26608 45240
rect 26660 45228 26666 45280
rect 1104 45178 28888 45200
rect 1104 45126 10982 45178
rect 11034 45126 11046 45178
rect 11098 45126 11110 45178
rect 11162 45126 11174 45178
rect 11226 45126 20982 45178
rect 21034 45126 21046 45178
rect 21098 45126 21110 45178
rect 21162 45126 21174 45178
rect 21226 45126 28888 45178
rect 1104 45104 28888 45126
rect 1673 45067 1731 45073
rect 1673 45033 1685 45067
rect 1719 45064 1731 45067
rect 1762 45064 1768 45076
rect 1719 45036 1768 45064
rect 1719 45033 1731 45036
rect 1673 45027 1731 45033
rect 1762 45024 1768 45036
rect 1820 45024 1826 45076
rect 1946 45064 1952 45076
rect 1907 45036 1952 45064
rect 1946 45024 1952 45036
rect 2004 45024 2010 45076
rect 12529 45067 12587 45073
rect 12529 45033 12541 45067
rect 12575 45064 12587 45067
rect 12618 45064 12624 45076
rect 12575 45036 12624 45064
rect 12575 45033 12587 45036
rect 12529 45027 12587 45033
rect 12618 45024 12624 45036
rect 12676 45024 12682 45076
rect 14550 45064 14556 45076
rect 14511 45036 14556 45064
rect 14550 45024 14556 45036
rect 14608 45024 14614 45076
rect 15565 45067 15623 45073
rect 15565 45033 15577 45067
rect 15611 45064 15623 45067
rect 15746 45064 15752 45076
rect 15611 45036 15752 45064
rect 15611 45033 15623 45036
rect 15565 45027 15623 45033
rect 15746 45024 15752 45036
rect 15804 45064 15810 45076
rect 16025 45067 16083 45073
rect 16025 45064 16037 45067
rect 15804 45036 16037 45064
rect 15804 45024 15810 45036
rect 16025 45033 16037 45036
rect 16071 45033 16083 45067
rect 16850 45064 16856 45076
rect 16811 45036 16856 45064
rect 16025 45027 16083 45033
rect 16850 45024 16856 45036
rect 16908 45024 16914 45076
rect 17034 45024 17040 45076
rect 17092 45064 17098 45076
rect 17221 45067 17279 45073
rect 17221 45064 17233 45067
rect 17092 45036 17233 45064
rect 17092 45024 17098 45036
rect 17221 45033 17233 45036
rect 17267 45033 17279 45067
rect 18138 45064 18144 45076
rect 18099 45036 18144 45064
rect 17221 45027 17279 45033
rect 18138 45024 18144 45036
rect 18196 45024 18202 45076
rect 18785 45067 18843 45073
rect 18785 45033 18797 45067
rect 18831 45064 18843 45067
rect 20346 45064 20352 45076
rect 18831 45036 20352 45064
rect 18831 45033 18843 45036
rect 18785 45027 18843 45033
rect 20346 45024 20352 45036
rect 20404 45024 20410 45076
rect 21542 45024 21548 45076
rect 21600 45064 21606 45076
rect 22002 45064 22008 45076
rect 21600 45036 22008 45064
rect 21600 45024 21606 45036
rect 22002 45024 22008 45036
rect 22060 45024 22066 45076
rect 23290 45064 23296 45076
rect 23251 45036 23296 45064
rect 23290 45024 23296 45036
rect 23348 45024 23354 45076
rect 23658 45064 23664 45076
rect 23619 45036 23664 45064
rect 23658 45024 23664 45036
rect 23716 45024 23722 45076
rect 24854 45064 24860 45076
rect 24815 45036 24860 45064
rect 24854 45024 24860 45036
rect 24912 45024 24918 45076
rect 25593 45067 25651 45073
rect 25593 45033 25605 45067
rect 25639 45064 25651 45067
rect 25774 45064 25780 45076
rect 25639 45036 25780 45064
rect 25639 45033 25651 45036
rect 25593 45027 25651 45033
rect 25774 45024 25780 45036
rect 25832 45064 25838 45076
rect 26694 45064 26700 45076
rect 25832 45036 26700 45064
rect 25832 45024 25838 45036
rect 26694 45024 26700 45036
rect 26752 45024 26758 45076
rect 13630 44996 13636 45008
rect 13591 44968 13636 44996
rect 13630 44956 13636 44968
rect 13688 44956 13694 45008
rect 19058 44956 19064 45008
rect 19116 44996 19122 45008
rect 19153 44999 19211 45005
rect 19153 44996 19165 44999
rect 19116 44968 19165 44996
rect 19116 44956 19122 44968
rect 19153 44965 19165 44968
rect 19199 44996 19211 44999
rect 19978 44996 19984 45008
rect 19199 44968 19984 44996
rect 19199 44965 19211 44968
rect 19153 44959 19211 44965
rect 19978 44956 19984 44968
rect 20036 44956 20042 45008
rect 21266 44956 21272 45008
rect 21324 44996 21330 45008
rect 21821 44999 21879 45005
rect 21821 44996 21833 44999
rect 21324 44968 21833 44996
rect 21324 44956 21330 44968
rect 21821 44965 21833 44968
rect 21867 44965 21879 44999
rect 23106 44996 23112 45008
rect 21821 44959 21879 44965
rect 22480 44968 23112 44996
rect 11790 44928 11796 44940
rect 11751 44900 11796 44928
rect 11790 44888 11796 44900
rect 11848 44888 11854 44940
rect 13446 44928 13452 44940
rect 13407 44900 13452 44928
rect 13446 44888 13452 44900
rect 13504 44888 13510 44940
rect 16666 44928 16672 44940
rect 16627 44900 16672 44928
rect 16666 44888 16672 44900
rect 16724 44888 16730 44940
rect 17678 44928 17684 44940
rect 17639 44900 17684 44928
rect 17678 44888 17684 44900
rect 17736 44888 17742 44940
rect 17957 44931 18015 44937
rect 17957 44897 17969 44931
rect 18003 44928 18015 44931
rect 18046 44928 18052 44940
rect 18003 44900 18052 44928
rect 18003 44897 18015 44900
rect 17957 44891 18015 44897
rect 18046 44888 18052 44900
rect 18104 44888 18110 44940
rect 18598 44888 18604 44940
rect 18656 44928 18662 44940
rect 19245 44931 19303 44937
rect 19245 44928 19257 44931
rect 18656 44900 19257 44928
rect 18656 44888 18662 44900
rect 19245 44897 19257 44900
rect 19291 44928 19303 44931
rect 19426 44928 19432 44940
rect 19291 44900 19432 44928
rect 19291 44897 19303 44900
rect 19245 44891 19303 44897
rect 19426 44888 19432 44900
rect 19484 44888 19490 44940
rect 21542 44888 21548 44940
rect 21600 44928 21606 44940
rect 22186 44928 22192 44940
rect 21600 44900 22192 44928
rect 21600 44888 21606 44900
rect 22186 44888 22192 44900
rect 22244 44888 22250 44940
rect 22480 44937 22508 44968
rect 23106 44956 23112 44968
rect 23164 44956 23170 45008
rect 25225 44999 25283 45005
rect 25225 44996 25237 44999
rect 23400 44968 25237 44996
rect 22465 44931 22523 44937
rect 22465 44897 22477 44931
rect 22511 44897 22523 44931
rect 22465 44891 22523 44897
rect 22554 44888 22560 44940
rect 22612 44928 22618 44940
rect 22833 44931 22891 44937
rect 22833 44928 22845 44931
rect 22612 44900 22845 44928
rect 22612 44888 22618 44900
rect 22833 44897 22845 44900
rect 22879 44928 22891 44931
rect 23400 44928 23428 44968
rect 25225 44965 25237 44968
rect 25271 44996 25283 44999
rect 26237 44999 26295 45005
rect 26237 44996 26249 44999
rect 25271 44968 26249 44996
rect 25271 44965 25283 44968
rect 25225 44959 25283 44965
rect 26237 44965 26249 44968
rect 26283 44965 26295 44999
rect 26237 44959 26295 44965
rect 26602 44956 26608 45008
rect 26660 44996 26666 45008
rect 26881 44999 26939 45005
rect 26881 44996 26893 44999
rect 26660 44968 26893 44996
rect 26660 44956 26666 44968
rect 26881 44965 26893 44968
rect 26927 44965 26939 44999
rect 26881 44959 26939 44965
rect 22879 44900 23428 44928
rect 22879 44897 22891 44900
rect 22833 44891 22891 44897
rect 23566 44888 23572 44940
rect 23624 44928 23630 44940
rect 23937 44931 23995 44937
rect 23937 44928 23949 44931
rect 23624 44900 23949 44928
rect 23624 44888 23630 44900
rect 23937 44897 23949 44900
rect 23983 44897 23995 44931
rect 25406 44928 25412 44940
rect 25367 44900 25412 44928
rect 23937 44891 23995 44897
rect 25406 44888 25412 44900
rect 25464 44888 25470 44940
rect 25961 44931 26019 44937
rect 25961 44897 25973 44931
rect 26007 44928 26019 44931
rect 26050 44928 26056 44940
rect 26007 44900 26056 44928
rect 26007 44897 26019 44900
rect 25961 44891 26019 44897
rect 26050 44888 26056 44900
rect 26108 44928 26114 44940
rect 26786 44928 26792 44940
rect 26108 44900 26792 44928
rect 26108 44888 26114 44900
rect 26786 44888 26792 44900
rect 26844 44888 26850 44940
rect 11885 44863 11943 44869
rect 11885 44829 11897 44863
rect 11931 44860 11943 44863
rect 11974 44860 11980 44872
rect 11931 44832 11980 44860
rect 11931 44829 11943 44832
rect 11885 44823 11943 44829
rect 11974 44820 11980 44832
rect 12032 44820 12038 44872
rect 18322 44820 18328 44872
rect 18380 44860 18386 44872
rect 19613 44863 19671 44869
rect 19613 44860 19625 44863
rect 18380 44832 19625 44860
rect 18380 44820 18386 44832
rect 19613 44829 19625 44832
rect 19659 44829 19671 44863
rect 19613 44823 19671 44829
rect 19702 44820 19708 44872
rect 19760 44860 19766 44872
rect 19760 44832 19805 44860
rect 19760 44820 19766 44832
rect 20346 44820 20352 44872
rect 20404 44860 20410 44872
rect 20625 44863 20683 44869
rect 20625 44860 20637 44863
rect 20404 44832 20637 44860
rect 20404 44820 20410 44832
rect 20625 44829 20637 44832
rect 20671 44860 20683 44863
rect 20898 44860 20904 44872
rect 20671 44832 20904 44860
rect 20671 44829 20683 44832
rect 20625 44823 20683 44829
rect 20898 44820 20904 44832
rect 20956 44820 20962 44872
rect 21174 44860 21180 44872
rect 21135 44832 21180 44860
rect 21174 44820 21180 44832
rect 21232 44820 21238 44872
rect 22094 44820 22100 44872
rect 22152 44860 22158 44872
rect 22373 44863 22431 44869
rect 22373 44860 22385 44863
rect 22152 44832 22385 44860
rect 22152 44820 22158 44832
rect 22373 44829 22385 44832
rect 22419 44829 22431 44863
rect 22373 44823 22431 44829
rect 22925 44863 22983 44869
rect 22925 44829 22937 44863
rect 22971 44829 22983 44863
rect 22925 44823 22983 44829
rect 16577 44795 16635 44801
rect 16577 44761 16589 44795
rect 16623 44792 16635 44795
rect 17770 44792 17776 44804
rect 16623 44764 17776 44792
rect 16623 44761 16635 44764
rect 16577 44755 16635 44761
rect 17770 44752 17776 44764
rect 17828 44752 17834 44804
rect 19521 44795 19579 44801
rect 19521 44761 19533 44795
rect 19567 44792 19579 44795
rect 19794 44792 19800 44804
rect 19567 44764 19800 44792
rect 19567 44761 19579 44764
rect 19521 44755 19579 44761
rect 19794 44752 19800 44764
rect 19852 44792 19858 44804
rect 20714 44792 20720 44804
rect 19852 44764 20720 44792
rect 19852 44752 19858 44764
rect 20714 44752 20720 44764
rect 20772 44752 20778 44804
rect 22462 44752 22468 44804
rect 22520 44792 22526 44804
rect 22940 44792 22968 44823
rect 23658 44820 23664 44872
rect 23716 44860 23722 44872
rect 23845 44863 23903 44869
rect 23845 44860 23857 44863
rect 23716 44832 23857 44860
rect 23716 44820 23722 44832
rect 23845 44829 23857 44832
rect 23891 44829 23903 44863
rect 23845 44823 23903 44829
rect 25130 44820 25136 44872
rect 25188 44860 25194 44872
rect 26510 44860 26516 44872
rect 25188 44832 26516 44860
rect 25188 44820 25194 44832
rect 26510 44820 26516 44832
rect 26568 44820 26574 44872
rect 27062 44820 27068 44872
rect 27120 44860 27126 44872
rect 27249 44863 27307 44869
rect 27249 44860 27261 44863
rect 27120 44832 27261 44860
rect 27120 44820 27126 44832
rect 27249 44829 27261 44832
rect 27295 44829 27307 44863
rect 27249 44823 27307 44829
rect 22520 44764 22968 44792
rect 22520 44752 22526 44764
rect 1578 44684 1584 44736
rect 1636 44724 1642 44736
rect 2317 44727 2375 44733
rect 2317 44724 2329 44727
rect 1636 44696 2329 44724
rect 1636 44684 1642 44696
rect 2317 44693 2329 44696
rect 2363 44693 2375 44727
rect 2317 44687 2375 44693
rect 19150 44684 19156 44736
rect 19208 44724 19214 44736
rect 19383 44727 19441 44733
rect 19383 44724 19395 44727
rect 19208 44696 19395 44724
rect 19208 44684 19214 44696
rect 19383 44693 19395 44696
rect 19429 44693 19441 44727
rect 19383 44687 19441 44693
rect 19978 44684 19984 44736
rect 20036 44724 20042 44736
rect 20257 44727 20315 44733
rect 20257 44724 20269 44727
rect 20036 44696 20269 44724
rect 20036 44684 20042 44696
rect 20257 44693 20269 44696
rect 20303 44693 20315 44727
rect 20257 44687 20315 44693
rect 21729 44727 21787 44733
rect 21729 44693 21741 44727
rect 21775 44724 21787 44727
rect 22278 44724 22284 44736
rect 21775 44696 22284 44724
rect 21775 44693 21787 44696
rect 21729 44687 21787 44693
rect 22278 44684 22284 44696
rect 22336 44684 22342 44736
rect 26878 44684 26884 44736
rect 26936 44724 26942 44736
rect 27525 44727 27583 44733
rect 27525 44724 27537 44727
rect 26936 44696 27537 44724
rect 26936 44684 26942 44696
rect 27525 44693 27537 44696
rect 27571 44693 27583 44727
rect 27525 44687 27583 44693
rect 1104 44634 28888 44656
rect 1104 44582 5982 44634
rect 6034 44582 6046 44634
rect 6098 44582 6110 44634
rect 6162 44582 6174 44634
rect 6226 44582 15982 44634
rect 16034 44582 16046 44634
rect 16098 44582 16110 44634
rect 16162 44582 16174 44634
rect 16226 44582 25982 44634
rect 26034 44582 26046 44634
rect 26098 44582 26110 44634
rect 26162 44582 26174 44634
rect 26226 44582 28888 44634
rect 1104 44560 28888 44582
rect 2958 44520 2964 44532
rect 2919 44492 2964 44520
rect 2958 44480 2964 44492
rect 3016 44480 3022 44532
rect 11790 44480 11796 44532
rect 11848 44520 11854 44532
rect 14185 44523 14243 44529
rect 14185 44520 14197 44523
rect 11848 44492 14197 44520
rect 11848 44480 11854 44492
rect 14185 44489 14197 44492
rect 14231 44489 14243 44523
rect 14185 44483 14243 44489
rect 15562 44480 15568 44532
rect 15620 44520 15626 44532
rect 15749 44523 15807 44529
rect 15749 44520 15761 44523
rect 15620 44492 15761 44520
rect 15620 44480 15626 44492
rect 15749 44489 15761 44492
rect 15795 44489 15807 44523
rect 15749 44483 15807 44489
rect 19705 44523 19763 44529
rect 19705 44489 19717 44523
rect 19751 44520 19763 44523
rect 19794 44520 19800 44532
rect 19751 44492 19800 44520
rect 19751 44489 19763 44492
rect 19705 44483 19763 44489
rect 12253 44455 12311 44461
rect 12253 44421 12265 44455
rect 12299 44452 12311 44455
rect 12618 44452 12624 44464
rect 12299 44424 12624 44452
rect 12299 44421 12311 44424
rect 12253 44415 12311 44421
rect 12618 44412 12624 44424
rect 12676 44452 12682 44464
rect 12713 44455 12771 44461
rect 12713 44452 12725 44455
rect 12676 44424 12725 44452
rect 12676 44412 12682 44424
rect 12713 44421 12725 44424
rect 12759 44421 12771 44455
rect 12713 44415 12771 44421
rect 1397 44387 1455 44393
rect 1397 44353 1409 44387
rect 1443 44384 1455 44387
rect 1578 44384 1584 44396
rect 1443 44356 1584 44384
rect 1443 44353 1455 44356
rect 1397 44347 1455 44353
rect 1578 44344 1584 44356
rect 1636 44344 1642 44396
rect 12805 44387 12863 44393
rect 12805 44353 12817 44387
rect 12851 44384 12863 44387
rect 12851 44356 13584 44384
rect 12851 44353 12863 44356
rect 12805 44347 12863 44353
rect 1673 44319 1731 44325
rect 1673 44285 1685 44319
rect 1719 44316 1731 44319
rect 1946 44316 1952 44328
rect 1719 44288 1952 44316
rect 1719 44285 1731 44288
rect 1673 44279 1731 44285
rect 1946 44276 1952 44288
rect 2004 44276 2010 44328
rect 10229 44319 10287 44325
rect 10229 44285 10241 44319
rect 10275 44316 10287 44319
rect 10965 44319 11023 44325
rect 10965 44316 10977 44319
rect 10275 44288 10977 44316
rect 10275 44285 10287 44288
rect 10229 44279 10287 44285
rect 10965 44285 10977 44288
rect 11011 44316 11023 44319
rect 11514 44316 11520 44328
rect 11011 44288 11520 44316
rect 11011 44285 11023 44288
rect 10965 44279 11023 44285
rect 11514 44276 11520 44288
rect 11572 44276 11578 44328
rect 12618 44325 12624 44328
rect 12584 44319 12624 44325
rect 12584 44285 12596 44319
rect 12584 44279 12624 44285
rect 12618 44276 12624 44279
rect 12676 44276 12682 44328
rect 11885 44251 11943 44257
rect 11885 44217 11897 44251
rect 11931 44248 11943 44251
rect 12437 44251 12495 44257
rect 12437 44248 12449 44251
rect 11931 44220 12449 44248
rect 11931 44217 11943 44220
rect 11885 44211 11943 44217
rect 12437 44217 12449 44220
rect 12483 44248 12495 44251
rect 12483 44220 13492 44248
rect 12483 44217 12495 44220
rect 12437 44211 12495 44217
rect 13464 44192 13492 44220
rect 10778 44180 10784 44192
rect 10739 44152 10784 44180
rect 10778 44140 10784 44152
rect 10836 44140 10842 44192
rect 11425 44183 11483 44189
rect 11425 44149 11437 44183
rect 11471 44180 11483 44183
rect 11790 44180 11796 44192
rect 11471 44152 11796 44180
rect 11471 44149 11483 44152
rect 11425 44143 11483 44149
rect 11790 44140 11796 44152
rect 11848 44140 11854 44192
rect 13078 44180 13084 44192
rect 13039 44152 13084 44180
rect 13078 44140 13084 44152
rect 13136 44140 13142 44192
rect 13446 44180 13452 44192
rect 13407 44152 13452 44180
rect 13446 44140 13452 44152
rect 13504 44140 13510 44192
rect 13556 44180 13584 44356
rect 13814 44276 13820 44328
rect 13872 44316 13878 44328
rect 14001 44319 14059 44325
rect 14001 44316 14013 44319
rect 13872 44288 14013 44316
rect 13872 44276 13878 44288
rect 14001 44285 14013 44288
rect 14047 44316 14059 44319
rect 14461 44319 14519 44325
rect 14461 44316 14473 44319
rect 14047 44288 14473 44316
rect 14047 44285 14059 44288
rect 14001 44279 14059 44285
rect 14461 44285 14473 44288
rect 14507 44285 14519 44319
rect 15764 44316 15792 44483
rect 19794 44480 19800 44492
rect 19852 44480 19858 44532
rect 20898 44520 20904 44532
rect 20180 44492 20904 44520
rect 17129 44455 17187 44461
rect 17129 44421 17141 44455
rect 17175 44452 17187 44455
rect 17954 44452 17960 44464
rect 17175 44424 17960 44452
rect 17175 44421 17187 44424
rect 17129 44415 17187 44421
rect 17954 44412 17960 44424
rect 18012 44412 18018 44464
rect 16666 44344 16672 44396
rect 16724 44384 16730 44396
rect 16761 44387 16819 44393
rect 16761 44384 16773 44387
rect 16724 44356 16773 44384
rect 16724 44344 16730 44356
rect 16761 44353 16773 44356
rect 16807 44384 16819 44387
rect 17494 44384 17500 44396
rect 16807 44356 17500 44384
rect 16807 44353 16819 44356
rect 16761 44347 16819 44353
rect 17494 44344 17500 44356
rect 17552 44344 17558 44396
rect 18322 44344 18328 44396
rect 18380 44384 18386 44396
rect 20180 44393 20208 44492
rect 20898 44480 20904 44492
rect 20956 44480 20962 44532
rect 21637 44523 21695 44529
rect 21637 44489 21649 44523
rect 21683 44520 21695 44523
rect 22462 44520 22468 44532
rect 21683 44492 22468 44520
rect 21683 44489 21695 44492
rect 21637 44483 21695 44489
rect 22462 44480 22468 44492
rect 22520 44480 22526 44532
rect 23106 44520 23112 44532
rect 23067 44492 23112 44520
rect 23106 44480 23112 44492
rect 23164 44480 23170 44532
rect 25130 44480 25136 44532
rect 25188 44520 25194 44532
rect 25593 44523 25651 44529
rect 25593 44520 25605 44523
rect 25188 44492 25605 44520
rect 25188 44480 25194 44492
rect 25593 44489 25605 44492
rect 25639 44489 25651 44523
rect 25593 44483 25651 44489
rect 20346 44452 20352 44464
rect 20272 44424 20352 44452
rect 18601 44387 18659 44393
rect 18601 44384 18613 44387
rect 18380 44356 18613 44384
rect 18380 44344 18386 44356
rect 18601 44353 18613 44356
rect 18647 44384 18659 44387
rect 19981 44387 20039 44393
rect 19981 44384 19993 44387
rect 18647 44356 19993 44384
rect 18647 44353 18659 44356
rect 18601 44347 18659 44353
rect 19981 44353 19993 44356
rect 20027 44353 20039 44387
rect 19981 44347 20039 44353
rect 20165 44387 20223 44393
rect 20165 44353 20177 44387
rect 20211 44353 20223 44387
rect 20165 44347 20223 44353
rect 15933 44319 15991 44325
rect 15933 44316 15945 44319
rect 15764 44288 15945 44316
rect 14461 44279 14519 44285
rect 15933 44285 15945 44288
rect 15979 44316 15991 44319
rect 16482 44316 16488 44328
rect 15979 44288 16488 44316
rect 15979 44285 15991 44288
rect 15933 44279 15991 44285
rect 16482 44276 16488 44288
rect 16540 44276 16546 44328
rect 16574 44276 16580 44328
rect 16632 44316 16638 44328
rect 16945 44319 17003 44325
rect 16945 44316 16957 44319
rect 16632 44288 16957 44316
rect 16632 44276 16638 44288
rect 16945 44285 16957 44288
rect 16991 44316 17003 44319
rect 18506 44316 18512 44328
rect 16991 44288 17540 44316
rect 18419 44288 18512 44316
rect 16991 44285 17003 44288
rect 16945 44279 17003 44285
rect 13909 44183 13967 44189
rect 13909 44180 13921 44183
rect 13556 44152 13921 44180
rect 13909 44149 13921 44152
rect 13955 44180 13967 44183
rect 13998 44180 14004 44192
rect 13955 44152 14004 44180
rect 13955 44149 13967 44152
rect 13909 44143 13967 44149
rect 13998 44140 14004 44152
rect 14056 44140 14062 44192
rect 16114 44180 16120 44192
rect 16075 44152 16120 44180
rect 16114 44140 16120 44152
rect 16172 44140 16178 44192
rect 16666 44140 16672 44192
rect 16724 44180 16730 44192
rect 16942 44180 16948 44192
rect 16724 44152 16948 44180
rect 16724 44140 16730 44152
rect 16942 44140 16948 44152
rect 17000 44140 17006 44192
rect 17512 44189 17540 44288
rect 18506 44276 18512 44288
rect 18564 44316 18570 44328
rect 19245 44319 19303 44325
rect 19245 44316 19257 44319
rect 18564 44288 19257 44316
rect 18564 44276 18570 44288
rect 19245 44285 19257 44288
rect 19291 44316 19303 44319
rect 19334 44316 19340 44328
rect 19291 44288 19340 44316
rect 19291 44285 19303 44288
rect 19245 44279 19303 44285
rect 19334 44276 19340 44288
rect 19392 44276 19398 44328
rect 20272 44248 20300 44424
rect 20346 44412 20352 44424
rect 20404 44412 20410 44464
rect 20438 44412 20444 44464
rect 20496 44412 20502 44464
rect 24670 44412 24676 44464
rect 24728 44412 24734 44464
rect 24762 44412 24768 44464
rect 24820 44452 24826 44464
rect 25038 44452 25044 44464
rect 24820 44424 25044 44452
rect 24820 44412 24826 44424
rect 25038 44412 25044 44424
rect 25096 44412 25102 44464
rect 20456 44384 20484 44412
rect 21174 44384 21180 44396
rect 20364 44356 21180 44384
rect 20364 44325 20392 44356
rect 21174 44344 21180 44356
rect 21232 44344 21238 44396
rect 24026 44344 24032 44396
rect 24084 44384 24090 44396
rect 24210 44384 24216 44396
rect 24084 44356 24216 44384
rect 24084 44344 24090 44356
rect 24210 44344 24216 44356
rect 24268 44344 24274 44396
rect 24688 44384 24716 44412
rect 24854 44384 24860 44396
rect 24688 44356 24860 44384
rect 24854 44344 24860 44356
rect 24912 44384 24918 44396
rect 25225 44387 25283 44393
rect 25225 44384 25237 44387
rect 24912 44356 25237 44384
rect 24912 44344 24918 44356
rect 25225 44353 25237 44356
rect 25271 44353 25283 44387
rect 25225 44347 25283 44353
rect 26053 44387 26111 44393
rect 26053 44353 26065 44387
rect 26099 44384 26111 44387
rect 26418 44384 26424 44396
rect 26099 44356 26424 44384
rect 26099 44353 26111 44356
rect 26053 44347 26111 44353
rect 26418 44344 26424 44356
rect 26476 44344 26482 44396
rect 26602 44384 26608 44396
rect 26515 44356 26608 44384
rect 20349 44319 20407 44325
rect 20349 44285 20361 44319
rect 20395 44285 20407 44319
rect 20349 44279 20407 44285
rect 20438 44276 20444 44328
rect 20496 44316 20502 44328
rect 20901 44319 20959 44325
rect 20901 44316 20913 44319
rect 20496 44288 20913 44316
rect 20496 44276 20502 44288
rect 20901 44285 20913 44288
rect 20947 44285 20959 44319
rect 20901 44279 20959 44285
rect 21269 44319 21327 44325
rect 21269 44285 21281 44319
rect 21315 44316 21327 44319
rect 22094 44316 22100 44328
rect 21315 44288 22100 44316
rect 21315 44285 21327 44288
rect 21269 44279 21327 44285
rect 22094 44276 22100 44288
rect 22152 44316 22158 44328
rect 22189 44319 22247 44325
rect 22189 44316 22201 44319
rect 22152 44288 22201 44316
rect 22152 44276 22158 44288
rect 22189 44285 22201 44288
rect 22235 44285 22247 44319
rect 22189 44279 22247 44285
rect 22278 44276 22284 44328
rect 22336 44316 22342 44328
rect 22373 44319 22431 44325
rect 22373 44316 22385 44319
rect 22336 44288 22385 44316
rect 22336 44276 22342 44288
rect 22373 44285 22385 44288
rect 22419 44285 22431 44319
rect 22554 44316 22560 44328
rect 22515 44288 22560 44316
rect 22373 44279 22431 44285
rect 22554 44276 22560 44288
rect 22612 44276 22618 44328
rect 22646 44276 22652 44328
rect 22704 44316 22710 44328
rect 23842 44316 23848 44328
rect 22704 44288 23848 44316
rect 22704 44276 22710 44288
rect 23842 44276 23848 44288
rect 23900 44316 23906 44328
rect 23937 44319 23995 44325
rect 23937 44316 23949 44319
rect 23900 44288 23949 44316
rect 23900 44276 23906 44288
rect 23937 44285 23949 44288
rect 23983 44285 23995 44319
rect 23937 44279 23995 44285
rect 24670 44276 24676 44328
rect 24728 44316 24734 44328
rect 24765 44319 24823 44325
rect 24765 44316 24777 44319
rect 24728 44288 24777 44316
rect 24728 44276 24734 44288
rect 24765 44285 24777 44288
rect 24811 44285 24823 44319
rect 24765 44279 24823 44285
rect 26145 44319 26203 44325
rect 26145 44285 26157 44319
rect 26191 44316 26203 44319
rect 26528 44316 26556 44356
rect 26602 44344 26608 44356
rect 26660 44384 26666 44396
rect 26878 44384 26884 44396
rect 26660 44356 26884 44384
rect 26660 44344 26666 44356
rect 26878 44344 26884 44356
rect 26936 44344 26942 44396
rect 26191 44288 26556 44316
rect 26191 44285 26203 44288
rect 26145 44279 26203 44285
rect 26694 44276 26700 44328
rect 26752 44316 26758 44328
rect 28077 44319 28135 44325
rect 28077 44316 28089 44319
rect 26752 44288 28089 44316
rect 26752 44276 26758 44288
rect 28077 44285 28089 44288
rect 28123 44285 28135 44319
rect 28077 44279 28135 44285
rect 20533 44251 20591 44257
rect 20533 44248 20545 44251
rect 20272 44220 20545 44248
rect 20533 44217 20545 44220
rect 20579 44217 20591 44251
rect 20533 44211 20591 44217
rect 21729 44251 21787 44257
rect 21729 44217 21741 44251
rect 21775 44248 21787 44251
rect 21818 44248 21824 44260
rect 21775 44220 21824 44248
rect 21775 44217 21787 44220
rect 21729 44211 21787 44217
rect 21818 44208 21824 44220
rect 21876 44208 21882 44260
rect 24029 44251 24087 44257
rect 24029 44217 24041 44251
rect 24075 44248 24087 44251
rect 25130 44248 25136 44260
rect 24075 44220 25136 44248
rect 24075 44217 24087 44220
rect 24029 44211 24087 44217
rect 25130 44208 25136 44220
rect 25188 44208 25194 44260
rect 17497 44183 17555 44189
rect 17497 44149 17509 44183
rect 17543 44180 17555 44183
rect 17678 44180 17684 44192
rect 17543 44152 17684 44180
rect 17543 44149 17555 44152
rect 17497 44143 17555 44149
rect 17678 44140 17684 44152
rect 17736 44180 17742 44192
rect 17773 44183 17831 44189
rect 17773 44180 17785 44183
rect 17736 44152 17785 44180
rect 17736 44140 17742 44152
rect 17773 44149 17785 44152
rect 17819 44149 17831 44183
rect 17773 44143 17831 44149
rect 20070 44140 20076 44192
rect 20128 44180 20134 44192
rect 20441 44183 20499 44189
rect 20441 44180 20453 44183
rect 20128 44152 20453 44180
rect 20128 44140 20134 44152
rect 20441 44149 20453 44152
rect 20487 44149 20499 44183
rect 20441 44143 20499 44149
rect 22462 44140 22468 44192
rect 22520 44180 22526 44192
rect 22646 44180 22652 44192
rect 22520 44152 22652 44180
rect 22520 44140 22526 44152
rect 22646 44140 22652 44152
rect 22704 44140 22710 44192
rect 23477 44183 23535 44189
rect 23477 44149 23489 44183
rect 23523 44180 23535 44183
rect 23566 44180 23572 44192
rect 23523 44152 23572 44180
rect 23523 44149 23535 44152
rect 23477 44143 23535 44149
rect 23566 44140 23572 44152
rect 23624 44140 23630 44192
rect 27706 44180 27712 44192
rect 27667 44152 27712 44180
rect 27706 44140 27712 44152
rect 27764 44140 27770 44192
rect 1104 44090 28888 44112
rect 1104 44038 10982 44090
rect 11034 44038 11046 44090
rect 11098 44038 11110 44090
rect 11162 44038 11174 44090
rect 11226 44038 20982 44090
rect 21034 44038 21046 44090
rect 21098 44038 21110 44090
rect 21162 44038 21174 44090
rect 21226 44038 28888 44090
rect 1104 44016 28888 44038
rect 16482 43936 16488 43988
rect 16540 43976 16546 43988
rect 17129 43979 17187 43985
rect 17129 43976 17141 43979
rect 16540 43948 17141 43976
rect 16540 43936 16546 43948
rect 17129 43945 17141 43948
rect 17175 43976 17187 43979
rect 17494 43976 17500 43988
rect 17175 43948 17500 43976
rect 17175 43945 17187 43948
rect 17129 43939 17187 43945
rect 17494 43936 17500 43948
rect 17552 43976 17558 43988
rect 17552 43948 17908 43976
rect 17552 43936 17558 43948
rect 12250 43908 12256 43920
rect 11808 43880 12256 43908
rect 1489 43843 1547 43849
rect 1489 43809 1501 43843
rect 1535 43840 1547 43843
rect 1578 43840 1584 43852
rect 1535 43812 1584 43840
rect 1535 43809 1547 43812
rect 1489 43803 1547 43809
rect 1578 43800 1584 43812
rect 1636 43800 1642 43852
rect 7558 43800 7564 43852
rect 7616 43840 7622 43852
rect 7837 43843 7895 43849
rect 7837 43840 7849 43843
rect 7616 43812 7849 43840
rect 7616 43800 7622 43812
rect 7837 43809 7849 43812
rect 7883 43809 7895 43843
rect 8570 43840 8576 43852
rect 8531 43812 8576 43840
rect 7837 43803 7895 43809
rect 8570 43800 8576 43812
rect 8628 43800 8634 43852
rect 8665 43843 8723 43849
rect 8665 43809 8677 43843
rect 8711 43840 8723 43843
rect 8754 43840 8760 43852
rect 8711 43812 8760 43840
rect 8711 43809 8723 43812
rect 8665 43803 8723 43809
rect 8754 43800 8760 43812
rect 8812 43800 8818 43852
rect 11606 43800 11612 43852
rect 11664 43840 11670 43852
rect 11808 43849 11836 43880
rect 12250 43868 12256 43880
rect 12308 43868 12314 43920
rect 16853 43911 16911 43917
rect 16853 43877 16865 43911
rect 16899 43908 16911 43911
rect 17586 43908 17592 43920
rect 16899 43880 17592 43908
rect 16899 43877 16911 43880
rect 16853 43871 16911 43877
rect 17586 43868 17592 43880
rect 17644 43868 17650 43920
rect 17880 43908 17908 43948
rect 17954 43936 17960 43988
rect 18012 43976 18018 43988
rect 19061 43979 19119 43985
rect 19061 43976 19073 43979
rect 18012 43948 19073 43976
rect 18012 43936 18018 43948
rect 19061 43945 19073 43948
rect 19107 43976 19119 43979
rect 19150 43976 19156 43988
rect 19107 43948 19156 43976
rect 19107 43945 19119 43948
rect 19061 43939 19119 43945
rect 19150 43936 19156 43948
rect 19208 43936 19214 43988
rect 19705 43979 19763 43985
rect 19705 43945 19717 43979
rect 19751 43976 19763 43979
rect 19886 43976 19892 43988
rect 19751 43948 19892 43976
rect 19751 43945 19763 43948
rect 19705 43939 19763 43945
rect 19886 43936 19892 43948
rect 19944 43936 19950 43988
rect 21269 43979 21327 43985
rect 21269 43945 21281 43979
rect 21315 43945 21327 43979
rect 23842 43976 23848 43988
rect 23803 43948 23848 43976
rect 21269 43939 21327 43945
rect 18046 43908 18052 43920
rect 17880 43880 18052 43908
rect 11793 43843 11851 43849
rect 11793 43840 11805 43843
rect 11664 43812 11805 43840
rect 11664 43800 11670 43812
rect 11793 43809 11805 43812
rect 11839 43809 11851 43843
rect 12066 43840 12072 43852
rect 12027 43812 12072 43840
rect 11793 43803 11851 43809
rect 12066 43800 12072 43812
rect 12124 43800 12130 43852
rect 13078 43840 13084 43852
rect 13039 43812 13084 43840
rect 13078 43800 13084 43812
rect 13136 43800 13142 43852
rect 16298 43840 16304 43852
rect 16259 43812 16304 43840
rect 16298 43800 16304 43812
rect 16356 43800 16362 43852
rect 16393 43843 16451 43849
rect 16393 43809 16405 43843
rect 16439 43840 16451 43843
rect 16482 43840 16488 43852
rect 16439 43812 16488 43840
rect 16439 43809 16451 43812
rect 16393 43803 16451 43809
rect 16482 43800 16488 43812
rect 16540 43800 16546 43852
rect 17678 43840 17684 43852
rect 17639 43812 17684 43840
rect 17678 43800 17684 43812
rect 17736 43800 17742 43852
rect 17770 43800 17776 43852
rect 17828 43840 17834 43852
rect 17972 43849 18000 43880
rect 18046 43868 18052 43880
rect 18104 43868 18110 43920
rect 18690 43868 18696 43920
rect 18748 43908 18754 43920
rect 21284 43908 21312 43939
rect 23842 43936 23848 43948
rect 23900 43936 23906 43988
rect 25406 43936 25412 43988
rect 25464 43976 25470 43988
rect 25869 43979 25927 43985
rect 25869 43976 25881 43979
rect 25464 43948 25881 43976
rect 25464 43936 25470 43948
rect 25869 43945 25881 43948
rect 25915 43945 25927 43979
rect 26694 43976 26700 43988
rect 26655 43948 26700 43976
rect 25869 43939 25927 43945
rect 26694 43936 26700 43948
rect 26752 43936 26758 43988
rect 26786 43936 26792 43988
rect 26844 43976 26850 43988
rect 26844 43948 26889 43976
rect 26844 43936 26850 43948
rect 21634 43908 21640 43920
rect 18748 43880 21640 43908
rect 18748 43868 18754 43880
rect 21634 43868 21640 43880
rect 21692 43868 21698 43920
rect 23474 43908 23480 43920
rect 22572 43880 23480 43908
rect 17957 43843 18015 43849
rect 17828 43812 17873 43840
rect 17828 43800 17834 43812
rect 17957 43809 17969 43843
rect 18003 43809 18015 43843
rect 19886 43840 19892 43852
rect 19847 43812 19892 43840
rect 17957 43803 18015 43809
rect 19886 43800 19892 43812
rect 19944 43800 19950 43852
rect 21082 43840 21088 43852
rect 21043 43812 21088 43840
rect 21082 43800 21088 43812
rect 21140 43800 21146 43852
rect 22572 43849 22600 43880
rect 23474 43868 23480 43880
rect 23532 43868 23538 43920
rect 26510 43908 26516 43920
rect 26471 43880 26516 43908
rect 26510 43868 26516 43880
rect 26568 43868 26574 43920
rect 26878 43908 26884 43920
rect 26839 43880 26884 43908
rect 26878 43868 26884 43880
rect 26936 43868 26942 43920
rect 22557 43843 22615 43849
rect 22557 43809 22569 43843
rect 22603 43809 22615 43843
rect 22738 43840 22744 43852
rect 22699 43812 22744 43840
rect 22557 43803 22615 43809
rect 22738 43800 22744 43812
rect 22796 43800 22802 43852
rect 22925 43843 22983 43849
rect 22925 43809 22937 43843
rect 22971 43840 22983 43843
rect 23106 43840 23112 43852
rect 22971 43812 23112 43840
rect 22971 43809 22983 43812
rect 22925 43803 22983 43809
rect 23106 43800 23112 43812
rect 23164 43800 23170 43852
rect 26329 43843 26387 43849
rect 26329 43809 26341 43843
rect 26375 43840 26387 43843
rect 26786 43840 26792 43852
rect 26375 43812 26792 43840
rect 26375 43809 26387 43812
rect 26329 43803 26387 43809
rect 26786 43800 26792 43812
rect 26844 43800 26850 43852
rect 1765 43775 1823 43781
rect 1765 43741 1777 43775
rect 1811 43772 1823 43775
rect 2222 43772 2228 43784
rect 1811 43744 2228 43772
rect 1811 43741 1823 43744
rect 1765 43735 1823 43741
rect 2222 43732 2228 43744
rect 2280 43732 2286 43784
rect 3142 43772 3148 43784
rect 3103 43744 3148 43772
rect 3142 43732 3148 43744
rect 3200 43732 3206 43784
rect 7742 43772 7748 43784
rect 7703 43744 7748 43772
rect 7742 43732 7748 43744
rect 7800 43732 7806 43784
rect 11241 43775 11299 43781
rect 11241 43741 11253 43775
rect 11287 43772 11299 43775
rect 11330 43772 11336 43784
rect 11287 43744 11336 43772
rect 11287 43741 11299 43744
rect 11241 43735 11299 43741
rect 11330 43732 11336 43744
rect 11388 43732 11394 43784
rect 12253 43775 12311 43781
rect 12253 43741 12265 43775
rect 12299 43741 12311 43775
rect 12618 43772 12624 43784
rect 12531 43744 12624 43772
rect 12253 43735 12311 43741
rect 10594 43664 10600 43716
rect 10652 43704 10658 43716
rect 12268 43704 12296 43735
rect 12618 43732 12624 43744
rect 12676 43772 12682 43784
rect 13170 43772 13176 43784
rect 12676 43744 13176 43772
rect 12676 43732 12682 43744
rect 13170 43732 13176 43744
rect 13228 43732 13234 43784
rect 18414 43772 18420 43784
rect 18375 43744 18420 43772
rect 18414 43732 18420 43744
rect 18472 43732 18478 43784
rect 22186 43732 22192 43784
rect 22244 43772 22250 43784
rect 23842 43772 23848 43784
rect 22244 43744 23848 43772
rect 22244 43732 22250 43744
rect 23842 43732 23848 43744
rect 23900 43772 23906 43784
rect 23937 43775 23995 43781
rect 23937 43772 23949 43775
rect 23900 43744 23949 43772
rect 23900 43732 23906 43744
rect 23937 43741 23949 43744
rect 23983 43741 23995 43775
rect 23937 43735 23995 43741
rect 24118 43732 24124 43784
rect 24176 43772 24182 43784
rect 24213 43775 24271 43781
rect 24213 43772 24225 43775
rect 24176 43744 24225 43772
rect 24176 43732 24182 43744
rect 24213 43741 24225 43744
rect 24259 43741 24271 43775
rect 24213 43735 24271 43741
rect 25593 43775 25651 43781
rect 25593 43741 25605 43775
rect 25639 43772 25651 43775
rect 25866 43772 25872 43784
rect 25639 43744 25872 43772
rect 25639 43741 25651 43744
rect 25593 43735 25651 43741
rect 25866 43732 25872 43744
rect 25924 43732 25930 43784
rect 27246 43772 27252 43784
rect 27207 43744 27252 43772
rect 27246 43732 27252 43744
rect 27304 43732 27310 43784
rect 10652 43676 12296 43704
rect 12989 43707 13047 43713
rect 10652 43664 10658 43676
rect 12989 43673 13001 43707
rect 13035 43704 13047 43707
rect 13354 43704 13360 43716
rect 13035 43676 13360 43704
rect 13035 43673 13047 43676
rect 12989 43667 13047 43673
rect 13354 43664 13360 43676
rect 13412 43664 13418 43716
rect 15746 43664 15752 43716
rect 15804 43704 15810 43716
rect 16114 43704 16120 43716
rect 15804 43676 16120 43704
rect 15804 43664 15810 43676
rect 16114 43664 16120 43676
rect 16172 43664 16178 43716
rect 22370 43704 22376 43716
rect 22331 43676 22376 43704
rect 22370 43664 22376 43676
rect 22428 43664 22434 43716
rect 13262 43636 13268 43648
rect 13223 43608 13268 43636
rect 13262 43596 13268 43608
rect 13320 43596 13326 43648
rect 17589 43639 17647 43645
rect 17589 43605 17601 43639
rect 17635 43636 17647 43639
rect 18598 43636 18604 43648
rect 17635 43608 18604 43636
rect 17635 43605 17647 43608
rect 17589 43599 17647 43605
rect 18598 43596 18604 43608
rect 18656 43636 18662 43648
rect 18693 43639 18751 43645
rect 18693 43636 18705 43639
rect 18656 43608 18705 43636
rect 18656 43596 18662 43608
rect 18693 43605 18705 43608
rect 18739 43605 18751 43639
rect 18693 43599 18751 43605
rect 19978 43596 19984 43648
rect 20036 43636 20042 43648
rect 20533 43639 20591 43645
rect 20533 43636 20545 43639
rect 20036 43608 20545 43636
rect 20036 43596 20042 43608
rect 20533 43605 20545 43608
rect 20579 43605 20591 43639
rect 20533 43599 20591 43605
rect 21821 43639 21879 43645
rect 21821 43605 21833 43639
rect 21867 43636 21879 43639
rect 22094 43636 22100 43648
rect 21867 43608 22100 43636
rect 21867 43605 21879 43608
rect 21821 43599 21879 43605
rect 22094 43596 22100 43608
rect 22152 43636 22158 43648
rect 22462 43636 22468 43648
rect 22152 43608 22468 43636
rect 22152 43596 22158 43608
rect 22462 43596 22468 43608
rect 22520 43596 22526 43648
rect 23477 43639 23535 43645
rect 23477 43605 23489 43639
rect 23523 43636 23535 43639
rect 24670 43636 24676 43648
rect 23523 43608 24676 43636
rect 23523 43605 23535 43608
rect 23477 43599 23535 43605
rect 24670 43596 24676 43608
rect 24728 43596 24734 43648
rect 27522 43636 27528 43648
rect 27483 43608 27528 43636
rect 27522 43596 27528 43608
rect 27580 43596 27586 43648
rect 1104 43546 28888 43568
rect 1104 43494 5982 43546
rect 6034 43494 6046 43546
rect 6098 43494 6110 43546
rect 6162 43494 6174 43546
rect 6226 43494 15982 43546
rect 16034 43494 16046 43546
rect 16098 43494 16110 43546
rect 16162 43494 16174 43546
rect 16226 43494 25982 43546
rect 26034 43494 26046 43546
rect 26098 43494 26110 43546
rect 26162 43494 26174 43546
rect 26226 43494 28888 43546
rect 1104 43472 28888 43494
rect 7742 43432 7748 43444
rect 7703 43404 7748 43432
rect 7742 43392 7748 43404
rect 7800 43392 7806 43444
rect 8481 43435 8539 43441
rect 8481 43401 8493 43435
rect 8527 43432 8539 43435
rect 8570 43432 8576 43444
rect 8527 43404 8576 43432
rect 8527 43401 8539 43404
rect 8481 43395 8539 43401
rect 8570 43392 8576 43404
rect 8628 43392 8634 43444
rect 11333 43435 11391 43441
rect 11333 43401 11345 43435
rect 11379 43432 11391 43435
rect 11514 43432 11520 43444
rect 11379 43404 11520 43432
rect 11379 43401 11391 43404
rect 11333 43395 11391 43401
rect 8113 43367 8171 43373
rect 8113 43333 8125 43367
rect 8159 43364 8171 43367
rect 8754 43364 8760 43376
rect 8159 43336 8760 43364
rect 8159 43333 8171 43336
rect 8113 43327 8171 43333
rect 8754 43324 8760 43336
rect 8812 43324 8818 43376
rect 9674 43324 9680 43376
rect 9732 43364 9738 43376
rect 10965 43367 11023 43373
rect 10965 43364 10977 43367
rect 9732 43336 10977 43364
rect 9732 43324 9738 43336
rect 10965 43333 10977 43336
rect 11011 43333 11023 43367
rect 10965 43327 11023 43333
rect 1762 43296 1768 43308
rect 1723 43268 1768 43296
rect 1762 43256 1768 43268
rect 1820 43256 1826 43308
rect 1489 43231 1547 43237
rect 1489 43197 1501 43231
rect 1535 43228 1547 43231
rect 1578 43228 1584 43240
rect 1535 43200 1584 43228
rect 1535 43197 1547 43200
rect 1489 43191 1547 43197
rect 1578 43188 1584 43200
rect 1636 43188 1642 43240
rect 3142 43228 3148 43240
rect 3103 43200 3148 43228
rect 3142 43188 3148 43200
rect 3200 43188 3206 43240
rect 10781 43231 10839 43237
rect 10781 43197 10793 43231
rect 10827 43228 10839 43231
rect 11348 43228 11376 43395
rect 11514 43392 11520 43404
rect 11572 43392 11578 43444
rect 12805 43435 12863 43441
rect 12805 43401 12817 43435
rect 12851 43432 12863 43435
rect 13078 43432 13084 43444
rect 12851 43404 13084 43432
rect 12851 43401 12863 43404
rect 12805 43395 12863 43401
rect 13078 43392 13084 43404
rect 13136 43392 13142 43444
rect 15746 43392 15752 43444
rect 15804 43432 15810 43444
rect 16117 43435 16175 43441
rect 16117 43432 16129 43435
rect 15804 43404 16129 43432
rect 15804 43392 15810 43404
rect 16117 43401 16129 43404
rect 16163 43401 16175 43435
rect 16117 43395 16175 43401
rect 16298 43392 16304 43444
rect 16356 43432 16362 43444
rect 16577 43435 16635 43441
rect 16577 43432 16589 43435
rect 16356 43404 16589 43432
rect 16356 43392 16362 43404
rect 16577 43401 16589 43404
rect 16623 43432 16635 43435
rect 17129 43435 17187 43441
rect 17129 43432 17141 43435
rect 16623 43404 17141 43432
rect 16623 43401 16635 43404
rect 16577 43395 16635 43401
rect 17129 43401 17141 43404
rect 17175 43432 17187 43435
rect 17402 43432 17408 43444
rect 17175 43404 17408 43432
rect 17175 43401 17187 43404
rect 17129 43395 17187 43401
rect 17402 43392 17408 43404
rect 17460 43392 17466 43444
rect 17678 43432 17684 43444
rect 17639 43404 17684 43432
rect 17678 43392 17684 43404
rect 17736 43392 17742 43444
rect 19426 43432 19432 43444
rect 19387 43404 19432 43432
rect 19426 43392 19432 43404
rect 19484 43392 19490 43444
rect 21082 43392 21088 43444
rect 21140 43432 21146 43444
rect 21821 43435 21879 43441
rect 21821 43432 21833 43435
rect 21140 43404 21833 43432
rect 21140 43392 21146 43404
rect 21821 43401 21833 43404
rect 21867 43432 21879 43435
rect 22465 43435 22523 43441
rect 22465 43432 22477 43435
rect 21867 43404 22477 43432
rect 21867 43401 21879 43404
rect 21821 43395 21879 43401
rect 22465 43401 22477 43404
rect 22511 43401 22523 43435
rect 22465 43395 22523 43401
rect 22741 43435 22799 43441
rect 22741 43401 22753 43435
rect 22787 43432 22799 43435
rect 22922 43432 22928 43444
rect 22787 43404 22928 43432
rect 22787 43401 22799 43404
rect 22741 43395 22799 43401
rect 22922 43392 22928 43404
rect 22980 43392 22986 43444
rect 23109 43435 23167 43441
rect 23109 43401 23121 43435
rect 23155 43432 23167 43435
rect 23658 43432 23664 43444
rect 23155 43404 23664 43432
rect 23155 43401 23167 43404
rect 23109 43395 23167 43401
rect 15841 43367 15899 43373
rect 15841 43333 15853 43367
rect 15887 43364 15899 43367
rect 16482 43364 16488 43376
rect 15887 43336 16488 43364
rect 15887 43333 15899 43336
rect 15841 43327 15899 43333
rect 16482 43324 16488 43336
rect 16540 43324 16546 43376
rect 19150 43324 19156 43376
rect 19208 43364 19214 43376
rect 20070 43364 20076 43376
rect 19208 43336 20076 43364
rect 19208 43324 19214 43336
rect 20070 43324 20076 43336
rect 20128 43324 20134 43376
rect 13814 43296 13820 43308
rect 13775 43268 13820 43296
rect 13814 43256 13820 43268
rect 13872 43256 13878 43308
rect 17678 43256 17684 43308
rect 17736 43296 17742 43308
rect 18046 43296 18052 43308
rect 17736 43268 18052 43296
rect 17736 43256 17742 43268
rect 18046 43256 18052 43268
rect 18104 43256 18110 43308
rect 20714 43256 20720 43308
rect 20772 43296 20778 43308
rect 21266 43296 21272 43308
rect 20772 43268 21272 43296
rect 20772 43256 20778 43268
rect 21266 43256 21272 43268
rect 21324 43296 21330 43308
rect 22281 43299 22339 43305
rect 21324 43268 21404 43296
rect 21324 43256 21330 43268
rect 10827 43200 11376 43228
rect 11701 43231 11759 43237
rect 10827 43197 10839 43200
rect 10781 43191 10839 43197
rect 11701 43197 11713 43231
rect 11747 43228 11759 43231
rect 12066 43228 12072 43240
rect 11747 43200 12072 43228
rect 11747 43197 11759 43200
rect 11701 43191 11759 43197
rect 12066 43188 12072 43200
rect 12124 43228 12130 43240
rect 12161 43231 12219 43237
rect 12161 43228 12173 43231
rect 12124 43200 12173 43228
rect 12124 43188 12130 43200
rect 12161 43197 12173 43200
rect 12207 43197 12219 43231
rect 12986 43228 12992 43240
rect 12947 43200 12992 43228
rect 12161 43191 12219 43197
rect 12176 43160 12204 43191
rect 12986 43188 12992 43200
rect 13044 43188 13050 43240
rect 13354 43228 13360 43240
rect 13315 43200 13360 43228
rect 13354 43188 13360 43200
rect 13412 43188 13418 43240
rect 13722 43228 13728 43240
rect 13683 43200 13728 43228
rect 13722 43188 13728 43200
rect 13780 43188 13786 43240
rect 16945 43231 17003 43237
rect 16945 43197 16957 43231
rect 16991 43228 17003 43231
rect 17034 43228 17040 43240
rect 16991 43200 17040 43228
rect 16991 43197 17003 43200
rect 16945 43191 17003 43197
rect 17034 43188 17040 43200
rect 17092 43228 17098 43240
rect 17770 43228 17776 43240
rect 17092 43200 17776 43228
rect 17092 43188 17098 43200
rect 17770 43188 17776 43200
rect 17828 43188 17834 43240
rect 18325 43231 18383 43237
rect 18325 43197 18337 43231
rect 18371 43228 18383 43231
rect 18966 43228 18972 43240
rect 18371 43200 18972 43228
rect 18371 43197 18383 43200
rect 18325 43191 18383 43197
rect 18966 43188 18972 43200
rect 19024 43188 19030 43240
rect 19978 43188 19984 43240
rect 20036 43228 20042 43240
rect 21376 43237 21404 43268
rect 22281 43265 22293 43299
rect 22327 43296 22339 43299
rect 22738 43296 22744 43308
rect 22327 43268 22744 43296
rect 22327 43265 22339 43268
rect 22281 43259 22339 43265
rect 22738 43256 22744 43268
rect 22796 43256 22802 43308
rect 21085 43231 21143 43237
rect 21085 43228 21097 43231
rect 20036 43200 21097 43228
rect 20036 43188 20042 43200
rect 21085 43197 21097 43200
rect 21131 43197 21143 43231
rect 21085 43191 21143 43197
rect 21361 43231 21419 43237
rect 21361 43197 21373 43231
rect 21407 43197 21419 43231
rect 21361 43191 21419 43197
rect 21545 43231 21603 43237
rect 21545 43197 21557 43231
rect 21591 43197 21603 43231
rect 21545 43191 21603 43197
rect 22557 43231 22615 43237
rect 22557 43197 22569 43231
rect 22603 43228 22615 43231
rect 23124 43228 23152 43395
rect 23658 43392 23664 43404
rect 23716 43392 23722 43444
rect 24029 43435 24087 43441
rect 24029 43401 24041 43435
rect 24075 43432 24087 43435
rect 24118 43432 24124 43444
rect 24075 43404 24124 43432
rect 24075 43401 24087 43404
rect 24029 43395 24087 43401
rect 24118 43392 24124 43404
rect 24176 43392 24182 43444
rect 25774 43392 25780 43444
rect 25832 43432 25838 43444
rect 25961 43435 26019 43441
rect 25961 43432 25973 43435
rect 25832 43404 25973 43432
rect 25832 43392 25838 43404
rect 25961 43401 25973 43404
rect 26007 43401 26019 43435
rect 26510 43432 26516 43444
rect 26471 43404 26516 43432
rect 25961 43395 26019 43401
rect 26510 43392 26516 43404
rect 26568 43392 26574 43444
rect 26694 43392 26700 43444
rect 26752 43432 26758 43444
rect 26973 43435 27031 43441
rect 26973 43432 26985 43435
rect 26752 43404 26985 43432
rect 26752 43392 26758 43404
rect 26973 43401 26985 43404
rect 27019 43401 27031 43435
rect 27338 43432 27344 43444
rect 27299 43404 27344 43432
rect 26973 43395 27031 43401
rect 27338 43392 27344 43404
rect 27396 43392 27402 43444
rect 23474 43364 23480 43376
rect 23435 43336 23480 43364
rect 23474 43324 23480 43336
rect 23532 43324 23538 43376
rect 26878 43324 26884 43376
rect 26936 43364 26942 43376
rect 28261 43367 28319 43373
rect 28261 43364 28273 43367
rect 26936 43336 28273 43364
rect 26936 43324 26942 43336
rect 28261 43333 28273 43336
rect 28307 43333 28319 43367
rect 28261 43327 28319 43333
rect 24489 43299 24547 43305
rect 24489 43265 24501 43299
rect 24535 43296 24547 43299
rect 27065 43299 27123 43305
rect 24535 43268 24900 43296
rect 24535 43265 24547 43268
rect 24489 43259 24547 43265
rect 24872 43240 24900 43268
rect 27065 43265 27077 43299
rect 27111 43296 27123 43299
rect 27522 43296 27528 43308
rect 27111 43268 27528 43296
rect 27111 43265 27123 43268
rect 27065 43259 27123 43265
rect 27522 43256 27528 43268
rect 27580 43256 27586 43308
rect 22603 43200 23152 43228
rect 22603 43197 22615 43200
rect 22557 43191 22615 43197
rect 13740 43160 13768 43188
rect 12176 43132 13768 43160
rect 19426 43120 19432 43172
rect 19484 43160 19490 43172
rect 20349 43163 20407 43169
rect 20349 43160 20361 43163
rect 19484 43132 20361 43160
rect 19484 43120 19490 43132
rect 20349 43129 20361 43132
rect 20395 43129 20407 43163
rect 20349 43123 20407 43129
rect 20533 43163 20591 43169
rect 20533 43129 20545 43163
rect 20579 43160 20591 43163
rect 20714 43160 20720 43172
rect 20579 43132 20720 43160
rect 20579 43129 20591 43132
rect 20533 43123 20591 43129
rect 10594 43092 10600 43104
rect 10555 43064 10600 43092
rect 10594 43052 10600 43064
rect 10652 43052 10658 43104
rect 20364 43092 20392 43123
rect 20714 43120 20720 43132
rect 20772 43120 20778 43172
rect 21560 43092 21588 43191
rect 23842 43188 23848 43240
rect 23900 43228 23906 43240
rect 24581 43231 24639 43237
rect 24581 43228 24593 43231
rect 23900 43200 24593 43228
rect 23900 43188 23906 43200
rect 24581 43197 24593 43200
rect 24627 43197 24639 43231
rect 24854 43228 24860 43240
rect 24815 43200 24860 43228
rect 24581 43191 24639 43197
rect 24854 43188 24860 43200
rect 24912 43188 24918 43240
rect 26326 43228 26332 43240
rect 25516 43200 26332 43228
rect 20364 43064 21588 43092
rect 22465 43095 22523 43101
rect 22465 43061 22477 43095
rect 22511 43092 22523 43095
rect 25516 43092 25544 43200
rect 26326 43188 26332 43200
rect 26384 43228 26390 43240
rect 27157 43231 27215 43237
rect 27157 43228 27169 43231
rect 26384 43200 27169 43228
rect 26384 43188 26390 43200
rect 27157 43197 27169 43200
rect 27203 43228 27215 43231
rect 27893 43231 27951 43237
rect 27893 43228 27905 43231
rect 27203 43200 27905 43228
rect 27203 43197 27215 43200
rect 27157 43191 27215 43197
rect 27893 43197 27905 43200
rect 27939 43197 27951 43231
rect 27893 43191 27951 43197
rect 22511 43064 25544 43092
rect 22511 43061 22523 43064
rect 22465 43055 22523 43061
rect 1104 43002 28888 43024
rect 1104 42950 10982 43002
rect 11034 42950 11046 43002
rect 11098 42950 11110 43002
rect 11162 42950 11174 43002
rect 11226 42950 20982 43002
rect 21034 42950 21046 43002
rect 21098 42950 21110 43002
rect 21162 42950 21174 43002
rect 21226 42950 28888 43002
rect 1104 42928 28888 42950
rect 1673 42891 1731 42897
rect 1673 42857 1685 42891
rect 1719 42888 1731 42891
rect 1762 42888 1768 42900
rect 1719 42860 1768 42888
rect 1719 42857 1731 42860
rect 1673 42851 1731 42857
rect 1762 42848 1768 42860
rect 1820 42848 1826 42900
rect 11330 42848 11336 42900
rect 11388 42888 11394 42900
rect 17034 42888 17040 42900
rect 11388 42860 12388 42888
rect 16995 42860 17040 42888
rect 11388 42848 11394 42860
rect 1578 42780 1584 42832
rect 1636 42820 1642 42832
rect 2317 42823 2375 42829
rect 2317 42820 2329 42823
rect 1636 42792 2329 42820
rect 1636 42780 1642 42792
rect 2317 42789 2329 42792
rect 2363 42789 2375 42823
rect 11425 42823 11483 42829
rect 11425 42820 11437 42823
rect 2317 42783 2375 42789
rect 10980 42792 11437 42820
rect 10226 42712 10232 42764
rect 10284 42752 10290 42764
rect 10980 42752 11008 42792
rect 11425 42789 11437 42792
rect 11471 42789 11483 42823
rect 11425 42783 11483 42789
rect 10284 42724 11008 42752
rect 11333 42755 11391 42761
rect 10284 42712 10290 42724
rect 11333 42721 11345 42755
rect 11379 42752 11391 42755
rect 11606 42752 11612 42764
rect 11379 42724 11612 42752
rect 11379 42721 11391 42724
rect 11333 42715 11391 42721
rect 11606 42712 11612 42724
rect 11664 42712 11670 42764
rect 12066 42752 12072 42764
rect 12027 42724 12072 42752
rect 12066 42712 12072 42724
rect 12124 42712 12130 42764
rect 11974 42684 11980 42696
rect 11935 42656 11980 42684
rect 11974 42644 11980 42656
rect 12032 42644 12038 42696
rect 12360 42684 12388 42860
rect 17034 42848 17040 42860
rect 17092 42848 17098 42900
rect 17494 42888 17500 42900
rect 17455 42860 17500 42888
rect 17494 42848 17500 42860
rect 17552 42848 17558 42900
rect 20625 42891 20683 42897
rect 20625 42857 20637 42891
rect 20671 42888 20683 42891
rect 21266 42888 21272 42900
rect 20671 42860 21272 42888
rect 20671 42857 20683 42860
rect 20625 42851 20683 42857
rect 21266 42848 21272 42860
rect 21324 42848 21330 42900
rect 26786 42848 26792 42900
rect 26844 42888 26850 42900
rect 27341 42891 27399 42897
rect 27341 42888 27353 42891
rect 26844 42860 27353 42888
rect 26844 42848 26850 42860
rect 27341 42857 27353 42860
rect 27387 42857 27399 42891
rect 27341 42851 27399 42857
rect 13814 42820 13820 42832
rect 13740 42792 13820 42820
rect 12434 42712 12440 42764
rect 12492 42752 12498 42764
rect 13740 42752 13768 42792
rect 13814 42780 13820 42792
rect 13872 42780 13878 42832
rect 21637 42823 21695 42829
rect 21637 42789 21649 42823
rect 21683 42820 21695 42823
rect 21726 42820 21732 42832
rect 21683 42792 21732 42820
rect 21683 42789 21695 42792
rect 21637 42783 21695 42789
rect 21726 42780 21732 42792
rect 21784 42780 21790 42832
rect 22922 42780 22928 42832
rect 22980 42820 22986 42832
rect 23106 42820 23112 42832
rect 22980 42792 23112 42820
rect 22980 42780 22986 42792
rect 23106 42780 23112 42792
rect 23164 42780 23170 42832
rect 12492 42724 13768 42752
rect 17589 42755 17647 42761
rect 12492 42712 12498 42724
rect 17589 42721 17601 42755
rect 17635 42752 17647 42755
rect 17678 42752 17684 42764
rect 17635 42724 17684 42752
rect 17635 42721 17647 42724
rect 17589 42715 17647 42721
rect 17678 42712 17684 42724
rect 17736 42712 17742 42764
rect 19150 42712 19156 42764
rect 19208 42752 19214 42764
rect 19702 42752 19708 42764
rect 19208 42724 19708 42752
rect 19208 42712 19214 42724
rect 19702 42712 19708 42724
rect 19760 42712 19766 42764
rect 19797 42755 19855 42761
rect 19797 42721 19809 42755
rect 19843 42752 19855 42755
rect 20070 42752 20076 42764
rect 19843 42724 20076 42752
rect 19843 42721 19855 42724
rect 19797 42715 19855 42721
rect 20070 42712 20076 42724
rect 20128 42752 20134 42764
rect 20438 42752 20444 42764
rect 20128 42724 20444 42752
rect 20128 42712 20134 42724
rect 20438 42712 20444 42724
rect 20496 42712 20502 42764
rect 21545 42755 21603 42761
rect 21545 42721 21557 42755
rect 21591 42752 21603 42755
rect 22278 42752 22284 42764
rect 21591 42724 22284 42752
rect 21591 42721 21603 42724
rect 21545 42715 21603 42721
rect 22278 42712 22284 42724
rect 22336 42712 22342 42764
rect 22646 42752 22652 42764
rect 22607 42724 22652 42752
rect 22646 42712 22652 42724
rect 22704 42712 22710 42764
rect 22738 42712 22744 42764
rect 22796 42752 22802 42764
rect 22796 42724 22841 42752
rect 22796 42712 22802 42724
rect 23842 42712 23848 42764
rect 23900 42752 23906 42764
rect 23937 42755 23995 42761
rect 23937 42752 23949 42755
rect 23900 42724 23949 42752
rect 23900 42712 23906 42724
rect 23937 42721 23949 42724
rect 23983 42721 23995 42755
rect 23937 42715 23995 42721
rect 24213 42755 24271 42761
rect 24213 42721 24225 42755
rect 24259 42752 24271 42755
rect 24578 42752 24584 42764
rect 24259 42724 24584 42752
rect 24259 42721 24271 42724
rect 24213 42715 24271 42721
rect 12529 42687 12587 42693
rect 12529 42684 12541 42687
rect 12360 42656 12541 42684
rect 12529 42653 12541 42656
rect 12575 42653 12587 42687
rect 12529 42647 12587 42653
rect 17865 42687 17923 42693
rect 17865 42653 17877 42687
rect 17911 42684 17923 42687
rect 18322 42684 18328 42696
rect 17911 42656 18328 42684
rect 17911 42653 17923 42656
rect 17865 42647 17923 42653
rect 18322 42644 18328 42656
rect 18380 42644 18386 42696
rect 21177 42687 21235 42693
rect 21177 42653 21189 42687
rect 21223 42684 21235 42687
rect 22186 42684 22192 42696
rect 21223 42656 22192 42684
rect 21223 42653 21235 42656
rect 21177 42647 21235 42653
rect 22186 42644 22192 42656
rect 22244 42644 22250 42696
rect 22373 42687 22431 42693
rect 22373 42653 22385 42687
rect 22419 42684 22431 42687
rect 22462 42684 22468 42696
rect 22419 42656 22468 42684
rect 22419 42653 22431 42656
rect 22373 42647 22431 42653
rect 22462 42644 22468 42656
rect 22520 42644 22526 42696
rect 23952 42684 23980 42715
rect 24578 42712 24584 42724
rect 24636 42712 24642 42764
rect 25590 42712 25596 42764
rect 25648 42752 25654 42764
rect 26513 42755 26571 42761
rect 26513 42752 26525 42755
rect 25648 42724 26525 42752
rect 25648 42712 25654 42724
rect 26513 42721 26525 42724
rect 26559 42721 26571 42755
rect 26513 42715 26571 42721
rect 26602 42712 26608 42764
rect 26660 42752 26666 42764
rect 26660 42724 26705 42752
rect 26660 42712 26666 42724
rect 25774 42684 25780 42696
rect 23952 42656 25780 42684
rect 25774 42644 25780 42656
rect 25832 42684 25838 42696
rect 25869 42687 25927 42693
rect 25869 42684 25881 42687
rect 25832 42656 25881 42684
rect 25832 42644 25838 42656
rect 25869 42653 25881 42656
rect 25915 42684 25927 42687
rect 26237 42687 26295 42693
rect 26237 42684 26249 42687
rect 25915 42656 26249 42684
rect 25915 42653 25927 42656
rect 25869 42647 25927 42653
rect 26237 42653 26249 42656
rect 26283 42653 26295 42687
rect 26237 42647 26295 42653
rect 19886 42576 19892 42628
rect 19944 42616 19950 42628
rect 20165 42619 20223 42625
rect 20165 42616 20177 42619
rect 19944 42588 20177 42616
rect 19944 42576 19950 42588
rect 20165 42585 20177 42588
rect 20211 42616 20223 42619
rect 20438 42616 20444 42628
rect 20211 42588 20444 42616
rect 20211 42585 20223 42588
rect 20165 42579 20223 42585
rect 20438 42576 20444 42588
rect 20496 42576 20502 42628
rect 2041 42551 2099 42557
rect 2041 42517 2053 42551
rect 2087 42548 2099 42551
rect 2222 42548 2228 42560
rect 2087 42520 2228 42548
rect 2087 42517 2099 42520
rect 2041 42511 2099 42517
rect 2222 42508 2228 42520
rect 2280 42508 2286 42560
rect 8665 42551 8723 42557
rect 8665 42517 8677 42551
rect 8711 42548 8723 42551
rect 10226 42548 10232 42560
rect 8711 42520 10232 42548
rect 8711 42517 8723 42520
rect 8665 42511 8723 42517
rect 10226 42508 10232 42520
rect 10284 42508 10290 42560
rect 12986 42548 12992 42560
rect 12947 42520 12992 42548
rect 12986 42508 12992 42520
rect 13044 42508 13050 42560
rect 18966 42548 18972 42560
rect 18927 42520 18972 42548
rect 18966 42508 18972 42520
rect 19024 42508 19030 42560
rect 22278 42508 22284 42560
rect 22336 42548 22342 42560
rect 22554 42548 22560 42560
rect 22336 42520 22560 42548
rect 22336 42508 22342 42520
rect 22554 42508 22560 42520
rect 22612 42548 22618 42560
rect 23109 42551 23167 42557
rect 23109 42548 23121 42551
rect 22612 42520 23121 42548
rect 22612 42508 22618 42520
rect 23109 42517 23121 42520
rect 23155 42517 23167 42551
rect 23109 42511 23167 42517
rect 23566 42508 23572 42560
rect 23624 42548 23630 42560
rect 23753 42551 23811 42557
rect 23753 42548 23765 42551
rect 23624 42520 23765 42548
rect 23624 42508 23630 42520
rect 23753 42517 23765 42520
rect 23799 42548 23811 42551
rect 24302 42548 24308 42560
rect 23799 42520 24308 42548
rect 23799 42517 23811 42520
rect 23753 42511 23811 42517
rect 24302 42508 24308 42520
rect 24360 42508 24366 42560
rect 25130 42508 25136 42560
rect 25188 42548 25194 42560
rect 25317 42551 25375 42557
rect 25317 42548 25329 42551
rect 25188 42520 25329 42548
rect 25188 42508 25194 42520
rect 25317 42517 25329 42520
rect 25363 42517 25375 42551
rect 26786 42548 26792 42560
rect 26747 42520 26792 42548
rect 25317 42511 25375 42517
rect 26786 42508 26792 42520
rect 26844 42508 26850 42560
rect 1104 42458 28888 42480
rect 1104 42406 5982 42458
rect 6034 42406 6046 42458
rect 6098 42406 6110 42458
rect 6162 42406 6174 42458
rect 6226 42406 15982 42458
rect 16034 42406 16046 42458
rect 16098 42406 16110 42458
rect 16162 42406 16174 42458
rect 16226 42406 25982 42458
rect 26034 42406 26046 42458
rect 26098 42406 26110 42458
rect 26162 42406 26174 42458
rect 26226 42406 28888 42458
rect 1104 42384 28888 42406
rect 1578 42344 1584 42356
rect 1539 42316 1584 42344
rect 1578 42304 1584 42316
rect 1636 42304 1642 42356
rect 10873 42347 10931 42353
rect 10873 42313 10885 42347
rect 10919 42344 10931 42347
rect 11330 42344 11336 42356
rect 10919 42316 11336 42344
rect 10919 42313 10931 42316
rect 10873 42307 10931 42313
rect 11330 42304 11336 42316
rect 11388 42304 11394 42356
rect 11885 42347 11943 42353
rect 11885 42313 11897 42347
rect 11931 42344 11943 42347
rect 11974 42344 11980 42356
rect 11931 42316 11980 42344
rect 11931 42313 11943 42316
rect 11885 42307 11943 42313
rect 8481 42211 8539 42217
rect 8481 42177 8493 42211
rect 8527 42208 8539 42211
rect 8527 42180 9628 42208
rect 8527 42177 8539 42180
rect 8481 42171 8539 42177
rect 9600 42152 9628 42180
rect 8757 42143 8815 42149
rect 8757 42109 8769 42143
rect 8803 42109 8815 42143
rect 8938 42140 8944 42152
rect 8899 42112 8944 42140
rect 8757 42103 8815 42109
rect 8772 42072 8800 42103
rect 8938 42100 8944 42112
rect 8996 42100 9002 42152
rect 9214 42140 9220 42152
rect 9175 42112 9220 42140
rect 9214 42100 9220 42112
rect 9272 42100 9278 42152
rect 9582 42140 9588 42152
rect 9543 42112 9588 42140
rect 9582 42100 9588 42112
rect 9640 42100 9646 42152
rect 10042 42140 10048 42152
rect 10003 42112 10048 42140
rect 10042 42100 10048 42112
rect 10100 42100 10106 42152
rect 10226 42140 10232 42152
rect 10187 42112 10232 42140
rect 10226 42100 10232 42112
rect 10284 42100 10290 42152
rect 11333 42143 11391 42149
rect 11333 42109 11345 42143
rect 11379 42140 11391 42143
rect 11900 42140 11928 42307
rect 11974 42304 11980 42316
rect 12032 42344 12038 42356
rect 12161 42347 12219 42353
rect 12161 42344 12173 42347
rect 12032 42316 12173 42344
rect 12032 42304 12038 42316
rect 12161 42313 12173 42316
rect 12207 42313 12219 42347
rect 12161 42307 12219 42313
rect 12986 42304 12992 42356
rect 13044 42344 13050 42356
rect 14461 42347 14519 42353
rect 14461 42344 14473 42347
rect 13044 42316 14473 42344
rect 13044 42304 13050 42316
rect 14461 42313 14473 42316
rect 14507 42313 14519 42347
rect 17770 42344 17776 42356
rect 17731 42316 17776 42344
rect 14461 42307 14519 42313
rect 17770 42304 17776 42316
rect 17828 42304 17834 42356
rect 18322 42344 18328 42356
rect 18235 42316 18328 42344
rect 18322 42304 18328 42316
rect 18380 42344 18386 42356
rect 19702 42344 19708 42356
rect 18380 42316 19708 42344
rect 18380 42304 18386 42316
rect 19702 42304 19708 42316
rect 19760 42304 19766 42356
rect 20714 42304 20720 42356
rect 20772 42344 20778 42356
rect 20993 42347 21051 42353
rect 20993 42344 21005 42347
rect 20772 42316 21005 42344
rect 20772 42304 20778 42316
rect 20993 42313 21005 42316
rect 21039 42313 21051 42347
rect 20993 42307 21051 42313
rect 17405 42279 17463 42285
rect 17405 42245 17417 42279
rect 17451 42276 17463 42279
rect 17678 42276 17684 42288
rect 17451 42248 17684 42276
rect 17451 42245 17463 42248
rect 17405 42239 17463 42245
rect 17678 42236 17684 42248
rect 17736 42236 17742 42288
rect 18874 42276 18880 42288
rect 18835 42248 18880 42276
rect 18874 42236 18880 42248
rect 18932 42236 18938 42288
rect 19613 42279 19671 42285
rect 19613 42245 19625 42279
rect 19659 42276 19671 42279
rect 19886 42276 19892 42288
rect 19659 42248 19892 42276
rect 19659 42245 19671 42248
rect 19613 42239 19671 42245
rect 19886 42236 19892 42248
rect 19944 42236 19950 42288
rect 19981 42279 20039 42285
rect 19981 42245 19993 42279
rect 20027 42276 20039 42279
rect 20438 42276 20444 42288
rect 20027 42248 20444 42276
rect 20027 42245 20039 42248
rect 19981 42239 20039 42245
rect 20438 42236 20444 42248
rect 20496 42236 20502 42288
rect 14185 42211 14243 42217
rect 14185 42177 14197 42211
rect 14231 42208 14243 42211
rect 19904 42208 19932 42236
rect 21008 42208 21036 42307
rect 21266 42304 21272 42356
rect 21324 42344 21330 42356
rect 21634 42344 21640 42356
rect 21324 42316 21640 42344
rect 21324 42304 21330 42316
rect 21634 42304 21640 42316
rect 21692 42304 21698 42356
rect 25041 42347 25099 42353
rect 25041 42313 25053 42347
rect 25087 42344 25099 42347
rect 26786 42344 26792 42356
rect 25087 42316 26792 42344
rect 25087 42313 25099 42316
rect 25041 42307 25099 42313
rect 22186 42236 22192 42288
rect 22244 42276 22250 42288
rect 23014 42276 23020 42288
rect 22244 42248 23020 42276
rect 22244 42236 22250 42248
rect 23014 42236 23020 42248
rect 23072 42236 23078 42288
rect 23937 42279 23995 42285
rect 23937 42245 23949 42279
rect 23983 42276 23995 42279
rect 24762 42276 24768 42288
rect 23983 42248 24768 42276
rect 23983 42245 23995 42248
rect 23937 42239 23995 42245
rect 24762 42236 24768 42248
rect 24820 42236 24826 42288
rect 21634 42208 21640 42220
rect 14231 42180 15148 42208
rect 19904 42180 20944 42208
rect 21008 42180 21640 42208
rect 14231 42177 14243 42180
rect 14185 42171 14243 42177
rect 11379 42112 11928 42140
rect 14277 42143 14335 42149
rect 11379 42109 11391 42112
rect 11333 42103 11391 42109
rect 14277 42109 14289 42143
rect 14323 42109 14335 42143
rect 14277 42103 14335 42109
rect 9030 42072 9036 42084
rect 8772 42044 9036 42072
rect 9030 42032 9036 42044
rect 9088 42032 9094 42084
rect 8113 42007 8171 42013
rect 8113 41973 8125 42007
rect 8159 42004 8171 42007
rect 9232 42004 9260 42100
rect 11241 42075 11299 42081
rect 11241 42041 11253 42075
rect 11287 42072 11299 42075
rect 12434 42072 12440 42084
rect 11287 42044 12440 42072
rect 11287 42041 11299 42044
rect 11241 42035 11299 42041
rect 12434 42032 12440 42044
rect 12492 42032 12498 42084
rect 14292 42072 14320 42103
rect 15120 42084 15148 42180
rect 18414 42100 18420 42152
rect 18472 42140 18478 42152
rect 18693 42143 18751 42149
rect 18693 42140 18705 42143
rect 18472 42112 18705 42140
rect 18472 42100 18478 42112
rect 18693 42109 18705 42112
rect 18739 42140 18751 42143
rect 19153 42143 19211 42149
rect 19153 42140 19165 42143
rect 18739 42112 19165 42140
rect 18739 42109 18751 42112
rect 18693 42103 18751 42109
rect 19153 42109 19165 42112
rect 19199 42109 19211 42143
rect 19153 42103 19211 42109
rect 20070 42100 20076 42152
rect 20128 42140 20134 42152
rect 20364 42149 20392 42180
rect 20165 42143 20223 42149
rect 20165 42140 20177 42143
rect 20128 42112 20177 42140
rect 20128 42100 20134 42112
rect 20165 42109 20177 42112
rect 20211 42109 20223 42143
rect 20165 42103 20223 42109
rect 20349 42143 20407 42149
rect 20349 42109 20361 42143
rect 20395 42109 20407 42143
rect 20349 42103 20407 42109
rect 20533 42143 20591 42149
rect 20533 42109 20545 42143
rect 20579 42109 20591 42143
rect 20533 42103 20591 42109
rect 15102 42072 15108 42084
rect 14016 42044 14320 42072
rect 15063 42044 15108 42072
rect 14016 42016 14044 42044
rect 15102 42032 15108 42044
rect 15160 42032 15166 42084
rect 19334 42032 19340 42084
rect 19392 42072 19398 42084
rect 20548 42072 20576 42103
rect 19392 42044 20576 42072
rect 19392 42032 19398 42044
rect 11514 42004 11520 42016
rect 8159 41976 9260 42004
rect 11475 41976 11520 42004
rect 8159 41973 8171 41976
rect 8113 41967 8171 41973
rect 11514 41964 11520 41976
rect 11572 41964 11578 42016
rect 11606 41964 11612 42016
rect 11664 42004 11670 42016
rect 12066 42004 12072 42016
rect 11664 41976 12072 42004
rect 11664 41964 11670 41976
rect 12066 41964 12072 41976
rect 12124 42004 12130 42016
rect 12621 42007 12679 42013
rect 12621 42004 12633 42007
rect 12124 41976 12633 42004
rect 12124 41964 12130 41976
rect 12621 41973 12633 41976
rect 12667 41973 12679 42007
rect 13998 42004 14004 42016
rect 13959 41976 14004 42004
rect 12621 41967 12679 41973
rect 13998 41964 14004 41976
rect 14056 41964 14062 42016
rect 20916 42004 20944 42180
rect 21634 42168 21640 42180
rect 21692 42208 21698 42220
rect 22557 42211 22615 42217
rect 22557 42208 22569 42211
rect 21692 42180 22569 42208
rect 21692 42168 21698 42180
rect 22557 42177 22569 42180
rect 22603 42177 22615 42211
rect 25056 42208 25084 42307
rect 26786 42304 26792 42316
rect 26844 42304 26850 42356
rect 25590 42276 25596 42288
rect 25551 42248 25596 42276
rect 25590 42236 25596 42248
rect 25648 42236 25654 42288
rect 25958 42276 25964 42288
rect 25919 42248 25964 42276
rect 25958 42236 25964 42248
rect 26016 42236 26022 42288
rect 22557 42171 22615 42177
rect 24136 42180 25084 42208
rect 21453 42143 21511 42149
rect 21453 42109 21465 42143
rect 21499 42140 21511 42143
rect 21818 42140 21824 42152
rect 21499 42112 21824 42140
rect 21499 42109 21511 42112
rect 21453 42103 21511 42109
rect 21818 42100 21824 42112
rect 21876 42140 21882 42152
rect 22097 42143 22155 42149
rect 22097 42140 22109 42143
rect 21876 42112 22109 42140
rect 21876 42100 21882 42112
rect 22097 42109 22109 42112
rect 22143 42140 22155 42143
rect 22143 42112 22324 42140
rect 22143 42109 22155 42112
rect 22097 42103 22155 42109
rect 21545 42075 21603 42081
rect 21545 42041 21557 42075
rect 21591 42072 21603 42075
rect 22186 42072 22192 42084
rect 21591 42044 22192 42072
rect 21591 42041 21603 42044
rect 21545 42035 21603 42041
rect 22186 42032 22192 42044
rect 22244 42032 22250 42084
rect 22296 42072 22324 42112
rect 22370 42100 22376 42152
rect 22428 42140 22434 42152
rect 24136 42149 24164 42180
rect 25866 42168 25872 42220
rect 25924 42208 25930 42220
rect 26326 42208 26332 42220
rect 25924 42180 26332 42208
rect 25924 42168 25930 42180
rect 26326 42168 26332 42180
rect 26384 42208 26390 42220
rect 26421 42211 26479 42217
rect 26421 42208 26433 42211
rect 26384 42180 26433 42208
rect 26384 42168 26390 42180
rect 26421 42177 26433 42180
rect 26467 42177 26479 42211
rect 26421 42171 26479 42177
rect 26510 42168 26516 42220
rect 26568 42168 26574 42220
rect 24121 42143 24179 42149
rect 22428 42112 22473 42140
rect 22428 42100 22434 42112
rect 24121 42109 24133 42143
rect 24167 42109 24179 42143
rect 24302 42140 24308 42152
rect 24263 42112 24308 42140
rect 24121 42103 24179 42109
rect 24302 42100 24308 42112
rect 24360 42100 24366 42152
rect 24489 42143 24547 42149
rect 24489 42109 24501 42143
rect 24535 42109 24547 42143
rect 24489 42103 24547 42109
rect 26145 42143 26203 42149
rect 26145 42109 26157 42143
rect 26191 42140 26203 42143
rect 26528 42140 26556 42168
rect 27522 42140 27528 42152
rect 26191 42112 27528 42140
rect 26191 42109 26203 42112
rect 26145 42103 26203 42109
rect 22646 42072 22652 42084
rect 22296 42044 22652 42072
rect 22646 42032 22652 42044
rect 22704 42072 22710 42084
rect 23477 42075 23535 42081
rect 23477 42072 23489 42075
rect 22704 42044 23489 42072
rect 22704 42032 22710 42044
rect 23477 42041 23489 42044
rect 23523 42072 23535 42075
rect 24504 42072 24532 42103
rect 23523 42044 24532 42072
rect 23523 42041 23535 42044
rect 23477 42035 23535 42041
rect 25866 42032 25872 42084
rect 25924 42072 25930 42084
rect 26160 42072 26188 42103
rect 27522 42100 27528 42112
rect 27580 42100 27586 42152
rect 25924 42044 26188 42072
rect 25924 42032 25930 42044
rect 22094 42004 22100 42016
rect 20916 41976 22100 42004
rect 22094 41964 22100 41976
rect 22152 41964 22158 42016
rect 22462 41964 22468 42016
rect 22520 42004 22526 42016
rect 22925 42007 22983 42013
rect 22925 42004 22937 42007
rect 22520 41976 22937 42004
rect 22520 41964 22526 41976
rect 22925 41973 22937 41976
rect 22971 42004 22983 42007
rect 23290 42004 23296 42016
rect 22971 41976 23296 42004
rect 22971 41973 22983 41976
rect 22925 41967 22983 41973
rect 23290 41964 23296 41976
rect 23348 41964 23354 42016
rect 27154 41964 27160 42016
rect 27212 42004 27218 42016
rect 27525 42007 27583 42013
rect 27525 42004 27537 42007
rect 27212 41976 27537 42004
rect 27212 41964 27218 41976
rect 27525 41973 27537 41976
rect 27571 41973 27583 42007
rect 27525 41967 27583 41973
rect 1104 41914 28888 41936
rect 1104 41862 10982 41914
rect 11034 41862 11046 41914
rect 11098 41862 11110 41914
rect 11162 41862 11174 41914
rect 11226 41862 20982 41914
rect 21034 41862 21046 41914
rect 21098 41862 21110 41914
rect 21162 41862 21174 41914
rect 21226 41862 28888 41914
rect 1104 41840 28888 41862
rect 8665 41803 8723 41809
rect 8665 41769 8677 41803
rect 8711 41800 8723 41803
rect 10042 41800 10048 41812
rect 8711 41772 10048 41800
rect 8711 41769 8723 41772
rect 8665 41763 8723 41769
rect 10042 41760 10048 41772
rect 10100 41760 10106 41812
rect 17402 41760 17408 41812
rect 17460 41800 17466 41812
rect 17678 41800 17684 41812
rect 17460 41772 17684 41800
rect 17460 41760 17466 41772
rect 17678 41760 17684 41772
rect 17736 41760 17742 41812
rect 18141 41803 18199 41809
rect 18141 41769 18153 41803
rect 18187 41800 18199 41803
rect 18966 41800 18972 41812
rect 18187 41772 18972 41800
rect 18187 41769 18199 41772
rect 18141 41763 18199 41769
rect 18966 41760 18972 41772
rect 19024 41760 19030 41812
rect 19334 41760 19340 41812
rect 19392 41800 19398 41812
rect 19613 41803 19671 41809
rect 19613 41800 19625 41803
rect 19392 41772 19625 41800
rect 19392 41760 19398 41772
rect 19613 41769 19625 41772
rect 19659 41769 19671 41803
rect 19613 41763 19671 41769
rect 19886 41760 19892 41812
rect 19944 41800 19950 41812
rect 20346 41800 20352 41812
rect 19944 41772 20352 41800
rect 19944 41760 19950 41772
rect 20346 41760 20352 41772
rect 20404 41760 20410 41812
rect 21818 41800 21824 41812
rect 21779 41772 21824 41800
rect 21818 41760 21824 41772
rect 21876 41760 21882 41812
rect 22189 41803 22247 41809
rect 22189 41769 22201 41803
rect 22235 41800 22247 41803
rect 22462 41800 22468 41812
rect 22235 41772 22468 41800
rect 22235 41769 22247 41772
rect 22189 41763 22247 41769
rect 22462 41760 22468 41772
rect 22520 41800 22526 41812
rect 22738 41800 22744 41812
rect 22520 41772 22744 41800
rect 22520 41760 22526 41772
rect 22738 41760 22744 41772
rect 22796 41760 22802 41812
rect 24029 41803 24087 41809
rect 24029 41769 24041 41803
rect 24075 41800 24087 41803
rect 24578 41800 24584 41812
rect 24075 41772 24584 41800
rect 24075 41769 24087 41772
rect 24029 41763 24087 41769
rect 24578 41760 24584 41772
rect 24636 41760 24642 41812
rect 25685 41803 25743 41809
rect 25685 41769 25697 41803
rect 25731 41800 25743 41803
rect 25774 41800 25780 41812
rect 25731 41772 25780 41800
rect 25731 41769 25743 41772
rect 25685 41763 25743 41769
rect 25774 41760 25780 41772
rect 25832 41760 25838 41812
rect 26237 41803 26295 41809
rect 26237 41769 26249 41803
rect 26283 41800 26295 41803
rect 26326 41800 26332 41812
rect 26283 41772 26332 41800
rect 26283 41769 26295 41772
rect 26237 41763 26295 41769
rect 26326 41760 26332 41772
rect 26384 41760 26390 41812
rect 27522 41800 27528 41812
rect 27483 41772 27528 41800
rect 27522 41760 27528 41772
rect 27580 41760 27586 41812
rect 10781 41735 10839 41741
rect 10781 41701 10793 41735
rect 10827 41732 10839 41735
rect 11422 41732 11428 41744
rect 10827 41704 11428 41732
rect 10827 41701 10839 41704
rect 10781 41695 10839 41701
rect 11422 41692 11428 41704
rect 11480 41732 11486 41744
rect 20714 41732 20720 41744
rect 11480 41704 11928 41732
rect 20675 41704 20720 41732
rect 11480 41692 11486 41704
rect 11900 41673 11928 41704
rect 20714 41692 20720 41704
rect 20772 41692 20778 41744
rect 21453 41735 21511 41741
rect 21453 41701 21465 41735
rect 21499 41732 21511 41735
rect 22370 41732 22376 41744
rect 21499 41704 22376 41732
rect 21499 41701 21511 41704
rect 21453 41695 21511 41701
rect 22370 41692 22376 41704
rect 22428 41692 22434 41744
rect 26510 41732 26516 41744
rect 26471 41704 26516 41732
rect 26510 41692 26516 41704
rect 26568 41692 26574 41744
rect 11517 41667 11575 41673
rect 11517 41633 11529 41667
rect 11563 41633 11575 41667
rect 11517 41627 11575 41633
rect 11885 41667 11943 41673
rect 11885 41633 11897 41667
rect 11931 41633 11943 41667
rect 11885 41627 11943 41633
rect 10778 41556 10784 41608
rect 10836 41596 10842 41608
rect 11425 41599 11483 41605
rect 11425 41596 11437 41599
rect 10836 41568 11437 41596
rect 10836 41556 10842 41568
rect 11425 41565 11437 41568
rect 11471 41565 11483 41599
rect 11425 41559 11483 41565
rect 10413 41531 10471 41537
rect 10413 41497 10425 41531
rect 10459 41528 10471 41531
rect 10870 41528 10876 41540
rect 10459 41500 10876 41528
rect 10459 41497 10471 41500
rect 10413 41491 10471 41497
rect 10870 41488 10876 41500
rect 10928 41488 10934 41540
rect 11532 41528 11560 41627
rect 19426 41624 19432 41676
rect 19484 41664 19490 41676
rect 19797 41667 19855 41673
rect 19797 41664 19809 41667
rect 19484 41636 19809 41664
rect 19484 41624 19490 41636
rect 19797 41633 19809 41636
rect 19843 41664 19855 41667
rect 19978 41664 19984 41676
rect 19843 41636 19984 41664
rect 19843 41633 19855 41636
rect 19797 41627 19855 41633
rect 19978 41624 19984 41636
rect 20036 41624 20042 41676
rect 20901 41667 20959 41673
rect 20901 41633 20913 41667
rect 20947 41633 20959 41667
rect 20901 41627 20959 41633
rect 21085 41667 21143 41673
rect 21085 41633 21097 41667
rect 21131 41664 21143 41667
rect 21266 41664 21272 41676
rect 21131 41636 21272 41664
rect 21131 41633 21143 41636
rect 21085 41627 21143 41633
rect 11790 41556 11796 41608
rect 11848 41596 11854 41608
rect 11977 41599 12035 41605
rect 11977 41596 11989 41599
rect 11848 41568 11989 41596
rect 11848 41556 11854 41568
rect 11977 41565 11989 41568
rect 12023 41565 12035 41599
rect 11977 41559 12035 41565
rect 12342 41528 12348 41540
rect 11532 41500 12348 41528
rect 12342 41488 12348 41500
rect 12400 41488 12406 41540
rect 19150 41488 19156 41540
rect 19208 41528 19214 41540
rect 19981 41531 20039 41537
rect 19981 41528 19993 41531
rect 19208 41500 19993 41528
rect 19208 41488 19214 41500
rect 19981 41497 19993 41500
rect 20027 41497 20039 41531
rect 20916 41528 20944 41627
rect 21266 41624 21272 41636
rect 21324 41624 21330 41676
rect 22554 41664 22560 41676
rect 22515 41636 22560 41664
rect 22554 41624 22560 41636
rect 22612 41624 22618 41676
rect 23014 41624 23020 41676
rect 23072 41664 23078 41676
rect 23109 41667 23167 41673
rect 23109 41664 23121 41667
rect 23072 41636 23121 41664
rect 23072 41624 23078 41636
rect 23109 41633 23121 41636
rect 23155 41633 23167 41667
rect 23109 41627 23167 41633
rect 24578 41624 24584 41676
rect 24636 41664 24642 41676
rect 25133 41667 25191 41673
rect 25133 41664 25145 41667
rect 24636 41636 25145 41664
rect 24636 41624 24642 41636
rect 25133 41633 25145 41636
rect 25179 41633 25191 41667
rect 27154 41664 27160 41676
rect 27115 41636 27160 41664
rect 25133 41627 25191 41633
rect 27154 41624 27160 41636
rect 27212 41624 27218 41676
rect 22002 41556 22008 41608
rect 22060 41596 22066 41608
rect 23198 41596 23204 41608
rect 22060 41568 23204 41596
rect 22060 41556 22066 41568
rect 23198 41556 23204 41568
rect 23256 41556 23262 41608
rect 24305 41599 24363 41605
rect 24305 41596 24317 41599
rect 23584 41568 24317 41596
rect 22462 41528 22468 41540
rect 20916 41500 22468 41528
rect 19981 41491 20039 41497
rect 22462 41488 22468 41500
rect 22520 41488 22526 41540
rect 23584 41472 23612 41568
rect 24305 41565 24317 41568
rect 24351 41565 24363 41599
rect 24305 41559 24363 41565
rect 24320 41528 24348 41559
rect 24394 41556 24400 41608
rect 24452 41596 24458 41608
rect 24452 41568 24497 41596
rect 24452 41556 24458 41568
rect 24670 41556 24676 41608
rect 24728 41596 24734 41608
rect 25225 41599 25283 41605
rect 25225 41596 25237 41599
rect 24728 41568 25237 41596
rect 24728 41556 24734 41568
rect 25225 41565 25237 41568
rect 25271 41565 25283 41599
rect 25225 41559 25283 41565
rect 25038 41528 25044 41540
rect 24320 41500 25044 41528
rect 25038 41488 25044 41500
rect 25096 41488 25102 41540
rect 9030 41460 9036 41472
rect 8991 41432 9036 41460
rect 9030 41420 9036 41432
rect 9088 41420 9094 41472
rect 10965 41463 11023 41469
rect 10965 41429 10977 41463
rect 11011 41460 11023 41463
rect 11330 41460 11336 41472
rect 11011 41432 11336 41460
rect 11011 41429 11023 41432
rect 10965 41423 11023 41429
rect 11330 41420 11336 41432
rect 11388 41420 11394 41472
rect 15654 41420 15660 41472
rect 15712 41460 15718 41472
rect 16117 41463 16175 41469
rect 16117 41460 16129 41463
rect 15712 41432 16129 41460
rect 15712 41420 15718 41432
rect 16117 41429 16129 41432
rect 16163 41429 16175 41463
rect 16117 41423 16175 41429
rect 23385 41463 23443 41469
rect 23385 41429 23397 41463
rect 23431 41460 23443 41463
rect 23566 41460 23572 41472
rect 23431 41432 23572 41460
rect 23431 41429 23443 41432
rect 23385 41423 23443 41429
rect 23566 41420 23572 41432
rect 23624 41420 23630 41472
rect 1104 41370 28888 41392
rect 1104 41318 5982 41370
rect 6034 41318 6046 41370
rect 6098 41318 6110 41370
rect 6162 41318 6174 41370
rect 6226 41318 15982 41370
rect 16034 41318 16046 41370
rect 16098 41318 16110 41370
rect 16162 41318 16174 41370
rect 16226 41318 25982 41370
rect 26034 41318 26046 41370
rect 26098 41318 26110 41370
rect 26162 41318 26174 41370
rect 26226 41318 28888 41370
rect 1104 41296 28888 41318
rect 11790 41256 11796 41268
rect 11751 41228 11796 41256
rect 11790 41216 11796 41228
rect 11848 41256 11854 41268
rect 12526 41256 12532 41268
rect 11848 41228 12532 41256
rect 11848 41216 11854 41228
rect 12526 41216 12532 41228
rect 12584 41216 12590 41268
rect 19794 41256 19800 41268
rect 19755 41228 19800 41256
rect 19794 41216 19800 41228
rect 19852 41216 19858 41268
rect 19978 41216 19984 41268
rect 20036 41256 20042 41268
rect 20073 41259 20131 41265
rect 20073 41256 20085 41259
rect 20036 41228 20085 41256
rect 20036 41216 20042 41228
rect 20073 41225 20085 41228
rect 20119 41225 20131 41259
rect 22462 41256 22468 41268
rect 22423 41228 22468 41256
rect 20073 41219 20131 41225
rect 22462 41216 22468 41228
rect 22520 41216 22526 41268
rect 22833 41259 22891 41265
rect 22833 41225 22845 41259
rect 22879 41256 22891 41259
rect 23014 41256 23020 41268
rect 22879 41228 23020 41256
rect 22879 41225 22891 41228
rect 22833 41219 22891 41225
rect 23014 41216 23020 41228
rect 23072 41216 23078 41268
rect 26329 41259 26387 41265
rect 26329 41225 26341 41259
rect 26375 41256 26387 41259
rect 26878 41256 26884 41268
rect 26375 41228 26884 41256
rect 26375 41225 26387 41228
rect 26329 41219 26387 41225
rect 26878 41216 26884 41228
rect 26936 41216 26942 41268
rect 10042 41148 10048 41200
rect 10100 41188 10106 41200
rect 11149 41191 11207 41197
rect 11149 41188 11161 41191
rect 10100 41160 11161 41188
rect 10100 41148 10106 41160
rect 11149 41157 11161 41160
rect 11195 41157 11207 41191
rect 11149 41151 11207 41157
rect 16393 41191 16451 41197
rect 16393 41157 16405 41191
rect 16439 41188 16451 41191
rect 16482 41188 16488 41200
rect 16439 41160 16488 41188
rect 16439 41157 16451 41160
rect 16393 41151 16451 41157
rect 16482 41148 16488 41160
rect 16540 41148 16546 41200
rect 19521 41191 19579 41197
rect 19521 41157 19533 41191
rect 19567 41188 19579 41191
rect 19702 41188 19708 41200
rect 19567 41160 19708 41188
rect 19567 41157 19579 41160
rect 19521 41151 19579 41157
rect 9861 41123 9919 41129
rect 9861 41089 9873 41123
rect 9907 41120 9919 41123
rect 9907 41092 11284 41120
rect 9907 41089 9919 41092
rect 9861 41083 9919 41089
rect 10321 41055 10379 41061
rect 10321 41052 10333 41055
rect 10152 41024 10333 41052
rect 10152 40928 10180 41024
rect 10321 41021 10333 41024
rect 10367 41021 10379 41055
rect 10686 41052 10692 41064
rect 10647 41024 10692 41052
rect 10321 41015 10379 41021
rect 10686 41012 10692 41024
rect 10744 41052 10750 41064
rect 10870 41052 10876 41064
rect 10744 41024 10876 41052
rect 10744 41012 10750 41024
rect 10870 41012 10876 41024
rect 10928 41012 10934 41064
rect 11256 41061 11284 41092
rect 15654 41080 15660 41132
rect 15712 41120 15718 41132
rect 15712 41092 16804 41120
rect 15712 41080 15718 41092
rect 11241 41055 11299 41061
rect 11241 41021 11253 41055
rect 11287 41052 11299 41055
rect 11514 41052 11520 41064
rect 11287 41024 11520 41052
rect 11287 41021 11299 41024
rect 11241 41015 11299 41021
rect 11514 41012 11520 41024
rect 11572 41052 11578 41064
rect 11698 41052 11704 41064
rect 11572 41024 11704 41052
rect 11572 41012 11578 41024
rect 11698 41012 11704 41024
rect 11756 41012 11762 41064
rect 16574 41052 16580 41064
rect 16535 41024 16580 41052
rect 16574 41012 16580 41024
rect 16632 41012 16638 41064
rect 16776 41061 16804 41092
rect 16761 41055 16819 41061
rect 16761 41021 16773 41055
rect 16807 41021 16819 41055
rect 16942 41052 16948 41064
rect 16903 41024 16948 41052
rect 16761 41015 16819 41021
rect 16942 41012 16948 41024
rect 17000 41012 17006 41064
rect 19628 41061 19656 41160
rect 19702 41148 19708 41160
rect 19760 41148 19766 41200
rect 20533 41191 20591 41197
rect 20533 41157 20545 41191
rect 20579 41188 20591 41191
rect 21634 41188 21640 41200
rect 20579 41160 21640 41188
rect 20579 41157 20591 41160
rect 20533 41151 20591 41157
rect 21634 41148 21640 41160
rect 21692 41188 21698 41200
rect 21910 41188 21916 41200
rect 21692 41160 21916 41188
rect 21692 41148 21698 41160
rect 21910 41148 21916 41160
rect 21968 41188 21974 41200
rect 26789 41191 26847 41197
rect 21968 41160 22048 41188
rect 21968 41148 21974 41160
rect 21174 41120 21180 41132
rect 21135 41092 21180 41120
rect 21174 41080 21180 41092
rect 21232 41080 21238 41132
rect 22020 41129 22048 41160
rect 26789 41157 26801 41191
rect 26835 41188 26847 41191
rect 27154 41188 27160 41200
rect 26835 41160 27160 41188
rect 26835 41157 26847 41160
rect 26789 41151 26847 41157
rect 27154 41148 27160 41160
rect 27212 41148 27218 41200
rect 22005 41123 22063 41129
rect 22005 41089 22017 41123
rect 22051 41089 22063 41123
rect 22005 41083 22063 41089
rect 24673 41123 24731 41129
rect 24673 41089 24685 41123
rect 24719 41120 24731 41123
rect 24719 41092 25084 41120
rect 24719 41089 24731 41092
rect 24673 41083 24731 41089
rect 19613 41055 19671 41061
rect 19613 41021 19625 41055
rect 19659 41021 19671 41055
rect 19613 41015 19671 41021
rect 21085 41055 21143 41061
rect 21085 41021 21097 41055
rect 21131 41052 21143 41055
rect 21542 41052 21548 41064
rect 21131 41024 21548 41052
rect 21131 41021 21143 41024
rect 21085 41015 21143 41021
rect 21542 41012 21548 41024
rect 21600 41012 21606 41064
rect 21634 41012 21640 41064
rect 21692 41052 21698 41064
rect 21818 41052 21824 41064
rect 21692 41024 21824 41052
rect 21692 41012 21698 41024
rect 21818 41012 21824 41024
rect 21876 41052 21882 41064
rect 21913 41055 21971 41061
rect 21913 41052 21925 41055
rect 21876 41024 21925 41052
rect 21876 41012 21882 41024
rect 21913 41021 21925 41024
rect 21959 41021 21971 41055
rect 21913 41015 21971 41021
rect 23658 41012 23664 41064
rect 23716 41052 23722 41064
rect 25056 41061 25084 41092
rect 23753 41055 23811 41061
rect 23753 41052 23765 41055
rect 23716 41024 23765 41052
rect 23716 41012 23722 41024
rect 23753 41021 23765 41024
rect 23799 41052 23811 41055
rect 24213 41055 24271 41061
rect 24213 41052 24225 41055
rect 23799 41024 24225 41052
rect 23799 41021 23811 41024
rect 23753 41015 23811 41021
rect 24213 41021 24225 41024
rect 24259 41021 24271 41055
rect 24213 41015 24271 41021
rect 24765 41055 24823 41061
rect 24765 41021 24777 41055
rect 24811 41052 24823 41055
rect 25041 41055 25099 41061
rect 24811 41024 24900 41052
rect 24811 41021 24823 41024
rect 24765 41015 24823 41021
rect 15746 40944 15752 40996
rect 15804 40984 15810 40996
rect 16025 40987 16083 40993
rect 16025 40984 16037 40987
rect 15804 40956 16037 40984
rect 15804 40944 15810 40956
rect 16025 40953 16037 40956
rect 16071 40984 16083 40987
rect 16960 40984 16988 41012
rect 16071 40956 16988 40984
rect 20901 40987 20959 40993
rect 16071 40953 16083 40956
rect 16025 40947 16083 40953
rect 20901 40953 20913 40987
rect 20947 40984 20959 40987
rect 21652 40984 21680 41012
rect 20947 40956 21680 40984
rect 23477 40987 23535 40993
rect 20947 40953 20959 40956
rect 20901 40947 20959 40953
rect 23477 40953 23489 40987
rect 23523 40984 23535 40987
rect 24302 40984 24308 40996
rect 23523 40956 24308 40984
rect 23523 40953 23535 40956
rect 23477 40947 23535 40953
rect 24302 40944 24308 40956
rect 24360 40984 24366 40996
rect 24670 40984 24676 40996
rect 24360 40956 24676 40984
rect 24360 40944 24366 40956
rect 24670 40944 24676 40956
rect 24728 40944 24734 40996
rect 10134 40916 10140 40928
rect 10095 40888 10140 40916
rect 10134 40876 10140 40888
rect 10192 40876 10198 40928
rect 12066 40916 12072 40928
rect 12027 40888 12072 40916
rect 12066 40876 12072 40888
rect 12124 40876 12130 40928
rect 12434 40876 12440 40928
rect 12492 40916 12498 40928
rect 12713 40919 12771 40925
rect 12713 40916 12725 40919
rect 12492 40888 12725 40916
rect 12492 40876 12498 40888
rect 12713 40885 12725 40888
rect 12759 40916 12771 40919
rect 12802 40916 12808 40928
rect 12759 40888 12808 40916
rect 12759 40885 12771 40888
rect 12713 40879 12771 40885
rect 12802 40876 12808 40888
rect 12860 40876 12866 40928
rect 13078 40916 13084 40928
rect 13039 40888 13084 40916
rect 13078 40876 13084 40888
rect 13136 40876 13142 40928
rect 23934 40916 23940 40928
rect 23895 40888 23940 40916
rect 23934 40876 23940 40888
rect 23992 40876 23998 40928
rect 24872 40916 24900 41024
rect 25041 41021 25053 41055
rect 25087 41052 25099 41055
rect 25314 41052 25320 41064
rect 25087 41024 25320 41052
rect 25087 41021 25099 41024
rect 25041 41015 25099 41021
rect 25314 41012 25320 41024
rect 25372 41012 25378 41064
rect 25866 40916 25872 40928
rect 24872 40888 25872 40916
rect 25866 40876 25872 40888
rect 25924 40876 25930 40928
rect 1104 40826 28888 40848
rect 1104 40774 10982 40826
rect 11034 40774 11046 40826
rect 11098 40774 11110 40826
rect 11162 40774 11174 40826
rect 11226 40774 20982 40826
rect 21034 40774 21046 40826
rect 21098 40774 21110 40826
rect 21162 40774 21174 40826
rect 21226 40774 28888 40826
rect 1104 40752 28888 40774
rect 10778 40672 10784 40724
rect 10836 40712 10842 40724
rect 10873 40715 10931 40721
rect 10873 40712 10885 40715
rect 10836 40684 10885 40712
rect 10836 40672 10842 40684
rect 10873 40681 10885 40684
rect 10919 40681 10931 40715
rect 10873 40675 10931 40681
rect 20717 40715 20775 40721
rect 20717 40681 20729 40715
rect 20763 40712 20775 40715
rect 21266 40712 21272 40724
rect 20763 40684 21272 40712
rect 20763 40681 20775 40684
rect 20717 40675 20775 40681
rect 21266 40672 21272 40684
rect 21324 40672 21330 40724
rect 21542 40712 21548 40724
rect 21503 40684 21548 40712
rect 21542 40672 21548 40684
rect 21600 40672 21606 40724
rect 21913 40715 21971 40721
rect 21913 40681 21925 40715
rect 21959 40712 21971 40715
rect 22002 40712 22008 40724
rect 21959 40684 22008 40712
rect 21959 40681 21971 40684
rect 21913 40675 21971 40681
rect 22002 40672 22008 40684
rect 22060 40672 22066 40724
rect 23198 40672 23204 40724
rect 23256 40712 23262 40724
rect 23385 40715 23443 40721
rect 23385 40712 23397 40715
rect 23256 40684 23397 40712
rect 23256 40672 23262 40684
rect 23385 40681 23397 40684
rect 23431 40681 23443 40715
rect 25038 40712 25044 40724
rect 24999 40684 25044 40712
rect 23385 40675 23443 40681
rect 25038 40672 25044 40684
rect 25096 40672 25102 40724
rect 25501 40715 25559 40721
rect 25501 40681 25513 40715
rect 25547 40712 25559 40715
rect 25866 40712 25872 40724
rect 25547 40684 25872 40712
rect 25547 40681 25559 40684
rect 25501 40675 25559 40681
rect 25866 40672 25872 40684
rect 25924 40672 25930 40724
rect 10413 40579 10471 40585
rect 10413 40545 10425 40579
rect 10459 40576 10471 40579
rect 10502 40576 10508 40588
rect 10459 40548 10508 40576
rect 10459 40545 10471 40548
rect 10413 40539 10471 40545
rect 10502 40536 10508 40548
rect 10560 40576 10566 40588
rect 10796 40576 10824 40672
rect 13078 40644 13084 40656
rect 12452 40616 13084 40644
rect 12066 40576 12072 40588
rect 10560 40548 10824 40576
rect 12027 40548 12072 40576
rect 10560 40536 10566 40548
rect 12066 40536 12072 40548
rect 12124 40576 12130 40588
rect 12342 40576 12348 40588
rect 12124 40548 12348 40576
rect 12124 40536 12130 40548
rect 12342 40536 12348 40548
rect 12400 40536 12406 40588
rect 12452 40585 12480 40616
rect 13078 40604 13084 40616
rect 13136 40604 13142 40656
rect 16758 40604 16764 40656
rect 16816 40604 16822 40656
rect 22554 40644 22560 40656
rect 22515 40616 22560 40644
rect 22554 40604 22560 40616
rect 22612 40644 22618 40656
rect 22833 40647 22891 40653
rect 22833 40644 22845 40647
rect 22612 40616 22845 40644
rect 22612 40604 22618 40616
rect 22833 40613 22845 40616
rect 22879 40613 22891 40647
rect 22833 40607 22891 40613
rect 12437 40579 12495 40585
rect 12437 40545 12449 40579
rect 12483 40545 12495 40579
rect 12437 40539 12495 40545
rect 14001 40579 14059 40585
rect 14001 40545 14013 40579
rect 14047 40576 14059 40579
rect 14182 40576 14188 40588
rect 14047 40548 14188 40576
rect 14047 40545 14059 40548
rect 14001 40539 14059 40545
rect 14182 40536 14188 40548
rect 14240 40536 14246 40588
rect 16577 40579 16635 40585
rect 16577 40545 16589 40579
rect 16623 40545 16635 40579
rect 16776 40576 16804 40604
rect 17037 40579 17095 40585
rect 17037 40576 17049 40579
rect 16776 40548 17049 40576
rect 16577 40539 16635 40545
rect 17037 40545 17049 40548
rect 17083 40545 17095 40579
rect 20990 40576 20996 40588
rect 20951 40548 20996 40576
rect 17037 40539 17095 40545
rect 10045 40511 10103 40517
rect 10045 40477 10057 40511
rect 10091 40508 10103 40511
rect 10226 40508 10232 40520
rect 10091 40480 10232 40508
rect 10091 40477 10103 40480
rect 10045 40471 10103 40477
rect 10226 40468 10232 40480
rect 10284 40468 10290 40520
rect 11974 40508 11980 40520
rect 10612 40480 11980 40508
rect 1486 40332 1492 40384
rect 1544 40372 1550 40384
rect 1581 40375 1639 40381
rect 1581 40372 1593 40375
rect 1544 40344 1593 40372
rect 1544 40332 1550 40344
rect 1581 40341 1593 40344
rect 1627 40341 1639 40375
rect 1581 40335 1639 40341
rect 10042 40332 10048 40384
rect 10100 40372 10106 40384
rect 10612 40381 10640 40480
rect 11974 40468 11980 40480
rect 12032 40468 12038 40520
rect 12526 40508 12532 40520
rect 12487 40480 12532 40508
rect 12526 40468 12532 40480
rect 12584 40468 12590 40520
rect 16592 40508 16620 40539
rect 20990 40536 20996 40548
rect 21048 40536 21054 40588
rect 21634 40536 21640 40588
rect 21692 40576 21698 40588
rect 22005 40579 22063 40585
rect 22005 40576 22017 40579
rect 21692 40548 22017 40576
rect 21692 40536 21698 40548
rect 22005 40545 22017 40548
rect 22051 40545 22063 40579
rect 22005 40539 22063 40545
rect 22097 40579 22155 40585
rect 22097 40545 22109 40579
rect 22143 40576 22155 40579
rect 22186 40576 22192 40588
rect 22143 40548 22192 40576
rect 22143 40545 22155 40548
rect 22097 40539 22155 40545
rect 22186 40536 22192 40548
rect 22244 40536 22250 40588
rect 24213 40579 24271 40585
rect 24213 40545 24225 40579
rect 24259 40576 24271 40579
rect 24486 40576 24492 40588
rect 24259 40548 24492 40576
rect 24259 40545 24271 40548
rect 24213 40539 24271 40545
rect 24486 40536 24492 40548
rect 24544 40536 24550 40588
rect 24581 40579 24639 40585
rect 24581 40545 24593 40579
rect 24627 40576 24639 40579
rect 25130 40576 25136 40588
rect 24627 40548 25136 40576
rect 24627 40545 24639 40548
rect 24581 40539 24639 40545
rect 25130 40536 25136 40548
rect 25188 40536 25194 40588
rect 16761 40511 16819 40517
rect 16761 40508 16773 40511
rect 16592 40480 16773 40508
rect 16761 40477 16773 40480
rect 16807 40508 16819 40511
rect 17218 40508 17224 40520
rect 16807 40480 17224 40508
rect 16807 40477 16819 40480
rect 16761 40471 16819 40477
rect 17218 40468 17224 40480
rect 17276 40508 17282 40520
rect 17402 40508 17408 40520
rect 17276 40480 17408 40508
rect 17276 40468 17282 40480
rect 17402 40468 17408 40480
rect 17460 40468 17466 40520
rect 11333 40443 11391 40449
rect 11333 40409 11345 40443
rect 11379 40440 11391 40443
rect 11790 40440 11796 40452
rect 11379 40412 11796 40440
rect 11379 40409 11391 40412
rect 11333 40403 11391 40409
rect 11790 40400 11796 40412
rect 11848 40400 11854 40452
rect 16209 40443 16267 40449
rect 16209 40409 16221 40443
rect 16255 40440 16267 40443
rect 16574 40440 16580 40452
rect 16255 40412 16580 40440
rect 16255 40409 16267 40412
rect 16209 40403 16267 40409
rect 16574 40400 16580 40412
rect 16632 40400 16638 40452
rect 21177 40443 21235 40449
rect 21177 40409 21189 40443
rect 21223 40440 21235 40443
rect 21652 40440 21680 40536
rect 23290 40468 23296 40520
rect 23348 40508 23354 40520
rect 24121 40511 24179 40517
rect 24121 40508 24133 40511
rect 23348 40480 24133 40508
rect 23348 40468 23354 40480
rect 24121 40477 24133 40480
rect 24167 40477 24179 40511
rect 24121 40471 24179 40477
rect 24673 40511 24731 40517
rect 24673 40477 24685 40511
rect 24719 40477 24731 40511
rect 24673 40471 24731 40477
rect 21223 40412 21680 40440
rect 21223 40409 21235 40412
rect 21177 40403 21235 40409
rect 24578 40400 24584 40452
rect 24636 40440 24642 40452
rect 24688 40440 24716 40471
rect 24636 40412 24716 40440
rect 24636 40400 24642 40412
rect 10597 40375 10655 40381
rect 10597 40372 10609 40375
rect 10100 40344 10609 40372
rect 10100 40332 10106 40344
rect 10597 40341 10609 40344
rect 10643 40341 10655 40375
rect 11514 40372 11520 40384
rect 11475 40344 11520 40372
rect 10597 40335 10655 40341
rect 11514 40332 11520 40344
rect 11572 40332 11578 40384
rect 12894 40372 12900 40384
rect 12855 40344 12900 40372
rect 12894 40332 12900 40344
rect 12952 40332 12958 40384
rect 12986 40332 12992 40384
rect 13044 40372 13050 40384
rect 13265 40375 13323 40381
rect 13265 40372 13277 40375
rect 13044 40344 13277 40372
rect 13044 40332 13050 40344
rect 13265 40341 13277 40344
rect 13311 40341 13323 40375
rect 13265 40335 13323 40341
rect 13906 40332 13912 40384
rect 13964 40372 13970 40384
rect 14185 40375 14243 40381
rect 14185 40372 14197 40375
rect 13964 40344 14197 40372
rect 13964 40332 13970 40344
rect 14185 40341 14197 40344
rect 14231 40341 14243 40375
rect 15654 40372 15660 40384
rect 15615 40344 15660 40372
rect 14185 40335 14243 40341
rect 15654 40332 15660 40344
rect 15712 40332 15718 40384
rect 18138 40372 18144 40384
rect 18099 40344 18144 40372
rect 18138 40332 18144 40344
rect 18196 40332 18202 40384
rect 23661 40375 23719 40381
rect 23661 40341 23673 40375
rect 23707 40372 23719 40375
rect 24118 40372 24124 40384
rect 23707 40344 24124 40372
rect 23707 40341 23719 40344
rect 23661 40335 23719 40341
rect 24118 40332 24124 40344
rect 24176 40332 24182 40384
rect 1104 40282 28888 40304
rect 1104 40230 5982 40282
rect 6034 40230 6046 40282
rect 6098 40230 6110 40282
rect 6162 40230 6174 40282
rect 6226 40230 15982 40282
rect 16034 40230 16046 40282
rect 16098 40230 16110 40282
rect 16162 40230 16174 40282
rect 16226 40230 25982 40282
rect 26034 40230 26046 40282
rect 26098 40230 26110 40282
rect 26162 40230 26174 40282
rect 26226 40230 28888 40282
rect 1104 40208 28888 40230
rect 11698 40128 11704 40180
rect 11756 40128 11762 40180
rect 11793 40171 11851 40177
rect 11793 40137 11805 40171
rect 11839 40168 11851 40171
rect 12526 40168 12532 40180
rect 11839 40140 12532 40168
rect 11839 40137 11851 40140
rect 11793 40131 11851 40137
rect 12526 40128 12532 40140
rect 12584 40128 12590 40180
rect 15102 40168 15108 40180
rect 15063 40140 15108 40168
rect 15102 40128 15108 40140
rect 15160 40128 15166 40180
rect 16758 40128 16764 40180
rect 16816 40168 16822 40180
rect 17589 40171 17647 40177
rect 17589 40168 17601 40171
rect 16816 40140 17601 40168
rect 16816 40128 16822 40140
rect 17589 40137 17601 40140
rect 17635 40137 17647 40171
rect 17589 40131 17647 40137
rect 21634 40128 21640 40180
rect 21692 40168 21698 40180
rect 22373 40171 22431 40177
rect 22373 40168 22385 40171
rect 21692 40140 22385 40168
rect 21692 40128 21698 40140
rect 22373 40137 22385 40140
rect 22419 40137 22431 40171
rect 22373 40131 22431 40137
rect 10226 40060 10232 40112
rect 10284 40100 10290 40112
rect 11716 40100 11744 40128
rect 11885 40103 11943 40109
rect 11885 40100 11897 40103
rect 10284 40072 11100 40100
rect 11716 40072 11897 40100
rect 10284 40060 10290 40072
rect 1762 40032 1768 40044
rect 1723 40004 1768 40032
rect 1762 39992 1768 40004
rect 1820 39992 1826 40044
rect 9950 40032 9956 40044
rect 9911 40004 9956 40032
rect 9950 39992 9956 40004
rect 10008 39992 10014 40044
rect 10962 40032 10968 40044
rect 10520 40004 10968 40032
rect 1486 39964 1492 39976
rect 1447 39936 1492 39964
rect 1486 39924 1492 39936
rect 1544 39924 1550 39976
rect 10520 39973 10548 40004
rect 10962 39992 10968 40004
rect 11020 39992 11026 40044
rect 11072 40032 11100 40072
rect 11885 40069 11897 40072
rect 11931 40069 11943 40103
rect 11885 40063 11943 40069
rect 11974 40060 11980 40112
rect 12032 40100 12038 40112
rect 12069 40103 12127 40109
rect 12069 40100 12081 40103
rect 12032 40072 12081 40100
rect 12032 40060 12038 40072
rect 12069 40069 12081 40072
rect 12115 40069 12127 40103
rect 12069 40063 12127 40069
rect 23750 40060 23756 40112
rect 23808 40100 23814 40112
rect 25409 40103 25467 40109
rect 25409 40100 25421 40103
rect 23808 40072 25421 40100
rect 23808 40060 23814 40072
rect 25409 40069 25421 40072
rect 25455 40069 25467 40103
rect 25409 40063 25467 40069
rect 11241 40035 11299 40041
rect 11241 40032 11253 40035
rect 11072 40004 11253 40032
rect 11241 40001 11253 40004
rect 11287 40032 11299 40035
rect 11698 40032 11704 40044
rect 11287 40004 11704 40032
rect 11287 40001 11299 40004
rect 11241 39995 11299 40001
rect 11698 39992 11704 40004
rect 11756 39992 11762 40044
rect 15930 40032 15936 40044
rect 15891 40004 15936 40032
rect 15930 39992 15936 40004
rect 15988 39992 15994 40044
rect 24578 40032 24584 40044
rect 24228 40004 24584 40032
rect 9125 39967 9183 39973
rect 9125 39933 9137 39967
rect 9171 39964 9183 39967
rect 10505 39967 10563 39973
rect 10505 39964 10517 39967
rect 9171 39936 10517 39964
rect 9171 39933 9183 39936
rect 9125 39927 9183 39933
rect 10505 39933 10517 39936
rect 10551 39933 10563 39967
rect 10505 39927 10563 39933
rect 10597 39967 10655 39973
rect 10597 39933 10609 39967
rect 10643 39933 10655 39967
rect 10870 39964 10876 39976
rect 10831 39936 10876 39964
rect 10597 39927 10655 39933
rect 3142 39896 3148 39908
rect 3103 39868 3148 39896
rect 3142 39856 3148 39868
rect 3200 39856 3206 39908
rect 9493 39899 9551 39905
rect 9493 39865 9505 39899
rect 9539 39896 9551 39899
rect 9674 39896 9680 39908
rect 9539 39868 9680 39896
rect 9539 39865 9551 39868
rect 9493 39859 9551 39865
rect 9674 39856 9680 39868
rect 9732 39896 9738 39908
rect 10612 39896 10640 39927
rect 10870 39924 10876 39936
rect 10928 39924 10934 39976
rect 11425 39967 11483 39973
rect 11425 39933 11437 39967
rect 11471 39964 11483 39967
rect 12066 39964 12072 39976
rect 11471 39936 12072 39964
rect 11471 39933 11483 39936
rect 11425 39927 11483 39933
rect 9732 39868 10640 39896
rect 9732 39856 9738 39868
rect 9861 39831 9919 39837
rect 9861 39797 9873 39831
rect 9907 39828 9919 39831
rect 11440 39828 11468 39927
rect 12066 39924 12072 39936
rect 12124 39924 12130 39976
rect 13357 39967 13415 39973
rect 13357 39933 13369 39967
rect 13403 39964 13415 39967
rect 14182 39964 14188 39976
rect 13403 39936 14188 39964
rect 13403 39933 13415 39936
rect 13357 39927 13415 39933
rect 14182 39924 14188 39936
rect 14240 39924 14246 39976
rect 15657 39967 15715 39973
rect 15657 39933 15669 39967
rect 15703 39964 15715 39967
rect 17218 39964 17224 39976
rect 15703 39936 17224 39964
rect 15703 39933 15715 39936
rect 15657 39927 15715 39933
rect 17218 39924 17224 39936
rect 17276 39924 17282 39976
rect 22002 39964 22008 39976
rect 21963 39936 22008 39964
rect 22002 39924 22008 39936
rect 22060 39964 22066 39976
rect 22278 39964 22284 39976
rect 22060 39936 22284 39964
rect 22060 39924 22066 39936
rect 22278 39924 22284 39936
rect 22336 39924 22342 39976
rect 24228 39973 24256 40004
rect 24578 39992 24584 40004
rect 24636 39992 24642 40044
rect 25130 40032 25136 40044
rect 25091 40004 25136 40032
rect 25130 39992 25136 40004
rect 25188 39992 25194 40044
rect 23661 39967 23719 39973
rect 23661 39933 23673 39967
rect 23707 39933 23719 39967
rect 23661 39927 23719 39933
rect 24213 39967 24271 39973
rect 24213 39933 24225 39967
rect 24259 39933 24271 39967
rect 25225 39967 25283 39973
rect 25225 39964 25237 39967
rect 24213 39927 24271 39933
rect 24320 39936 25237 39964
rect 13817 39899 13875 39905
rect 13817 39865 13829 39899
rect 13863 39865 13875 39899
rect 13817 39859 13875 39865
rect 9907 39800 11468 39828
rect 11885 39831 11943 39837
rect 9907 39797 9919 39800
rect 9861 39791 9919 39797
rect 11885 39797 11897 39831
rect 11931 39828 11943 39831
rect 11974 39828 11980 39840
rect 11931 39800 11980 39828
rect 11931 39797 11943 39800
rect 11885 39791 11943 39797
rect 11974 39788 11980 39800
rect 12032 39788 12038 39840
rect 12618 39828 12624 39840
rect 12579 39800 12624 39828
rect 12618 39788 12624 39800
rect 12676 39788 12682 39840
rect 13630 39828 13636 39840
rect 13591 39800 13636 39828
rect 13630 39788 13636 39800
rect 13688 39828 13694 39840
rect 13832 39828 13860 39859
rect 20990 39856 20996 39908
rect 21048 39896 21054 39908
rect 21085 39899 21143 39905
rect 21085 39896 21097 39899
rect 21048 39868 21097 39896
rect 21048 39856 21054 39868
rect 21085 39865 21097 39868
rect 21131 39896 21143 39899
rect 22370 39896 22376 39908
rect 21131 39868 22376 39896
rect 21131 39865 21143 39868
rect 21085 39859 21143 39865
rect 22370 39856 22376 39868
rect 22428 39856 22434 39908
rect 23474 39896 23480 39908
rect 23435 39868 23480 39896
rect 23474 39856 23480 39868
rect 23532 39896 23538 39908
rect 23676 39896 23704 39927
rect 23532 39868 23704 39896
rect 23532 39856 23538 39868
rect 13688 39800 13860 39828
rect 13688 39788 13694 39800
rect 16758 39788 16764 39840
rect 16816 39828 16822 39840
rect 17037 39831 17095 39837
rect 17037 39828 17049 39831
rect 16816 39800 17049 39828
rect 16816 39788 16822 39800
rect 17037 39797 17049 39800
rect 17083 39797 17095 39831
rect 17037 39791 17095 39797
rect 21726 39788 21732 39840
rect 21784 39828 21790 39840
rect 21821 39831 21879 39837
rect 21821 39828 21833 39831
rect 21784 39800 21833 39828
rect 21784 39788 21790 39800
rect 21821 39797 21833 39800
rect 21867 39797 21879 39831
rect 21821 39791 21879 39797
rect 22554 39788 22560 39840
rect 22612 39828 22618 39840
rect 23017 39831 23075 39837
rect 23017 39828 23029 39831
rect 22612 39800 23029 39828
rect 22612 39788 22618 39800
rect 23017 39797 23029 39800
rect 23063 39828 23075 39831
rect 23290 39828 23296 39840
rect 23063 39800 23296 39828
rect 23063 39797 23075 39800
rect 23017 39791 23075 39797
rect 23290 39788 23296 39800
rect 23348 39788 23354 39840
rect 23658 39788 23664 39840
rect 23716 39828 23722 39840
rect 24320 39828 24348 39936
rect 25225 39933 25237 39936
rect 25271 39964 25283 39967
rect 25685 39967 25743 39973
rect 25685 39964 25697 39967
rect 25271 39936 25697 39964
rect 25271 39933 25283 39936
rect 25225 39927 25283 39933
rect 25685 39933 25697 39936
rect 25731 39933 25743 39967
rect 25685 39927 25743 39933
rect 24397 39899 24455 39905
rect 24397 39865 24409 39899
rect 24443 39896 24455 39899
rect 24486 39896 24492 39908
rect 24443 39868 24492 39896
rect 24443 39865 24455 39868
rect 24397 39859 24455 39865
rect 24486 39856 24492 39868
rect 24544 39856 24550 39908
rect 23716 39800 24348 39828
rect 23716 39788 23722 39800
rect 24578 39788 24584 39840
rect 24636 39828 24642 39840
rect 24673 39831 24731 39837
rect 24673 39828 24685 39831
rect 24636 39800 24685 39828
rect 24636 39788 24642 39800
rect 24673 39797 24685 39800
rect 24719 39797 24731 39831
rect 24673 39791 24731 39797
rect 1104 39738 28888 39760
rect 1104 39686 10982 39738
rect 11034 39686 11046 39738
rect 11098 39686 11110 39738
rect 11162 39686 11174 39738
rect 11226 39686 20982 39738
rect 21034 39686 21046 39738
rect 21098 39686 21110 39738
rect 21162 39686 21174 39738
rect 21226 39686 28888 39738
rect 1104 39664 28888 39686
rect 1673 39627 1731 39633
rect 1673 39593 1685 39627
rect 1719 39624 1731 39627
rect 1762 39624 1768 39636
rect 1719 39596 1768 39624
rect 1719 39593 1731 39596
rect 1673 39587 1731 39593
rect 1762 39584 1768 39596
rect 1820 39584 1826 39636
rect 10502 39624 10508 39636
rect 10463 39596 10508 39624
rect 10502 39584 10508 39596
rect 10560 39584 10566 39636
rect 16577 39627 16635 39633
rect 16577 39593 16589 39627
rect 16623 39624 16635 39627
rect 16850 39624 16856 39636
rect 16623 39596 16856 39624
rect 16623 39593 16635 39596
rect 16577 39587 16635 39593
rect 16850 39584 16856 39596
rect 16908 39624 16914 39636
rect 17310 39624 17316 39636
rect 16908 39596 17316 39624
rect 16908 39584 16914 39596
rect 17310 39584 17316 39596
rect 17368 39584 17374 39636
rect 19426 39624 19432 39636
rect 19387 39596 19432 39624
rect 19426 39584 19432 39596
rect 19484 39584 19490 39636
rect 21542 39584 21548 39636
rect 21600 39624 21606 39636
rect 21821 39627 21879 39633
rect 21821 39624 21833 39627
rect 21600 39596 21833 39624
rect 21600 39584 21606 39596
rect 21821 39593 21833 39596
rect 21867 39593 21879 39627
rect 21821 39587 21879 39593
rect 22186 39584 22192 39636
rect 22244 39624 22250 39636
rect 22373 39627 22431 39633
rect 22373 39624 22385 39627
rect 22244 39596 22385 39624
rect 22244 39584 22250 39596
rect 22373 39593 22385 39596
rect 22419 39593 22431 39627
rect 24486 39624 24492 39636
rect 24447 39596 24492 39624
rect 22373 39587 22431 39593
rect 24486 39584 24492 39596
rect 24544 39584 24550 39636
rect 24670 39584 24676 39636
rect 24728 39624 24734 39636
rect 24765 39627 24823 39633
rect 24765 39624 24777 39627
rect 24728 39596 24777 39624
rect 24728 39584 24734 39596
rect 24765 39593 24777 39596
rect 24811 39593 24823 39627
rect 24765 39587 24823 39593
rect 11149 39559 11207 39565
rect 11149 39525 11161 39559
rect 11195 39556 11207 39559
rect 12158 39556 12164 39568
rect 11195 39528 12164 39556
rect 11195 39525 11207 39528
rect 11149 39519 11207 39525
rect 12158 39516 12164 39528
rect 12216 39516 12222 39568
rect 21910 39556 21916 39568
rect 21560 39528 21916 39556
rect 21560 39500 21588 39528
rect 21910 39516 21916 39528
rect 21968 39516 21974 39568
rect 9493 39491 9551 39497
rect 9493 39457 9505 39491
rect 9539 39488 9551 39491
rect 11514 39488 11520 39500
rect 9539 39460 11520 39488
rect 9539 39457 9551 39460
rect 9493 39451 9551 39457
rect 11514 39448 11520 39460
rect 11572 39488 11578 39500
rect 11609 39491 11667 39497
rect 11609 39488 11621 39491
rect 11572 39460 11621 39488
rect 11572 39448 11578 39460
rect 11609 39457 11621 39460
rect 11655 39457 11667 39491
rect 11790 39488 11796 39500
rect 11751 39460 11796 39488
rect 11609 39451 11667 39457
rect 11790 39448 11796 39460
rect 11848 39448 11854 39500
rect 11977 39491 12035 39497
rect 11977 39457 11989 39491
rect 12023 39457 12035 39491
rect 11977 39451 12035 39457
rect 12897 39491 12955 39497
rect 12897 39457 12909 39491
rect 12943 39457 12955 39491
rect 12897 39451 12955 39457
rect 10870 39380 10876 39432
rect 10928 39420 10934 39432
rect 11992 39420 12020 39451
rect 10928 39392 12020 39420
rect 12253 39423 12311 39429
rect 10928 39380 10934 39392
rect 12253 39389 12265 39423
rect 12299 39389 12311 39423
rect 12253 39383 12311 39389
rect 9125 39355 9183 39361
rect 9125 39321 9137 39355
rect 9171 39352 9183 39355
rect 12268 39352 12296 39383
rect 12342 39380 12348 39432
rect 12400 39420 12406 39432
rect 12529 39423 12587 39429
rect 12529 39420 12541 39423
rect 12400 39392 12541 39420
rect 12400 39380 12406 39392
rect 12529 39389 12541 39392
rect 12575 39389 12587 39423
rect 12912 39420 12940 39451
rect 12986 39448 12992 39500
rect 13044 39488 13050 39500
rect 13538 39488 13544 39500
rect 13044 39460 13089 39488
rect 13499 39460 13544 39488
rect 13044 39448 13050 39460
rect 13538 39448 13544 39460
rect 13596 39448 13602 39500
rect 13722 39488 13728 39500
rect 13683 39460 13728 39488
rect 13722 39448 13728 39460
rect 13780 39488 13786 39500
rect 14737 39491 14795 39497
rect 14737 39488 14749 39491
rect 13780 39460 14749 39488
rect 13780 39448 13786 39460
rect 14737 39457 14749 39460
rect 14783 39457 14795 39491
rect 15286 39488 15292 39500
rect 15247 39460 15292 39488
rect 14737 39451 14795 39457
rect 15286 39448 15292 39460
rect 15344 39448 15350 39500
rect 16758 39488 16764 39500
rect 16719 39460 16764 39488
rect 16758 39448 16764 39460
rect 16816 39448 16822 39500
rect 21542 39488 21548 39500
rect 21455 39460 21548 39488
rect 21542 39448 21548 39460
rect 21600 39448 21606 39500
rect 21726 39488 21732 39500
rect 21687 39460 21732 39488
rect 21726 39448 21732 39460
rect 21784 39448 21790 39500
rect 23569 39491 23627 39497
rect 23569 39457 23581 39491
rect 23615 39488 23627 39491
rect 23658 39488 23664 39500
rect 23615 39460 23664 39488
rect 23615 39457 23627 39460
rect 23569 39451 23627 39457
rect 23658 39448 23664 39460
rect 23716 39448 23722 39500
rect 24578 39488 24584 39500
rect 24044 39460 24584 39488
rect 14090 39420 14096 39432
rect 12912 39392 14096 39420
rect 12529 39383 12587 39389
rect 14090 39380 14096 39392
rect 14148 39380 14154 39432
rect 16666 39420 16672 39432
rect 16579 39392 16672 39420
rect 16666 39380 16672 39392
rect 16724 39420 16730 39432
rect 17034 39420 17040 39432
rect 16724 39392 17040 39420
rect 16724 39380 16730 39392
rect 17034 39380 17040 39392
rect 17092 39380 17098 39432
rect 17218 39380 17224 39432
rect 17276 39420 17282 39432
rect 17589 39423 17647 39429
rect 17589 39420 17601 39423
rect 17276 39392 17601 39420
rect 17276 39380 17282 39392
rect 17589 39389 17601 39392
rect 17635 39420 17647 39423
rect 18046 39420 18052 39432
rect 17635 39392 18052 39420
rect 17635 39389 17647 39392
rect 17589 39383 17647 39389
rect 18046 39380 18052 39392
rect 18104 39380 18110 39432
rect 18322 39420 18328 39432
rect 18283 39392 18328 39420
rect 18322 39380 18328 39392
rect 18380 39380 18386 39432
rect 13078 39352 13084 39364
rect 9171 39324 13084 39352
rect 9171 39321 9183 39324
rect 9125 39315 9183 39321
rect 13078 39312 13084 39324
rect 13136 39312 13142 39364
rect 10042 39284 10048 39296
rect 10003 39256 10048 39284
rect 10042 39244 10048 39256
rect 10100 39244 10106 39296
rect 10778 39284 10784 39296
rect 10739 39256 10784 39284
rect 10778 39244 10784 39256
rect 10836 39244 10842 39296
rect 11974 39244 11980 39296
rect 12032 39284 12038 39296
rect 12158 39284 12164 39296
rect 12032 39256 12164 39284
rect 12032 39244 12038 39256
rect 12158 39244 12164 39256
rect 12216 39284 12222 39296
rect 12713 39287 12771 39293
rect 12713 39284 12725 39287
rect 12216 39256 12725 39284
rect 12216 39244 12222 39256
rect 12713 39253 12725 39256
rect 12759 39253 12771 39287
rect 12713 39247 12771 39253
rect 12802 39244 12808 39296
rect 12860 39284 12866 39296
rect 13173 39287 13231 39293
rect 13173 39284 13185 39287
rect 12860 39256 13185 39284
rect 12860 39244 12866 39256
rect 13173 39253 13185 39256
rect 13219 39253 13231 39287
rect 13173 39247 13231 39253
rect 13814 39244 13820 39296
rect 13872 39284 13878 39296
rect 14369 39287 14427 39293
rect 14369 39284 14381 39287
rect 13872 39256 14381 39284
rect 13872 39244 13878 39256
rect 14369 39253 14381 39256
rect 14415 39253 14427 39287
rect 14369 39247 14427 39253
rect 15010 39244 15016 39296
rect 15068 39284 15074 39296
rect 15473 39287 15531 39293
rect 15473 39284 15485 39287
rect 15068 39256 15485 39284
rect 15068 39244 15074 39256
rect 15473 39253 15485 39256
rect 15519 39253 15531 39287
rect 15746 39284 15752 39296
rect 15707 39256 15752 39284
rect 15473 39247 15531 39253
rect 15746 39244 15752 39256
rect 15804 39244 15810 39296
rect 16209 39287 16267 39293
rect 16209 39253 16221 39287
rect 16255 39284 16267 39287
rect 16390 39284 16396 39296
rect 16255 39256 16396 39284
rect 16255 39253 16267 39256
rect 16209 39247 16267 39253
rect 16390 39244 16396 39256
rect 16448 39244 16454 39296
rect 16574 39244 16580 39296
rect 16632 39284 16638 39296
rect 16945 39287 17003 39293
rect 16945 39284 16957 39287
rect 16632 39256 16957 39284
rect 16632 39244 16638 39256
rect 16945 39253 16957 39256
rect 16991 39253 17003 39287
rect 16945 39247 17003 39253
rect 21453 39287 21511 39293
rect 21453 39253 21465 39287
rect 21499 39284 21511 39287
rect 22002 39284 22008 39296
rect 21499 39256 22008 39284
rect 21499 39253 21511 39256
rect 21453 39247 21511 39253
rect 22002 39244 22008 39256
rect 22060 39244 22066 39296
rect 23474 39244 23480 39296
rect 23532 39284 23538 39296
rect 24044 39293 24072 39460
rect 24578 39448 24584 39460
rect 24636 39448 24642 39500
rect 23753 39287 23811 39293
rect 23753 39284 23765 39287
rect 23532 39256 23765 39284
rect 23532 39244 23538 39256
rect 23753 39253 23765 39256
rect 23799 39284 23811 39287
rect 24029 39287 24087 39293
rect 24029 39284 24041 39287
rect 23799 39256 24041 39284
rect 23799 39253 23811 39256
rect 23753 39247 23811 39253
rect 24029 39253 24041 39256
rect 24075 39253 24087 39287
rect 24029 39247 24087 39253
rect 1104 39194 28888 39216
rect 1104 39142 5982 39194
rect 6034 39142 6046 39194
rect 6098 39142 6110 39194
rect 6162 39142 6174 39194
rect 6226 39142 15982 39194
rect 16034 39142 16046 39194
rect 16098 39142 16110 39194
rect 16162 39142 16174 39194
rect 16226 39142 25982 39194
rect 26034 39142 26046 39194
rect 26098 39142 26110 39194
rect 26162 39142 26174 39194
rect 26226 39142 28888 39194
rect 1104 39120 28888 39142
rect 3145 39083 3203 39089
rect 3145 39049 3157 39083
rect 3191 39080 3203 39083
rect 3326 39080 3332 39092
rect 3191 39052 3332 39080
rect 3191 39049 3203 39052
rect 3145 39043 3203 39049
rect 3326 39040 3332 39052
rect 3384 39040 3390 39092
rect 12434 39040 12440 39092
rect 12492 39080 12498 39092
rect 12897 39083 12955 39089
rect 12897 39080 12909 39083
rect 12492 39052 12909 39080
rect 12492 39040 12498 39052
rect 12897 39049 12909 39052
rect 12943 39049 12955 39083
rect 12897 39043 12955 39049
rect 14090 39040 14096 39092
rect 14148 39080 14154 39092
rect 15197 39083 15255 39089
rect 15197 39080 15209 39083
rect 14148 39052 15209 39080
rect 14148 39040 14154 39052
rect 15197 39049 15209 39052
rect 15243 39049 15255 39083
rect 15197 39043 15255 39049
rect 16758 39040 16764 39092
rect 16816 39080 16822 39092
rect 17037 39083 17095 39089
rect 17037 39080 17049 39083
rect 16816 39052 17049 39080
rect 16816 39040 16822 39052
rect 17037 39049 17049 39052
rect 17083 39049 17095 39083
rect 17037 39043 17095 39049
rect 18322 39040 18328 39092
rect 18380 39080 18386 39092
rect 19429 39083 19487 39089
rect 19429 39080 19441 39083
rect 18380 39052 19441 39080
rect 18380 39040 18386 39052
rect 19429 39049 19441 39052
rect 19475 39049 19487 39083
rect 19429 39043 19487 39049
rect 21177 39083 21235 39089
rect 21177 39049 21189 39083
rect 21223 39080 21235 39083
rect 21726 39080 21732 39092
rect 21223 39052 21732 39080
rect 21223 39049 21235 39052
rect 21177 39043 21235 39049
rect 21726 39040 21732 39052
rect 21784 39040 21790 39092
rect 23658 39040 23664 39092
rect 23716 39080 23722 39092
rect 23845 39083 23903 39089
rect 23845 39080 23857 39083
rect 23716 39052 23857 39080
rect 23716 39040 23722 39052
rect 23845 39049 23857 39052
rect 23891 39049 23903 39083
rect 23845 39043 23903 39049
rect 24486 39040 24492 39092
rect 24544 39080 24550 39092
rect 27525 39083 27583 39089
rect 27525 39080 27537 39083
rect 24544 39052 27537 39080
rect 24544 39040 24550 39052
rect 27525 39049 27537 39052
rect 27571 39049 27583 39083
rect 27525 39043 27583 39049
rect 10413 39015 10471 39021
rect 10413 39012 10425 39015
rect 9600 38984 10425 39012
rect 1486 38904 1492 38956
rect 1544 38944 1550 38956
rect 1581 38947 1639 38953
rect 1581 38944 1593 38947
rect 1544 38916 1593 38944
rect 1544 38904 1550 38916
rect 1581 38913 1593 38916
rect 1627 38944 1639 38947
rect 1762 38944 1768 38956
rect 1627 38916 1768 38944
rect 1627 38913 1639 38916
rect 1581 38907 1639 38913
rect 1762 38904 1768 38916
rect 1820 38904 1826 38956
rect 1670 38836 1676 38888
rect 1728 38876 1734 38888
rect 1857 38879 1915 38885
rect 1857 38876 1869 38879
rect 1728 38848 1869 38876
rect 1728 38836 1734 38848
rect 1857 38845 1869 38848
rect 1903 38845 1915 38879
rect 1857 38839 1915 38845
rect 8846 38836 8852 38888
rect 8904 38876 8910 38888
rect 9600 38885 9628 38984
rect 10413 38981 10425 38984
rect 10459 38981 10471 39015
rect 21542 39012 21548 39024
rect 21503 38984 21548 39012
rect 10413 38975 10471 38981
rect 21542 38972 21548 38984
rect 21600 39012 21606 39024
rect 21637 39015 21695 39021
rect 21637 39012 21649 39015
rect 21600 38984 21649 39012
rect 21600 38972 21606 38984
rect 21637 38981 21649 38984
rect 21683 39012 21695 39015
rect 21821 39015 21879 39021
rect 21821 39012 21833 39015
rect 21683 38984 21833 39012
rect 21683 38981 21695 38984
rect 21637 38975 21695 38981
rect 21821 38981 21833 38984
rect 21867 38981 21879 39015
rect 21821 38975 21879 38981
rect 10134 38944 10140 38956
rect 10095 38916 10140 38944
rect 10134 38904 10140 38916
rect 10192 38904 10198 38956
rect 11517 38947 11575 38953
rect 11517 38913 11529 38947
rect 11563 38944 11575 38947
rect 15286 38944 15292 38956
rect 11563 38916 12664 38944
rect 11563 38913 11575 38916
rect 11517 38907 11575 38913
rect 12636 38888 12664 38916
rect 14016 38916 15292 38944
rect 9585 38879 9643 38885
rect 9585 38876 9597 38879
rect 8904 38848 9597 38876
rect 8904 38836 8910 38848
rect 9585 38845 9597 38848
rect 9631 38845 9643 38879
rect 9585 38839 9643 38845
rect 9677 38879 9735 38885
rect 9677 38845 9689 38879
rect 9723 38876 9735 38879
rect 11149 38879 11207 38885
rect 9723 38848 9904 38876
rect 9723 38845 9735 38848
rect 9677 38839 9735 38845
rect 9125 38811 9183 38817
rect 9125 38777 9137 38811
rect 9171 38808 9183 38811
rect 9766 38808 9772 38820
rect 9171 38780 9772 38808
rect 9171 38777 9183 38780
rect 9125 38771 9183 38777
rect 9766 38768 9772 38780
rect 9824 38768 9830 38820
rect 8757 38743 8815 38749
rect 8757 38709 8769 38743
rect 8803 38740 8815 38743
rect 9306 38740 9312 38752
rect 8803 38712 9312 38740
rect 8803 38709 8815 38712
rect 8757 38703 8815 38709
rect 9306 38700 9312 38712
rect 9364 38700 9370 38752
rect 9490 38740 9496 38752
rect 9451 38712 9496 38740
rect 9490 38700 9496 38712
rect 9548 38740 9554 38752
rect 9876 38740 9904 38848
rect 11149 38845 11161 38879
rect 11195 38876 11207 38879
rect 11330 38876 11336 38888
rect 11195 38848 11336 38876
rect 11195 38845 11207 38848
rect 11149 38839 11207 38845
rect 11330 38836 11336 38848
rect 11388 38836 11394 38888
rect 12158 38836 12164 38888
rect 12216 38876 12222 38888
rect 12437 38879 12495 38885
rect 12437 38876 12449 38879
rect 12216 38848 12449 38876
rect 12216 38836 12222 38848
rect 12437 38845 12449 38848
rect 12483 38845 12495 38879
rect 12618 38876 12624 38888
rect 12579 38848 12624 38876
rect 12437 38839 12495 38845
rect 12618 38836 12624 38848
rect 12676 38836 12682 38888
rect 12710 38836 12716 38888
rect 12768 38876 12774 38888
rect 12894 38876 12900 38888
rect 12768 38848 12900 38876
rect 12768 38836 12774 38848
rect 12894 38836 12900 38848
rect 12952 38836 12958 38888
rect 13538 38876 13544 38888
rect 13499 38848 13544 38876
rect 13538 38836 13544 38848
rect 13596 38836 13602 38888
rect 14016 38885 14044 38916
rect 15286 38904 15292 38916
rect 15344 38944 15350 38956
rect 15654 38944 15660 38956
rect 15344 38916 15660 38944
rect 15344 38904 15350 38916
rect 15654 38904 15660 38916
rect 15712 38904 15718 38956
rect 17770 38904 17776 38956
rect 17828 38944 17834 38956
rect 17865 38947 17923 38953
rect 17865 38944 17877 38947
rect 17828 38916 17877 38944
rect 17828 38904 17834 38916
rect 17865 38913 17877 38916
rect 17911 38944 17923 38947
rect 22370 38944 22376 38956
rect 17911 38916 18368 38944
rect 17911 38913 17923 38916
rect 17865 38907 17923 38913
rect 13909 38879 13967 38885
rect 13909 38845 13921 38879
rect 13955 38876 13967 38879
rect 14001 38879 14059 38885
rect 14001 38876 14013 38879
rect 13955 38848 14013 38876
rect 13955 38845 13967 38848
rect 13909 38839 13967 38845
rect 14001 38845 14013 38848
rect 14047 38845 14059 38879
rect 14001 38839 14059 38845
rect 14185 38879 14243 38885
rect 14185 38845 14197 38879
rect 14231 38845 14243 38879
rect 14185 38839 14243 38845
rect 10965 38811 11023 38817
rect 10965 38777 10977 38811
rect 11011 38808 11023 38811
rect 11793 38811 11851 38817
rect 11793 38808 11805 38811
rect 11011 38780 11805 38808
rect 11011 38777 11023 38780
rect 10965 38771 11023 38777
rect 11793 38777 11805 38780
rect 11839 38808 11851 38811
rect 13556 38808 13584 38836
rect 11839 38780 13584 38808
rect 11839 38777 11851 38780
rect 11793 38771 11851 38777
rect 14200 38752 14228 38839
rect 14918 38836 14924 38888
rect 14976 38876 14982 38888
rect 15381 38879 15439 38885
rect 15381 38876 15393 38879
rect 14976 38848 15393 38876
rect 14976 38836 14982 38848
rect 15381 38845 15393 38848
rect 15427 38876 15439 38879
rect 16390 38876 16396 38888
rect 15427 38848 16396 38876
rect 15427 38845 15439 38848
rect 15381 38839 15439 38845
rect 16390 38836 16396 38848
rect 16448 38836 16454 38888
rect 17497 38879 17555 38885
rect 17497 38845 17509 38879
rect 17543 38876 17555 38879
rect 18046 38876 18052 38888
rect 17543 38848 18052 38876
rect 17543 38845 17555 38848
rect 17497 38839 17555 38845
rect 18046 38836 18052 38848
rect 18104 38836 18110 38888
rect 18340 38885 18368 38916
rect 22020 38916 22376 38944
rect 18325 38879 18383 38885
rect 18325 38845 18337 38879
rect 18371 38876 18383 38879
rect 18414 38876 18420 38888
rect 18371 38848 18420 38876
rect 18371 38845 18383 38848
rect 18325 38839 18383 38845
rect 18414 38836 18420 38848
rect 18472 38836 18478 38888
rect 21174 38836 21180 38888
rect 21232 38876 21238 38888
rect 21542 38876 21548 38888
rect 21232 38848 21548 38876
rect 21232 38836 21238 38848
rect 21542 38836 21548 38848
rect 21600 38836 21606 38888
rect 21910 38836 21916 38888
rect 21968 38876 21974 38888
rect 22020 38885 22048 38916
rect 22370 38904 22376 38916
rect 22428 38944 22434 38956
rect 22833 38947 22891 38953
rect 22833 38944 22845 38947
rect 22428 38916 22845 38944
rect 22428 38904 22434 38916
rect 22833 38913 22845 38916
rect 22879 38913 22891 38947
rect 22833 38907 22891 38913
rect 26053 38947 26111 38953
rect 26053 38913 26065 38947
rect 26099 38944 26111 38947
rect 26099 38916 26464 38944
rect 26099 38913 26111 38916
rect 26053 38907 26111 38913
rect 26436 38888 26464 38916
rect 22005 38879 22063 38885
rect 22005 38876 22017 38879
rect 21968 38848 22017 38876
rect 21968 38836 21974 38848
rect 22005 38845 22017 38848
rect 22051 38845 22063 38879
rect 22005 38839 22063 38845
rect 22097 38879 22155 38885
rect 22097 38845 22109 38879
rect 22143 38845 22155 38879
rect 22554 38876 22560 38888
rect 22515 38848 22560 38876
rect 22097 38839 22155 38845
rect 14553 38811 14611 38817
rect 14553 38777 14565 38811
rect 14599 38808 14611 38811
rect 15102 38808 15108 38820
rect 14599 38780 15108 38808
rect 14599 38777 14611 38780
rect 14553 38771 14611 38777
rect 15102 38768 15108 38780
rect 15160 38768 15166 38820
rect 15286 38768 15292 38820
rect 15344 38808 15350 38820
rect 16209 38811 16267 38817
rect 16209 38808 16221 38811
rect 15344 38780 16221 38808
rect 15344 38768 15350 38780
rect 16209 38777 16221 38780
rect 16255 38777 16267 38811
rect 16209 38771 16267 38777
rect 21637 38811 21695 38817
rect 21637 38777 21649 38811
rect 21683 38808 21695 38811
rect 22112 38808 22140 38839
rect 22554 38836 22560 38848
rect 22612 38836 22618 38888
rect 25774 38836 25780 38888
rect 25832 38876 25838 38888
rect 26142 38876 26148 38888
rect 25832 38848 26148 38876
rect 25832 38836 25838 38848
rect 26142 38836 26148 38848
rect 26200 38836 26206 38888
rect 26418 38876 26424 38888
rect 26379 38848 26424 38876
rect 26418 38836 26424 38848
rect 26476 38836 26482 38888
rect 21683 38780 22140 38808
rect 21683 38777 21695 38780
rect 21637 38771 21695 38777
rect 9548 38712 9904 38740
rect 9548 38700 9554 38712
rect 10042 38700 10048 38752
rect 10100 38740 10106 38752
rect 10781 38743 10839 38749
rect 10781 38740 10793 38743
rect 10100 38712 10793 38740
rect 10100 38700 10106 38712
rect 10781 38709 10793 38712
rect 10827 38740 10839 38743
rect 10870 38740 10876 38752
rect 10827 38712 10876 38740
rect 10827 38709 10839 38712
rect 10781 38703 10839 38709
rect 10870 38700 10876 38712
rect 10928 38700 10934 38752
rect 12158 38740 12164 38752
rect 12119 38712 12164 38740
rect 12158 38700 12164 38712
rect 12216 38700 12222 38752
rect 14182 38700 14188 38752
rect 14240 38740 14246 38752
rect 14829 38743 14887 38749
rect 14829 38740 14841 38743
rect 14240 38712 14841 38740
rect 14240 38700 14246 38712
rect 14829 38709 14841 38712
rect 14875 38709 14887 38743
rect 14829 38703 14887 38709
rect 15470 38700 15476 38752
rect 15528 38740 15534 38752
rect 15565 38743 15623 38749
rect 15565 38740 15577 38743
rect 15528 38712 15577 38740
rect 15528 38700 15534 38712
rect 15565 38709 15577 38712
rect 15611 38709 15623 38743
rect 15565 38703 15623 38709
rect 15654 38700 15660 38752
rect 15712 38740 15718 38752
rect 15841 38743 15899 38749
rect 15841 38740 15853 38743
rect 15712 38712 15853 38740
rect 15712 38700 15718 38712
rect 15841 38709 15853 38712
rect 15887 38709 15899 38743
rect 15841 38703 15899 38709
rect 16761 38743 16819 38749
rect 16761 38709 16773 38743
rect 16807 38740 16819 38743
rect 17034 38740 17040 38752
rect 16807 38712 17040 38740
rect 16807 38709 16819 38712
rect 16761 38703 16819 38709
rect 17034 38700 17040 38712
rect 17092 38700 17098 38752
rect 23474 38700 23480 38752
rect 23532 38740 23538 38752
rect 24581 38743 24639 38749
rect 24581 38740 24593 38743
rect 23532 38712 24593 38740
rect 23532 38700 23538 38712
rect 24581 38709 24593 38712
rect 24627 38709 24639 38743
rect 24581 38703 24639 38709
rect 1104 38650 28888 38672
rect 1104 38598 10982 38650
rect 11034 38598 11046 38650
rect 11098 38598 11110 38650
rect 11162 38598 11174 38650
rect 11226 38598 20982 38650
rect 21034 38598 21046 38650
rect 21098 38598 21110 38650
rect 21162 38598 21174 38650
rect 21226 38598 28888 38650
rect 1104 38576 28888 38598
rect 8757 38539 8815 38545
rect 8757 38505 8769 38539
rect 8803 38536 8815 38539
rect 9493 38539 9551 38545
rect 9493 38536 9505 38539
rect 8803 38508 9505 38536
rect 8803 38505 8815 38508
rect 8757 38499 8815 38505
rect 9493 38505 9505 38508
rect 9539 38536 9551 38539
rect 9539 38508 10548 38536
rect 9539 38505 9551 38508
rect 9493 38499 9551 38505
rect 8113 38471 8171 38477
rect 8113 38437 8125 38471
rect 8159 38468 8171 38471
rect 9306 38468 9312 38480
rect 8159 38440 9312 38468
rect 8159 38437 8171 38440
rect 8113 38431 8171 38437
rect 9306 38428 9312 38440
rect 9364 38428 9370 38480
rect 9674 38468 9680 38480
rect 9635 38440 9680 38468
rect 9674 38428 9680 38440
rect 9732 38428 9738 38480
rect 10520 38412 10548 38508
rect 11330 38496 11336 38548
rect 11388 38536 11394 38548
rect 15565 38539 15623 38545
rect 15565 38536 15577 38539
rect 11388 38508 15577 38536
rect 11388 38496 11394 38508
rect 15565 38505 15577 38508
rect 15611 38505 15623 38539
rect 16482 38536 16488 38548
rect 16443 38508 16488 38536
rect 15565 38499 15623 38505
rect 16482 38496 16488 38508
rect 16540 38496 16546 38548
rect 18141 38539 18199 38545
rect 18141 38505 18153 38539
rect 18187 38536 18199 38539
rect 18322 38536 18328 38548
rect 18187 38508 18328 38536
rect 18187 38505 18199 38508
rect 18141 38499 18199 38505
rect 18322 38496 18328 38508
rect 18380 38496 18386 38548
rect 20257 38539 20315 38545
rect 20257 38505 20269 38539
rect 20303 38536 20315 38539
rect 20714 38536 20720 38548
rect 20303 38508 20720 38536
rect 20303 38505 20315 38508
rect 20257 38499 20315 38505
rect 20714 38496 20720 38508
rect 20772 38496 20778 38548
rect 26142 38536 26148 38548
rect 26103 38508 26148 38536
rect 26142 38496 26148 38508
rect 26200 38496 26206 38548
rect 12069 38471 12127 38477
rect 12069 38437 12081 38471
rect 12115 38468 12127 38471
rect 12158 38468 12164 38480
rect 12115 38440 12164 38468
rect 12115 38437 12127 38440
rect 12069 38431 12127 38437
rect 12158 38428 12164 38440
rect 12216 38428 12222 38480
rect 15102 38428 15108 38480
rect 15160 38468 15166 38480
rect 15160 38440 16344 38468
rect 15160 38428 15166 38440
rect 8570 38400 8576 38412
rect 8531 38372 8576 38400
rect 8570 38360 8576 38372
rect 8628 38360 8634 38412
rect 8754 38360 8760 38412
rect 8812 38400 8818 38412
rect 9398 38400 9404 38412
rect 8812 38372 9404 38400
rect 8812 38360 8818 38372
rect 9398 38360 9404 38372
rect 9456 38360 9462 38412
rect 10226 38360 10232 38412
rect 10284 38400 10290 38412
rect 10321 38403 10379 38409
rect 10321 38400 10333 38403
rect 10284 38372 10333 38400
rect 10284 38360 10290 38372
rect 10321 38369 10333 38372
rect 10367 38369 10379 38403
rect 10321 38363 10379 38369
rect 10502 38360 10508 38412
rect 10560 38400 10566 38412
rect 10689 38403 10747 38409
rect 10689 38400 10701 38403
rect 10560 38372 10701 38400
rect 10560 38360 10566 38372
rect 10689 38369 10701 38372
rect 10735 38369 10747 38403
rect 10870 38400 10876 38412
rect 10831 38372 10876 38400
rect 10689 38363 10747 38369
rect 10870 38360 10876 38372
rect 10928 38360 10934 38412
rect 12802 38360 12808 38412
rect 12860 38400 12866 38412
rect 13173 38403 13231 38409
rect 13173 38400 13185 38403
rect 12860 38372 13185 38400
rect 12860 38360 12866 38372
rect 13173 38369 13185 38372
rect 13219 38400 13231 38403
rect 13538 38400 13544 38412
rect 13219 38372 13544 38400
rect 13219 38369 13231 38372
rect 13173 38363 13231 38369
rect 13538 38360 13544 38372
rect 13596 38360 13602 38412
rect 14185 38403 14243 38409
rect 14185 38369 14197 38403
rect 14231 38400 14243 38403
rect 14642 38400 14648 38412
rect 14231 38372 14648 38400
rect 14231 38369 14243 38372
rect 14185 38363 14243 38369
rect 14642 38360 14648 38372
rect 14700 38360 14706 38412
rect 16316 38409 16344 38440
rect 16390 38428 16396 38480
rect 16448 38468 16454 38480
rect 16448 38440 17264 38468
rect 16448 38428 16454 38440
rect 15289 38403 15347 38409
rect 15289 38369 15301 38403
rect 15335 38369 15347 38403
rect 15289 38363 15347 38369
rect 16301 38403 16359 38409
rect 16301 38369 16313 38403
rect 16347 38400 16359 38403
rect 16574 38400 16580 38412
rect 16347 38372 16580 38400
rect 16347 38369 16359 38372
rect 16301 38363 16359 38369
rect 8481 38335 8539 38341
rect 8481 38301 8493 38335
rect 8527 38332 8539 38335
rect 9674 38332 9680 38344
rect 8527 38304 9680 38332
rect 8527 38301 8539 38304
rect 8481 38295 8539 38301
rect 9674 38292 9680 38304
rect 9732 38292 9738 38344
rect 10413 38335 10471 38341
rect 10413 38301 10425 38335
rect 10459 38332 10471 38335
rect 10594 38332 10600 38344
rect 10459 38304 10600 38332
rect 10459 38301 10471 38304
rect 10413 38295 10471 38301
rect 10594 38292 10600 38304
rect 10652 38292 10658 38344
rect 12526 38332 12532 38344
rect 12487 38304 12532 38332
rect 12526 38292 12532 38304
rect 12584 38292 12590 38344
rect 15010 38292 15016 38344
rect 15068 38292 15074 38344
rect 15304 38332 15332 38363
rect 16574 38360 16580 38372
rect 16632 38360 16638 38412
rect 16482 38332 16488 38344
rect 15304 38304 16488 38332
rect 16482 38292 16488 38304
rect 16540 38332 16546 38344
rect 16850 38332 16856 38344
rect 16540 38304 16856 38332
rect 16540 38292 16546 38304
rect 16850 38292 16856 38304
rect 16908 38292 16914 38344
rect 1394 38224 1400 38276
rect 1452 38264 1458 38276
rect 1854 38264 1860 38276
rect 1452 38236 1860 38264
rect 1452 38224 1458 38236
rect 1854 38224 1860 38236
rect 1912 38264 1918 38276
rect 1949 38267 2007 38273
rect 1949 38264 1961 38267
rect 1912 38236 1961 38264
rect 1912 38224 1918 38236
rect 1949 38233 1961 38236
rect 1995 38233 2007 38267
rect 1949 38227 2007 38233
rect 8294 38224 8300 38276
rect 8352 38264 8358 38276
rect 9033 38267 9091 38273
rect 9033 38264 9045 38267
rect 8352 38236 9045 38264
rect 8352 38224 8358 38236
rect 9033 38233 9045 38236
rect 9079 38233 9091 38267
rect 9033 38227 9091 38233
rect 11241 38267 11299 38273
rect 11241 38233 11253 38267
rect 11287 38264 11299 38267
rect 11422 38264 11428 38276
rect 11287 38236 11428 38264
rect 11287 38233 11299 38236
rect 11241 38227 11299 38233
rect 11422 38224 11428 38236
rect 11480 38264 11486 38276
rect 12342 38264 12348 38276
rect 11480 38236 12348 38264
rect 11480 38224 11486 38236
rect 12342 38224 12348 38236
rect 12400 38224 12406 38276
rect 14093 38267 14151 38273
rect 14093 38233 14105 38267
rect 14139 38264 14151 38267
rect 14458 38264 14464 38276
rect 14139 38236 14464 38264
rect 14139 38233 14151 38236
rect 14093 38227 14151 38233
rect 14458 38224 14464 38236
rect 14516 38264 14522 38276
rect 15028 38264 15056 38292
rect 14516 38236 15056 38264
rect 14516 38224 14522 38236
rect 15102 38224 15108 38276
rect 15160 38264 15166 38276
rect 15746 38264 15752 38276
rect 15160 38236 15752 38264
rect 15160 38224 15166 38236
rect 15746 38224 15752 38236
rect 15804 38224 15810 38276
rect 15841 38267 15899 38273
rect 15841 38233 15853 38267
rect 15887 38264 15899 38267
rect 16298 38264 16304 38276
rect 15887 38236 16304 38264
rect 15887 38233 15899 38236
rect 15841 38227 15899 38233
rect 16298 38224 16304 38236
rect 16356 38224 16362 38276
rect 1578 38196 1584 38208
rect 1539 38168 1584 38196
rect 1578 38156 1584 38168
rect 1636 38156 1642 38208
rect 11514 38196 11520 38208
rect 11475 38168 11520 38196
rect 11514 38156 11520 38168
rect 11572 38156 11578 38208
rect 12437 38199 12495 38205
rect 12437 38165 12449 38199
rect 12483 38196 12495 38199
rect 12894 38196 12900 38208
rect 12483 38168 12900 38196
rect 12483 38165 12495 38168
rect 12437 38159 12495 38165
rect 12894 38156 12900 38168
rect 12952 38156 12958 38208
rect 13354 38156 13360 38208
rect 13412 38196 13418 38208
rect 13541 38199 13599 38205
rect 13541 38196 13553 38199
rect 13412 38168 13553 38196
rect 13412 38156 13418 38168
rect 13541 38165 13553 38168
rect 13587 38165 13599 38199
rect 14366 38196 14372 38208
rect 14327 38168 14372 38196
rect 13541 38159 13599 38165
rect 14366 38156 14372 38168
rect 14424 38156 14430 38208
rect 15010 38196 15016 38208
rect 14971 38168 15016 38196
rect 15010 38156 15016 38168
rect 15068 38156 15074 38208
rect 15378 38156 15384 38208
rect 15436 38196 15442 38208
rect 15473 38199 15531 38205
rect 15473 38196 15485 38199
rect 15436 38168 15485 38196
rect 15436 38156 15442 38168
rect 15473 38165 15485 38168
rect 15519 38165 15531 38199
rect 15473 38159 15531 38165
rect 15565 38199 15623 38205
rect 15565 38165 15577 38199
rect 15611 38196 15623 38199
rect 16209 38199 16267 38205
rect 16209 38196 16221 38199
rect 15611 38168 16221 38196
rect 15611 38165 15623 38168
rect 15565 38159 15623 38165
rect 16209 38165 16221 38168
rect 16255 38196 16267 38199
rect 16390 38196 16396 38208
rect 16255 38168 16396 38196
rect 16255 38165 16267 38168
rect 16209 38159 16267 38165
rect 16390 38156 16396 38168
rect 16448 38156 16454 38208
rect 16758 38196 16764 38208
rect 16719 38168 16764 38196
rect 16758 38156 16764 38168
rect 16816 38156 16822 38208
rect 17236 38205 17264 38440
rect 18046 38428 18052 38480
rect 18104 38468 18110 38480
rect 18417 38471 18475 38477
rect 18417 38468 18429 38471
rect 18104 38440 18429 38468
rect 18104 38428 18110 38440
rect 18417 38437 18429 38440
rect 18463 38437 18475 38471
rect 18417 38431 18475 38437
rect 23658 38400 23664 38412
rect 23619 38372 23664 38400
rect 23658 38360 23664 38372
rect 23716 38360 23722 38412
rect 21726 38292 21732 38344
rect 21784 38332 21790 38344
rect 22646 38332 22652 38344
rect 21784 38304 22652 38332
rect 21784 38292 21790 38304
rect 22646 38292 22652 38304
rect 22704 38292 22710 38344
rect 17221 38199 17279 38205
rect 17221 38165 17233 38199
rect 17267 38196 17279 38199
rect 17402 38196 17408 38208
rect 17267 38168 17408 38196
rect 17267 38165 17279 38168
rect 17221 38159 17279 38165
rect 17402 38156 17408 38168
rect 17460 38156 17466 38208
rect 17589 38199 17647 38205
rect 17589 38165 17601 38199
rect 17635 38196 17647 38199
rect 19426 38196 19432 38208
rect 17635 38168 19432 38196
rect 17635 38165 17647 38168
rect 17589 38159 17647 38165
rect 19426 38156 19432 38168
rect 19484 38156 19490 38208
rect 1104 38106 28888 38128
rect 1104 38054 5982 38106
rect 6034 38054 6046 38106
rect 6098 38054 6110 38106
rect 6162 38054 6174 38106
rect 6226 38054 15982 38106
rect 16034 38054 16046 38106
rect 16098 38054 16110 38106
rect 16162 38054 16174 38106
rect 16226 38054 25982 38106
rect 26034 38054 26046 38106
rect 26098 38054 26110 38106
rect 26162 38054 26174 38106
rect 26226 38054 28888 38106
rect 1104 38032 28888 38054
rect 8941 37995 8999 38001
rect 8941 37961 8953 37995
rect 8987 37992 8999 37995
rect 9030 37992 9036 38004
rect 8987 37964 9036 37992
rect 8987 37961 8999 37964
rect 8941 37955 8999 37961
rect 7561 37859 7619 37865
rect 7561 37825 7573 37859
rect 7607 37856 7619 37859
rect 8662 37856 8668 37868
rect 7607 37828 8668 37856
rect 7607 37825 7619 37828
rect 7561 37819 7619 37825
rect 8662 37816 8668 37828
rect 8720 37816 8726 37868
rect 7929 37791 7987 37797
rect 7929 37757 7941 37791
rect 7975 37788 7987 37791
rect 8202 37788 8208 37800
rect 7975 37760 8208 37788
rect 7975 37757 7987 37760
rect 7929 37751 7987 37757
rect 8202 37748 8208 37760
rect 8260 37748 8266 37800
rect 8389 37791 8447 37797
rect 8389 37757 8401 37791
rect 8435 37788 8447 37791
rect 8956 37788 8984 37955
rect 9030 37952 9036 37964
rect 9088 37952 9094 38004
rect 9677 37995 9735 38001
rect 9677 37961 9689 37995
rect 9723 37992 9735 37995
rect 11057 37995 11115 38001
rect 11057 37992 11069 37995
rect 9723 37964 11069 37992
rect 9723 37961 9735 37964
rect 9677 37955 9735 37961
rect 11057 37961 11069 37964
rect 11103 37992 11115 37995
rect 11514 37992 11520 38004
rect 11103 37964 11520 37992
rect 11103 37961 11115 37964
rect 11057 37955 11115 37961
rect 11514 37952 11520 37964
rect 11572 37952 11578 38004
rect 12342 37952 12348 38004
rect 12400 37992 12406 38004
rect 13170 37992 13176 38004
rect 12400 37964 13176 37992
rect 12400 37952 12406 37964
rect 13170 37952 13176 37964
rect 13228 37952 13234 38004
rect 14642 37952 14648 38004
rect 14700 37992 14706 38004
rect 15013 37995 15071 38001
rect 15013 37992 15025 37995
rect 14700 37964 15025 37992
rect 14700 37952 14706 37964
rect 15013 37961 15025 37964
rect 15059 37992 15071 37995
rect 15746 37992 15752 38004
rect 15059 37964 15752 37992
rect 15059 37961 15071 37964
rect 15013 37955 15071 37961
rect 15746 37952 15752 37964
rect 15804 37952 15810 38004
rect 16574 37992 16580 38004
rect 16535 37964 16580 37992
rect 16574 37952 16580 37964
rect 16632 37952 16638 38004
rect 18506 37952 18512 38004
rect 18564 37992 18570 38004
rect 18601 37995 18659 38001
rect 18601 37992 18613 37995
rect 18564 37964 18613 37992
rect 18564 37952 18570 37964
rect 18601 37961 18613 37964
rect 18647 37992 18659 37995
rect 18969 37995 19027 38001
rect 18969 37992 18981 37995
rect 18647 37964 18981 37992
rect 18647 37961 18659 37964
rect 18601 37955 18659 37961
rect 18969 37961 18981 37964
rect 19015 37992 19027 37995
rect 19518 37992 19524 38004
rect 19015 37964 19524 37992
rect 19015 37961 19027 37964
rect 18969 37955 19027 37961
rect 19518 37952 19524 37964
rect 19576 37952 19582 38004
rect 23477 37995 23535 38001
rect 23477 37961 23489 37995
rect 23523 37992 23535 37995
rect 23566 37992 23572 38004
rect 23523 37964 23572 37992
rect 23523 37961 23535 37964
rect 23477 37955 23535 37961
rect 23566 37952 23572 37964
rect 23624 37952 23630 38004
rect 23750 37952 23756 38004
rect 23808 37952 23814 38004
rect 23934 37952 23940 38004
rect 23992 37992 23998 38004
rect 23992 37964 24716 37992
rect 23992 37952 23998 37964
rect 9398 37884 9404 37936
rect 9456 37884 9462 37936
rect 10594 37924 10600 37936
rect 10507 37896 10600 37924
rect 10594 37884 10600 37896
rect 10652 37924 10658 37936
rect 10919 37927 10977 37933
rect 10919 37924 10931 37927
rect 10652 37896 10931 37924
rect 10652 37884 10658 37896
rect 10919 37893 10931 37896
rect 10965 37893 10977 37927
rect 10919 37887 10977 37893
rect 15289 37927 15347 37933
rect 15289 37893 15301 37927
rect 15335 37924 15347 37927
rect 15654 37924 15660 37936
rect 15335 37896 15660 37924
rect 15335 37893 15347 37896
rect 15289 37887 15347 37893
rect 15654 37884 15660 37896
rect 15712 37884 15718 37936
rect 16114 37884 16120 37936
rect 16172 37924 16178 37936
rect 16390 37924 16396 37936
rect 16172 37896 16396 37924
rect 16172 37884 16178 37896
rect 16390 37884 16396 37896
rect 16448 37884 16454 37936
rect 23768 37924 23796 37952
rect 21192 37896 23796 37924
rect 9416 37856 9444 37884
rect 9416 37828 9536 37856
rect 9508 37797 9536 37828
rect 8435 37760 8984 37788
rect 9401 37791 9459 37797
rect 8435 37757 8447 37760
rect 8389 37751 8447 37757
rect 9401 37757 9413 37791
rect 9447 37757 9459 37791
rect 9401 37751 9459 37757
rect 9493 37791 9551 37797
rect 9493 37757 9505 37791
rect 9539 37757 9551 37791
rect 9493 37751 9551 37757
rect 4890 37680 4896 37732
rect 4948 37720 4954 37732
rect 8297 37723 8355 37729
rect 8297 37720 8309 37723
rect 4948 37692 8309 37720
rect 4948 37680 4954 37692
rect 8297 37689 8309 37692
rect 8343 37720 8355 37723
rect 8478 37720 8484 37732
rect 8343 37692 8484 37720
rect 8343 37689 8355 37692
rect 8297 37683 8355 37689
rect 8478 37680 8484 37692
rect 8536 37720 8542 37732
rect 9217 37723 9275 37729
rect 9217 37720 9229 37723
rect 8536 37692 9229 37720
rect 8536 37680 8542 37692
rect 9217 37689 9229 37692
rect 9263 37720 9275 37723
rect 9416 37720 9444 37751
rect 10134 37720 10140 37732
rect 9263 37692 9444 37720
rect 9600 37692 10140 37720
rect 9263 37689 9275 37692
rect 9217 37683 9275 37689
rect 7193 37655 7251 37661
rect 7193 37621 7205 37655
rect 7239 37652 7251 37655
rect 7834 37652 7840 37664
rect 7239 37624 7840 37652
rect 7239 37621 7251 37624
rect 7193 37615 7251 37621
rect 7834 37612 7840 37624
rect 7892 37612 7898 37664
rect 8573 37655 8631 37661
rect 8573 37621 8585 37655
rect 8619 37652 8631 37655
rect 9490 37652 9496 37664
rect 8619 37624 9496 37652
rect 8619 37621 8631 37624
rect 8573 37615 8631 37621
rect 9490 37612 9496 37624
rect 9548 37652 9554 37664
rect 9600 37652 9628 37692
rect 10134 37680 10140 37692
rect 10192 37680 10198 37732
rect 9548 37624 9628 37652
rect 9548 37612 9554 37624
rect 9858 37612 9864 37664
rect 9916 37652 9922 37664
rect 10612 37661 10640 37884
rect 11149 37859 11207 37865
rect 11149 37856 11161 37859
rect 10888 37828 11161 37856
rect 10888 37800 10916 37828
rect 11149 37825 11161 37828
rect 11195 37825 11207 37859
rect 11149 37819 11207 37825
rect 11517 37859 11575 37865
rect 11517 37825 11529 37859
rect 11563 37856 11575 37859
rect 11790 37856 11796 37868
rect 11563 37828 11796 37856
rect 11563 37825 11575 37828
rect 11517 37819 11575 37825
rect 11790 37816 11796 37828
rect 11848 37816 11854 37868
rect 11885 37859 11943 37865
rect 11885 37825 11897 37859
rect 11931 37856 11943 37859
rect 12437 37859 12495 37865
rect 12437 37856 12449 37859
rect 11931 37828 12449 37856
rect 11931 37825 11943 37828
rect 11885 37819 11943 37825
rect 12437 37825 12449 37828
rect 12483 37856 12495 37859
rect 13170 37856 13176 37868
rect 12483 37828 13176 37856
rect 12483 37825 12495 37828
rect 12437 37819 12495 37825
rect 13170 37816 13176 37828
rect 13228 37816 13234 37868
rect 13998 37816 14004 37868
rect 14056 37856 14062 37868
rect 14737 37859 14795 37865
rect 14737 37856 14749 37859
rect 14056 37828 14749 37856
rect 14056 37816 14062 37828
rect 14737 37825 14749 37828
rect 14783 37825 14795 37859
rect 14737 37819 14795 37825
rect 15378 37816 15384 37868
rect 15436 37856 15442 37868
rect 15436 37828 16436 37856
rect 15436 37816 15442 37828
rect 16408 37800 16436 37828
rect 16574 37816 16580 37868
rect 16632 37856 16638 37868
rect 17405 37859 17463 37865
rect 17405 37856 17417 37859
rect 16632 37828 17417 37856
rect 16632 37816 16638 37828
rect 17405 37825 17417 37828
rect 17451 37856 17463 37859
rect 18506 37856 18512 37868
rect 17451 37828 18512 37856
rect 17451 37825 17463 37828
rect 17405 37819 17463 37825
rect 18506 37816 18512 37828
rect 18564 37816 18570 37868
rect 20073 37859 20131 37865
rect 20073 37825 20085 37859
rect 20119 37856 20131 37859
rect 20806 37856 20812 37868
rect 20119 37828 20812 37856
rect 20119 37825 20131 37828
rect 20073 37819 20131 37825
rect 20806 37816 20812 37828
rect 20864 37856 20870 37868
rect 21192 37865 21220 37896
rect 21177 37859 21235 37865
rect 21177 37856 21189 37859
rect 20864 37828 21189 37856
rect 20864 37816 20870 37828
rect 21177 37825 21189 37828
rect 21223 37825 21235 37859
rect 21177 37819 21235 37825
rect 23658 37816 23664 37868
rect 23716 37856 23722 37868
rect 23716 37828 24624 37856
rect 23716 37816 23722 37828
rect 10778 37788 10784 37800
rect 10739 37760 10784 37788
rect 10778 37748 10784 37760
rect 10836 37748 10842 37800
rect 10870 37748 10876 37800
rect 10928 37748 10934 37800
rect 12253 37791 12311 37797
rect 12253 37757 12265 37791
rect 12299 37788 12311 37791
rect 12621 37791 12679 37797
rect 12621 37788 12633 37791
rect 12299 37760 12633 37788
rect 12299 37757 12311 37760
rect 12253 37751 12311 37757
rect 12621 37757 12633 37760
rect 12667 37788 12679 37791
rect 12986 37788 12992 37800
rect 12667 37760 12992 37788
rect 12667 37757 12679 37760
rect 12621 37751 12679 37757
rect 12986 37748 12992 37760
rect 13044 37748 13050 37800
rect 14274 37788 14280 37800
rect 14187 37760 14280 37788
rect 14274 37748 14280 37760
rect 14332 37788 14338 37800
rect 15286 37788 15292 37800
rect 14332 37760 15292 37788
rect 14332 37748 14338 37760
rect 15286 37748 15292 37760
rect 15344 37748 15350 37800
rect 15654 37748 15660 37800
rect 15712 37788 15718 37800
rect 16301 37791 16359 37797
rect 16301 37788 16313 37791
rect 15712 37760 16313 37788
rect 15712 37748 15718 37760
rect 16301 37757 16313 37760
rect 16347 37757 16359 37791
rect 16301 37751 16359 37757
rect 16390 37748 16396 37800
rect 16448 37748 16454 37800
rect 17310 37748 17316 37800
rect 17368 37788 17374 37800
rect 17681 37791 17739 37797
rect 17681 37788 17693 37791
rect 17368 37760 17693 37788
rect 17368 37748 17374 37760
rect 17681 37757 17693 37760
rect 17727 37757 17739 37791
rect 20254 37788 20260 37800
rect 20215 37760 20260 37788
rect 17681 37751 17739 37757
rect 20254 37748 20260 37760
rect 20312 37748 20318 37800
rect 20714 37748 20720 37800
rect 20772 37788 20778 37800
rect 21085 37791 21143 37797
rect 21085 37788 21097 37791
rect 20772 37760 21097 37788
rect 20772 37748 20778 37760
rect 21085 37757 21097 37760
rect 21131 37757 21143 37791
rect 21085 37751 21143 37757
rect 23566 37748 23572 37800
rect 23624 37788 23630 37800
rect 24596 37797 24624 37828
rect 24688 37797 24716 37964
rect 25406 37952 25412 38004
rect 25464 37992 25470 38004
rect 25961 37995 26019 38001
rect 25961 37992 25973 37995
rect 25464 37964 25973 37992
rect 25464 37952 25470 37964
rect 25961 37961 25973 37964
rect 26007 37961 26019 37995
rect 25961 37955 26019 37961
rect 25976 37856 26004 37955
rect 26421 37859 26479 37865
rect 26421 37856 26433 37859
rect 25976 37828 26433 37856
rect 26421 37825 26433 37828
rect 26467 37825 26479 37859
rect 26421 37819 26479 37825
rect 23753 37791 23811 37797
rect 23753 37788 23765 37791
rect 23624 37760 23765 37788
rect 23624 37748 23630 37760
rect 23753 37757 23765 37760
rect 23799 37757 23811 37791
rect 23753 37751 23811 37757
rect 24581 37791 24639 37797
rect 24581 37757 24593 37791
rect 24627 37757 24639 37791
rect 24581 37751 24639 37757
rect 24673 37791 24731 37797
rect 24673 37757 24685 37791
rect 24719 37757 24731 37791
rect 24673 37751 24731 37757
rect 12805 37723 12863 37729
rect 12805 37689 12817 37723
rect 12851 37720 12863 37723
rect 12894 37720 12900 37732
rect 12851 37692 12900 37720
rect 12851 37689 12863 37692
rect 12805 37683 12863 37689
rect 12894 37680 12900 37692
rect 12952 37680 12958 37732
rect 13170 37720 13176 37732
rect 13131 37692 13176 37720
rect 13170 37680 13176 37692
rect 13228 37680 13234 37732
rect 14001 37723 14059 37729
rect 14001 37689 14013 37723
rect 14047 37720 14059 37723
rect 14369 37723 14427 37729
rect 14047 37692 14320 37720
rect 14047 37689 14059 37692
rect 14001 37683 14059 37689
rect 10229 37655 10287 37661
rect 10229 37652 10241 37655
rect 9916 37624 10241 37652
rect 9916 37612 9922 37624
rect 10229 37621 10241 37624
rect 10275 37652 10287 37655
rect 10597 37655 10655 37661
rect 10597 37652 10609 37655
rect 10275 37624 10609 37652
rect 10275 37621 10287 37624
rect 10229 37615 10287 37621
rect 10597 37621 10609 37624
rect 10643 37621 10655 37655
rect 12710 37652 12716 37664
rect 12671 37624 12716 37652
rect 10597 37615 10655 37621
rect 12710 37612 12716 37624
rect 12768 37652 12774 37664
rect 13449 37655 13507 37661
rect 13449 37652 13461 37655
rect 12768 37624 13461 37652
rect 12768 37612 12774 37624
rect 13449 37621 13461 37624
rect 13495 37621 13507 37655
rect 13449 37615 13507 37621
rect 13909 37655 13967 37661
rect 13909 37621 13921 37655
rect 13955 37652 13967 37655
rect 14182 37652 14188 37664
rect 13955 37624 14188 37652
rect 13955 37621 13967 37624
rect 13909 37615 13967 37621
rect 14182 37612 14188 37624
rect 14240 37612 14246 37664
rect 14292 37652 14320 37692
rect 14369 37689 14381 37723
rect 14415 37720 14427 37723
rect 14458 37720 14464 37732
rect 14415 37692 14464 37720
rect 14415 37689 14427 37692
rect 14369 37683 14427 37689
rect 14458 37680 14464 37692
rect 14516 37680 14522 37732
rect 15565 37723 15623 37729
rect 15565 37720 15577 37723
rect 15396 37692 15577 37720
rect 14918 37652 14924 37664
rect 14292 37624 14924 37652
rect 14918 37612 14924 37624
rect 14976 37612 14982 37664
rect 15286 37652 15292 37664
rect 15199 37624 15292 37652
rect 15286 37612 15292 37624
rect 15344 37652 15350 37664
rect 15396 37661 15424 37692
rect 15565 37689 15577 37692
rect 15611 37689 15623 37723
rect 15746 37720 15752 37732
rect 15707 37692 15752 37720
rect 15565 37683 15623 37689
rect 15746 37680 15752 37692
rect 15804 37680 15810 37732
rect 15930 37720 15936 37732
rect 15843 37692 15936 37720
rect 15930 37680 15936 37692
rect 15988 37720 15994 37732
rect 16758 37720 16764 37732
rect 15988 37692 16764 37720
rect 15988 37680 15994 37692
rect 16758 37680 16764 37692
rect 16816 37680 16822 37732
rect 17037 37723 17095 37729
rect 17037 37689 17049 37723
rect 17083 37720 17095 37723
rect 17494 37720 17500 37732
rect 17083 37692 17500 37720
rect 17083 37689 17095 37692
rect 17037 37683 17095 37689
rect 17494 37680 17500 37692
rect 17552 37680 17558 37732
rect 20346 37720 20352 37732
rect 20307 37692 20352 37720
rect 20346 37680 20352 37692
rect 20404 37680 20410 37732
rect 23842 37720 23848 37732
rect 23803 37692 23848 37720
rect 23842 37680 23848 37692
rect 23900 37680 23906 37732
rect 24688 37720 24716 37751
rect 24762 37748 24768 37800
rect 24820 37788 24826 37800
rect 26145 37791 26203 37797
rect 26145 37788 26157 37791
rect 24820 37760 26157 37788
rect 24820 37748 24826 37760
rect 26145 37757 26157 37760
rect 26191 37788 26203 37791
rect 26234 37788 26240 37800
rect 26191 37760 26240 37788
rect 26191 37757 26203 37760
rect 26145 37751 26203 37757
rect 26234 37748 26240 37760
rect 26292 37748 26298 37800
rect 24596 37692 24716 37720
rect 15381 37655 15439 37661
rect 15381 37652 15393 37655
rect 15344 37624 15393 37652
rect 15344 37612 15350 37624
rect 15381 37621 15393 37624
rect 15427 37621 15439 37655
rect 15381 37615 15439 37621
rect 15841 37655 15899 37661
rect 15841 37621 15853 37655
rect 15887 37652 15899 37655
rect 16298 37652 16304 37664
rect 15887 37624 16304 37652
rect 15887 37621 15899 37624
rect 15841 37615 15899 37621
rect 16298 37612 16304 37624
rect 16356 37612 16362 37664
rect 17402 37612 17408 37664
rect 17460 37652 17466 37664
rect 18325 37655 18383 37661
rect 18325 37652 18337 37655
rect 17460 37624 18337 37652
rect 17460 37612 17466 37624
rect 18325 37621 18337 37624
rect 18371 37652 18383 37655
rect 18874 37652 18880 37664
rect 18371 37624 18880 37652
rect 18371 37621 18383 37624
rect 18325 37615 18383 37621
rect 18874 37612 18880 37624
rect 18932 37612 18938 37664
rect 23658 37612 23664 37664
rect 23716 37652 23722 37664
rect 24596 37652 24624 37692
rect 27522 37652 27528 37664
rect 23716 37624 24624 37652
rect 27483 37624 27528 37652
rect 23716 37612 23722 37624
rect 27522 37612 27528 37624
rect 27580 37612 27586 37664
rect 1104 37562 28888 37584
rect 1104 37510 10982 37562
rect 11034 37510 11046 37562
rect 11098 37510 11110 37562
rect 11162 37510 11174 37562
rect 11226 37510 20982 37562
rect 21034 37510 21046 37562
rect 21098 37510 21110 37562
rect 21162 37510 21174 37562
rect 21226 37510 28888 37562
rect 1104 37488 28888 37510
rect 6917 37451 6975 37457
rect 6917 37417 6929 37451
rect 6963 37448 6975 37451
rect 7742 37448 7748 37460
rect 6963 37420 7748 37448
rect 6963 37417 6975 37420
rect 6917 37411 6975 37417
rect 7742 37408 7748 37420
rect 7800 37408 7806 37460
rect 8938 37408 8944 37460
rect 8996 37448 9002 37460
rect 9398 37448 9404 37460
rect 8996 37420 9404 37448
rect 8996 37408 9002 37420
rect 9398 37408 9404 37420
rect 9456 37408 9462 37460
rect 12621 37451 12679 37457
rect 9784 37420 11560 37448
rect 3053 37383 3111 37389
rect 3053 37349 3065 37383
rect 3099 37380 3111 37383
rect 3142 37380 3148 37392
rect 3099 37352 3148 37380
rect 3099 37349 3111 37352
rect 3053 37343 3111 37349
rect 3142 37340 3148 37352
rect 3200 37340 3206 37392
rect 8662 37380 8668 37392
rect 8623 37352 8668 37380
rect 8662 37340 8668 37352
rect 8720 37340 8726 37392
rect 1670 37312 1676 37324
rect 1631 37284 1676 37312
rect 1670 37272 1676 37284
rect 1728 37272 1734 37324
rect 7285 37315 7343 37321
rect 7285 37312 7297 37315
rect 6840 37284 7297 37312
rect 1394 37244 1400 37256
rect 1355 37216 1400 37244
rect 1394 37204 1400 37216
rect 1452 37204 1458 37256
rect 6546 37204 6552 37256
rect 6604 37244 6610 37256
rect 6840 37244 6868 37284
rect 7285 37281 7297 37284
rect 7331 37281 7343 37315
rect 7285 37275 7343 37281
rect 9490 37272 9496 37324
rect 9548 37312 9554 37324
rect 9784 37321 9812 37420
rect 10321 37383 10379 37389
rect 10321 37349 10333 37383
rect 10367 37380 10379 37383
rect 10778 37380 10784 37392
rect 10367 37352 10784 37380
rect 10367 37349 10379 37352
rect 10321 37343 10379 37349
rect 10778 37340 10784 37352
rect 10836 37340 10842 37392
rect 10870 37340 10876 37392
rect 10928 37380 10934 37392
rect 11532 37389 11560 37420
rect 12621 37417 12633 37451
rect 12667 37448 12679 37451
rect 12802 37448 12808 37460
rect 12667 37420 12808 37448
rect 12667 37417 12679 37420
rect 12621 37411 12679 37417
rect 12802 37408 12808 37420
rect 12860 37408 12866 37460
rect 13630 37408 13636 37460
rect 13688 37448 13694 37460
rect 14185 37451 14243 37457
rect 14185 37448 14197 37451
rect 13688 37420 14197 37448
rect 13688 37408 13694 37420
rect 14185 37417 14197 37420
rect 14231 37448 14243 37451
rect 14918 37448 14924 37460
rect 14231 37420 14924 37448
rect 14231 37417 14243 37420
rect 14185 37411 14243 37417
rect 14918 37408 14924 37420
rect 14976 37408 14982 37460
rect 15378 37408 15384 37460
rect 15436 37448 15442 37460
rect 15933 37451 15991 37457
rect 15933 37448 15945 37451
rect 15436 37420 15945 37448
rect 15436 37408 15442 37420
rect 15933 37417 15945 37420
rect 15979 37417 15991 37451
rect 15933 37411 15991 37417
rect 19518 37408 19524 37460
rect 19576 37448 19582 37460
rect 19613 37451 19671 37457
rect 19613 37448 19625 37451
rect 19576 37420 19625 37448
rect 19576 37408 19582 37420
rect 19613 37417 19625 37420
rect 19659 37417 19671 37451
rect 20254 37448 20260 37460
rect 20215 37420 20260 37448
rect 19613 37411 19671 37417
rect 20254 37408 20260 37420
rect 20312 37408 20318 37460
rect 22094 37448 22100 37460
rect 21928 37420 22100 37448
rect 11517 37383 11575 37389
rect 10928 37352 10973 37380
rect 10928 37340 10934 37352
rect 11517 37349 11529 37383
rect 11563 37380 11575 37383
rect 11790 37380 11796 37392
rect 11563 37352 11796 37380
rect 11563 37349 11575 37352
rect 11517 37343 11575 37349
rect 11790 37340 11796 37352
rect 11848 37340 11854 37392
rect 12434 37340 12440 37392
rect 12492 37380 12498 37392
rect 13357 37383 13415 37389
rect 13357 37380 13369 37383
rect 12492 37352 13369 37380
rect 12492 37340 12498 37352
rect 13357 37349 13369 37352
rect 13403 37349 13415 37383
rect 13357 37343 13415 37349
rect 13449 37383 13507 37389
rect 13449 37349 13461 37383
rect 13495 37380 13507 37383
rect 13538 37380 13544 37392
rect 13495 37352 13544 37380
rect 13495 37349 13507 37352
rect 13449 37343 13507 37349
rect 13538 37340 13544 37352
rect 13596 37340 13602 37392
rect 13722 37340 13728 37392
rect 13780 37380 13786 37392
rect 13817 37383 13875 37389
rect 13817 37380 13829 37383
rect 13780 37352 13829 37380
rect 13780 37340 13786 37352
rect 13817 37349 13829 37352
rect 13863 37380 13875 37383
rect 15010 37380 15016 37392
rect 13863 37352 15016 37380
rect 13863 37349 13875 37352
rect 13817 37343 13875 37349
rect 15010 37340 15016 37352
rect 15068 37340 15074 37392
rect 15105 37383 15163 37389
rect 15105 37349 15117 37383
rect 15151 37380 15163 37383
rect 15654 37380 15660 37392
rect 15151 37352 15660 37380
rect 15151 37349 15163 37352
rect 15105 37343 15163 37349
rect 15654 37340 15660 37352
rect 15712 37340 15718 37392
rect 9769 37315 9827 37321
rect 9769 37312 9781 37315
rect 9548 37284 9781 37312
rect 9548 37272 9554 37284
rect 9769 37281 9781 37284
rect 9815 37281 9827 37315
rect 9769 37275 9827 37281
rect 9861 37315 9919 37321
rect 9861 37281 9873 37315
rect 9907 37281 9919 37315
rect 11330 37312 11336 37324
rect 11291 37284 11336 37312
rect 9861 37275 9919 37281
rect 7006 37244 7012 37256
rect 6604 37216 6868 37244
rect 6967 37216 7012 37244
rect 6604 37204 6610 37216
rect 7006 37204 7012 37216
rect 7064 37204 7070 37256
rect 9214 37204 9220 37256
rect 9272 37244 9278 37256
rect 9876 37244 9904 37275
rect 11330 37272 11336 37284
rect 11388 37272 11394 37324
rect 11422 37272 11428 37324
rect 11480 37312 11486 37324
rect 12161 37315 12219 37321
rect 12161 37312 12173 37315
rect 11480 37284 12173 37312
rect 11480 37272 11486 37284
rect 12161 37281 12173 37284
rect 12207 37281 12219 37315
rect 12161 37275 12219 37281
rect 12802 37272 12808 37324
rect 12860 37312 12866 37324
rect 12986 37312 12992 37324
rect 12860 37284 12992 37312
rect 12860 37272 12866 37284
rect 12986 37272 12992 37284
rect 13044 37312 13050 37324
rect 13265 37315 13323 37321
rect 13265 37312 13277 37315
rect 13044 37284 13277 37312
rect 13044 37272 13050 37284
rect 13265 37281 13277 37284
rect 13311 37281 13323 37315
rect 13265 37275 13323 37281
rect 15289 37315 15347 37321
rect 15289 37281 15301 37315
rect 15335 37312 15347 37315
rect 16669 37315 16727 37321
rect 16669 37312 16681 37315
rect 15335 37284 16681 37312
rect 15335 37281 15347 37284
rect 15289 37275 15347 37281
rect 16669 37281 16681 37284
rect 16715 37312 16727 37315
rect 16758 37312 16764 37324
rect 16715 37284 16764 37312
rect 16715 37281 16727 37284
rect 16669 37275 16727 37281
rect 16758 37272 16764 37284
rect 16816 37272 16822 37324
rect 16850 37272 16856 37324
rect 16908 37312 16914 37324
rect 16908 37284 16953 37312
rect 16908 37272 16914 37284
rect 17402 37272 17408 37324
rect 17460 37312 17466 37324
rect 17589 37315 17647 37321
rect 17589 37312 17601 37315
rect 17460 37284 17601 37312
rect 17460 37272 17466 37284
rect 17589 37281 17601 37284
rect 17635 37281 17647 37315
rect 18138 37312 18144 37324
rect 17589 37275 17647 37281
rect 17880 37284 18144 37312
rect 9272 37216 9904 37244
rect 9272 37204 9278 37216
rect 10594 37204 10600 37256
rect 10652 37244 10658 37256
rect 11149 37247 11207 37253
rect 11149 37244 11161 37247
rect 10652 37216 11161 37244
rect 10652 37204 10658 37216
rect 11149 37213 11161 37216
rect 11195 37213 11207 37247
rect 11149 37207 11207 37213
rect 11885 37247 11943 37253
rect 11885 37213 11897 37247
rect 11931 37213 11943 37247
rect 11885 37207 11943 37213
rect 13081 37247 13139 37253
rect 13081 37213 13093 37247
rect 13127 37213 13139 37247
rect 15654 37244 15660 37256
rect 15615 37216 15660 37244
rect 13081 37207 13139 37213
rect 11054 37136 11060 37188
rect 11112 37176 11118 37188
rect 11900 37176 11928 37207
rect 11112 37148 11928 37176
rect 11112 37136 11118 37148
rect 6181 37111 6239 37117
rect 6181 37077 6193 37111
rect 6227 37108 6239 37111
rect 6362 37108 6368 37120
rect 6227 37080 6368 37108
rect 6227 37077 6239 37080
rect 6181 37071 6239 37077
rect 6362 37068 6368 37080
rect 6420 37108 6426 37120
rect 6457 37111 6515 37117
rect 6457 37108 6469 37111
rect 6420 37080 6469 37108
rect 6420 37068 6426 37080
rect 6457 37077 6469 37080
rect 6503 37077 6515 37111
rect 9030 37108 9036 37120
rect 8991 37080 9036 37108
rect 6457 37071 6515 37077
rect 9030 37068 9036 37080
rect 9088 37068 9094 37120
rect 11238 37068 11244 37120
rect 11296 37108 11302 37120
rect 12897 37111 12955 37117
rect 12897 37108 12909 37111
rect 11296 37080 12909 37108
rect 11296 37068 11302 37080
rect 12897 37077 12909 37080
rect 12943 37108 12955 37111
rect 13096 37108 13124 37207
rect 15654 37204 15660 37216
rect 15712 37204 15718 37256
rect 17221 37247 17279 37253
rect 17221 37213 17233 37247
rect 17267 37244 17279 37247
rect 17267 37216 17724 37244
rect 17267 37213 17279 37216
rect 17221 37207 17279 37213
rect 17696 37188 17724 37216
rect 17770 37204 17776 37256
rect 17828 37244 17834 37256
rect 17880 37244 17908 37284
rect 18138 37272 18144 37284
rect 18196 37312 18202 37324
rect 18233 37315 18291 37321
rect 18233 37312 18245 37315
rect 18196 37284 18245 37312
rect 18196 37272 18202 37284
rect 18233 37281 18245 37284
rect 18279 37281 18291 37315
rect 18414 37312 18420 37324
rect 18375 37284 18420 37312
rect 18233 37275 18291 37281
rect 18414 37272 18420 37284
rect 18472 37272 18478 37324
rect 20272 37312 20300 37408
rect 21928 37321 21956 37420
rect 22094 37408 22100 37420
rect 22152 37408 22158 37460
rect 25498 37448 25504 37460
rect 25459 37420 25504 37448
rect 25498 37408 25504 37420
rect 25556 37408 25562 37460
rect 26234 37448 26240 37460
rect 26195 37420 26240 37448
rect 26234 37408 26240 37420
rect 26292 37408 26298 37460
rect 21913 37315 21971 37321
rect 21913 37312 21925 37315
rect 20272 37284 21925 37312
rect 21913 37281 21925 37284
rect 21959 37281 21971 37315
rect 21913 37275 21971 37281
rect 22005 37315 22063 37321
rect 22005 37281 22017 37315
rect 22051 37312 22063 37315
rect 22554 37312 22560 37324
rect 22051 37284 22560 37312
rect 22051 37281 22063 37284
rect 22005 37275 22063 37281
rect 22554 37272 22560 37284
rect 22612 37272 22618 37324
rect 22738 37312 22744 37324
rect 22699 37284 22744 37312
rect 22738 37272 22744 37284
rect 22796 37272 22802 37324
rect 23658 37312 23664 37324
rect 23619 37284 23664 37312
rect 23658 37272 23664 37284
rect 23716 37272 23722 37324
rect 24026 37272 24032 37324
rect 24084 37312 24090 37324
rect 24213 37315 24271 37321
rect 24213 37312 24225 37315
rect 24084 37284 24225 37312
rect 24084 37272 24090 37284
rect 24213 37281 24225 37284
rect 24259 37281 24271 37315
rect 24213 37275 24271 37281
rect 17828 37216 17908 37244
rect 17828 37204 17834 37216
rect 22462 37204 22468 37256
rect 22520 37244 22526 37256
rect 22833 37247 22891 37253
rect 22833 37244 22845 37247
rect 22520 37216 22845 37244
rect 22520 37204 22526 37216
rect 22833 37213 22845 37216
rect 22879 37244 22891 37247
rect 23474 37244 23480 37256
rect 22879 37216 23480 37244
rect 22879 37213 22891 37216
rect 22833 37207 22891 37213
rect 23474 37204 23480 37216
rect 23532 37204 23538 37256
rect 23937 37247 23995 37253
rect 23937 37213 23949 37247
rect 23983 37244 23995 37247
rect 24670 37244 24676 37256
rect 23983 37216 24676 37244
rect 23983 37213 23995 37216
rect 23937 37207 23995 37213
rect 24670 37204 24676 37216
rect 24728 37204 24734 37256
rect 15454 37179 15512 37185
rect 15454 37145 15466 37179
rect 15500 37176 15512 37179
rect 16393 37179 16451 37185
rect 16393 37176 16405 37179
rect 15500 37148 16405 37176
rect 15500 37145 15512 37148
rect 15454 37139 15512 37145
rect 16393 37145 16405 37148
rect 16439 37176 16451 37179
rect 17586 37176 17592 37188
rect 16439 37148 17592 37176
rect 16439 37145 16451 37148
rect 16393 37139 16451 37145
rect 17586 37136 17592 37148
rect 17644 37136 17650 37188
rect 17678 37136 17684 37188
rect 17736 37176 17742 37188
rect 18601 37179 18659 37185
rect 18601 37176 18613 37179
rect 17736 37148 18613 37176
rect 17736 37136 17742 37148
rect 18601 37145 18613 37148
rect 18647 37145 18659 37179
rect 18601 37139 18659 37145
rect 14461 37111 14519 37117
rect 14461 37108 14473 37111
rect 12943 37080 14473 37108
rect 12943 37077 12955 37080
rect 12897 37071 12955 37077
rect 14461 37077 14473 37080
rect 14507 37108 14519 37111
rect 14734 37108 14740 37120
rect 14507 37080 14740 37108
rect 14507 37077 14519 37080
rect 14461 37071 14519 37077
rect 14734 37068 14740 37080
rect 14792 37068 14798 37120
rect 15565 37111 15623 37117
rect 15565 37077 15577 37111
rect 15611 37108 15623 37111
rect 15654 37108 15660 37120
rect 15611 37080 15660 37108
rect 15611 37077 15623 37080
rect 15565 37071 15623 37077
rect 15654 37068 15660 37080
rect 15712 37068 15718 37120
rect 15746 37068 15752 37120
rect 15804 37108 15810 37120
rect 16666 37108 16672 37120
rect 15804 37080 16672 37108
rect 15804 37068 15810 37080
rect 16666 37068 16672 37080
rect 16724 37108 16730 37120
rect 16991 37111 17049 37117
rect 16991 37108 17003 37111
rect 16724 37080 17003 37108
rect 16724 37068 16730 37080
rect 16991 37077 17003 37080
rect 17037 37077 17049 37111
rect 16991 37071 17049 37077
rect 17129 37111 17187 37117
rect 17129 37077 17141 37111
rect 17175 37108 17187 37111
rect 17218 37108 17224 37120
rect 17175 37080 17224 37108
rect 17175 37077 17187 37080
rect 17129 37071 17187 37077
rect 17218 37068 17224 37080
rect 17276 37068 17282 37120
rect 17957 37111 18015 37117
rect 17957 37077 17969 37111
rect 18003 37108 18015 37111
rect 18782 37108 18788 37120
rect 18003 37080 18788 37108
rect 18003 37077 18015 37080
rect 17957 37071 18015 37077
rect 18782 37068 18788 37080
rect 18840 37068 18846 37120
rect 18969 37111 19027 37117
rect 18969 37077 18981 37111
rect 19015 37108 19027 37111
rect 19058 37108 19064 37120
rect 19015 37080 19064 37108
rect 19015 37077 19027 37080
rect 18969 37071 19027 37077
rect 19058 37068 19064 37080
rect 19116 37068 19122 37120
rect 19337 37111 19395 37117
rect 19337 37077 19349 37111
rect 19383 37108 19395 37111
rect 19426 37108 19432 37120
rect 19383 37080 19432 37108
rect 19383 37077 19395 37080
rect 19337 37071 19395 37077
rect 19426 37068 19432 37080
rect 19484 37068 19490 37120
rect 1104 37018 28888 37040
rect 1104 36966 5982 37018
rect 6034 36966 6046 37018
rect 6098 36966 6110 37018
rect 6162 36966 6174 37018
rect 6226 36966 15982 37018
rect 16034 36966 16046 37018
rect 16098 36966 16110 37018
rect 16162 36966 16174 37018
rect 16226 36966 25982 37018
rect 26034 36966 26046 37018
rect 26098 36966 26110 37018
rect 26162 36966 26174 37018
rect 26226 36966 28888 37018
rect 1104 36944 28888 36966
rect 1670 36904 1676 36916
rect 1631 36876 1676 36904
rect 1670 36864 1676 36876
rect 1728 36864 1734 36916
rect 6273 36907 6331 36913
rect 6273 36873 6285 36907
rect 6319 36904 6331 36907
rect 6822 36904 6828 36916
rect 6319 36876 6828 36904
rect 6319 36873 6331 36876
rect 6273 36867 6331 36873
rect 6822 36864 6828 36876
rect 6880 36864 6886 36916
rect 8941 36907 8999 36913
rect 8941 36873 8953 36907
rect 8987 36904 8999 36907
rect 9490 36904 9496 36916
rect 8987 36876 9496 36904
rect 8987 36873 8999 36876
rect 8941 36867 8999 36873
rect 9490 36864 9496 36876
rect 9548 36864 9554 36916
rect 9766 36864 9772 36916
rect 9824 36904 9830 36916
rect 10919 36907 10977 36913
rect 10919 36904 10931 36907
rect 9824 36876 10931 36904
rect 9824 36864 9830 36876
rect 10919 36873 10931 36876
rect 10965 36873 10977 36907
rect 11054 36904 11060 36916
rect 11015 36876 11060 36904
rect 10919 36867 10977 36873
rect 11054 36864 11060 36876
rect 11112 36864 11118 36916
rect 11330 36864 11336 36916
rect 11388 36904 11394 36916
rect 11793 36907 11851 36913
rect 11793 36904 11805 36907
rect 11388 36876 11805 36904
rect 11388 36864 11394 36876
rect 11793 36873 11805 36876
rect 11839 36904 11851 36907
rect 12342 36904 12348 36916
rect 11839 36876 12348 36904
rect 11839 36873 11851 36876
rect 11793 36867 11851 36873
rect 12342 36864 12348 36876
rect 12400 36864 12406 36916
rect 12526 36864 12532 36916
rect 12584 36904 12590 36916
rect 12713 36907 12771 36913
rect 12713 36904 12725 36907
rect 12584 36876 12725 36904
rect 12584 36864 12590 36876
rect 12713 36873 12725 36876
rect 12759 36873 12771 36907
rect 12713 36867 12771 36873
rect 13062 36907 13120 36913
rect 13062 36873 13074 36907
rect 13108 36904 13120 36907
rect 13722 36904 13728 36916
rect 13108 36876 13728 36904
rect 13108 36873 13120 36876
rect 13062 36867 13120 36873
rect 6546 36836 6552 36848
rect 6507 36808 6552 36836
rect 6546 36796 6552 36808
rect 6604 36796 6610 36848
rect 10594 36836 10600 36848
rect 9508 36808 10600 36836
rect 9508 36780 9536 36808
rect 10594 36796 10600 36808
rect 10652 36796 10658 36848
rect 2130 36768 2136 36780
rect 2091 36740 2136 36768
rect 2130 36728 2136 36740
rect 2188 36728 2194 36780
rect 7098 36768 7104 36780
rect 7011 36740 7104 36768
rect 7098 36728 7104 36740
rect 7156 36768 7162 36780
rect 7926 36768 7932 36780
rect 7156 36740 7932 36768
rect 7156 36728 7162 36740
rect 7926 36728 7932 36740
rect 7984 36728 7990 36780
rect 8846 36728 8852 36780
rect 8904 36768 8910 36780
rect 9306 36768 9312 36780
rect 8904 36740 9312 36768
rect 8904 36728 8910 36740
rect 9306 36728 9312 36740
rect 9364 36728 9370 36780
rect 9490 36728 9496 36780
rect 9548 36728 9554 36780
rect 10229 36771 10287 36777
rect 10229 36768 10241 36771
rect 9600 36740 10241 36768
rect 1394 36660 1400 36712
rect 1452 36700 1458 36712
rect 1857 36703 1915 36709
rect 1857 36700 1869 36703
rect 1452 36672 1869 36700
rect 1452 36660 1458 36672
rect 1857 36669 1869 36672
rect 1903 36700 1915 36703
rect 2406 36700 2412 36712
rect 1903 36672 2412 36700
rect 1903 36669 1915 36672
rect 1857 36663 1915 36669
rect 2406 36660 2412 36672
rect 2464 36660 2470 36712
rect 5537 36703 5595 36709
rect 5537 36669 5549 36703
rect 5583 36700 5595 36703
rect 6362 36700 6368 36712
rect 5583 36672 6368 36700
rect 5583 36669 5595 36672
rect 5537 36663 5595 36669
rect 6362 36660 6368 36672
rect 6420 36700 6426 36712
rect 6825 36703 6883 36709
rect 6825 36700 6837 36703
rect 6420 36672 6837 36700
rect 6420 36660 6426 36672
rect 6825 36669 6837 36672
rect 6871 36700 6883 36703
rect 6914 36700 6920 36712
rect 6871 36672 6920 36700
rect 6871 36669 6883 36672
rect 6825 36663 6883 36669
rect 6914 36660 6920 36672
rect 6972 36660 6978 36712
rect 9398 36700 9404 36712
rect 9359 36672 9404 36700
rect 9398 36660 9404 36672
rect 9456 36660 9462 36712
rect 9600 36709 9628 36740
rect 10229 36737 10241 36740
rect 10275 36737 10287 36771
rect 11146 36768 11152 36780
rect 11107 36740 11152 36768
rect 10229 36731 10287 36737
rect 11146 36728 11152 36740
rect 11204 36728 11210 36780
rect 11517 36771 11575 36777
rect 11517 36737 11529 36771
rect 11563 36768 11575 36771
rect 12618 36768 12624 36780
rect 11563 36740 12624 36768
rect 11563 36737 11575 36740
rect 11517 36731 11575 36737
rect 12618 36728 12624 36740
rect 12676 36728 12682 36780
rect 12728 36768 12756 36867
rect 13722 36864 13728 36876
rect 13780 36864 13786 36916
rect 15654 36864 15660 36916
rect 15712 36904 15718 36916
rect 16390 36904 16396 36916
rect 15712 36876 16396 36904
rect 15712 36864 15718 36876
rect 16390 36864 16396 36876
rect 16448 36864 16454 36916
rect 17405 36907 17463 36913
rect 17405 36904 17417 36907
rect 16592 36876 17417 36904
rect 16592 36848 16620 36876
rect 17405 36873 17417 36876
rect 17451 36904 17463 36907
rect 17678 36904 17684 36916
rect 17451 36876 17684 36904
rect 17451 36873 17463 36876
rect 17405 36867 17463 36873
rect 17678 36864 17684 36876
rect 17736 36864 17742 36916
rect 18414 36864 18420 36916
rect 18472 36904 18478 36916
rect 18509 36907 18567 36913
rect 18509 36904 18521 36907
rect 18472 36876 18521 36904
rect 18472 36864 18478 36876
rect 18509 36873 18521 36876
rect 18555 36873 18567 36907
rect 18509 36867 18567 36873
rect 22094 36864 22100 36916
rect 22152 36904 22158 36916
rect 22189 36907 22247 36913
rect 22189 36904 22201 36907
rect 22152 36876 22201 36904
rect 22152 36864 22158 36876
rect 22189 36873 22201 36876
rect 22235 36873 22247 36907
rect 22189 36867 22247 36873
rect 22649 36907 22707 36913
rect 22649 36873 22661 36907
rect 22695 36904 22707 36907
rect 22738 36904 22744 36916
rect 22695 36876 22744 36904
rect 22695 36873 22707 36876
rect 22649 36867 22707 36873
rect 22738 36864 22744 36876
rect 22796 36864 22802 36916
rect 23934 36904 23940 36916
rect 23895 36876 23940 36904
rect 23934 36864 23940 36876
rect 23992 36864 23998 36916
rect 24397 36907 24455 36913
rect 24397 36873 24409 36907
rect 24443 36904 24455 36907
rect 24762 36904 24768 36916
rect 24443 36876 24768 36904
rect 24443 36873 24455 36876
rect 24397 36867 24455 36873
rect 24762 36864 24768 36876
rect 24820 36864 24826 36916
rect 13173 36839 13231 36845
rect 13173 36805 13185 36839
rect 13219 36836 13231 36839
rect 13354 36836 13360 36848
rect 13219 36808 13360 36836
rect 13219 36805 13231 36808
rect 13173 36799 13231 36805
rect 13354 36796 13360 36808
rect 13412 36796 13418 36848
rect 15010 36836 15016 36848
rect 14476 36808 15016 36836
rect 14476 36777 14504 36808
rect 15010 36796 15016 36808
rect 15068 36836 15074 36848
rect 15286 36836 15292 36848
rect 15068 36808 15292 36836
rect 15068 36796 15074 36808
rect 15286 36796 15292 36808
rect 15344 36796 15350 36848
rect 15749 36839 15807 36845
rect 15749 36805 15761 36839
rect 15795 36836 15807 36839
rect 15933 36839 15991 36845
rect 15933 36836 15945 36839
rect 15795 36808 15945 36836
rect 15795 36805 15807 36808
rect 15749 36799 15807 36805
rect 15933 36805 15945 36808
rect 15979 36836 15991 36839
rect 16574 36836 16580 36848
rect 15979 36808 16580 36836
rect 15979 36805 15991 36808
rect 15933 36799 15991 36805
rect 16574 36796 16580 36808
rect 16632 36796 16638 36848
rect 17218 36796 17224 36848
rect 17276 36836 17282 36848
rect 18233 36839 18291 36845
rect 18233 36836 18245 36839
rect 17276 36808 18245 36836
rect 17276 36796 17282 36808
rect 18233 36805 18245 36808
rect 18279 36805 18291 36839
rect 18233 36799 18291 36805
rect 19245 36839 19303 36845
rect 19245 36805 19257 36839
rect 19291 36805 19303 36839
rect 19245 36799 19303 36805
rect 13265 36771 13323 36777
rect 13265 36768 13277 36771
rect 12728 36740 13277 36768
rect 13265 36737 13277 36740
rect 13311 36737 13323 36771
rect 13265 36731 13323 36737
rect 14461 36771 14519 36777
rect 14461 36737 14473 36771
rect 14507 36737 14519 36771
rect 14461 36731 14519 36737
rect 14550 36728 14556 36780
rect 14608 36768 14614 36780
rect 15197 36771 15255 36777
rect 15197 36768 15209 36771
rect 14608 36740 15209 36768
rect 14608 36728 14614 36740
rect 15197 36737 15209 36740
rect 15243 36737 15255 36771
rect 16758 36768 16764 36780
rect 15197 36731 15255 36737
rect 15396 36740 16620 36768
rect 16719 36740 16764 36768
rect 9585 36703 9643 36709
rect 9585 36669 9597 36703
rect 9631 36669 9643 36703
rect 9585 36663 9643 36669
rect 6454 36592 6460 36644
rect 6512 36632 6518 36644
rect 8481 36635 8539 36641
rect 6512 36604 6960 36632
rect 6512 36592 6518 36604
rect 3234 36564 3240 36576
rect 3195 36536 3240 36564
rect 3234 36524 3240 36536
rect 3292 36524 3298 36576
rect 5905 36567 5963 36573
rect 5905 36533 5917 36567
rect 5951 36564 5963 36567
rect 6638 36564 6644 36576
rect 5951 36536 6644 36564
rect 5951 36533 5963 36536
rect 5905 36527 5963 36533
rect 6638 36524 6644 36536
rect 6696 36524 6702 36576
rect 6932 36564 6960 36604
rect 8481 36601 8493 36635
rect 8527 36632 8539 36635
rect 8846 36632 8852 36644
rect 8527 36604 8852 36632
rect 8527 36601 8539 36604
rect 8481 36595 8539 36601
rect 8846 36592 8852 36604
rect 8904 36592 8910 36644
rect 9600 36632 9628 36663
rect 9674 36660 9680 36712
rect 9732 36700 9738 36712
rect 10781 36703 10839 36709
rect 10781 36700 10793 36703
rect 9732 36672 10793 36700
rect 9732 36660 9738 36672
rect 10781 36669 10793 36672
rect 10827 36669 10839 36703
rect 10781 36663 10839 36669
rect 12897 36703 12955 36709
rect 12897 36669 12909 36703
rect 12943 36700 12955 36703
rect 13078 36700 13084 36712
rect 12943 36672 13084 36700
rect 12943 36669 12955 36672
rect 12897 36663 12955 36669
rect 9048 36604 9628 36632
rect 9048 36564 9076 36604
rect 9214 36564 9220 36576
rect 6932 36536 9076 36564
rect 9175 36536 9220 36564
rect 9214 36524 9220 36536
rect 9272 36524 9278 36576
rect 9674 36564 9680 36576
rect 9635 36536 9680 36564
rect 9674 36524 9680 36536
rect 9732 36524 9738 36576
rect 10796 36564 10824 36663
rect 13078 36660 13084 36672
rect 13136 36700 13142 36712
rect 13722 36700 13728 36712
rect 13136 36672 13728 36700
rect 13136 36660 13142 36672
rect 13722 36660 13728 36672
rect 13780 36660 13786 36712
rect 14182 36660 14188 36712
rect 14240 36700 14246 36712
rect 14369 36703 14427 36709
rect 14369 36700 14381 36703
rect 14240 36672 14381 36700
rect 14240 36660 14246 36672
rect 14369 36669 14381 36672
rect 14415 36700 14427 36703
rect 15396 36700 15424 36740
rect 16298 36700 16304 36712
rect 14415 36672 15424 36700
rect 15580 36672 16304 36700
rect 14415 36669 14427 36672
rect 14369 36663 14427 36669
rect 12253 36635 12311 36641
rect 12253 36601 12265 36635
rect 12299 36632 12311 36635
rect 12434 36632 12440 36644
rect 12299 36604 12440 36632
rect 12299 36601 12311 36604
rect 12253 36595 12311 36601
rect 12434 36592 12440 36604
rect 12492 36592 12498 36644
rect 14734 36632 14740 36644
rect 14695 36604 14740 36632
rect 14734 36592 14740 36604
rect 14792 36592 14798 36644
rect 14844 36641 14872 36672
rect 14829 36635 14887 36641
rect 14829 36601 14841 36635
rect 14875 36601 14887 36635
rect 14829 36595 14887 36601
rect 13541 36567 13599 36573
rect 13541 36564 13553 36567
rect 10796 36536 13553 36564
rect 13541 36533 13553 36536
rect 13587 36533 13599 36567
rect 13541 36527 13599 36533
rect 14001 36567 14059 36573
rect 14001 36533 14013 36567
rect 14047 36564 14059 36567
rect 14274 36564 14280 36576
rect 14047 36536 14280 36564
rect 14047 36533 14059 36536
rect 14001 36527 14059 36533
rect 14274 36524 14280 36536
rect 14332 36524 14338 36576
rect 14550 36524 14556 36576
rect 14608 36564 14614 36576
rect 14645 36567 14703 36573
rect 14645 36564 14657 36567
rect 14608 36536 14657 36564
rect 14608 36524 14614 36536
rect 14645 36533 14657 36536
rect 14691 36533 14703 36567
rect 14645 36527 14703 36533
rect 15286 36524 15292 36576
rect 15344 36564 15350 36576
rect 15580 36573 15608 36672
rect 16298 36660 16304 36672
rect 16356 36660 16362 36712
rect 16592 36700 16620 36740
rect 16758 36728 16764 36740
rect 16816 36728 16822 36780
rect 16850 36728 16856 36780
rect 16908 36768 16914 36780
rect 17129 36771 17187 36777
rect 17129 36768 17141 36771
rect 16908 36740 17141 36768
rect 16908 36728 16914 36740
rect 17129 36737 17141 36740
rect 17175 36768 17187 36771
rect 19260 36768 19288 36799
rect 17175 36740 19288 36768
rect 20533 36771 20591 36777
rect 17175 36737 17187 36740
rect 17129 36731 17187 36737
rect 20533 36737 20545 36771
rect 20579 36768 20591 36771
rect 21634 36768 21640 36780
rect 20579 36740 21640 36768
rect 20579 36737 20591 36740
rect 20533 36731 20591 36737
rect 16868 36700 16896 36728
rect 18046 36700 18052 36712
rect 16592 36672 16896 36700
rect 17959 36672 18052 36700
rect 18046 36660 18052 36672
rect 18104 36700 18110 36712
rect 18877 36703 18935 36709
rect 18877 36700 18889 36703
rect 18104 36672 18889 36700
rect 18104 36660 18110 36672
rect 18877 36669 18889 36672
rect 18923 36669 18935 36703
rect 19058 36700 19064 36712
rect 19019 36672 19064 36700
rect 18877 36663 18935 36669
rect 19058 36660 19064 36672
rect 19116 36700 19122 36712
rect 20640 36709 20668 36740
rect 21634 36728 21640 36740
rect 21692 36728 21698 36780
rect 25866 36728 25872 36780
rect 25924 36768 25930 36780
rect 26053 36771 26111 36777
rect 26053 36768 26065 36771
rect 25924 36740 26065 36768
rect 25924 36728 25930 36740
rect 26053 36737 26065 36740
rect 26099 36737 26111 36771
rect 26053 36731 26111 36737
rect 26145 36771 26203 36777
rect 26145 36737 26157 36771
rect 26191 36768 26203 36771
rect 26326 36768 26332 36780
rect 26191 36740 26332 36768
rect 26191 36737 26203 36740
rect 26145 36731 26203 36737
rect 19521 36703 19579 36709
rect 19521 36700 19533 36703
rect 19116 36672 19533 36700
rect 19116 36660 19122 36672
rect 19521 36669 19533 36672
rect 19567 36700 19579 36703
rect 19889 36703 19947 36709
rect 19889 36700 19901 36703
rect 19567 36672 19901 36700
rect 19567 36669 19579 36672
rect 19521 36663 19579 36669
rect 19889 36669 19901 36672
rect 19935 36669 19947 36703
rect 19889 36663 19947 36669
rect 20625 36703 20683 36709
rect 20625 36669 20637 36703
rect 20671 36669 20683 36703
rect 20625 36663 20683 36669
rect 20714 36660 20720 36712
rect 20772 36700 20778 36712
rect 21085 36703 21143 36709
rect 21085 36700 21097 36703
rect 20772 36672 21097 36700
rect 20772 36660 20778 36672
rect 21085 36669 21097 36672
rect 21131 36669 21143 36703
rect 26068 36700 26096 36731
rect 26326 36728 26332 36740
rect 26384 36728 26390 36780
rect 26421 36703 26479 36709
rect 26421 36700 26433 36703
rect 26068 36672 26433 36700
rect 21085 36663 21143 36669
rect 26421 36669 26433 36672
rect 26467 36669 26479 36703
rect 26421 36663 26479 36669
rect 15749 36635 15807 36641
rect 15749 36601 15761 36635
rect 15795 36632 15807 36635
rect 16025 36635 16083 36641
rect 16025 36632 16037 36635
rect 15795 36604 16037 36632
rect 15795 36601 15807 36604
rect 15749 36595 15807 36601
rect 16025 36601 16037 36604
rect 16071 36601 16083 36635
rect 16025 36595 16083 36601
rect 16114 36592 16120 36644
rect 16172 36632 16178 36644
rect 16393 36635 16451 36641
rect 16393 36632 16405 36635
rect 16172 36604 16405 36632
rect 16172 36592 16178 36604
rect 16393 36601 16405 36604
rect 16439 36601 16451 36635
rect 16393 36595 16451 36601
rect 16666 36592 16672 36644
rect 16724 36632 16730 36644
rect 17773 36635 17831 36641
rect 17773 36632 17785 36635
rect 16724 36604 17785 36632
rect 16724 36592 16730 36604
rect 17773 36601 17785 36604
rect 17819 36601 17831 36635
rect 17773 36595 17831 36601
rect 21361 36635 21419 36641
rect 21361 36601 21373 36635
rect 21407 36632 21419 36635
rect 21542 36632 21548 36644
rect 21407 36604 21548 36632
rect 21407 36601 21419 36604
rect 21361 36595 21419 36601
rect 21542 36592 21548 36604
rect 21600 36592 21606 36644
rect 21913 36635 21971 36641
rect 21913 36601 21925 36635
rect 21959 36632 21971 36635
rect 22462 36632 22468 36644
rect 21959 36604 22468 36632
rect 21959 36601 21971 36604
rect 21913 36595 21971 36601
rect 22462 36592 22468 36604
rect 22520 36592 22526 36644
rect 15565 36567 15623 36573
rect 15565 36564 15577 36567
rect 15344 36536 15577 36564
rect 15344 36524 15350 36536
rect 15565 36533 15577 36536
rect 15611 36533 15623 36567
rect 15565 36527 15623 36533
rect 15930 36524 15936 36576
rect 15988 36564 15994 36576
rect 16209 36567 16267 36573
rect 16209 36564 16221 36567
rect 15988 36536 16221 36564
rect 15988 36524 15994 36536
rect 16209 36533 16221 36536
rect 16255 36564 16267 36567
rect 16482 36564 16488 36576
rect 16255 36536 16488 36564
rect 16255 36533 16267 36536
rect 16209 36527 16267 36533
rect 16482 36524 16488 36536
rect 16540 36524 16546 36576
rect 27706 36564 27712 36576
rect 27667 36536 27712 36564
rect 27706 36524 27712 36536
rect 27764 36524 27770 36576
rect 1104 36474 28888 36496
rect 1104 36422 10982 36474
rect 11034 36422 11046 36474
rect 11098 36422 11110 36474
rect 11162 36422 11174 36474
rect 11226 36422 20982 36474
rect 21034 36422 21046 36474
rect 21098 36422 21110 36474
rect 21162 36422 21174 36474
rect 21226 36422 28888 36474
rect 1104 36400 28888 36422
rect 1949 36363 2007 36369
rect 1949 36329 1961 36363
rect 1995 36360 2007 36363
rect 2130 36360 2136 36372
rect 1995 36332 2136 36360
rect 1995 36329 2007 36332
rect 1949 36323 2007 36329
rect 2130 36320 2136 36332
rect 2188 36320 2194 36372
rect 6917 36363 6975 36369
rect 6917 36329 6929 36363
rect 6963 36360 6975 36363
rect 7098 36360 7104 36372
rect 6963 36332 7104 36360
rect 6963 36329 6975 36332
rect 6917 36323 6975 36329
rect 7098 36320 7104 36332
rect 7156 36320 7162 36372
rect 7561 36363 7619 36369
rect 7561 36329 7573 36363
rect 7607 36360 7619 36363
rect 7834 36360 7840 36372
rect 7607 36332 7840 36360
rect 7607 36329 7619 36332
rect 7561 36323 7619 36329
rect 7834 36320 7840 36332
rect 7892 36360 7898 36372
rect 8294 36360 8300 36372
rect 7892 36332 8300 36360
rect 7892 36320 7898 36332
rect 8294 36320 8300 36332
rect 8352 36320 8358 36372
rect 10137 36363 10195 36369
rect 10137 36329 10149 36363
rect 10183 36360 10195 36363
rect 10686 36360 10692 36372
rect 10183 36332 10692 36360
rect 10183 36329 10195 36332
rect 10137 36323 10195 36329
rect 10686 36320 10692 36332
rect 10744 36320 10750 36372
rect 13538 36320 13544 36372
rect 13596 36360 13602 36372
rect 14553 36363 14611 36369
rect 14553 36360 14565 36363
rect 13596 36332 14565 36360
rect 13596 36320 13602 36332
rect 14553 36329 14565 36332
rect 14599 36360 14611 36363
rect 15010 36360 15016 36372
rect 14599 36332 15016 36360
rect 14599 36329 14611 36332
rect 14553 36323 14611 36329
rect 15010 36320 15016 36332
rect 15068 36320 15074 36372
rect 19610 36360 19616 36372
rect 19571 36332 19616 36360
rect 19610 36320 19616 36332
rect 19668 36320 19674 36372
rect 19978 36360 19984 36372
rect 19939 36332 19984 36360
rect 19978 36320 19984 36332
rect 20036 36320 20042 36372
rect 20438 36320 20444 36372
rect 20496 36360 20502 36372
rect 20714 36360 20720 36372
rect 20496 36332 20720 36360
rect 20496 36320 20502 36332
rect 20714 36320 20720 36332
rect 20772 36320 20778 36372
rect 8389 36295 8447 36301
rect 8389 36261 8401 36295
rect 8435 36292 8447 36295
rect 8570 36292 8576 36304
rect 8435 36264 8576 36292
rect 8435 36261 8447 36264
rect 8389 36255 8447 36261
rect 8570 36252 8576 36264
rect 8628 36252 8634 36304
rect 8757 36295 8815 36301
rect 8757 36261 8769 36295
rect 8803 36292 8815 36295
rect 8803 36264 10640 36292
rect 8803 36261 8815 36264
rect 8757 36255 8815 36261
rect 10612 36236 10640 36264
rect 10870 36252 10876 36304
rect 10928 36292 10934 36304
rect 11698 36292 11704 36304
rect 10928 36264 11704 36292
rect 10928 36252 10934 36264
rect 11698 36252 11704 36264
rect 11756 36292 11762 36304
rect 13265 36295 13323 36301
rect 13265 36292 13277 36295
rect 11756 36264 13277 36292
rect 11756 36252 11762 36264
rect 13265 36261 13277 36264
rect 13311 36292 13323 36295
rect 13630 36292 13636 36304
rect 13311 36264 13636 36292
rect 13311 36261 13323 36264
rect 13265 36255 13323 36261
rect 13630 36252 13636 36264
rect 13688 36252 13694 36304
rect 14001 36295 14059 36301
rect 14001 36261 14013 36295
rect 14047 36292 14059 36295
rect 14090 36292 14096 36304
rect 14047 36264 14096 36292
rect 14047 36261 14059 36264
rect 14001 36255 14059 36261
rect 3694 36184 3700 36236
rect 3752 36224 3758 36236
rect 4893 36227 4951 36233
rect 4893 36224 4905 36227
rect 3752 36196 4905 36224
rect 3752 36184 3758 36196
rect 4893 36193 4905 36196
rect 4939 36224 4951 36227
rect 5166 36224 5172 36236
rect 4939 36196 5172 36224
rect 4939 36193 4951 36196
rect 4893 36187 4951 36193
rect 5166 36184 5172 36196
rect 5224 36184 5230 36236
rect 8205 36227 8263 36233
rect 8205 36224 8217 36227
rect 7852 36196 8217 36224
rect 4154 36116 4160 36168
rect 4212 36156 4218 36168
rect 4617 36159 4675 36165
rect 4617 36156 4629 36159
rect 4212 36128 4629 36156
rect 4212 36116 4218 36128
rect 4617 36125 4629 36128
rect 4663 36125 4675 36159
rect 4617 36119 4675 36125
rect 2317 36023 2375 36029
rect 2317 35989 2329 36023
rect 2363 36020 2375 36023
rect 2406 36020 2412 36032
rect 2363 35992 2412 36020
rect 2363 35989 2375 35992
rect 2317 35983 2375 35989
rect 2406 35980 2412 35992
rect 2464 35980 2470 36032
rect 5350 35980 5356 36032
rect 5408 36020 5414 36032
rect 5997 36023 6055 36029
rect 5997 36020 6009 36023
rect 5408 35992 6009 36020
rect 5408 35980 5414 35992
rect 5997 35989 6009 35992
rect 6043 35989 6055 36023
rect 5997 35983 6055 35989
rect 7650 35980 7656 36032
rect 7708 36020 7714 36032
rect 7852 36029 7880 36196
rect 8205 36193 8217 36196
rect 8251 36193 8263 36227
rect 10134 36224 10140 36236
rect 10095 36196 10140 36224
rect 8205 36187 8263 36193
rect 10134 36184 10140 36196
rect 10192 36184 10198 36236
rect 10594 36224 10600 36236
rect 10555 36196 10600 36224
rect 10594 36184 10600 36196
rect 10652 36184 10658 36236
rect 10686 36184 10692 36236
rect 10744 36224 10750 36236
rect 11241 36227 11299 36233
rect 10744 36196 10789 36224
rect 10744 36184 10750 36196
rect 11241 36193 11253 36227
rect 11287 36224 11299 36227
rect 12618 36224 12624 36236
rect 11287 36196 12624 36224
rect 11287 36193 11299 36196
rect 11241 36187 11299 36193
rect 8021 36159 8079 36165
rect 8021 36125 8033 36159
rect 8067 36156 8079 36159
rect 8570 36156 8576 36168
rect 8067 36128 8576 36156
rect 8067 36125 8079 36128
rect 8021 36119 8079 36125
rect 8570 36116 8576 36128
rect 8628 36116 8634 36168
rect 9493 36159 9551 36165
rect 9493 36125 9505 36159
rect 9539 36156 9551 36159
rect 11256 36156 11284 36187
rect 12618 36184 12624 36196
rect 12676 36184 12682 36236
rect 12802 36184 12808 36236
rect 12860 36224 12866 36236
rect 13081 36227 13139 36233
rect 13081 36224 13093 36227
rect 12860 36196 13093 36224
rect 12860 36184 12866 36196
rect 13081 36193 13093 36196
rect 13127 36193 13139 36227
rect 13081 36187 13139 36193
rect 13173 36227 13231 36233
rect 13173 36193 13185 36227
rect 13219 36224 13231 36227
rect 13354 36224 13360 36236
rect 13219 36196 13360 36224
rect 13219 36193 13231 36196
rect 13173 36187 13231 36193
rect 13354 36184 13360 36196
rect 13412 36184 13418 36236
rect 14016 36224 14044 36255
rect 14090 36252 14096 36264
rect 14148 36292 14154 36304
rect 14734 36292 14740 36304
rect 14148 36264 14740 36292
rect 14148 36252 14154 36264
rect 14734 36252 14740 36264
rect 14792 36252 14798 36304
rect 16298 36252 16304 36304
rect 16356 36292 16362 36304
rect 17129 36295 17187 36301
rect 17129 36292 17141 36295
rect 16356 36264 17141 36292
rect 16356 36252 16362 36264
rect 17129 36261 17141 36264
rect 17175 36261 17187 36295
rect 17129 36255 17187 36261
rect 17221 36295 17279 36301
rect 17221 36261 17233 36295
rect 17267 36261 17279 36295
rect 17586 36292 17592 36304
rect 17547 36264 17592 36292
rect 17221 36255 17279 36261
rect 13464 36196 14044 36224
rect 9539 36128 11284 36156
rect 12897 36159 12955 36165
rect 9539 36125 9551 36128
rect 9493 36119 9551 36125
rect 12897 36125 12909 36159
rect 12943 36156 12955 36159
rect 13464 36156 13492 36196
rect 14550 36184 14556 36236
rect 14608 36224 14614 36236
rect 15930 36224 15936 36236
rect 14608 36196 15936 36224
rect 14608 36184 14614 36196
rect 15930 36184 15936 36196
rect 15988 36184 15994 36236
rect 17037 36227 17095 36233
rect 17037 36193 17049 36227
rect 17083 36193 17095 36227
rect 17236 36224 17264 36255
rect 17586 36252 17592 36264
rect 17644 36252 17650 36304
rect 21818 36292 21824 36304
rect 21779 36264 21824 36292
rect 21818 36252 21824 36264
rect 21876 36252 21882 36304
rect 17770 36224 17776 36236
rect 17236 36196 17776 36224
rect 17037 36187 17095 36193
rect 13630 36156 13636 36168
rect 12943 36128 13492 36156
rect 13591 36128 13636 36156
rect 12943 36125 12955 36128
rect 12897 36119 12955 36125
rect 13630 36116 13636 36128
rect 13688 36116 13694 36168
rect 16025 36159 16083 36165
rect 16025 36125 16037 36159
rect 16071 36156 16083 36159
rect 16482 36156 16488 36168
rect 16071 36128 16488 36156
rect 16071 36125 16083 36128
rect 16025 36119 16083 36125
rect 16482 36116 16488 36128
rect 16540 36116 16546 36168
rect 16850 36156 16856 36168
rect 16811 36128 16856 36156
rect 16850 36116 16856 36128
rect 16908 36116 16914 36168
rect 7926 36048 7932 36100
rect 7984 36088 7990 36100
rect 9122 36088 9128 36100
rect 7984 36060 9128 36088
rect 7984 36048 7990 36060
rect 9122 36048 9128 36060
rect 9180 36088 9186 36100
rect 11054 36088 11060 36100
rect 9180 36060 11060 36088
rect 9180 36048 9186 36060
rect 11054 36048 11060 36060
rect 11112 36048 11118 36100
rect 12161 36091 12219 36097
rect 12161 36057 12173 36091
rect 12207 36088 12219 36091
rect 12434 36088 12440 36100
rect 12207 36060 12440 36088
rect 12207 36057 12219 36060
rect 12161 36051 12219 36057
rect 12434 36048 12440 36060
rect 12492 36048 12498 36100
rect 15010 36048 15016 36100
rect 15068 36088 15074 36100
rect 16114 36088 16120 36100
rect 15068 36060 16120 36088
rect 15068 36048 15074 36060
rect 16114 36048 16120 36060
rect 16172 36048 16178 36100
rect 16206 36048 16212 36100
rect 16264 36048 16270 36100
rect 16761 36091 16819 36097
rect 16761 36057 16773 36091
rect 16807 36088 16819 36091
rect 17052 36088 17080 36187
rect 17604 36168 17632 36196
rect 17770 36184 17776 36196
rect 17828 36184 17834 36236
rect 18509 36227 18567 36233
rect 18509 36193 18521 36227
rect 18555 36224 18567 36227
rect 19058 36224 19064 36236
rect 18555 36196 19064 36224
rect 18555 36193 18567 36196
rect 18509 36187 18567 36193
rect 19058 36184 19064 36196
rect 19116 36184 19122 36236
rect 19426 36184 19432 36236
rect 19484 36224 19490 36236
rect 19797 36227 19855 36233
rect 19797 36224 19809 36227
rect 19484 36196 19809 36224
rect 19484 36184 19490 36196
rect 19797 36193 19809 36196
rect 19843 36224 19855 36227
rect 21174 36224 21180 36236
rect 19843 36196 21180 36224
rect 19843 36193 19855 36196
rect 19797 36187 19855 36193
rect 21174 36184 21180 36196
rect 21232 36184 21238 36236
rect 22557 36227 22615 36233
rect 22557 36193 22569 36227
rect 22603 36224 22615 36227
rect 22830 36224 22836 36236
rect 22603 36196 22836 36224
rect 22603 36193 22615 36196
rect 22557 36187 22615 36193
rect 22830 36184 22836 36196
rect 22888 36184 22894 36236
rect 17586 36116 17592 36168
rect 17644 36116 17650 36168
rect 18230 36116 18236 36168
rect 18288 36156 18294 36168
rect 18417 36159 18475 36165
rect 18417 36156 18429 36159
rect 18288 36128 18429 36156
rect 18288 36116 18294 36128
rect 18417 36125 18429 36128
rect 18463 36125 18475 36159
rect 18417 36119 18475 36125
rect 20714 36116 20720 36168
rect 20772 36156 20778 36168
rect 21542 36156 21548 36168
rect 20772 36128 21548 36156
rect 20772 36116 20778 36128
rect 21542 36116 21548 36128
rect 21600 36156 21606 36168
rect 21729 36159 21787 36165
rect 21729 36156 21741 36159
rect 21600 36128 21741 36156
rect 21600 36116 21606 36128
rect 21729 36125 21741 36128
rect 21775 36125 21787 36159
rect 21729 36119 21787 36125
rect 21818 36116 21824 36168
rect 21876 36156 21882 36168
rect 22002 36156 22008 36168
rect 21876 36128 22008 36156
rect 21876 36116 21882 36128
rect 22002 36116 22008 36128
rect 22060 36116 22066 36168
rect 22462 36116 22468 36168
rect 22520 36156 22526 36168
rect 22649 36159 22707 36165
rect 22649 36156 22661 36159
rect 22520 36128 22661 36156
rect 22520 36116 22526 36128
rect 22649 36125 22661 36128
rect 22695 36125 22707 36159
rect 22649 36119 22707 36125
rect 17218 36088 17224 36100
rect 16807 36060 17224 36088
rect 16807 36057 16819 36060
rect 16761 36051 16819 36057
rect 17218 36048 17224 36060
rect 17276 36048 17282 36100
rect 20254 36088 20260 36100
rect 20215 36060 20260 36088
rect 20254 36048 20260 36060
rect 20312 36048 20318 36100
rect 7837 36023 7895 36029
rect 7837 36020 7849 36023
rect 7708 35992 7849 36020
rect 7708 35980 7714 35992
rect 7837 35989 7849 35992
rect 7883 35989 7895 36023
rect 9030 36020 9036 36032
rect 8991 35992 9036 36020
rect 7837 35983 7895 35989
rect 9030 35980 9036 35992
rect 9088 35980 9094 36032
rect 11701 36023 11759 36029
rect 11701 35989 11713 36023
rect 11747 36020 11759 36023
rect 11790 36020 11796 36032
rect 11747 35992 11796 36020
rect 11747 35989 11759 35992
rect 11701 35983 11759 35989
rect 11790 35980 11796 35992
rect 11848 35980 11854 36032
rect 12526 36020 12532 36032
rect 12487 35992 12532 36020
rect 12526 35980 12532 35992
rect 12584 36020 12590 36032
rect 13906 36020 13912 36032
rect 12584 35992 13912 36020
rect 12584 35980 12590 35992
rect 13906 35980 13912 35992
rect 13964 35980 13970 36032
rect 14826 36020 14832 36032
rect 14787 35992 14832 36020
rect 14826 35980 14832 35992
rect 14884 36020 14890 36032
rect 16224 36020 16252 36048
rect 16390 36020 16396 36032
rect 14884 35992 16252 36020
rect 16351 35992 16396 36020
rect 14884 35980 14890 35992
rect 16390 35980 16396 35992
rect 16448 35980 16454 36032
rect 16666 35980 16672 36032
rect 16724 36020 16730 36032
rect 17494 36020 17500 36032
rect 16724 35992 17500 36020
rect 16724 35980 16730 35992
rect 17494 35980 17500 35992
rect 17552 35980 17558 36032
rect 17954 35980 17960 36032
rect 18012 36020 18018 36032
rect 18049 36023 18107 36029
rect 18049 36020 18061 36023
rect 18012 35992 18061 36020
rect 18012 35980 18018 35992
rect 18049 35989 18061 35992
rect 18095 36020 18107 36023
rect 18693 36023 18751 36029
rect 18693 36020 18705 36023
rect 18095 35992 18705 36020
rect 18095 35989 18107 35992
rect 18049 35983 18107 35989
rect 18693 35989 18705 35992
rect 18739 35989 18751 36023
rect 18693 35983 18751 35989
rect 19150 35980 19156 36032
rect 19208 36020 19214 36032
rect 19337 36023 19395 36029
rect 19337 36020 19349 36023
rect 19208 35992 19349 36020
rect 19208 35980 19214 35992
rect 19337 35989 19349 35992
rect 19383 35989 19395 36023
rect 21174 36020 21180 36032
rect 21135 35992 21180 36020
rect 19337 35983 19395 35989
rect 21174 35980 21180 35992
rect 21232 35980 21238 36032
rect 23566 35980 23572 36032
rect 23624 36020 23630 36032
rect 23661 36023 23719 36029
rect 23661 36020 23673 36023
rect 23624 35992 23673 36020
rect 23624 35980 23630 35992
rect 23661 35989 23673 35992
rect 23707 35989 23719 36023
rect 23661 35983 23719 35989
rect 26237 36023 26295 36029
rect 26237 35989 26249 36023
rect 26283 36020 26295 36023
rect 26326 36020 26332 36032
rect 26283 35992 26332 36020
rect 26283 35989 26295 35992
rect 26237 35983 26295 35989
rect 26326 35980 26332 35992
rect 26384 35980 26390 36032
rect 1104 35930 28888 35952
rect 1104 35878 5982 35930
rect 6034 35878 6046 35930
rect 6098 35878 6110 35930
rect 6162 35878 6174 35930
rect 6226 35878 15982 35930
rect 16034 35878 16046 35930
rect 16098 35878 16110 35930
rect 16162 35878 16174 35930
rect 16226 35878 25982 35930
rect 26034 35878 26046 35930
rect 26098 35878 26110 35930
rect 26162 35878 26174 35930
rect 26226 35878 28888 35930
rect 1104 35856 28888 35878
rect 4614 35816 4620 35828
rect 4575 35788 4620 35816
rect 4614 35776 4620 35788
rect 4672 35776 4678 35828
rect 4890 35816 4896 35828
rect 4851 35788 4896 35816
rect 4890 35776 4896 35788
rect 4948 35776 4954 35828
rect 5166 35816 5172 35828
rect 5127 35788 5172 35816
rect 5166 35776 5172 35788
rect 5224 35776 5230 35828
rect 8570 35816 8576 35828
rect 8531 35788 8576 35816
rect 8570 35776 8576 35788
rect 8628 35776 8634 35828
rect 15102 35776 15108 35828
rect 15160 35816 15166 35828
rect 17218 35816 17224 35828
rect 15160 35788 17080 35816
rect 17179 35788 17224 35816
rect 15160 35776 15166 35788
rect 2406 35748 2412 35760
rect 1596 35720 2412 35748
rect 1394 35436 1400 35488
rect 1452 35476 1458 35488
rect 1596 35485 1624 35720
rect 2406 35708 2412 35720
rect 2464 35748 2470 35760
rect 4154 35748 4160 35760
rect 2464 35720 4160 35748
rect 2464 35708 2470 35720
rect 4154 35708 4160 35720
rect 4212 35708 4218 35760
rect 7650 35708 7656 35760
rect 7708 35748 7714 35760
rect 8849 35751 8907 35757
rect 8849 35748 8861 35751
rect 7708 35720 8861 35748
rect 7708 35708 7714 35720
rect 8849 35717 8861 35720
rect 8895 35748 8907 35751
rect 8941 35751 8999 35757
rect 8941 35748 8953 35751
rect 8895 35720 8953 35748
rect 8895 35717 8907 35720
rect 8849 35711 8907 35717
rect 8941 35717 8953 35720
rect 8987 35748 8999 35751
rect 10413 35751 10471 35757
rect 10413 35748 10425 35751
rect 8987 35720 10425 35748
rect 8987 35717 8999 35720
rect 8941 35711 8999 35717
rect 10413 35717 10425 35720
rect 10459 35748 10471 35751
rect 10505 35751 10563 35757
rect 10505 35748 10517 35751
rect 10459 35720 10517 35748
rect 10459 35717 10471 35720
rect 10413 35711 10471 35717
rect 10505 35717 10517 35720
rect 10551 35717 10563 35751
rect 10505 35711 10563 35717
rect 12802 35708 12808 35760
rect 12860 35748 12866 35760
rect 13541 35751 13599 35757
rect 13541 35748 13553 35751
rect 12860 35720 13553 35748
rect 12860 35708 12866 35720
rect 13541 35717 13553 35720
rect 13587 35748 13599 35751
rect 14274 35748 14280 35760
rect 13587 35720 14280 35748
rect 13587 35717 13599 35720
rect 13541 35711 13599 35717
rect 14274 35708 14280 35720
rect 14332 35708 14338 35760
rect 15841 35751 15899 35757
rect 15841 35717 15853 35751
rect 15887 35748 15899 35751
rect 16298 35748 16304 35760
rect 15887 35720 16304 35748
rect 15887 35717 15899 35720
rect 15841 35711 15899 35717
rect 2866 35680 2872 35692
rect 2827 35652 2872 35680
rect 2866 35640 2872 35652
rect 2924 35640 2930 35692
rect 6638 35640 6644 35692
rect 6696 35680 6702 35692
rect 7190 35680 7196 35692
rect 6696 35652 7196 35680
rect 6696 35640 6702 35652
rect 7190 35640 7196 35652
rect 7248 35680 7254 35692
rect 7248 35652 7972 35680
rect 7248 35640 7254 35652
rect 1854 35572 1860 35624
rect 1912 35612 1918 35624
rect 2501 35615 2559 35621
rect 2501 35612 2513 35615
rect 1912 35584 2513 35612
rect 1912 35572 1918 35584
rect 2501 35581 2513 35584
rect 2547 35612 2559 35615
rect 3145 35615 3203 35621
rect 3145 35612 3157 35615
rect 2547 35584 3157 35612
rect 2547 35581 2559 35584
rect 2501 35575 2559 35581
rect 3145 35581 3157 35584
rect 3191 35581 3203 35615
rect 3145 35575 3203 35581
rect 4709 35615 4767 35621
rect 4709 35581 4721 35615
rect 4755 35581 4767 35615
rect 4709 35575 4767 35581
rect 5721 35615 5779 35621
rect 5721 35581 5733 35615
rect 5767 35612 5779 35615
rect 6178 35612 6184 35624
rect 5767 35584 6184 35612
rect 5767 35581 5779 35584
rect 5721 35575 5779 35581
rect 2314 35544 2320 35556
rect 2227 35516 2320 35544
rect 2314 35504 2320 35516
rect 2372 35504 2378 35556
rect 4522 35504 4528 35556
rect 4580 35544 4586 35556
rect 4724 35544 4752 35575
rect 6178 35572 6184 35584
rect 6236 35572 6242 35624
rect 7101 35615 7159 35621
rect 7101 35581 7113 35615
rect 7147 35612 7159 35615
rect 7834 35612 7840 35624
rect 7147 35584 7840 35612
rect 7147 35581 7159 35584
rect 7101 35575 7159 35581
rect 7834 35572 7840 35584
rect 7892 35572 7898 35624
rect 7944 35553 7972 35652
rect 8202 35640 8208 35692
rect 8260 35680 8266 35692
rect 8297 35683 8355 35689
rect 8297 35680 8309 35683
rect 8260 35652 8309 35680
rect 8260 35640 8266 35652
rect 8297 35649 8309 35652
rect 8343 35649 8355 35683
rect 8297 35643 8355 35649
rect 9766 35640 9772 35692
rect 9824 35680 9830 35692
rect 9861 35683 9919 35689
rect 9861 35680 9873 35683
rect 9824 35652 9873 35680
rect 9824 35640 9830 35652
rect 9861 35649 9873 35652
rect 9907 35649 9919 35683
rect 9861 35643 9919 35649
rect 10045 35683 10103 35689
rect 10045 35649 10057 35683
rect 10091 35680 10103 35683
rect 11330 35680 11336 35692
rect 10091 35652 11336 35680
rect 10091 35649 10103 35652
rect 10045 35643 10103 35649
rect 11330 35640 11336 35652
rect 11388 35640 11394 35692
rect 12434 35640 12440 35692
rect 12492 35640 12498 35692
rect 13078 35640 13084 35692
rect 13136 35680 13142 35692
rect 13173 35683 13231 35689
rect 13173 35680 13185 35683
rect 13136 35652 13185 35680
rect 13136 35640 13142 35652
rect 13173 35649 13185 35652
rect 13219 35649 13231 35683
rect 13173 35643 13231 35649
rect 14001 35683 14059 35689
rect 14001 35649 14013 35683
rect 14047 35680 14059 35683
rect 14550 35680 14556 35692
rect 14047 35652 14556 35680
rect 14047 35649 14059 35652
rect 14001 35643 14059 35649
rect 14550 35640 14556 35652
rect 14608 35640 14614 35692
rect 15102 35640 15108 35692
rect 15160 35640 15166 35692
rect 15473 35683 15531 35689
rect 15473 35649 15485 35683
rect 15519 35680 15531 35683
rect 15856 35680 15884 35711
rect 16298 35708 16304 35720
rect 16356 35708 16362 35760
rect 17052 35748 17080 35788
rect 17218 35776 17224 35788
rect 17276 35776 17282 35828
rect 18138 35776 18144 35828
rect 18196 35816 18202 35828
rect 18877 35819 18935 35825
rect 18877 35816 18889 35819
rect 18196 35788 18889 35816
rect 18196 35776 18202 35788
rect 18877 35785 18889 35788
rect 18923 35785 18935 35819
rect 18877 35779 18935 35785
rect 19334 35776 19340 35828
rect 19392 35816 19398 35828
rect 19613 35819 19671 35825
rect 19613 35816 19625 35819
rect 19392 35788 19625 35816
rect 19392 35776 19398 35788
rect 19613 35785 19625 35788
rect 19659 35785 19671 35819
rect 19613 35779 19671 35785
rect 21269 35819 21327 35825
rect 21269 35785 21281 35819
rect 21315 35816 21327 35819
rect 21634 35816 21640 35828
rect 21315 35788 21640 35816
rect 21315 35785 21327 35788
rect 21269 35779 21327 35785
rect 17770 35748 17776 35760
rect 17052 35720 17776 35748
rect 17770 35708 17776 35720
rect 17828 35708 17834 35760
rect 18230 35708 18236 35760
rect 18288 35748 18294 35760
rect 19061 35751 19119 35757
rect 19061 35748 19073 35751
rect 18288 35720 19073 35748
rect 18288 35708 18294 35720
rect 19061 35717 19073 35720
rect 19107 35717 19119 35751
rect 19061 35711 19119 35717
rect 15519 35652 15884 35680
rect 15519 35649 15531 35652
rect 15473 35643 15531 35649
rect 15930 35640 15936 35692
rect 15988 35680 15994 35692
rect 15988 35652 16033 35680
rect 15988 35640 15994 35652
rect 16850 35640 16856 35692
rect 16908 35680 16914 35692
rect 16945 35683 17003 35689
rect 16945 35680 16957 35683
rect 16908 35652 16957 35680
rect 16908 35640 16914 35652
rect 16945 35649 16957 35652
rect 16991 35680 17003 35683
rect 17865 35683 17923 35689
rect 17865 35680 17877 35683
rect 16991 35652 17877 35680
rect 16991 35649 17003 35652
rect 16945 35643 17003 35649
rect 17865 35649 17877 35652
rect 17911 35680 17923 35683
rect 18049 35683 18107 35689
rect 18049 35680 18061 35683
rect 17911 35652 18061 35680
rect 17911 35649 17923 35652
rect 17865 35643 17923 35649
rect 18049 35649 18061 35652
rect 18095 35680 18107 35683
rect 18414 35680 18420 35692
rect 18095 35652 18420 35680
rect 18095 35649 18107 35652
rect 18049 35643 18107 35649
rect 18414 35640 18420 35652
rect 18472 35640 18478 35692
rect 18785 35683 18843 35689
rect 18785 35649 18797 35683
rect 18831 35680 18843 35683
rect 18877 35683 18935 35689
rect 18877 35680 18889 35683
rect 18831 35652 18889 35680
rect 18831 35649 18843 35652
rect 18785 35643 18843 35649
rect 18877 35649 18889 35652
rect 18923 35649 18935 35683
rect 18877 35643 18935 35649
rect 8478 35612 8484 35624
rect 8036 35584 8484 35612
rect 5629 35547 5687 35553
rect 5629 35544 5641 35547
rect 4580 35516 5641 35544
rect 4580 35504 4586 35516
rect 5629 35513 5641 35516
rect 5675 35544 5687 35547
rect 6641 35547 6699 35553
rect 6641 35544 6653 35547
rect 5675 35516 6653 35544
rect 5675 35513 5687 35516
rect 5629 35507 5687 35513
rect 6641 35513 6653 35516
rect 6687 35544 6699 35547
rect 7561 35547 7619 35553
rect 7561 35544 7573 35547
rect 6687 35516 7573 35544
rect 6687 35513 6699 35516
rect 6641 35507 6699 35513
rect 7561 35513 7573 35516
rect 7607 35544 7619 35547
rect 7929 35547 7987 35553
rect 7607 35516 7880 35544
rect 7607 35513 7619 35516
rect 7561 35507 7619 35513
rect 1581 35479 1639 35485
rect 1581 35476 1593 35479
rect 1452 35448 1593 35476
rect 1452 35436 1458 35448
rect 1581 35445 1593 35448
rect 1627 35445 1639 35479
rect 1581 35439 1639 35445
rect 1670 35436 1676 35488
rect 1728 35476 1734 35488
rect 2133 35479 2191 35485
rect 2133 35476 2145 35479
rect 1728 35448 2145 35476
rect 1728 35436 1734 35448
rect 2133 35445 2145 35448
rect 2179 35476 2191 35479
rect 2332 35476 2360 35504
rect 2179 35448 2360 35476
rect 5905 35479 5963 35485
rect 2179 35445 2191 35448
rect 2133 35439 2191 35445
rect 5905 35445 5917 35479
rect 5951 35476 5963 35479
rect 6914 35476 6920 35488
rect 5951 35448 6920 35476
rect 5951 35445 5963 35448
rect 5905 35439 5963 35445
rect 6914 35436 6920 35448
rect 6972 35436 6978 35488
rect 7098 35436 7104 35488
rect 7156 35476 7162 35488
rect 7377 35479 7435 35485
rect 7377 35476 7389 35479
rect 7156 35448 7389 35476
rect 7156 35436 7162 35448
rect 7377 35445 7389 35448
rect 7423 35476 7435 35479
rect 7650 35476 7656 35488
rect 7423 35448 7656 35476
rect 7423 35445 7435 35448
rect 7377 35439 7435 35445
rect 7650 35436 7656 35448
rect 7708 35476 7714 35488
rect 7745 35479 7803 35485
rect 7745 35476 7757 35479
rect 7708 35448 7757 35476
rect 7708 35436 7714 35448
rect 7745 35445 7757 35448
rect 7791 35445 7803 35479
rect 7852 35476 7880 35516
rect 7929 35513 7941 35547
rect 7975 35513 7987 35547
rect 7929 35507 7987 35513
rect 8036 35476 8064 35584
rect 8478 35572 8484 35584
rect 8536 35612 8542 35624
rect 9122 35612 9128 35624
rect 8536 35584 9128 35612
rect 8536 35572 8542 35584
rect 9122 35572 9128 35584
rect 9180 35612 9186 35624
rect 9180 35584 9628 35612
rect 9180 35572 9186 35584
rect 8849 35547 8907 35553
rect 8849 35513 8861 35547
rect 8895 35544 8907 35547
rect 9309 35547 9367 35553
rect 9309 35544 9321 35547
rect 8895 35516 9321 35544
rect 8895 35513 8907 35516
rect 8849 35507 8907 35513
rect 9309 35513 9321 35516
rect 9355 35513 9367 35547
rect 9490 35544 9496 35556
rect 9451 35516 9496 35544
rect 9309 35507 9367 35513
rect 9490 35504 9496 35516
rect 9548 35504 9554 35556
rect 9600 35544 9628 35584
rect 10134 35572 10140 35624
rect 10192 35612 10198 35624
rect 10229 35615 10287 35621
rect 10229 35612 10241 35615
rect 10192 35584 10241 35612
rect 10192 35572 10198 35584
rect 10229 35581 10241 35584
rect 10275 35612 10287 35615
rect 11698 35612 11704 35624
rect 10275 35584 11704 35612
rect 10275 35581 10287 35584
rect 10229 35575 10287 35581
rect 11698 35572 11704 35584
rect 11756 35572 11762 35624
rect 11885 35615 11943 35621
rect 11885 35581 11897 35615
rect 11931 35612 11943 35615
rect 12452 35612 12480 35640
rect 11931 35584 12848 35612
rect 11931 35581 11943 35584
rect 11885 35575 11943 35581
rect 10689 35547 10747 35553
rect 10689 35544 10701 35547
rect 9600 35516 10701 35544
rect 10689 35513 10701 35516
rect 10735 35544 10747 35547
rect 10778 35544 10784 35556
rect 10735 35516 10784 35544
rect 10735 35513 10747 35516
rect 10689 35507 10747 35513
rect 10778 35504 10784 35516
rect 10836 35504 10842 35556
rect 11054 35544 11060 35556
rect 11015 35516 11060 35544
rect 11054 35504 11060 35516
rect 11112 35504 11118 35556
rect 11422 35544 11428 35556
rect 11383 35516 11428 35544
rect 11422 35504 11428 35516
rect 11480 35504 11486 35556
rect 12158 35504 12164 35556
rect 12216 35544 12222 35556
rect 12253 35547 12311 35553
rect 12253 35544 12265 35547
rect 12216 35516 12265 35544
rect 12216 35504 12222 35516
rect 12253 35513 12265 35516
rect 12299 35544 12311 35547
rect 12434 35544 12440 35556
rect 12299 35516 12440 35544
rect 12299 35513 12311 35516
rect 12253 35507 12311 35513
rect 12434 35504 12440 35516
rect 12492 35504 12498 35556
rect 12820 35553 12848 35584
rect 14182 35572 14188 35624
rect 14240 35612 14246 35624
rect 14277 35615 14335 35621
rect 14277 35612 14289 35615
rect 14240 35584 14289 35612
rect 14240 35572 14246 35584
rect 14277 35581 14289 35584
rect 14323 35581 14335 35615
rect 15120 35612 15148 35640
rect 14277 35575 14335 35581
rect 14384 35584 15148 35612
rect 15712 35615 15770 35621
rect 12805 35547 12863 35553
rect 12805 35513 12817 35547
rect 12851 35544 12863 35547
rect 13354 35544 13360 35556
rect 12851 35516 13360 35544
rect 12851 35513 12863 35516
rect 12805 35507 12863 35513
rect 13354 35504 13360 35516
rect 13412 35504 13418 35556
rect 13814 35504 13820 35556
rect 13872 35544 13878 35556
rect 14384 35553 14412 35584
rect 15712 35581 15724 35615
rect 15758 35612 15770 35615
rect 16022 35612 16028 35624
rect 15758 35584 16028 35612
rect 15758 35581 15770 35584
rect 15712 35575 15770 35581
rect 16022 35572 16028 35584
rect 16080 35572 16086 35624
rect 17218 35572 17224 35624
rect 17276 35612 17282 35624
rect 18138 35612 18144 35624
rect 17276 35584 18144 35612
rect 17276 35572 17282 35584
rect 18138 35572 18144 35584
rect 18196 35612 18202 35624
rect 18233 35615 18291 35621
rect 18233 35612 18245 35615
rect 18196 35584 18245 35612
rect 18196 35572 18202 35584
rect 18233 35581 18245 35584
rect 18279 35581 18291 35615
rect 19628 35612 19656 35779
rect 21634 35776 21640 35788
rect 21692 35776 21698 35828
rect 22462 35816 22468 35828
rect 22423 35788 22468 35816
rect 22462 35776 22468 35788
rect 22520 35776 22526 35828
rect 23477 35683 23535 35689
rect 23477 35649 23489 35683
rect 23523 35680 23535 35683
rect 23934 35680 23940 35692
rect 23523 35652 23940 35680
rect 23523 35649 23535 35652
rect 23477 35643 23535 35649
rect 23934 35640 23940 35652
rect 23992 35640 23998 35692
rect 26145 35683 26203 35689
rect 26145 35649 26157 35683
rect 26191 35680 26203 35683
rect 26326 35680 26332 35692
rect 26191 35652 26332 35680
rect 26191 35649 26203 35652
rect 26145 35643 26203 35649
rect 26326 35640 26332 35652
rect 26384 35640 26390 35692
rect 26421 35683 26479 35689
rect 26421 35649 26433 35683
rect 26467 35680 26479 35683
rect 27798 35680 27804 35692
rect 26467 35652 27804 35680
rect 26467 35649 26479 35652
rect 26421 35643 26479 35649
rect 19889 35615 19947 35621
rect 19889 35612 19901 35615
rect 19628 35584 19901 35612
rect 18233 35575 18291 35581
rect 19889 35581 19901 35584
rect 19935 35581 19947 35615
rect 21634 35612 21640 35624
rect 21595 35584 21640 35612
rect 19889 35575 19947 35581
rect 21634 35572 21640 35584
rect 21692 35572 21698 35624
rect 23014 35572 23020 35624
rect 23072 35612 23078 35624
rect 23566 35612 23572 35624
rect 23072 35584 23572 35612
rect 23072 35572 23078 35584
rect 23566 35572 23572 35584
rect 23624 35612 23630 35624
rect 23661 35615 23719 35621
rect 23661 35612 23673 35615
rect 23624 35584 23673 35612
rect 23624 35572 23630 35584
rect 23661 35581 23673 35584
rect 23707 35581 23719 35615
rect 23661 35575 23719 35581
rect 26053 35615 26111 35621
rect 26053 35581 26065 35615
rect 26099 35612 26111 35615
rect 26436 35612 26464 35643
rect 27798 35640 27804 35652
rect 27856 35640 27862 35692
rect 26099 35584 26464 35612
rect 26099 35581 26111 35584
rect 26053 35575 26111 35581
rect 14369 35547 14427 35553
rect 14369 35544 14381 35547
rect 13872 35516 14381 35544
rect 13872 35504 13878 35516
rect 14369 35513 14381 35516
rect 14415 35513 14427 35547
rect 14734 35544 14740 35556
rect 14695 35516 14740 35544
rect 14369 35507 14427 35513
rect 14734 35504 14740 35516
rect 14792 35504 14798 35556
rect 15565 35547 15623 35553
rect 15565 35513 15577 35547
rect 15611 35544 15623 35547
rect 16482 35544 16488 35556
rect 15611 35516 16488 35544
rect 15611 35513 15623 35516
rect 15565 35507 15623 35513
rect 16482 35504 16488 35516
rect 16540 35504 16546 35556
rect 16758 35504 16764 35556
rect 16816 35544 16822 35556
rect 18417 35547 18475 35553
rect 18417 35544 18429 35547
rect 16816 35516 18429 35544
rect 16816 35504 16822 35516
rect 18417 35513 18429 35516
rect 18463 35544 18475 35547
rect 19150 35544 19156 35556
rect 18463 35516 19156 35544
rect 18463 35513 18475 35516
rect 18417 35507 18475 35513
rect 19150 35504 19156 35516
rect 19208 35504 19214 35556
rect 20530 35544 20536 35556
rect 20491 35516 20536 35544
rect 20530 35504 20536 35516
rect 20588 35504 20594 35556
rect 22097 35547 22155 35553
rect 22097 35513 22109 35547
rect 22143 35544 22155 35547
rect 22278 35544 22284 35556
rect 22143 35516 22284 35544
rect 22143 35513 22155 35516
rect 22097 35507 22155 35513
rect 22278 35504 22284 35516
rect 22336 35504 22342 35556
rect 25314 35544 25320 35556
rect 25275 35516 25320 35544
rect 25314 35504 25320 35516
rect 25372 35504 25378 35556
rect 27798 35544 27804 35556
rect 27759 35516 27804 35544
rect 27798 35504 27804 35516
rect 27856 35504 27862 35556
rect 7852 35448 8064 35476
rect 7745 35439 7803 35445
rect 8294 35436 8300 35488
rect 8352 35476 8358 35488
rect 9030 35476 9036 35488
rect 8352 35448 9036 35476
rect 8352 35436 8358 35448
rect 9030 35436 9036 35448
rect 9088 35476 9094 35488
rect 9401 35479 9459 35485
rect 9401 35476 9413 35479
rect 9088 35448 9413 35476
rect 9088 35436 9094 35448
rect 9401 35445 9413 35448
rect 9447 35476 9459 35479
rect 10045 35479 10103 35485
rect 10045 35476 10057 35479
rect 9447 35448 10057 35476
rect 9447 35445 9459 35448
rect 9401 35439 9459 35445
rect 10045 35445 10057 35448
rect 10091 35476 10103 35479
rect 10134 35476 10140 35488
rect 10091 35448 10140 35476
rect 10091 35445 10103 35448
rect 10045 35439 10103 35445
rect 10134 35436 10140 35448
rect 10192 35436 10198 35488
rect 10413 35479 10471 35485
rect 10413 35445 10425 35479
rect 10459 35476 10471 35479
rect 10873 35479 10931 35485
rect 10873 35476 10885 35479
rect 10459 35448 10885 35476
rect 10459 35445 10471 35448
rect 10413 35439 10471 35445
rect 10873 35445 10885 35448
rect 10919 35445 10931 35479
rect 10873 35439 10931 35445
rect 10965 35479 11023 35485
rect 10965 35445 10977 35479
rect 11011 35476 11023 35479
rect 11330 35476 11336 35488
rect 11011 35448 11336 35476
rect 11011 35445 11023 35448
rect 10965 35439 11023 35445
rect 11330 35436 11336 35448
rect 11388 35436 11394 35488
rect 12526 35436 12532 35488
rect 12584 35476 12590 35488
rect 12621 35479 12679 35485
rect 12621 35476 12633 35479
rect 12584 35448 12633 35476
rect 12584 35436 12590 35448
rect 12621 35445 12633 35448
rect 12667 35445 12679 35479
rect 12621 35439 12679 35445
rect 12713 35479 12771 35485
rect 12713 35445 12725 35479
rect 12759 35476 12771 35479
rect 12986 35476 12992 35488
rect 12759 35448 12992 35476
rect 12759 35445 12771 35448
rect 12713 35439 12771 35445
rect 12986 35436 12992 35448
rect 13044 35436 13050 35488
rect 13906 35476 13912 35488
rect 13867 35448 13912 35476
rect 13906 35436 13912 35448
rect 13964 35476 13970 35488
rect 14185 35479 14243 35485
rect 14185 35476 14197 35479
rect 13964 35448 14197 35476
rect 13964 35436 13970 35448
rect 14185 35445 14197 35448
rect 14231 35445 14243 35479
rect 14185 35439 14243 35445
rect 14918 35436 14924 35488
rect 14976 35476 14982 35488
rect 15013 35479 15071 35485
rect 15013 35476 15025 35479
rect 14976 35448 15025 35476
rect 14976 35436 14982 35448
rect 15013 35445 15025 35448
rect 15059 35445 15071 35479
rect 15013 35439 15071 35445
rect 15470 35436 15476 35488
rect 15528 35476 15534 35488
rect 16209 35479 16267 35485
rect 16209 35476 16221 35479
rect 15528 35448 16221 35476
rect 15528 35436 15534 35448
rect 16209 35445 16221 35448
rect 16255 35445 16267 35479
rect 16209 35439 16267 35445
rect 17954 35436 17960 35488
rect 18012 35476 18018 35488
rect 18230 35476 18236 35488
rect 18012 35448 18236 35476
rect 18012 35436 18018 35448
rect 18230 35436 18236 35448
rect 18288 35476 18294 35488
rect 18325 35479 18383 35485
rect 18325 35476 18337 35479
rect 18288 35448 18337 35476
rect 18288 35436 18294 35448
rect 18325 35445 18337 35448
rect 18371 35445 18383 35479
rect 18325 35439 18383 35445
rect 20714 35436 20720 35488
rect 20772 35476 20778 35488
rect 20809 35479 20867 35485
rect 20809 35476 20821 35479
rect 20772 35448 20821 35476
rect 20772 35436 20778 35448
rect 20809 35445 20821 35448
rect 20855 35445 20867 35479
rect 22830 35476 22836 35488
rect 22791 35448 22836 35476
rect 20809 35439 20867 35445
rect 22830 35436 22836 35448
rect 22888 35436 22894 35488
rect 1104 35386 28888 35408
rect 1104 35334 10982 35386
rect 11034 35334 11046 35386
rect 11098 35334 11110 35386
rect 11162 35334 11174 35386
rect 11226 35334 20982 35386
rect 21034 35334 21046 35386
rect 21098 35334 21110 35386
rect 21162 35334 21174 35386
rect 21226 35334 28888 35386
rect 1104 35312 28888 35334
rect 4614 35272 4620 35284
rect 4575 35244 4620 35272
rect 4614 35232 4620 35244
rect 4672 35232 4678 35284
rect 5629 35275 5687 35281
rect 5629 35241 5641 35275
rect 5675 35272 5687 35275
rect 9490 35272 9496 35284
rect 5675 35244 9496 35272
rect 5675 35241 5687 35244
rect 5629 35235 5687 35241
rect 9490 35232 9496 35244
rect 9548 35232 9554 35284
rect 9953 35275 10011 35281
rect 9953 35241 9965 35275
rect 9999 35272 10011 35275
rect 10134 35272 10140 35284
rect 9999 35244 10140 35272
rect 9999 35241 10011 35244
rect 9953 35235 10011 35241
rect 10134 35232 10140 35244
rect 10192 35232 10198 35284
rect 10594 35232 10600 35284
rect 10652 35272 10658 35284
rect 10689 35275 10747 35281
rect 10689 35272 10701 35275
rect 10652 35244 10701 35272
rect 10652 35232 10658 35244
rect 10689 35241 10701 35244
rect 10735 35241 10747 35275
rect 10689 35235 10747 35241
rect 10778 35232 10784 35284
rect 10836 35272 10842 35284
rect 11057 35275 11115 35281
rect 11057 35272 11069 35275
rect 10836 35244 11069 35272
rect 10836 35232 10842 35244
rect 11057 35241 11069 35244
rect 11103 35241 11115 35275
rect 13449 35275 13507 35281
rect 13449 35272 13461 35275
rect 11057 35235 11115 35241
rect 11256 35244 13461 35272
rect 11256 35216 11284 35244
rect 13449 35241 13461 35244
rect 13495 35241 13507 35275
rect 14182 35272 14188 35284
rect 14143 35244 14188 35272
rect 13449 35235 13507 35241
rect 14182 35232 14188 35244
rect 14240 35232 14246 35284
rect 14918 35232 14924 35284
rect 14976 35272 14982 35284
rect 15930 35272 15936 35284
rect 14976 35244 15936 35272
rect 14976 35232 14982 35244
rect 15930 35232 15936 35244
rect 15988 35232 15994 35284
rect 16393 35275 16451 35281
rect 16393 35241 16405 35275
rect 16439 35272 16451 35275
rect 16482 35272 16488 35284
rect 16439 35244 16488 35272
rect 16439 35241 16451 35244
rect 16393 35235 16451 35241
rect 16482 35232 16488 35244
rect 16540 35272 16546 35284
rect 18046 35272 18052 35284
rect 16540 35244 18052 35272
rect 16540 35232 16546 35244
rect 18046 35232 18052 35244
rect 18104 35232 18110 35284
rect 18138 35232 18144 35284
rect 18196 35272 18202 35284
rect 18196 35244 18241 35272
rect 18196 35232 18202 35244
rect 19334 35232 19340 35284
rect 19392 35272 19398 35284
rect 19429 35275 19487 35281
rect 19429 35272 19441 35275
rect 19392 35244 19441 35272
rect 19392 35232 19398 35244
rect 19429 35241 19441 35244
rect 19475 35241 19487 35275
rect 19886 35272 19892 35284
rect 19847 35244 19892 35272
rect 19429 35235 19487 35241
rect 19886 35232 19892 35244
rect 19944 35232 19950 35284
rect 20530 35272 20536 35284
rect 20443 35244 20536 35272
rect 20530 35232 20536 35244
rect 20588 35272 20594 35284
rect 22186 35272 22192 35284
rect 20588 35244 22192 35272
rect 20588 35232 20594 35244
rect 22186 35232 22192 35244
rect 22244 35232 22250 35284
rect 9122 35204 9128 35216
rect 9083 35176 9128 35204
rect 9122 35164 9128 35176
rect 9180 35164 9186 35216
rect 11238 35204 11244 35216
rect 11199 35176 11244 35204
rect 11238 35164 11244 35176
rect 11296 35164 11302 35216
rect 11974 35204 11980 35216
rect 11935 35176 11980 35204
rect 11974 35164 11980 35176
rect 12032 35164 12038 35216
rect 12526 35204 12532 35216
rect 12487 35176 12532 35204
rect 12526 35164 12532 35176
rect 12584 35204 12590 35216
rect 12710 35204 12716 35216
rect 12584 35176 12716 35204
rect 12584 35164 12590 35176
rect 12710 35164 12716 35176
rect 12768 35164 12774 35216
rect 13262 35204 13268 35216
rect 12967 35176 13268 35204
rect 5074 35136 5080 35148
rect 5035 35108 5080 35136
rect 5074 35096 5080 35108
rect 5132 35096 5138 35148
rect 6089 35139 6147 35145
rect 6089 35105 6101 35139
rect 6135 35136 6147 35139
rect 6638 35136 6644 35148
rect 6135 35108 6644 35136
rect 6135 35105 6147 35108
rect 6089 35099 6147 35105
rect 6638 35096 6644 35108
rect 6696 35096 6702 35148
rect 7006 35096 7012 35148
rect 7064 35136 7070 35148
rect 7101 35139 7159 35145
rect 7101 35136 7113 35139
rect 7064 35108 7113 35136
rect 7064 35096 7070 35108
rect 7101 35105 7113 35108
rect 7147 35105 7159 35139
rect 7101 35099 7159 35105
rect 7834 35096 7840 35148
rect 7892 35136 7898 35148
rect 8938 35136 8944 35148
rect 7892 35108 8944 35136
rect 7892 35096 7898 35108
rect 8938 35096 8944 35108
rect 8996 35096 9002 35148
rect 9858 35136 9864 35148
rect 9819 35108 9864 35136
rect 9858 35096 9864 35108
rect 9916 35096 9922 35148
rect 10029 35139 10087 35145
rect 10029 35105 10041 35139
rect 10075 35136 10087 35139
rect 10075 35105 10088 35136
rect 10029 35099 10088 35105
rect 3418 35028 3424 35080
rect 3476 35068 3482 35080
rect 5994 35068 6000 35080
rect 3476 35040 5856 35068
rect 5955 35040 6000 35068
rect 3476 35028 3482 35040
rect 3881 35003 3939 35009
rect 3881 34969 3893 35003
rect 3927 35000 3939 35003
rect 5350 35000 5356 35012
rect 3927 34972 5356 35000
rect 3927 34969 3939 34972
rect 3881 34963 3939 34969
rect 5350 34960 5356 34972
rect 5408 34960 5414 35012
rect 5828 35000 5856 35040
rect 5994 35028 6000 35040
rect 6052 35028 6058 35080
rect 7377 35071 7435 35077
rect 7377 35068 7389 35071
rect 6932 35040 7389 35068
rect 6932 35000 6960 35040
rect 7377 35037 7389 35040
rect 7423 35068 7435 35071
rect 9030 35068 9036 35080
rect 7423 35040 9036 35068
rect 7423 35037 7435 35040
rect 7377 35031 7435 35037
rect 9030 35028 9036 35040
rect 9088 35028 9094 35080
rect 9122 35028 9128 35080
rect 9180 35068 9186 35080
rect 9398 35068 9404 35080
rect 9180 35040 9404 35068
rect 9180 35028 9186 35040
rect 9398 35028 9404 35040
rect 9456 35068 9462 35080
rect 9677 35071 9735 35077
rect 9677 35068 9689 35071
rect 9456 35040 9689 35068
rect 9456 35028 9462 35040
rect 9677 35037 9689 35040
rect 9723 35037 9735 35071
rect 9677 35031 9735 35037
rect 9858 35000 9864 35012
rect 5828 34972 6960 35000
rect 8036 34972 9864 35000
rect 1394 34892 1400 34944
rect 1452 34932 1458 34944
rect 1581 34935 1639 34941
rect 1581 34932 1593 34935
rect 1452 34904 1593 34932
rect 1452 34892 1458 34904
rect 1581 34901 1593 34904
rect 1627 34901 1639 34935
rect 3418 34932 3424 34944
rect 3379 34904 3424 34932
rect 1581 34895 1639 34901
rect 3418 34892 3424 34904
rect 3476 34892 3482 34944
rect 4982 34932 4988 34944
rect 4943 34904 4988 34932
rect 4982 34892 4988 34904
rect 5040 34892 5046 34944
rect 5258 34932 5264 34944
rect 5219 34904 5264 34932
rect 5258 34892 5264 34904
rect 5316 34892 5322 34944
rect 6273 34935 6331 34941
rect 6273 34901 6285 34935
rect 6319 34932 6331 34935
rect 6362 34932 6368 34944
rect 6319 34904 6368 34932
rect 6319 34901 6331 34904
rect 6273 34895 6331 34901
rect 6362 34892 6368 34904
rect 6420 34892 6426 34944
rect 6546 34932 6552 34944
rect 6507 34904 6552 34932
rect 6546 34892 6552 34904
rect 6604 34892 6610 34944
rect 6822 34892 6828 34944
rect 6880 34932 6886 34944
rect 7009 34935 7067 34941
rect 7009 34932 7021 34935
rect 6880 34904 7021 34932
rect 6880 34892 6886 34904
rect 7009 34901 7021 34904
rect 7055 34932 7067 34935
rect 8036 34932 8064 34972
rect 9858 34960 9864 34972
rect 9916 34960 9922 35012
rect 9950 34960 9956 35012
rect 10008 35000 10014 35012
rect 10060 35000 10088 35099
rect 10134 35096 10140 35148
rect 10192 35136 10198 35148
rect 10413 35139 10471 35145
rect 10413 35136 10425 35139
rect 10192 35108 10425 35136
rect 10192 35096 10198 35108
rect 10413 35105 10425 35108
rect 10459 35136 10471 35139
rect 11471 35139 11529 35145
rect 11471 35136 11483 35139
rect 10459 35108 11483 35136
rect 10459 35105 10471 35108
rect 10413 35099 10471 35105
rect 11471 35105 11483 35108
rect 11517 35105 11529 35139
rect 12802 35136 12808 35148
rect 12763 35108 12808 35136
rect 11471 35099 11529 35105
rect 12802 35096 12808 35108
rect 12860 35096 12866 35148
rect 12967 35145 12995 35176
rect 13262 35164 13268 35176
rect 13320 35164 13326 35216
rect 14734 35204 14740 35216
rect 13372 35176 14740 35204
rect 12952 35139 13010 35145
rect 12952 35105 12964 35139
rect 12998 35105 13010 35139
rect 13372 35136 13400 35176
rect 14734 35164 14740 35176
rect 14792 35164 14798 35216
rect 15102 35164 15108 35216
rect 15160 35204 15166 35216
rect 15289 35207 15347 35213
rect 15289 35204 15301 35207
rect 15160 35176 15301 35204
rect 15160 35164 15166 35176
rect 15289 35173 15301 35176
rect 15335 35173 15347 35207
rect 15657 35207 15715 35213
rect 15657 35204 15669 35207
rect 15289 35167 15347 35173
rect 15396 35176 15669 35204
rect 12952 35099 13010 35105
rect 13077 35108 13400 35136
rect 14461 35139 14519 35145
rect 10594 35028 10600 35080
rect 10652 35068 10658 35080
rect 11609 35071 11667 35077
rect 11609 35068 11621 35071
rect 10652 35040 11621 35068
rect 10652 35028 10658 35040
rect 11609 35037 11621 35040
rect 11655 35068 11667 35071
rect 13077 35068 13105 35108
rect 14461 35105 14473 35139
rect 14507 35136 14519 35139
rect 14550 35136 14556 35148
rect 14507 35108 14556 35136
rect 14507 35105 14519 35108
rect 14461 35099 14519 35105
rect 14550 35096 14556 35108
rect 14608 35096 14614 35148
rect 11655 35040 13105 35068
rect 13173 35071 13231 35077
rect 11655 35037 11667 35040
rect 11609 35031 11667 35037
rect 13173 35037 13185 35071
rect 13219 35068 13231 35071
rect 13998 35068 14004 35080
rect 13219 35040 14004 35068
rect 13219 35037 13231 35040
rect 13173 35031 13231 35037
rect 13998 35028 14004 35040
rect 14056 35028 14062 35080
rect 14274 35028 14280 35080
rect 14332 35068 14338 35080
rect 15396 35068 15424 35176
rect 15657 35173 15669 35176
rect 15703 35204 15715 35207
rect 16666 35204 16672 35216
rect 15703 35176 16672 35204
rect 15703 35173 15715 35176
rect 15657 35167 15715 35173
rect 16666 35164 16672 35176
rect 16724 35164 16730 35216
rect 17218 35204 17224 35216
rect 17179 35176 17224 35204
rect 17218 35164 17224 35176
rect 17276 35164 17282 35216
rect 17586 35204 17592 35216
rect 17547 35176 17592 35204
rect 17586 35164 17592 35176
rect 17644 35164 17650 35216
rect 18414 35204 18420 35216
rect 18375 35176 18420 35204
rect 18414 35164 18420 35176
rect 18472 35164 18478 35216
rect 19904 35204 19932 35232
rect 20438 35204 20444 35216
rect 19904 35176 20444 35204
rect 20438 35164 20444 35176
rect 20496 35164 20502 35216
rect 22278 35204 22284 35216
rect 21744 35176 22284 35204
rect 15473 35139 15531 35145
rect 15473 35136 15485 35139
rect 14332 35040 15424 35068
rect 15469 35105 15485 35136
rect 15519 35105 15531 35139
rect 15469 35099 15531 35105
rect 15565 35139 15623 35145
rect 15565 35105 15577 35139
rect 15611 35136 15623 35139
rect 16390 35136 16396 35148
rect 15611 35108 16396 35136
rect 15611 35105 15623 35108
rect 15565 35099 15623 35105
rect 14332 35028 14338 35040
rect 10008 34972 10088 35000
rect 10008 34960 10014 34972
rect 12066 34960 12072 35012
rect 12124 35000 12130 35012
rect 12526 35000 12532 35012
rect 12124 34972 12532 35000
rect 12124 34960 12130 34972
rect 12526 34960 12532 34972
rect 12584 34960 12590 35012
rect 12710 34960 12716 35012
rect 12768 35000 12774 35012
rect 15469 35000 15497 35099
rect 16390 35096 16396 35108
rect 16448 35096 16454 35148
rect 17037 35139 17095 35145
rect 17037 35136 17049 35139
rect 16592 35108 17049 35136
rect 15654 35028 15660 35080
rect 15712 35068 15718 35080
rect 16025 35071 16083 35077
rect 16025 35068 16037 35071
rect 15712 35040 16037 35068
rect 15712 35028 15718 35040
rect 16025 35037 16037 35040
rect 16071 35037 16083 35071
rect 16025 35031 16083 35037
rect 16592 35012 16620 35108
rect 17037 35105 17049 35108
rect 17083 35105 17095 35139
rect 17037 35099 17095 35105
rect 17129 35139 17187 35145
rect 17129 35105 17141 35139
rect 17175 35105 17187 35139
rect 17129 35099 17187 35105
rect 19061 35139 19119 35145
rect 19061 35105 19073 35139
rect 19107 35136 19119 35139
rect 19426 35136 19432 35148
rect 19107 35108 19432 35136
rect 19107 35105 19119 35108
rect 19061 35099 19119 35105
rect 16850 35068 16856 35080
rect 16811 35040 16856 35068
rect 16850 35028 16856 35040
rect 16908 35028 16914 35080
rect 16574 35000 16580 35012
rect 12768 34972 16580 35000
rect 12768 34960 12774 34972
rect 16574 34960 16580 34972
rect 16632 34960 16638 35012
rect 16758 34960 16764 35012
rect 16816 35000 16822 35012
rect 17144 35000 17172 35099
rect 19426 35096 19432 35108
rect 19484 35096 19490 35148
rect 21744 35145 21772 35176
rect 22278 35164 22284 35176
rect 22336 35164 22342 35216
rect 21729 35139 21787 35145
rect 21729 35105 21741 35139
rect 21775 35105 21787 35139
rect 22002 35136 22008 35148
rect 21963 35108 22008 35136
rect 21729 35099 21787 35105
rect 22002 35096 22008 35108
rect 22060 35096 22066 35148
rect 23382 35136 23388 35148
rect 23343 35108 23388 35136
rect 23382 35096 23388 35108
rect 23440 35096 23446 35148
rect 21177 35071 21235 35077
rect 21177 35037 21189 35071
rect 21223 35068 21235 35071
rect 21634 35068 21640 35080
rect 21223 35040 21640 35068
rect 21223 35037 21235 35040
rect 21177 35031 21235 35037
rect 21634 35028 21640 35040
rect 21692 35028 21698 35080
rect 22186 35068 22192 35080
rect 22147 35040 22192 35068
rect 22186 35028 22192 35040
rect 22244 35028 22250 35080
rect 23109 35071 23167 35077
rect 23109 35068 23121 35071
rect 23032 35040 23121 35068
rect 16816 34972 17172 35000
rect 16816 34960 16822 34972
rect 23032 34944 23060 35040
rect 23109 35037 23121 35040
rect 23155 35037 23167 35071
rect 23109 35031 23167 35037
rect 8662 34932 8668 34944
rect 7055 34904 8064 34932
rect 8623 34904 8668 34932
rect 7055 34901 7067 34904
rect 7009 34895 7067 34901
rect 8662 34892 8668 34904
rect 8720 34892 8726 34944
rect 8938 34892 8944 34944
rect 8996 34932 9002 34944
rect 11422 34941 11428 34944
rect 9401 34935 9459 34941
rect 9401 34932 9413 34935
rect 8996 34904 9413 34932
rect 8996 34892 9002 34904
rect 9401 34901 9413 34904
rect 9447 34901 9459 34935
rect 9401 34895 9459 34901
rect 11406 34935 11428 34941
rect 11406 34901 11418 34935
rect 11406 34895 11428 34901
rect 11422 34892 11428 34895
rect 11480 34892 11486 34944
rect 11698 34892 11704 34944
rect 11756 34932 11762 34944
rect 12434 34932 12440 34944
rect 11756 34904 12440 34932
rect 11756 34892 11762 34904
rect 12434 34892 12440 34904
rect 12492 34932 12498 34944
rect 13081 34935 13139 34941
rect 13081 34932 13093 34935
rect 12492 34904 13093 34932
rect 12492 34892 12498 34904
rect 13081 34901 13093 34904
rect 13127 34901 13139 34935
rect 13081 34895 13139 34901
rect 13814 34892 13820 34944
rect 13872 34932 13878 34944
rect 14001 34935 14059 34941
rect 14001 34932 14013 34935
rect 13872 34904 14013 34932
rect 13872 34892 13878 34904
rect 14001 34901 14013 34904
rect 14047 34932 14059 34935
rect 14185 34935 14243 34941
rect 14185 34932 14197 34935
rect 14047 34904 14197 34932
rect 14047 34901 14059 34904
rect 14001 34895 14059 34901
rect 14185 34901 14197 34904
rect 14231 34901 14243 34935
rect 14185 34895 14243 34901
rect 15105 34935 15163 34941
rect 15105 34901 15117 34935
rect 15151 34932 15163 34935
rect 15286 34932 15292 34944
rect 15151 34904 15292 34932
rect 15151 34901 15163 34904
rect 15105 34895 15163 34901
rect 15286 34892 15292 34904
rect 15344 34932 15350 34944
rect 16666 34932 16672 34944
rect 15344 34904 16672 34932
rect 15344 34892 15350 34904
rect 16666 34892 16672 34904
rect 16724 34932 16730 34944
rect 17494 34932 17500 34944
rect 16724 34904 17500 34932
rect 16724 34892 16730 34904
rect 17494 34892 17500 34904
rect 17552 34892 17558 34944
rect 22462 34932 22468 34944
rect 22423 34904 22468 34932
rect 22462 34892 22468 34904
rect 22520 34892 22526 34944
rect 23014 34932 23020 34944
rect 22975 34904 23020 34932
rect 23014 34892 23020 34904
rect 23072 34892 23078 34944
rect 23474 34892 23480 34944
rect 23532 34932 23538 34944
rect 24489 34935 24547 34941
rect 24489 34932 24501 34935
rect 23532 34904 24501 34932
rect 23532 34892 23538 34904
rect 24489 34901 24501 34904
rect 24535 34901 24547 34935
rect 24489 34895 24547 34901
rect 24946 34892 24952 34944
rect 25004 34932 25010 34944
rect 25498 34932 25504 34944
rect 25004 34904 25504 34932
rect 25004 34892 25010 34904
rect 25498 34892 25504 34904
rect 25556 34892 25562 34944
rect 26237 34935 26295 34941
rect 26237 34901 26249 34935
rect 26283 34932 26295 34935
rect 26326 34932 26332 34944
rect 26283 34904 26332 34932
rect 26283 34901 26295 34904
rect 26237 34895 26295 34901
rect 26326 34892 26332 34904
rect 26384 34892 26390 34944
rect 1104 34842 28888 34864
rect 1104 34790 5982 34842
rect 6034 34790 6046 34842
rect 6098 34790 6110 34842
rect 6162 34790 6174 34842
rect 6226 34790 15982 34842
rect 16034 34790 16046 34842
rect 16098 34790 16110 34842
rect 16162 34790 16174 34842
rect 16226 34790 25982 34842
rect 26034 34790 26046 34842
rect 26098 34790 26110 34842
rect 26162 34790 26174 34842
rect 26226 34790 28888 34842
rect 1104 34768 28888 34790
rect 4522 34728 4528 34740
rect 4483 34700 4528 34728
rect 4522 34688 4528 34700
rect 4580 34688 4586 34740
rect 4982 34688 4988 34740
rect 5040 34728 5046 34740
rect 11238 34728 11244 34740
rect 5040 34700 11244 34728
rect 5040 34688 5046 34700
rect 11238 34688 11244 34700
rect 11296 34688 11302 34740
rect 12158 34728 12164 34740
rect 12119 34700 12164 34728
rect 12158 34688 12164 34700
rect 12216 34728 12222 34740
rect 12216 34700 12480 34728
rect 12216 34688 12222 34700
rect 5074 34660 5080 34672
rect 5035 34632 5080 34660
rect 5074 34620 5080 34632
rect 5132 34620 5138 34672
rect 5997 34663 6055 34669
rect 5997 34660 6009 34663
rect 5460 34632 6009 34660
rect 3878 34592 3884 34604
rect 3839 34564 3884 34592
rect 3878 34552 3884 34564
rect 3936 34552 3942 34604
rect 4982 34552 4988 34604
rect 5040 34592 5046 34604
rect 5350 34592 5356 34604
rect 5040 34564 5356 34592
rect 5040 34552 5046 34564
rect 5350 34552 5356 34564
rect 5408 34552 5414 34604
rect 1394 34524 1400 34536
rect 1355 34496 1400 34524
rect 1394 34484 1400 34496
rect 1452 34484 1458 34536
rect 1670 34524 1676 34536
rect 1631 34496 1676 34524
rect 1670 34484 1676 34496
rect 1728 34484 1734 34536
rect 3513 34527 3571 34533
rect 3513 34493 3525 34527
rect 3559 34524 3571 34527
rect 3970 34524 3976 34536
rect 3559 34496 3976 34524
rect 3559 34493 3571 34496
rect 3513 34487 3571 34493
rect 3970 34484 3976 34496
rect 4028 34484 4034 34536
rect 4249 34527 4307 34533
rect 4249 34493 4261 34527
rect 4295 34524 4307 34527
rect 4341 34527 4399 34533
rect 4341 34524 4353 34527
rect 4295 34496 4353 34524
rect 4295 34493 4307 34496
rect 4249 34487 4307 34493
rect 4341 34493 4353 34496
rect 4387 34524 4399 34527
rect 5258 34524 5264 34536
rect 4387 34496 5264 34524
rect 4387 34493 4399 34496
rect 4341 34487 4399 34493
rect 5258 34484 5264 34496
rect 5316 34484 5322 34536
rect 5460 34533 5488 34632
rect 5997 34629 6009 34632
rect 6043 34629 6055 34663
rect 6638 34660 6644 34672
rect 6599 34632 6644 34660
rect 5997 34623 6055 34629
rect 6638 34620 6644 34632
rect 6696 34620 6702 34672
rect 9769 34663 9827 34669
rect 6748 34632 8984 34660
rect 5902 34592 5908 34604
rect 5863 34564 5908 34592
rect 5902 34552 5908 34564
rect 5960 34552 5966 34604
rect 6546 34592 6552 34604
rect 6012 34564 6552 34592
rect 5445 34527 5503 34533
rect 5445 34493 5457 34527
rect 5491 34493 5503 34527
rect 6012 34524 6040 34564
rect 6546 34552 6552 34564
rect 6604 34592 6610 34604
rect 6748 34592 6776 34632
rect 8956 34604 8984 34632
rect 9769 34629 9781 34663
rect 9815 34660 9827 34663
rect 10042 34660 10048 34672
rect 9815 34632 10048 34660
rect 9815 34629 9827 34632
rect 9769 34623 9827 34629
rect 10042 34620 10048 34632
rect 10100 34660 10106 34672
rect 10100 34632 10824 34660
rect 10100 34620 10106 34632
rect 6604 34564 6776 34592
rect 6604 34552 6610 34564
rect 6914 34552 6920 34604
rect 6972 34592 6978 34604
rect 7837 34595 7895 34601
rect 7837 34592 7849 34595
rect 6972 34564 7849 34592
rect 6972 34552 6978 34564
rect 7837 34561 7849 34564
rect 7883 34561 7895 34595
rect 8110 34592 8116 34604
rect 8071 34564 8116 34592
rect 7837 34555 7895 34561
rect 5445 34487 5503 34493
rect 5552 34496 6040 34524
rect 4614 34416 4620 34468
rect 4672 34456 4678 34468
rect 5552 34456 5580 34496
rect 6362 34484 6368 34536
rect 6420 34524 6426 34536
rect 7009 34527 7067 34533
rect 7009 34524 7021 34527
rect 6420 34496 7021 34524
rect 6420 34484 6426 34496
rect 7009 34493 7021 34496
rect 7055 34524 7067 34527
rect 7561 34527 7619 34533
rect 7561 34524 7573 34527
rect 7055 34496 7573 34524
rect 7055 34493 7067 34496
rect 7009 34487 7067 34493
rect 7561 34493 7573 34496
rect 7607 34524 7619 34527
rect 7650 34524 7656 34536
rect 7607 34496 7656 34524
rect 7607 34493 7619 34496
rect 7561 34487 7619 34493
rect 7650 34484 7656 34496
rect 7708 34484 7714 34536
rect 7852 34524 7880 34555
rect 8110 34552 8116 34564
rect 8168 34552 8174 34604
rect 8938 34592 8944 34604
rect 8899 34564 8944 34592
rect 8938 34552 8944 34564
rect 8996 34552 9002 34604
rect 9490 34552 9496 34604
rect 9548 34592 9554 34604
rect 10134 34592 10140 34604
rect 9548 34564 10140 34592
rect 9548 34552 9554 34564
rect 10134 34552 10140 34564
rect 10192 34552 10198 34604
rect 10318 34552 10324 34604
rect 10376 34592 10382 34604
rect 10796 34592 10824 34632
rect 11330 34620 11336 34672
rect 11388 34660 11394 34672
rect 11606 34660 11612 34672
rect 11388 34632 11612 34660
rect 11388 34620 11394 34632
rect 11606 34620 11612 34632
rect 11664 34620 11670 34672
rect 11698 34620 11704 34672
rect 11756 34660 11762 34672
rect 11882 34660 11888 34672
rect 11756 34632 11888 34660
rect 11756 34620 11762 34632
rect 11882 34620 11888 34632
rect 11940 34620 11946 34672
rect 10376 34564 10732 34592
rect 10796 34564 12204 34592
rect 10376 34552 10382 34564
rect 8294 34524 8300 34536
rect 7852 34496 8300 34524
rect 8294 34484 8300 34496
rect 8352 34484 8358 34536
rect 8478 34524 8484 34536
rect 8439 34496 8484 34524
rect 8478 34484 8484 34496
rect 8536 34484 8542 34536
rect 8662 34524 8668 34536
rect 8623 34496 8668 34524
rect 8662 34484 8668 34496
rect 8720 34484 8726 34536
rect 9030 34524 9036 34536
rect 8991 34496 9036 34524
rect 9030 34484 9036 34496
rect 9088 34524 9094 34536
rect 10045 34527 10103 34533
rect 10045 34524 10057 34527
rect 9088 34496 10057 34524
rect 9088 34484 9094 34496
rect 10045 34493 10057 34496
rect 10091 34493 10103 34527
rect 10502 34524 10508 34536
rect 10463 34496 10508 34524
rect 10045 34487 10103 34493
rect 10502 34484 10508 34496
rect 10560 34484 10566 34536
rect 10704 34533 10732 34564
rect 10689 34527 10747 34533
rect 10689 34493 10701 34527
rect 10735 34493 10747 34527
rect 10689 34487 10747 34493
rect 10873 34527 10931 34533
rect 10873 34493 10885 34527
rect 10919 34493 10931 34527
rect 10873 34487 10931 34493
rect 7098 34456 7104 34468
rect 4672 34428 5580 34456
rect 5920 34428 7104 34456
rect 4672 34416 4678 34428
rect 2774 34348 2780 34400
rect 2832 34388 2838 34400
rect 2832 34360 2877 34388
rect 2832 34348 2838 34360
rect 5166 34348 5172 34400
rect 5224 34388 5230 34400
rect 5920 34388 5948 34428
rect 7098 34416 7104 34428
rect 7156 34456 7162 34468
rect 7156 34428 7236 34456
rect 7156 34416 7162 34428
rect 5224 34360 5948 34388
rect 5997 34391 6055 34397
rect 5224 34348 5230 34360
rect 5997 34357 6009 34391
rect 6043 34388 6055 34391
rect 6273 34391 6331 34397
rect 6273 34388 6285 34391
rect 6043 34360 6285 34388
rect 6043 34357 6055 34360
rect 5997 34351 6055 34357
rect 6273 34357 6285 34360
rect 6319 34388 6331 34391
rect 6546 34388 6552 34400
rect 6319 34360 6552 34388
rect 6319 34357 6331 34360
rect 6273 34351 6331 34357
rect 6546 34348 6552 34360
rect 6604 34348 6610 34400
rect 7208 34397 7236 34428
rect 10778 34416 10784 34468
rect 10836 34456 10842 34468
rect 10888 34456 10916 34487
rect 12176 34468 12204 34564
rect 12452 34524 12480 34700
rect 14182 34688 14188 34740
rect 14240 34688 14246 34740
rect 14550 34688 14556 34740
rect 14608 34728 14614 34740
rect 15010 34728 15016 34740
rect 14608 34700 15016 34728
rect 14608 34688 14614 34700
rect 15010 34688 15016 34700
rect 15068 34688 15074 34740
rect 15102 34688 15108 34740
rect 15160 34728 15166 34740
rect 15289 34731 15347 34737
rect 15289 34728 15301 34731
rect 15160 34700 15301 34728
rect 15160 34688 15166 34700
rect 15289 34697 15301 34700
rect 15335 34697 15347 34731
rect 15289 34691 15347 34697
rect 16574 34688 16580 34740
rect 16632 34728 16638 34740
rect 16761 34731 16819 34737
rect 16761 34728 16773 34731
rect 16632 34700 16773 34728
rect 16632 34688 16638 34700
rect 16761 34697 16773 34700
rect 16807 34728 16819 34731
rect 17129 34731 17187 34737
rect 17129 34728 17141 34731
rect 16807 34700 17141 34728
rect 16807 34697 16819 34700
rect 16761 34691 16819 34697
rect 17129 34697 17141 34700
rect 17175 34697 17187 34731
rect 17129 34691 17187 34697
rect 17865 34731 17923 34737
rect 17865 34697 17877 34731
rect 17911 34728 17923 34731
rect 18414 34728 18420 34740
rect 17911 34700 18420 34728
rect 17911 34697 17923 34700
rect 17865 34691 17923 34697
rect 18414 34688 18420 34700
rect 18472 34688 18478 34740
rect 19426 34728 19432 34740
rect 19387 34700 19432 34728
rect 19426 34688 19432 34700
rect 19484 34688 19490 34740
rect 20070 34688 20076 34740
rect 20128 34728 20134 34740
rect 20257 34731 20315 34737
rect 20257 34728 20269 34731
rect 20128 34700 20269 34728
rect 20128 34688 20134 34700
rect 20257 34697 20269 34700
rect 20303 34697 20315 34731
rect 20257 34691 20315 34697
rect 21913 34731 21971 34737
rect 21913 34697 21925 34731
rect 21959 34728 21971 34731
rect 22002 34728 22008 34740
rect 21959 34700 22008 34728
rect 21959 34697 21971 34700
rect 21913 34691 21971 34697
rect 22002 34688 22008 34700
rect 22060 34688 22066 34740
rect 22186 34688 22192 34740
rect 22244 34728 22250 34740
rect 22557 34731 22615 34737
rect 22557 34728 22569 34731
rect 22244 34700 22569 34728
rect 22244 34688 22250 34700
rect 22557 34697 22569 34700
rect 22603 34697 22615 34731
rect 22557 34691 22615 34697
rect 23109 34731 23167 34737
rect 23109 34697 23121 34731
rect 23155 34728 23167 34731
rect 23382 34728 23388 34740
rect 23155 34700 23388 34728
rect 23155 34697 23167 34700
rect 23109 34691 23167 34697
rect 23382 34688 23388 34700
rect 23440 34688 23446 34740
rect 24946 34728 24952 34740
rect 23492 34700 24952 34728
rect 12986 34620 12992 34672
rect 13044 34660 13050 34672
rect 14200 34660 14228 34688
rect 17770 34660 17776 34672
rect 13044 34632 17776 34660
rect 13044 34620 13050 34632
rect 17770 34620 17776 34632
rect 17828 34620 17834 34672
rect 18325 34663 18383 34669
rect 18325 34629 18337 34663
rect 18371 34629 18383 34663
rect 18325 34623 18383 34629
rect 13262 34592 13268 34604
rect 13223 34564 13268 34592
rect 13262 34552 13268 34564
rect 13320 34552 13326 34604
rect 14093 34595 14151 34601
rect 14093 34561 14105 34595
rect 14139 34592 14151 34595
rect 14185 34595 14243 34601
rect 14185 34592 14197 34595
rect 14139 34564 14197 34592
rect 14139 34561 14151 34564
rect 14093 34555 14151 34561
rect 14185 34561 14197 34564
rect 14231 34592 14243 34595
rect 14734 34592 14740 34604
rect 14231 34564 14740 34592
rect 14231 34561 14243 34564
rect 14185 34555 14243 34561
rect 14734 34552 14740 34564
rect 14792 34552 14798 34604
rect 16482 34592 16488 34604
rect 15948 34564 16488 34592
rect 15948 34536 15976 34564
rect 16482 34552 16488 34564
rect 16540 34552 16546 34604
rect 18046 34552 18052 34604
rect 18104 34592 18110 34604
rect 18340 34592 18368 34623
rect 18432 34601 18460 34688
rect 19981 34663 20039 34669
rect 19981 34629 19993 34663
rect 20027 34660 20039 34663
rect 22278 34660 22284 34672
rect 20027 34632 21404 34660
rect 22191 34632 22284 34660
rect 20027 34629 20039 34632
rect 19981 34623 20039 34629
rect 18104 34564 18368 34592
rect 18417 34595 18475 34601
rect 18104 34552 18110 34564
rect 18417 34561 18429 34595
rect 18463 34561 18475 34595
rect 19058 34592 19064 34604
rect 19019 34564 19064 34592
rect 18417 34555 18475 34561
rect 19058 34552 19064 34564
rect 19116 34552 19122 34604
rect 20530 34592 20536 34604
rect 20491 34564 20536 34592
rect 20530 34552 20536 34564
rect 20588 34552 20594 34604
rect 12529 34527 12587 34533
rect 12529 34524 12541 34527
rect 12452 34496 12541 34524
rect 12529 34493 12541 34496
rect 12575 34493 12587 34527
rect 12710 34524 12716 34536
rect 12671 34496 12716 34524
rect 12529 34487 12587 34493
rect 12710 34484 12716 34496
rect 12768 34484 12774 34536
rect 12881 34527 12939 34533
rect 12881 34493 12893 34527
rect 12927 34524 12939 34527
rect 13078 34524 13084 34536
rect 12927 34496 13084 34524
rect 12927 34493 12939 34496
rect 12881 34487 12939 34493
rect 13078 34484 13084 34496
rect 13136 34484 13142 34536
rect 14366 34524 14372 34536
rect 14327 34496 14372 34524
rect 14366 34484 14372 34496
rect 14424 34524 14430 34536
rect 14921 34527 14979 34533
rect 14424 34496 14688 34524
rect 14424 34484 14430 34496
rect 11974 34456 11980 34468
rect 10836 34428 11980 34456
rect 10836 34416 10842 34428
rect 11974 34416 11980 34428
rect 12032 34416 12038 34468
rect 12158 34416 12164 34468
rect 12216 34456 12222 34468
rect 12342 34456 12348 34468
rect 12216 34428 12348 34456
rect 12216 34416 12222 34428
rect 12342 34416 12348 34428
rect 12400 34416 12406 34468
rect 12434 34416 12440 34468
rect 12492 34456 12498 34468
rect 13541 34459 13599 34465
rect 13541 34456 13553 34459
rect 12492 34428 13553 34456
rect 12492 34416 12498 34428
rect 13541 34425 13553 34428
rect 13587 34425 13599 34459
rect 13541 34419 13599 34425
rect 13814 34416 13820 34468
rect 13872 34456 13878 34468
rect 14550 34456 14556 34468
rect 13872 34428 14556 34456
rect 13872 34416 13878 34428
rect 14550 34416 14556 34428
rect 14608 34416 14614 34468
rect 14660 34456 14688 34496
rect 14921 34493 14933 34527
rect 14967 34524 14979 34527
rect 15102 34524 15108 34536
rect 14967 34496 15108 34524
rect 14967 34493 14979 34496
rect 14921 34487 14979 34493
rect 15102 34484 15108 34496
rect 15160 34484 15166 34536
rect 15749 34527 15807 34533
rect 15749 34493 15761 34527
rect 15795 34524 15807 34527
rect 15930 34524 15936 34536
rect 15795 34496 15936 34524
rect 15795 34493 15807 34496
rect 15749 34487 15807 34493
rect 15930 34484 15936 34496
rect 15988 34484 15994 34536
rect 18196 34527 18254 34533
rect 18196 34493 18208 34527
rect 18242 34524 18254 34527
rect 18874 34524 18880 34536
rect 18242 34496 18880 34524
rect 18242 34493 18254 34496
rect 18196 34487 18254 34493
rect 18874 34484 18880 34496
rect 18932 34484 18938 34536
rect 20070 34484 20076 34536
rect 20128 34524 20134 34536
rect 20254 34524 20260 34536
rect 20128 34496 20260 34524
rect 20128 34484 20134 34496
rect 20254 34484 20260 34496
rect 20312 34524 20318 34536
rect 21376 34533 21404 34632
rect 22278 34620 22284 34632
rect 22336 34660 22342 34672
rect 23492 34660 23520 34700
rect 24946 34688 24952 34700
rect 25004 34688 25010 34740
rect 25314 34688 25320 34740
rect 25372 34728 25378 34740
rect 25961 34731 26019 34737
rect 25961 34728 25973 34731
rect 25372 34700 25973 34728
rect 25372 34688 25378 34700
rect 25961 34697 25973 34700
rect 26007 34697 26019 34731
rect 27706 34728 27712 34740
rect 27667 34700 27712 34728
rect 25961 34691 26019 34697
rect 22336 34632 23520 34660
rect 22336 34620 22342 34632
rect 21542 34592 21548 34604
rect 21503 34564 21548 34592
rect 21542 34552 21548 34564
rect 21600 34552 21606 34604
rect 23477 34595 23535 34601
rect 23477 34561 23489 34595
rect 23523 34592 23535 34595
rect 25038 34592 25044 34604
rect 23523 34564 23796 34592
rect 24999 34564 25044 34592
rect 23523 34561 23535 34564
rect 23477 34555 23535 34561
rect 23768 34536 23796 34564
rect 25038 34552 25044 34564
rect 25096 34552 25102 34604
rect 25976 34592 26004 34691
rect 27706 34688 27712 34700
rect 27764 34688 27770 34740
rect 26421 34595 26479 34601
rect 26421 34592 26433 34595
rect 25976 34564 26433 34592
rect 26421 34561 26433 34564
rect 26467 34561 26479 34595
rect 26421 34555 26479 34561
rect 20809 34527 20867 34533
rect 20809 34524 20821 34527
rect 20312 34496 20821 34524
rect 20312 34484 20318 34496
rect 20809 34493 20821 34496
rect 20855 34493 20867 34527
rect 20809 34487 20867 34493
rect 21361 34527 21419 34533
rect 21361 34493 21373 34527
rect 21407 34524 21419 34527
rect 21634 34524 21640 34536
rect 21407 34496 21640 34524
rect 21407 34493 21419 34496
rect 21361 34487 21419 34493
rect 21634 34484 21640 34496
rect 21692 34484 21698 34536
rect 23014 34484 23020 34536
rect 23072 34524 23078 34536
rect 23661 34527 23719 34533
rect 23661 34524 23673 34527
rect 23072 34496 23673 34524
rect 23072 34484 23078 34496
rect 23661 34493 23673 34496
rect 23707 34493 23719 34527
rect 23661 34487 23719 34493
rect 14660 34428 14964 34456
rect 7193 34391 7251 34397
rect 7193 34357 7205 34391
rect 7239 34357 7251 34391
rect 7193 34351 7251 34357
rect 9122 34348 9128 34400
rect 9180 34388 9186 34400
rect 10318 34388 10324 34400
rect 9180 34360 10324 34388
rect 9180 34348 9186 34360
rect 10318 34348 10324 34360
rect 10376 34388 10382 34400
rect 11333 34391 11391 34397
rect 11333 34388 11345 34391
rect 10376 34360 11345 34388
rect 10376 34348 10382 34360
rect 11333 34357 11345 34360
rect 11379 34357 11391 34391
rect 11333 34351 11391 34357
rect 11885 34391 11943 34397
rect 11885 34357 11897 34391
rect 11931 34388 11943 34391
rect 12802 34388 12808 34400
rect 11931 34360 12808 34388
rect 11931 34357 11943 34360
rect 11885 34351 11943 34357
rect 12802 34348 12808 34360
rect 12860 34348 12866 34400
rect 14461 34391 14519 34397
rect 14461 34357 14473 34391
rect 14507 34388 14519 34391
rect 14826 34388 14832 34400
rect 14507 34360 14832 34388
rect 14507 34357 14519 34360
rect 14461 34351 14519 34357
rect 14826 34348 14832 34360
rect 14884 34348 14890 34400
rect 14936 34388 14964 34428
rect 15010 34416 15016 34468
rect 15068 34456 15074 34468
rect 15562 34456 15568 34468
rect 15068 34428 15568 34456
rect 15068 34416 15074 34428
rect 15562 34416 15568 34428
rect 15620 34456 15626 34468
rect 16117 34459 16175 34465
rect 16117 34456 16129 34459
rect 15620 34428 16129 34456
rect 15620 34416 15626 34428
rect 16117 34425 16129 34428
rect 16163 34425 16175 34459
rect 16482 34456 16488 34468
rect 16443 34428 16488 34456
rect 16117 34419 16175 34425
rect 16482 34416 16488 34428
rect 16540 34416 16546 34468
rect 17954 34416 17960 34468
rect 18012 34456 18018 34468
rect 18049 34459 18107 34465
rect 18049 34456 18061 34459
rect 18012 34428 18061 34456
rect 18012 34416 18018 34428
rect 18049 34425 18061 34428
rect 18095 34425 18107 34459
rect 18049 34419 18107 34425
rect 19610 34416 19616 34468
rect 19668 34456 19674 34468
rect 20714 34456 20720 34468
rect 19668 34428 20720 34456
rect 19668 34416 19674 34428
rect 20714 34416 20720 34428
rect 20772 34416 20778 34468
rect 20898 34416 20904 34468
rect 20956 34456 20962 34468
rect 20956 34428 21680 34456
rect 20956 34416 20962 34428
rect 21652 34400 21680 34428
rect 15933 34391 15991 34397
rect 15933 34388 15945 34391
rect 14936 34360 15945 34388
rect 15933 34357 15945 34360
rect 15979 34357 15991 34391
rect 15933 34351 15991 34357
rect 16025 34391 16083 34397
rect 16025 34357 16037 34391
rect 16071 34388 16083 34391
rect 16666 34388 16672 34400
rect 16071 34360 16672 34388
rect 16071 34357 16083 34360
rect 16025 34351 16083 34357
rect 16666 34348 16672 34360
rect 16724 34348 16730 34400
rect 16942 34348 16948 34400
rect 17000 34388 17006 34400
rect 17218 34388 17224 34400
rect 17000 34360 17224 34388
rect 17000 34348 17006 34360
rect 17218 34348 17224 34360
rect 17276 34348 17282 34400
rect 18506 34348 18512 34400
rect 18564 34388 18570 34400
rect 18693 34391 18751 34397
rect 18693 34388 18705 34391
rect 18564 34360 18705 34388
rect 18564 34348 18570 34360
rect 18693 34357 18705 34360
rect 18739 34357 18751 34391
rect 18693 34351 18751 34357
rect 21634 34348 21640 34400
rect 21692 34348 21698 34400
rect 23676 34388 23704 34487
rect 23750 34484 23756 34536
rect 23808 34524 23814 34536
rect 23937 34527 23995 34533
rect 23937 34524 23949 34527
rect 23808 34496 23949 34524
rect 23808 34484 23814 34496
rect 23937 34493 23949 34496
rect 23983 34493 23995 34527
rect 23937 34487 23995 34493
rect 26145 34527 26203 34533
rect 26145 34493 26157 34527
rect 26191 34524 26203 34527
rect 26234 34524 26240 34536
rect 26191 34496 26240 34524
rect 26191 34493 26203 34496
rect 26145 34487 26203 34493
rect 26234 34484 26240 34496
rect 26292 34484 26298 34536
rect 24302 34388 24308 34400
rect 23676 34360 24308 34388
rect 24302 34348 24308 34360
rect 24360 34348 24366 34400
rect 1104 34298 28888 34320
rect 1104 34246 10982 34298
rect 11034 34246 11046 34298
rect 11098 34246 11110 34298
rect 11162 34246 11174 34298
rect 11226 34246 20982 34298
rect 21034 34246 21046 34298
rect 21098 34246 21110 34298
rect 21162 34246 21174 34298
rect 21226 34246 28888 34298
rect 1104 34224 28888 34246
rect 1670 34184 1676 34196
rect 1631 34156 1676 34184
rect 1670 34144 1676 34156
rect 1728 34144 1734 34196
rect 3418 34184 3424 34196
rect 3379 34156 3424 34184
rect 3418 34144 3424 34156
rect 3476 34144 3482 34196
rect 4338 34184 4344 34196
rect 4299 34156 4344 34184
rect 4338 34144 4344 34156
rect 4396 34144 4402 34196
rect 4614 34184 4620 34196
rect 4575 34156 4620 34184
rect 4614 34144 4620 34156
rect 4672 34144 4678 34196
rect 4985 34187 5043 34193
rect 4985 34153 4997 34187
rect 5031 34184 5043 34187
rect 5442 34184 5448 34196
rect 5031 34156 5448 34184
rect 5031 34153 5043 34156
rect 4985 34147 5043 34153
rect 5442 34144 5448 34156
rect 5500 34144 5506 34196
rect 5629 34187 5687 34193
rect 5629 34153 5641 34187
rect 5675 34184 5687 34187
rect 6362 34184 6368 34196
rect 5675 34156 6368 34184
rect 5675 34153 5687 34156
rect 5629 34147 5687 34153
rect 6362 34144 6368 34156
rect 6420 34144 6426 34196
rect 6549 34187 6607 34193
rect 6549 34153 6561 34187
rect 6595 34184 6607 34187
rect 6822 34184 6828 34196
rect 6595 34156 6828 34184
rect 6595 34153 6607 34156
rect 6549 34147 6607 34153
rect 6822 34144 6828 34156
rect 6880 34144 6886 34196
rect 10226 34184 10232 34196
rect 9692 34156 10232 34184
rect 5350 34116 5356 34128
rect 5311 34088 5356 34116
rect 5350 34076 5356 34088
rect 5408 34076 5414 34128
rect 5534 34076 5540 34128
rect 5592 34116 5598 34128
rect 5721 34119 5779 34125
rect 5721 34116 5733 34119
rect 5592 34088 5733 34116
rect 5592 34076 5598 34088
rect 5721 34085 5733 34088
rect 5767 34085 5779 34119
rect 5721 34079 5779 34085
rect 5810 34076 5816 34128
rect 5868 34116 5874 34128
rect 9692 34125 9720 34156
rect 10226 34144 10232 34156
rect 10284 34144 10290 34196
rect 10502 34144 10508 34196
rect 10560 34144 10566 34196
rect 12158 34184 12164 34196
rect 12119 34156 12164 34184
rect 12158 34144 12164 34156
rect 12216 34144 12222 34196
rect 13538 34144 13544 34196
rect 13596 34184 13602 34196
rect 13909 34187 13967 34193
rect 13596 34156 13676 34184
rect 13596 34144 13602 34156
rect 9677 34119 9735 34125
rect 5868 34088 6868 34116
rect 5868 34076 5874 34088
rect 6840 34060 6868 34088
rect 9677 34085 9689 34119
rect 9723 34085 9735 34119
rect 10520 34116 10548 34144
rect 10870 34116 10876 34128
rect 10520 34088 10876 34116
rect 9677 34079 9735 34085
rect 4430 34048 4436 34060
rect 4391 34020 4436 34048
rect 4430 34008 4436 34020
rect 4488 34008 4494 34060
rect 5258 34008 5264 34060
rect 5316 34048 5322 34060
rect 5445 34051 5503 34057
rect 5445 34048 5457 34051
rect 5316 34020 5457 34048
rect 5316 34008 5322 34020
rect 5445 34017 5457 34020
rect 5491 34048 5503 34051
rect 6638 34048 6644 34060
rect 5491 34020 6644 34048
rect 5491 34017 5503 34020
rect 5445 34011 5503 34017
rect 6638 34008 6644 34020
rect 6696 34008 6702 34060
rect 6822 34008 6828 34060
rect 6880 34008 6886 34060
rect 9858 34008 9864 34060
rect 9916 34048 9922 34060
rect 10796 34057 10824 34088
rect 10870 34076 10876 34088
rect 10928 34076 10934 34128
rect 11974 34076 11980 34128
rect 12032 34116 12038 34128
rect 13648 34125 13676 34156
rect 13909 34153 13921 34187
rect 13955 34184 13967 34187
rect 14366 34184 14372 34196
rect 13955 34156 14372 34184
rect 13955 34153 13967 34156
rect 13909 34147 13967 34153
rect 14366 34144 14372 34156
rect 14424 34144 14430 34196
rect 16758 34184 16764 34196
rect 16719 34156 16764 34184
rect 16758 34144 16764 34156
rect 16816 34144 16822 34196
rect 16850 34144 16856 34196
rect 16908 34184 16914 34196
rect 17681 34187 17739 34193
rect 17681 34184 17693 34187
rect 16908 34156 17693 34184
rect 16908 34144 16914 34156
rect 17681 34153 17693 34156
rect 17727 34153 17739 34187
rect 18046 34184 18052 34196
rect 18007 34156 18052 34184
rect 17681 34147 17739 34153
rect 18046 34144 18052 34156
rect 18104 34144 18110 34196
rect 20257 34187 20315 34193
rect 20257 34153 20269 34187
rect 20303 34184 20315 34187
rect 20806 34184 20812 34196
rect 20303 34156 20812 34184
rect 20303 34153 20315 34156
rect 20257 34147 20315 34153
rect 20806 34144 20812 34156
rect 20864 34184 20870 34196
rect 22370 34184 22376 34196
rect 20864 34156 22232 34184
rect 22331 34156 22376 34184
rect 20864 34144 20870 34156
rect 12345 34119 12403 34125
rect 12345 34116 12357 34119
rect 12032 34088 12357 34116
rect 12032 34076 12038 34088
rect 12345 34085 12357 34088
rect 12391 34085 12403 34119
rect 12345 34079 12403 34085
rect 13633 34119 13691 34125
rect 13633 34085 13645 34119
rect 13679 34085 13691 34119
rect 13633 34079 13691 34085
rect 14001 34119 14059 34125
rect 14001 34085 14013 34119
rect 14047 34116 14059 34119
rect 14182 34116 14188 34128
rect 14047 34088 14188 34116
rect 14047 34085 14059 34088
rect 14001 34079 14059 34085
rect 14182 34076 14188 34088
rect 14240 34076 14246 34128
rect 14274 34076 14280 34128
rect 14332 34116 14338 34128
rect 14645 34119 14703 34125
rect 14645 34116 14657 34119
rect 14332 34088 14657 34116
rect 14332 34076 14338 34088
rect 14645 34085 14657 34088
rect 14691 34116 14703 34119
rect 14734 34116 14740 34128
rect 14691 34088 14740 34116
rect 14691 34085 14703 34088
rect 14645 34079 14703 34085
rect 14734 34076 14740 34088
rect 14792 34116 14798 34128
rect 15013 34119 15071 34125
rect 15013 34116 15025 34119
rect 14792 34088 15025 34116
rect 14792 34076 14798 34088
rect 15013 34085 15025 34088
rect 15059 34085 15071 34119
rect 15013 34079 15071 34085
rect 15102 34076 15108 34128
rect 15160 34116 15166 34128
rect 17954 34116 17960 34128
rect 15160 34088 15479 34116
rect 15160 34076 15166 34088
rect 10137 34051 10195 34057
rect 10137 34048 10149 34051
rect 9916 34020 10149 34048
rect 9916 34008 9922 34020
rect 10137 34017 10149 34020
rect 10183 34017 10195 34051
rect 10137 34011 10195 34017
rect 10321 34051 10379 34057
rect 10321 34017 10333 34051
rect 10367 34017 10379 34051
rect 10321 34011 10379 34017
rect 10597 34051 10655 34057
rect 10597 34017 10609 34051
rect 10643 34048 10655 34051
rect 10781 34051 10839 34057
rect 10643 34020 10732 34048
rect 10643 34017 10655 34020
rect 10597 34011 10655 34017
rect 6178 33980 6184 33992
rect 6139 33952 6184 33980
rect 6178 33940 6184 33952
rect 6236 33940 6242 33992
rect 7006 33980 7012 33992
rect 6967 33952 7012 33980
rect 7006 33940 7012 33952
rect 7064 33940 7070 33992
rect 7285 33983 7343 33989
rect 7285 33949 7297 33983
rect 7331 33980 7343 33983
rect 8110 33980 8116 33992
rect 7331 33952 8116 33980
rect 7331 33949 7343 33952
rect 7285 33943 7343 33949
rect 4982 33872 4988 33924
rect 5040 33912 5046 33924
rect 5040 33884 7052 33912
rect 5040 33872 5046 33884
rect 3786 33844 3792 33856
rect 3747 33816 3792 33844
rect 3786 33804 3792 33816
rect 3844 33804 3850 33856
rect 4522 33804 4528 33856
rect 4580 33844 4586 33856
rect 6914 33844 6920 33856
rect 4580 33816 6920 33844
rect 4580 33804 4586 33816
rect 6914 33804 6920 33816
rect 6972 33804 6978 33856
rect 7024 33844 7052 33884
rect 7944 33844 7972 33952
rect 8110 33940 8116 33952
rect 8168 33940 8174 33992
rect 8294 33940 8300 33992
rect 8352 33980 8358 33992
rect 9493 33983 9551 33989
rect 9493 33980 9505 33983
rect 8352 33952 9505 33980
rect 8352 33940 8358 33952
rect 9493 33949 9505 33952
rect 9539 33980 9551 33983
rect 9539 33952 9904 33980
rect 9539 33949 9551 33952
rect 9493 33943 9551 33949
rect 9876 33912 9904 33952
rect 9950 33940 9956 33992
rect 10008 33980 10014 33992
rect 10336 33980 10364 34011
rect 10008 33952 10364 33980
rect 10704 33980 10732 34020
rect 10781 34017 10793 34051
rect 10827 34017 10839 34051
rect 10781 34011 10839 34017
rect 11422 34008 11428 34060
rect 11480 34048 11486 34060
rect 12253 34051 12311 34057
rect 12253 34048 12265 34051
rect 11480 34020 12265 34048
rect 11480 34008 11486 34020
rect 12253 34017 12265 34020
rect 12299 34017 12311 34051
rect 12253 34011 12311 34017
rect 13541 34051 13599 34057
rect 13541 34017 13553 34051
rect 13587 34048 13599 34051
rect 13817 34051 13875 34057
rect 13817 34048 13829 34051
rect 13587 34020 13829 34048
rect 13587 34017 13599 34020
rect 13541 34011 13599 34017
rect 13817 34017 13829 34020
rect 13863 34048 13875 34051
rect 14292 34048 14320 34076
rect 15286 34048 15292 34060
rect 13863 34020 14320 34048
rect 15247 34020 15292 34048
rect 13863 34017 13875 34020
rect 13817 34011 13875 34017
rect 15286 34008 15292 34020
rect 15344 34008 15350 34060
rect 15451 34057 15479 34088
rect 16868 34088 17960 34116
rect 16868 34060 16896 34088
rect 17954 34076 17960 34088
rect 18012 34076 18018 34128
rect 21269 34119 21327 34125
rect 21269 34085 21281 34119
rect 21315 34116 21327 34119
rect 21634 34116 21640 34128
rect 21315 34088 21640 34116
rect 21315 34085 21327 34088
rect 21269 34079 21327 34085
rect 21634 34076 21640 34088
rect 21692 34076 21698 34128
rect 22204 34116 22232 34156
rect 22370 34144 22376 34156
rect 22428 34144 22434 34196
rect 23198 34116 23204 34128
rect 22204 34088 23204 34116
rect 23198 34076 23204 34088
rect 23256 34116 23262 34128
rect 23256 34088 23520 34116
rect 23256 34076 23262 34088
rect 15436 34051 15494 34057
rect 15436 34017 15448 34051
rect 15482 34048 15494 34051
rect 16666 34048 16672 34060
rect 15482 34020 16672 34048
rect 15482 34017 15494 34020
rect 15436 34011 15494 34017
rect 16666 34008 16672 34020
rect 16724 34008 16730 34060
rect 16850 34048 16856 34060
rect 16811 34020 16856 34048
rect 16850 34008 16856 34020
rect 16908 34008 16914 34060
rect 16942 34008 16948 34060
rect 17000 34048 17006 34060
rect 17037 34051 17095 34057
rect 17037 34048 17049 34051
rect 17000 34020 17049 34048
rect 17000 34008 17006 34020
rect 17037 34017 17049 34020
rect 17083 34017 17095 34051
rect 17037 34011 17095 34017
rect 18509 34051 18567 34057
rect 18509 34017 18521 34051
rect 18555 34048 18567 34051
rect 19242 34048 19248 34060
rect 18555 34020 19248 34048
rect 18555 34017 18567 34020
rect 18509 34011 18567 34017
rect 19242 34008 19248 34020
rect 19300 34008 19306 34060
rect 20714 34008 20720 34060
rect 20772 34048 20778 34060
rect 21085 34051 21143 34057
rect 21085 34048 21097 34051
rect 20772 34020 21097 34048
rect 20772 34008 20778 34020
rect 21085 34017 21097 34020
rect 21131 34017 21143 34051
rect 21085 34011 21143 34017
rect 21177 34051 21235 34057
rect 21177 34017 21189 34051
rect 21223 34048 21235 34051
rect 21358 34048 21364 34060
rect 21223 34020 21364 34048
rect 21223 34017 21235 34020
rect 21177 34011 21235 34017
rect 21358 34008 21364 34020
rect 21416 34008 21422 34060
rect 23382 34048 23388 34060
rect 23343 34020 23388 34048
rect 23382 34008 23388 34020
rect 23440 34008 23446 34060
rect 23492 34057 23520 34088
rect 23477 34051 23535 34057
rect 23477 34017 23489 34051
rect 23523 34017 23535 34051
rect 23477 34011 23535 34017
rect 25225 34051 25283 34057
rect 25225 34017 25237 34051
rect 25271 34048 25283 34051
rect 25314 34048 25320 34060
rect 25271 34020 25320 34048
rect 25271 34017 25283 34020
rect 25225 34011 25283 34017
rect 25314 34008 25320 34020
rect 25372 34008 25378 34060
rect 10962 33980 10968 33992
rect 10704 33952 10968 33980
rect 10008 33940 10014 33952
rect 10962 33940 10968 33952
rect 11020 33940 11026 33992
rect 11057 33983 11115 33989
rect 11057 33949 11069 33983
rect 11103 33949 11115 33983
rect 11057 33943 11115 33949
rect 11885 33983 11943 33989
rect 11885 33949 11897 33983
rect 11931 33980 11943 33983
rect 11977 33983 12035 33989
rect 11977 33980 11989 33983
rect 11931 33952 11989 33980
rect 11931 33949 11943 33952
rect 11885 33943 11943 33949
rect 11977 33949 11989 33952
rect 12023 33980 12035 33983
rect 12066 33980 12072 33992
rect 12023 33952 12072 33980
rect 12023 33949 12035 33952
rect 11977 33943 12035 33949
rect 11072 33912 11100 33943
rect 12066 33940 12072 33952
rect 12124 33940 12130 33992
rect 12713 33983 12771 33989
rect 12713 33949 12725 33983
rect 12759 33980 12771 33983
rect 13262 33980 13268 33992
rect 12759 33952 13268 33980
rect 12759 33949 12771 33952
rect 12713 33943 12771 33949
rect 13262 33940 13268 33952
rect 13320 33940 13326 33992
rect 14369 33983 14427 33989
rect 14369 33949 14381 33983
rect 14415 33980 14427 33983
rect 15657 33983 15715 33989
rect 14415 33952 15608 33980
rect 14415 33949 14427 33952
rect 14369 33943 14427 33949
rect 9876 33884 11100 33912
rect 11517 33915 11575 33921
rect 11517 33881 11529 33915
rect 11563 33912 11575 33915
rect 12894 33912 12900 33924
rect 11563 33884 12900 33912
rect 11563 33881 11575 33884
rect 11517 33875 11575 33881
rect 12894 33872 12900 33884
rect 12952 33872 12958 33924
rect 15580 33856 15608 33952
rect 15657 33949 15669 33983
rect 15703 33980 15715 33983
rect 16482 33980 16488 33992
rect 15703 33952 16488 33980
rect 15703 33949 15715 33952
rect 15657 33943 15715 33949
rect 16482 33940 16488 33952
rect 16540 33940 16546 33992
rect 17310 33980 17316 33992
rect 17271 33952 17316 33980
rect 17310 33940 17316 33952
rect 17368 33940 17374 33992
rect 18230 33980 18236 33992
rect 18191 33952 18236 33980
rect 18230 33940 18236 33952
rect 18288 33940 18294 33992
rect 20806 33940 20812 33992
rect 20864 33980 20870 33992
rect 20901 33983 20959 33989
rect 20901 33980 20913 33983
rect 20864 33952 20913 33980
rect 20864 33940 20870 33952
rect 20901 33949 20913 33952
rect 20947 33949 20959 33983
rect 21634 33980 21640 33992
rect 21595 33952 21640 33980
rect 20901 33943 20959 33949
rect 15930 33872 15936 33924
rect 15988 33912 15994 33924
rect 20916 33912 20944 33943
rect 21634 33940 21640 33952
rect 21692 33940 21698 33992
rect 22557 33983 22615 33989
rect 22557 33949 22569 33983
rect 22603 33949 22615 33983
rect 22557 33943 22615 33949
rect 22649 33983 22707 33989
rect 22649 33949 22661 33983
rect 22695 33980 22707 33983
rect 22830 33980 22836 33992
rect 22695 33952 22836 33980
rect 22695 33949 22707 33952
rect 22649 33943 22707 33949
rect 21913 33915 21971 33921
rect 21913 33912 21925 33915
rect 15988 33884 16436 33912
rect 20916 33884 21925 33912
rect 15988 33872 15994 33884
rect 7024 33816 7972 33844
rect 8202 33804 8208 33856
rect 8260 33844 8266 33856
rect 8389 33847 8447 33853
rect 8389 33844 8401 33847
rect 8260 33816 8401 33844
rect 8260 33804 8266 33816
rect 8389 33813 8401 33816
rect 8435 33813 8447 33847
rect 8389 33807 8447 33813
rect 8662 33804 8668 33856
rect 8720 33844 8726 33856
rect 9033 33847 9091 33853
rect 9033 33844 9045 33847
rect 8720 33816 9045 33844
rect 8720 33804 8726 33816
rect 9033 33813 9045 33816
rect 9079 33813 9091 33847
rect 13078 33844 13084 33856
rect 12991 33816 13084 33844
rect 9033 33807 9091 33813
rect 13078 33804 13084 33816
rect 13136 33844 13142 33856
rect 13998 33844 14004 33856
rect 13136 33816 14004 33844
rect 13136 33804 13142 33816
rect 13998 33804 14004 33816
rect 14056 33804 14062 33856
rect 15562 33844 15568 33856
rect 15523 33816 15568 33844
rect 15562 33804 15568 33816
rect 15620 33804 15626 33856
rect 15654 33804 15660 33856
rect 15712 33844 15718 33856
rect 16408 33853 16436 33884
rect 21913 33881 21925 33884
rect 21959 33881 21971 33915
rect 22572 33912 22600 33943
rect 22830 33940 22836 33952
rect 22888 33940 22894 33992
rect 23014 33940 23020 33992
rect 23072 33980 23078 33992
rect 24397 33983 24455 33989
rect 24397 33980 24409 33983
rect 23072 33952 24409 33980
rect 23072 33940 23078 33952
rect 24397 33949 24409 33952
rect 24443 33949 24455 33983
rect 24946 33980 24952 33992
rect 24907 33952 24952 33980
rect 24397 33943 24455 33949
rect 24946 33940 24952 33952
rect 25004 33940 25010 33992
rect 25038 33940 25044 33992
rect 25096 33980 25102 33992
rect 25409 33983 25467 33989
rect 25409 33980 25421 33983
rect 25096 33952 25421 33980
rect 25096 33940 25102 33952
rect 25409 33949 25421 33952
rect 25455 33949 25467 33983
rect 25409 33943 25467 33949
rect 23032 33912 23060 33940
rect 22572 33884 23060 33912
rect 21913 33875 21971 33881
rect 15749 33847 15807 33853
rect 15749 33844 15761 33847
rect 15712 33816 15761 33844
rect 15712 33804 15718 33816
rect 15749 33813 15761 33816
rect 15795 33813 15807 33847
rect 15749 33807 15807 33813
rect 16393 33847 16451 33853
rect 16393 33813 16405 33847
rect 16439 33844 16451 33847
rect 16482 33844 16488 33856
rect 16439 33816 16488 33844
rect 16439 33813 16451 33816
rect 16393 33807 16451 33813
rect 16482 33804 16488 33816
rect 16540 33804 16546 33856
rect 19797 33847 19855 33853
rect 19797 33813 19809 33847
rect 19843 33844 19855 33847
rect 20070 33844 20076 33856
rect 19843 33816 20076 33844
rect 19843 33813 19855 33816
rect 19797 33807 19855 33813
rect 20070 33804 20076 33816
rect 20128 33804 20134 33856
rect 20714 33844 20720 33856
rect 20675 33816 20720 33844
rect 20714 33804 20720 33816
rect 20772 33804 20778 33856
rect 23474 33804 23480 33856
rect 23532 33844 23538 33856
rect 23845 33847 23903 33853
rect 23845 33844 23857 33847
rect 23532 33816 23857 33844
rect 23532 33804 23538 33816
rect 23845 33813 23857 33816
rect 23891 33813 23903 33847
rect 24302 33844 24308 33856
rect 24263 33816 24308 33844
rect 23845 33807 23903 33813
rect 24302 33804 24308 33816
rect 24360 33804 24366 33856
rect 26237 33847 26295 33853
rect 26237 33813 26249 33847
rect 26283 33844 26295 33847
rect 26326 33844 26332 33856
rect 26283 33816 26332 33844
rect 26283 33813 26295 33816
rect 26237 33807 26295 33813
rect 26326 33804 26332 33816
rect 26384 33804 26390 33856
rect 1104 33754 28888 33776
rect 1104 33702 5982 33754
rect 6034 33702 6046 33754
rect 6098 33702 6110 33754
rect 6162 33702 6174 33754
rect 6226 33702 15982 33754
rect 16034 33702 16046 33754
rect 16098 33702 16110 33754
rect 16162 33702 16174 33754
rect 16226 33702 25982 33754
rect 26034 33702 26046 33754
rect 26098 33702 26110 33754
rect 26162 33702 26174 33754
rect 26226 33702 28888 33754
rect 1104 33680 28888 33702
rect 4522 33640 4528 33652
rect 4483 33612 4528 33640
rect 4522 33600 4528 33612
rect 4580 33600 4586 33652
rect 6273 33643 6331 33649
rect 5184 33612 6224 33640
rect 3513 33575 3571 33581
rect 3513 33541 3525 33575
rect 3559 33572 3571 33575
rect 5184 33572 5212 33612
rect 3559 33544 5212 33572
rect 3559 33541 3571 33544
rect 3513 33535 3571 33541
rect 5258 33532 5264 33584
rect 5316 33572 5322 33584
rect 5810 33572 5816 33584
rect 5316 33544 5816 33572
rect 5316 33532 5322 33544
rect 5810 33532 5816 33544
rect 5868 33532 5874 33584
rect 6196 33572 6224 33612
rect 6273 33609 6285 33643
rect 6319 33640 6331 33643
rect 6362 33640 6368 33652
rect 6319 33612 6368 33640
rect 6319 33609 6331 33612
rect 6273 33603 6331 33609
rect 6362 33600 6368 33612
rect 6420 33600 6426 33652
rect 6638 33640 6644 33652
rect 6599 33612 6644 33640
rect 6638 33600 6644 33612
rect 6696 33600 6702 33652
rect 7098 33640 7104 33652
rect 7059 33612 7104 33640
rect 7098 33600 7104 33612
rect 7156 33600 7162 33652
rect 8110 33600 8116 33652
rect 8168 33600 8174 33652
rect 8570 33600 8576 33652
rect 8628 33640 8634 33652
rect 9033 33643 9091 33649
rect 9033 33640 9045 33643
rect 8628 33612 9045 33640
rect 8628 33600 8634 33612
rect 9033 33609 9045 33612
rect 9079 33640 9091 33643
rect 9079 33612 10272 33640
rect 9079 33609 9091 33612
rect 9033 33603 9091 33609
rect 7742 33572 7748 33584
rect 6196 33544 7748 33572
rect 7742 33532 7748 33544
rect 7800 33532 7806 33584
rect 8128 33572 8156 33600
rect 10134 33572 10140 33584
rect 7944 33544 10140 33572
rect 2777 33507 2835 33513
rect 2777 33473 2789 33507
rect 2823 33504 2835 33507
rect 3145 33507 3203 33513
rect 3145 33504 3157 33507
rect 2823 33476 3157 33504
rect 2823 33473 2835 33476
rect 2777 33467 2835 33473
rect 3145 33473 3157 33476
rect 3191 33504 3203 33507
rect 4982 33504 4988 33516
rect 3191 33476 4988 33504
rect 3191 33473 3203 33476
rect 3145 33467 3203 33473
rect 4982 33464 4988 33476
rect 5040 33464 5046 33516
rect 5350 33504 5356 33516
rect 5311 33476 5356 33504
rect 5350 33464 5356 33476
rect 5408 33464 5414 33516
rect 7282 33504 7288 33516
rect 7243 33476 7288 33504
rect 7282 33464 7288 33476
rect 7340 33464 7346 33516
rect 7944 33513 7972 33544
rect 7929 33507 7987 33513
rect 7929 33473 7941 33507
rect 7975 33473 7987 33507
rect 8110 33504 8116 33516
rect 8071 33476 8116 33504
rect 7929 33467 7987 33473
rect 8110 33464 8116 33476
rect 8168 33464 8174 33516
rect 4249 33439 4307 33445
rect 4249 33405 4261 33439
rect 4295 33436 4307 33439
rect 4338 33436 4344 33448
rect 4295 33408 4344 33436
rect 4295 33405 4307 33408
rect 4249 33399 4307 33405
rect 4338 33396 4344 33408
rect 4396 33396 4402 33448
rect 5442 33436 5448 33448
rect 5403 33408 5448 33436
rect 5442 33396 5448 33408
rect 5500 33396 5506 33448
rect 6914 33396 6920 33448
rect 6972 33436 6978 33448
rect 7837 33439 7895 33445
rect 7837 33436 7849 33439
rect 6972 33408 7849 33436
rect 6972 33396 6978 33408
rect 7300 33380 7328 33408
rect 7837 33405 7849 33408
rect 7883 33405 7895 33439
rect 8202 33436 8208 33448
rect 8163 33408 8208 33436
rect 7837 33399 7895 33405
rect 8202 33396 8208 33408
rect 8260 33396 8266 33448
rect 9692 33445 9720 33544
rect 10134 33532 10140 33544
rect 10192 33532 10198 33584
rect 10244 33504 10272 33612
rect 10870 33600 10876 33652
rect 10928 33640 10934 33652
rect 11701 33643 11759 33649
rect 11701 33640 11713 33643
rect 10928 33612 11713 33640
rect 10928 33600 10934 33612
rect 11701 33609 11713 33612
rect 11747 33640 11759 33643
rect 12158 33640 12164 33652
rect 11747 33612 12164 33640
rect 11747 33609 11759 33612
rect 11701 33603 11759 33609
rect 12158 33600 12164 33612
rect 12216 33600 12222 33652
rect 13538 33600 13544 33652
rect 13596 33640 13602 33652
rect 13633 33643 13691 33649
rect 13633 33640 13645 33643
rect 13596 33612 13645 33640
rect 13596 33600 13602 33612
rect 13633 33609 13645 33612
rect 13679 33609 13691 33643
rect 13633 33603 13691 33609
rect 15562 33600 15568 33652
rect 15620 33640 15626 33652
rect 17589 33643 17647 33649
rect 17589 33640 17601 33643
rect 15620 33612 17601 33640
rect 15620 33600 15626 33612
rect 17589 33609 17601 33612
rect 17635 33609 17647 33643
rect 17589 33603 17647 33609
rect 19153 33643 19211 33649
rect 19153 33609 19165 33643
rect 19199 33640 19211 33643
rect 19242 33640 19248 33652
rect 19199 33612 19248 33640
rect 19199 33609 19211 33612
rect 19153 33603 19211 33609
rect 19242 33600 19248 33612
rect 19300 33600 19306 33652
rect 20622 33600 20628 33652
rect 20680 33640 20686 33652
rect 22649 33643 22707 33649
rect 22649 33640 22661 33643
rect 20680 33612 22661 33640
rect 20680 33600 20686 33612
rect 22649 33609 22661 33612
rect 22695 33609 22707 33643
rect 22649 33603 22707 33609
rect 22925 33643 22983 33649
rect 22925 33609 22937 33643
rect 22971 33640 22983 33643
rect 23014 33640 23020 33652
rect 22971 33612 23020 33640
rect 22971 33609 22983 33612
rect 22925 33603 22983 33609
rect 23014 33600 23020 33612
rect 23072 33600 23078 33652
rect 23198 33640 23204 33652
rect 23159 33612 23204 33640
rect 23198 33600 23204 33612
rect 23256 33600 23262 33652
rect 23566 33600 23572 33652
rect 23624 33640 23630 33652
rect 23845 33643 23903 33649
rect 23845 33640 23857 33643
rect 23624 33612 23857 33640
rect 23624 33600 23630 33612
rect 23845 33609 23857 33612
rect 23891 33609 23903 33643
rect 23845 33603 23903 33609
rect 24489 33643 24547 33649
rect 24489 33609 24501 33643
rect 24535 33640 24547 33643
rect 25038 33640 25044 33652
rect 24535 33612 25044 33640
rect 24535 33609 24547 33612
rect 24489 33603 24547 33609
rect 10962 33572 10968 33584
rect 10923 33544 10968 33572
rect 10962 33532 10968 33544
rect 11020 33532 11026 33584
rect 12066 33532 12072 33584
rect 12124 33572 12130 33584
rect 12526 33572 12532 33584
rect 12124 33544 12532 33572
rect 12124 33532 12130 33544
rect 12526 33532 12532 33544
rect 12584 33532 12590 33584
rect 13078 33572 13084 33584
rect 12728 33544 13084 33572
rect 10980 33504 11008 33532
rect 12728 33504 12756 33544
rect 13078 33532 13084 33544
rect 13136 33532 13142 33584
rect 15010 33532 15016 33584
rect 15068 33572 15074 33584
rect 15378 33572 15384 33584
rect 15068 33544 15384 33572
rect 15068 33532 15074 33544
rect 15378 33532 15384 33544
rect 15436 33572 15442 33584
rect 15436 33544 16344 33572
rect 15436 33532 15442 33544
rect 10152 33476 11008 33504
rect 12636 33476 12756 33504
rect 9677 33439 9735 33445
rect 9677 33405 9689 33439
rect 9723 33405 9735 33439
rect 9950 33436 9956 33448
rect 9911 33408 9956 33436
rect 9677 33399 9735 33405
rect 9950 33396 9956 33408
rect 10008 33396 10014 33448
rect 10152 33445 10180 33476
rect 10137 33439 10195 33445
rect 10137 33405 10149 33439
rect 10183 33405 10195 33439
rect 10137 33399 10195 33405
rect 10226 33396 10232 33448
rect 10284 33436 10290 33448
rect 10321 33439 10379 33445
rect 10321 33436 10333 33439
rect 10284 33408 10333 33436
rect 10284 33396 10290 33408
rect 10321 33405 10333 33408
rect 10367 33436 10379 33439
rect 10502 33436 10508 33448
rect 10367 33408 10508 33436
rect 10367 33405 10379 33408
rect 10321 33399 10379 33405
rect 10502 33396 10508 33408
rect 10560 33396 10566 33448
rect 10689 33439 10747 33445
rect 10689 33405 10701 33439
rect 10735 33436 10747 33439
rect 10778 33436 10784 33448
rect 10735 33408 10784 33436
rect 10735 33405 10747 33408
rect 10689 33399 10747 33405
rect 10778 33396 10784 33408
rect 10836 33396 10842 33448
rect 12636 33445 12664 33476
rect 12802 33464 12808 33516
rect 12860 33504 12866 33516
rect 13538 33504 13544 33516
rect 12860 33476 13544 33504
rect 12860 33464 12866 33476
rect 13538 33464 13544 33476
rect 13596 33464 13602 33516
rect 14918 33464 14924 33516
rect 14976 33504 14982 33516
rect 16206 33504 16212 33516
rect 14976 33476 15424 33504
rect 14976 33464 14982 33476
rect 15396 33448 15424 33476
rect 15580 33476 16212 33504
rect 12437 33439 12495 33445
rect 12437 33436 12449 33439
rect 12268 33408 12449 33436
rect 3878 33368 3884 33380
rect 3839 33340 3884 33368
rect 3878 33328 3884 33340
rect 3936 33328 3942 33380
rect 4430 33328 4436 33380
rect 4488 33368 4494 33380
rect 4893 33371 4951 33377
rect 4893 33368 4905 33371
rect 4488 33340 4905 33368
rect 4488 33328 4494 33340
rect 4893 33337 4905 33340
rect 4939 33368 4951 33371
rect 4982 33368 4988 33380
rect 4939 33340 4988 33368
rect 4939 33337 4951 33340
rect 4893 33331 4951 33337
rect 4982 33328 4988 33340
rect 5040 33368 5046 33380
rect 5902 33368 5908 33380
rect 5040 33340 5672 33368
rect 5863 33340 5908 33368
rect 5040 33328 5046 33340
rect 5261 33303 5319 33309
rect 5261 33269 5273 33303
rect 5307 33300 5319 33303
rect 5534 33300 5540 33312
rect 5307 33272 5540 33300
rect 5307 33269 5319 33272
rect 5261 33263 5319 33269
rect 5534 33260 5540 33272
rect 5592 33260 5598 33312
rect 5644 33300 5672 33340
rect 5902 33328 5908 33340
rect 5960 33328 5966 33380
rect 7282 33328 7288 33380
rect 7340 33328 7346 33380
rect 8754 33368 8760 33380
rect 8036 33340 8760 33368
rect 8036 33300 8064 33340
rect 8754 33328 8760 33340
rect 8812 33328 8818 33380
rect 9214 33368 9220 33380
rect 9175 33340 9220 33368
rect 9214 33328 9220 33340
rect 9272 33328 9278 33380
rect 12158 33368 12164 33380
rect 10336 33340 12164 33368
rect 10336 33312 10364 33340
rect 12158 33328 12164 33340
rect 12216 33368 12222 33380
rect 12268 33368 12296 33408
rect 12437 33405 12449 33408
rect 12483 33405 12495 33439
rect 12437 33399 12495 33405
rect 12621 33439 12679 33445
rect 12621 33405 12633 33439
rect 12667 33405 12679 33439
rect 12621 33399 12679 33405
rect 13078 33396 13084 33448
rect 13136 33436 13142 33448
rect 13173 33439 13231 33445
rect 13173 33436 13185 33439
rect 13136 33408 13185 33436
rect 13136 33396 13142 33408
rect 13173 33405 13185 33408
rect 13219 33405 13231 33439
rect 15102 33436 15108 33448
rect 15063 33408 15108 33436
rect 13173 33399 13231 33405
rect 15102 33396 15108 33408
rect 15160 33396 15166 33448
rect 15378 33396 15384 33448
rect 15436 33396 15442 33448
rect 15580 33445 15608 33476
rect 16206 33464 16212 33476
rect 16264 33464 16270 33516
rect 15565 33439 15623 33445
rect 15565 33405 15577 33439
rect 15611 33405 15623 33439
rect 15565 33399 15623 33405
rect 15841 33439 15899 33445
rect 15841 33405 15853 33439
rect 15887 33436 15899 33439
rect 15930 33436 15936 33448
rect 15887 33408 15936 33436
rect 15887 33405 15899 33408
rect 15841 33399 15899 33405
rect 15930 33396 15936 33408
rect 15988 33396 15994 33448
rect 16117 33439 16175 33445
rect 16117 33405 16129 33439
rect 16163 33436 16175 33439
rect 16316 33436 16344 33544
rect 23106 33532 23112 33584
rect 23164 33572 23170 33584
rect 24504 33572 24532 33603
rect 25038 33600 25044 33612
rect 25096 33600 25102 33652
rect 25498 33600 25504 33652
rect 25556 33640 25562 33652
rect 25961 33643 26019 33649
rect 25961 33640 25973 33643
rect 25556 33612 25973 33640
rect 25556 33600 25562 33612
rect 25961 33609 25973 33612
rect 26007 33609 26019 33643
rect 25961 33603 26019 33609
rect 23164 33544 24532 33572
rect 23164 33532 23170 33544
rect 24946 33532 24952 33584
rect 25004 33572 25010 33584
rect 25133 33575 25191 33581
rect 25133 33572 25145 33575
rect 25004 33544 25145 33572
rect 25004 33532 25010 33544
rect 25133 33541 25145 33544
rect 25179 33541 25191 33575
rect 25133 33535 25191 33541
rect 20346 33464 20352 33516
rect 20404 33504 20410 33516
rect 20622 33504 20628 33516
rect 20404 33476 20628 33504
rect 20404 33464 20410 33476
rect 20622 33464 20628 33476
rect 20680 33464 20686 33516
rect 20898 33504 20904 33516
rect 20859 33476 20904 33504
rect 20898 33464 20904 33476
rect 20956 33464 20962 33516
rect 22554 33504 22560 33516
rect 22515 33476 22560 33504
rect 22554 33464 22560 33476
rect 22612 33464 22618 33516
rect 24857 33507 24915 33513
rect 24857 33473 24869 33507
rect 24903 33504 24915 33507
rect 25314 33504 25320 33516
rect 24903 33476 25320 33504
rect 24903 33473 24915 33476
rect 24857 33467 24915 33473
rect 25314 33464 25320 33476
rect 25372 33464 25378 33516
rect 16163 33408 16344 33436
rect 18693 33439 18751 33445
rect 16163 33405 16175 33408
rect 16117 33399 16175 33405
rect 18693 33405 18705 33439
rect 18739 33436 18751 33439
rect 18874 33436 18880 33448
rect 18739 33408 18880 33436
rect 18739 33405 18751 33408
rect 18693 33399 18751 33405
rect 18874 33396 18880 33408
rect 18932 33396 18938 33448
rect 19610 33396 19616 33448
rect 19668 33436 19674 33448
rect 19981 33439 20039 33445
rect 19981 33436 19993 33439
rect 19668 33408 19993 33436
rect 19668 33396 19674 33408
rect 19981 33405 19993 33408
rect 20027 33405 20039 33439
rect 19981 33399 20039 33405
rect 20438 33396 20444 33448
rect 20496 33436 20502 33448
rect 20809 33439 20867 33445
rect 20809 33436 20821 33439
rect 20496 33408 20821 33436
rect 20496 33396 20502 33408
rect 20809 33405 20821 33408
rect 20855 33405 20867 33439
rect 20809 33399 20867 33405
rect 22097 33439 22155 33445
rect 22097 33405 22109 33439
rect 22143 33436 22155 33439
rect 22278 33436 22284 33448
rect 22143 33408 22284 33436
rect 22143 33405 22155 33408
rect 22097 33399 22155 33405
rect 22278 33396 22284 33408
rect 22336 33396 22342 33448
rect 25976 33436 26004 33603
rect 26145 33507 26203 33513
rect 26145 33473 26157 33507
rect 26191 33504 26203 33507
rect 26326 33504 26332 33516
rect 26191 33476 26332 33504
rect 26191 33473 26203 33476
rect 26145 33467 26203 33473
rect 26326 33464 26332 33476
rect 26384 33464 26390 33516
rect 26421 33439 26479 33445
rect 26421 33436 26433 33439
rect 25976 33408 26433 33436
rect 26421 33405 26433 33408
rect 26467 33405 26479 33439
rect 26421 33399 26479 33405
rect 12216 33340 12296 33368
rect 12216 33328 12222 33340
rect 12342 33328 12348 33380
rect 12400 33368 12406 33380
rect 12805 33371 12863 33377
rect 12805 33368 12817 33371
rect 12400 33340 12817 33368
rect 12400 33328 12406 33340
rect 12805 33337 12817 33340
rect 12851 33337 12863 33371
rect 14001 33371 14059 33377
rect 14001 33368 14013 33371
rect 12805 33331 12863 33337
rect 12912 33340 14013 33368
rect 12912 33312 12940 33340
rect 14001 33337 14013 33340
rect 14047 33337 14059 33371
rect 16942 33368 16948 33380
rect 16855 33340 16948 33368
rect 14001 33331 14059 33337
rect 16942 33328 16948 33340
rect 17000 33368 17006 33380
rect 18782 33368 18788 33380
rect 17000 33340 18788 33368
rect 17000 33328 17006 33340
rect 18782 33328 18788 33340
rect 18840 33328 18846 33380
rect 20073 33371 20131 33377
rect 20073 33337 20085 33371
rect 20119 33368 20131 33371
rect 20346 33368 20352 33380
rect 20119 33340 20352 33368
rect 20119 33337 20131 33340
rect 20073 33331 20131 33337
rect 20346 33328 20352 33340
rect 20404 33328 20410 33380
rect 20898 33328 20904 33380
rect 20956 33368 20962 33380
rect 21821 33371 21879 33377
rect 21821 33368 21833 33371
rect 20956 33340 21833 33368
rect 20956 33328 20962 33340
rect 21821 33337 21833 33340
rect 21867 33337 21879 33371
rect 21821 33331 21879 33337
rect 22189 33371 22247 33377
rect 22189 33337 22201 33371
rect 22235 33368 22247 33371
rect 22370 33368 22376 33380
rect 22235 33340 22376 33368
rect 22235 33337 22247 33340
rect 22189 33331 22247 33337
rect 22370 33328 22376 33340
rect 22428 33368 22434 33380
rect 23290 33368 23296 33380
rect 22428 33340 23296 33368
rect 22428 33328 22434 33340
rect 23290 33328 23296 33340
rect 23348 33328 23354 33380
rect 8662 33300 8668 33312
rect 5644 33272 8064 33300
rect 8623 33272 8668 33300
rect 8662 33260 8668 33272
rect 8720 33260 8726 33312
rect 10318 33260 10324 33312
rect 10376 33260 10382 33312
rect 11974 33300 11980 33312
rect 11935 33272 11980 33300
rect 11974 33260 11980 33272
rect 12032 33260 12038 33312
rect 12713 33303 12771 33309
rect 12713 33269 12725 33303
rect 12759 33300 12771 33303
rect 12894 33300 12900 33312
rect 12759 33272 12900 33300
rect 12759 33269 12771 33272
rect 12713 33263 12771 33269
rect 12894 33260 12900 33272
rect 12952 33260 12958 33312
rect 14366 33300 14372 33312
rect 14327 33272 14372 33300
rect 14366 33260 14372 33272
rect 14424 33260 14430 33312
rect 14826 33260 14832 33312
rect 14884 33300 14890 33312
rect 14921 33303 14979 33309
rect 14921 33300 14933 33303
rect 14884 33272 14933 33300
rect 14884 33260 14890 33272
rect 14921 33269 14933 33272
rect 14967 33269 14979 33303
rect 14921 33263 14979 33269
rect 15930 33260 15936 33312
rect 15988 33300 15994 33312
rect 17313 33303 17371 33309
rect 17313 33300 17325 33303
rect 15988 33272 17325 33300
rect 15988 33260 15994 33272
rect 17313 33269 17325 33272
rect 17359 33300 17371 33303
rect 18046 33300 18052 33312
rect 17359 33272 18052 33300
rect 17359 33269 17371 33272
rect 17313 33263 17371 33269
rect 18046 33260 18052 33272
rect 18104 33260 18110 33312
rect 19426 33300 19432 33312
rect 19387 33272 19432 33300
rect 19426 33260 19432 33272
rect 19484 33260 19490 33312
rect 21358 33300 21364 33312
rect 21271 33272 21364 33300
rect 21358 33260 21364 33272
rect 21416 33300 21422 33312
rect 21637 33303 21695 33309
rect 21637 33300 21649 33303
rect 21416 33272 21649 33300
rect 21416 33260 21422 33272
rect 21637 33269 21649 33272
rect 21683 33300 21695 33303
rect 21910 33300 21916 33312
rect 21683 33272 21916 33300
rect 21683 33269 21695 33272
rect 21637 33263 21695 33269
rect 21910 33260 21916 33272
rect 21968 33300 21974 33312
rect 22005 33303 22063 33309
rect 22005 33300 22017 33303
rect 21968 33272 22017 33300
rect 21968 33260 21974 33272
rect 22005 33269 22017 33272
rect 22051 33269 22063 33303
rect 22005 33263 22063 33269
rect 22649 33303 22707 33309
rect 22649 33269 22661 33303
rect 22695 33300 22707 33303
rect 27525 33303 27583 33309
rect 27525 33300 27537 33303
rect 22695 33272 27537 33300
rect 22695 33269 22707 33272
rect 22649 33263 22707 33269
rect 27525 33269 27537 33272
rect 27571 33269 27583 33303
rect 27525 33263 27583 33269
rect 1104 33210 28888 33232
rect 1104 33158 10982 33210
rect 11034 33158 11046 33210
rect 11098 33158 11110 33210
rect 11162 33158 11174 33210
rect 11226 33158 20982 33210
rect 21034 33158 21046 33210
rect 21098 33158 21110 33210
rect 21162 33158 21174 33210
rect 21226 33158 28888 33210
rect 1104 33136 28888 33158
rect 4614 33096 4620 33108
rect 4575 33068 4620 33096
rect 4614 33056 4620 33068
rect 4672 33056 4678 33108
rect 4893 33099 4951 33105
rect 4893 33065 4905 33099
rect 4939 33096 4951 33099
rect 7745 33099 7803 33105
rect 4939 33068 7696 33096
rect 4939 33065 4951 33068
rect 4893 33059 4951 33065
rect 7006 33028 7012 33040
rect 6840 33000 7012 33028
rect 4709 32963 4767 32969
rect 4709 32929 4721 32963
rect 4755 32960 4767 32963
rect 5166 32960 5172 32972
rect 4755 32932 5172 32960
rect 4755 32929 4767 32932
rect 4709 32923 4767 32929
rect 5166 32920 5172 32932
rect 5224 32920 5230 32972
rect 6840 32960 6868 33000
rect 7006 32988 7012 33000
rect 7064 32988 7070 33040
rect 7668 33028 7696 33068
rect 7745 33065 7757 33099
rect 7791 33096 7803 33099
rect 7834 33096 7840 33108
rect 7791 33068 7840 33096
rect 7791 33065 7803 33068
rect 7745 33059 7803 33065
rect 7834 33056 7840 33068
rect 7892 33096 7898 33108
rect 8110 33096 8116 33108
rect 7892 33068 8116 33096
rect 7892 33056 7898 33068
rect 8110 33056 8116 33068
rect 8168 33056 8174 33108
rect 8386 33056 8392 33108
rect 8444 33096 8450 33108
rect 9217 33099 9275 33105
rect 9217 33096 9229 33099
rect 8444 33068 9229 33096
rect 8444 33056 8450 33068
rect 9217 33065 9229 33068
rect 9263 33096 9275 33099
rect 9490 33096 9496 33108
rect 9263 33068 9496 33096
rect 9263 33065 9275 33068
rect 9217 33059 9275 33065
rect 9490 33056 9496 33068
rect 9548 33056 9554 33108
rect 11609 33099 11667 33105
rect 11609 33065 11621 33099
rect 11655 33096 11667 33099
rect 11655 33068 14228 33096
rect 11655 33065 11667 33068
rect 11609 33059 11667 33065
rect 8021 33031 8079 33037
rect 8021 33028 8033 33031
rect 7668 33000 8033 33028
rect 8021 32997 8033 33000
rect 8067 33028 8079 33031
rect 8754 33028 8760 33040
rect 8067 33000 8760 33028
rect 8067 32997 8079 33000
rect 8021 32991 8079 32997
rect 8754 32988 8760 33000
rect 8812 32988 8818 33040
rect 9122 32988 9128 33040
rect 9180 33028 9186 33040
rect 9677 33031 9735 33037
rect 9180 33000 9628 33028
rect 9180 32988 9186 33000
rect 9600 32972 9628 33000
rect 9677 32997 9689 33031
rect 9723 33028 9735 33031
rect 10410 33028 10416 33040
rect 9723 33000 10416 33028
rect 9723 32997 9735 33000
rect 9677 32991 9735 32997
rect 10410 32988 10416 33000
rect 10468 32988 10474 33040
rect 10502 32988 10508 33040
rect 10560 32988 10566 33040
rect 8294 32960 8300 32972
rect 5736 32932 6868 32960
rect 8255 32932 8300 32960
rect 5736 32904 5764 32932
rect 8294 32920 8300 32932
rect 8352 32920 8358 32972
rect 9306 32920 9312 32972
rect 9364 32960 9370 32972
rect 9401 32963 9459 32969
rect 9401 32960 9413 32963
rect 9364 32932 9413 32960
rect 9364 32920 9370 32932
rect 9401 32929 9413 32932
rect 9447 32929 9459 32963
rect 9401 32923 9459 32929
rect 9582 32920 9588 32972
rect 9640 32920 9646 32972
rect 10318 32960 10324 32972
rect 10279 32932 10324 32960
rect 10318 32920 10324 32932
rect 10376 32920 10382 32972
rect 10520 32960 10548 32988
rect 11716 32969 11744 33068
rect 12158 32988 12164 33040
rect 12216 33028 12222 33040
rect 12437 33031 12495 33037
rect 12437 33028 12449 33031
rect 12216 33000 12449 33028
rect 12216 32988 12222 33000
rect 12437 32997 12449 33000
rect 12483 32997 12495 33031
rect 12710 33028 12716 33040
rect 12671 33000 12716 33028
rect 12437 32991 12495 32997
rect 10689 32963 10747 32969
rect 10689 32960 10701 32963
rect 10520 32932 10701 32960
rect 10689 32929 10701 32932
rect 10735 32929 10747 32963
rect 10689 32923 10747 32929
rect 11701 32963 11759 32969
rect 11701 32929 11713 32963
rect 11747 32929 11759 32963
rect 12452 32960 12480 32991
rect 12710 32988 12716 33000
rect 12768 32988 12774 33040
rect 12894 32988 12900 33040
rect 12952 33028 12958 33040
rect 14090 33028 14096 33040
rect 12952 33000 13584 33028
rect 12952 32988 12958 33000
rect 13078 32960 13084 32972
rect 12452 32932 13084 32960
rect 11701 32923 11759 32929
rect 13078 32920 13084 32932
rect 13136 32920 13142 32972
rect 13556 32969 13584 33000
rect 14016 33000 14096 33028
rect 13173 32963 13231 32969
rect 13173 32929 13185 32963
rect 13219 32929 13231 32963
rect 13173 32923 13231 32929
rect 13449 32963 13507 32969
rect 13449 32929 13461 32963
rect 13495 32929 13507 32963
rect 13449 32923 13507 32929
rect 13541 32963 13599 32969
rect 13541 32929 13553 32963
rect 13587 32929 13599 32963
rect 13541 32923 13599 32929
rect 3418 32852 3424 32904
rect 3476 32892 3482 32904
rect 3513 32895 3571 32901
rect 3513 32892 3525 32895
rect 3476 32864 3525 32892
rect 3476 32852 3482 32864
rect 3513 32861 3525 32864
rect 3559 32892 3571 32895
rect 5718 32892 5724 32904
rect 3559 32864 5724 32892
rect 3559 32861 3571 32864
rect 3513 32855 3571 32861
rect 5718 32852 5724 32864
rect 5776 32852 5782 32904
rect 5902 32852 5908 32904
rect 5960 32892 5966 32904
rect 5997 32895 6055 32901
rect 5997 32892 6009 32895
rect 5960 32864 6009 32892
rect 5960 32852 5966 32864
rect 5997 32861 6009 32864
rect 6043 32861 6055 32895
rect 5997 32855 6055 32861
rect 7377 32895 7435 32901
rect 7377 32861 7389 32895
rect 7423 32892 7435 32895
rect 7742 32892 7748 32904
rect 7423 32864 7748 32892
rect 7423 32861 7435 32864
rect 7377 32855 7435 32861
rect 7742 32852 7748 32864
rect 7800 32852 7806 32904
rect 8205 32895 8263 32901
rect 8205 32892 8217 32895
rect 8036 32864 8217 32892
rect 7006 32784 7012 32836
rect 7064 32824 7070 32836
rect 7650 32824 7656 32836
rect 7064 32796 7656 32824
rect 7064 32784 7070 32796
rect 7650 32784 7656 32796
rect 7708 32784 7714 32836
rect 3878 32756 3884 32768
rect 3839 32728 3884 32756
rect 3878 32716 3884 32728
rect 3936 32716 3942 32768
rect 5442 32756 5448 32768
rect 5403 32728 5448 32756
rect 5442 32716 5448 32728
rect 5500 32716 5506 32768
rect 6914 32716 6920 32768
rect 6972 32756 6978 32768
rect 8036 32756 8064 32864
rect 8205 32861 8217 32864
rect 8251 32861 8263 32895
rect 8205 32855 8263 32861
rect 8757 32895 8815 32901
rect 8757 32861 8769 32895
rect 8803 32892 8815 32895
rect 9122 32892 9128 32904
rect 8803 32864 9128 32892
rect 8803 32861 8815 32864
rect 8757 32855 8815 32861
rect 9122 32852 9128 32864
rect 9180 32892 9186 32904
rect 10229 32895 10287 32901
rect 10229 32892 10241 32895
rect 9180 32864 10241 32892
rect 9180 32852 9186 32864
rect 10229 32861 10241 32864
rect 10275 32861 10287 32895
rect 10778 32892 10784 32904
rect 10739 32864 10784 32892
rect 10229 32855 10287 32861
rect 10778 32852 10784 32864
rect 10836 32852 10842 32904
rect 12250 32852 12256 32904
rect 12308 32892 12314 32904
rect 12434 32892 12440 32904
rect 12308 32864 12440 32892
rect 12308 32852 12314 32864
rect 12434 32852 12440 32864
rect 12492 32852 12498 32904
rect 12986 32852 12992 32904
rect 13044 32892 13050 32904
rect 13188 32892 13216 32923
rect 13044 32864 13216 32892
rect 13464 32892 13492 32923
rect 13814 32892 13820 32904
rect 13464 32864 13584 32892
rect 13775 32864 13820 32892
rect 13044 32852 13050 32864
rect 8110 32784 8116 32836
rect 8168 32824 8174 32836
rect 9401 32827 9459 32833
rect 9401 32824 9413 32827
rect 8168 32796 9413 32824
rect 8168 32784 8174 32796
rect 9401 32793 9413 32796
rect 9447 32824 9459 32827
rect 13004 32824 13032 32852
rect 9447 32796 13032 32824
rect 13556 32824 13584 32864
rect 13814 32852 13820 32864
rect 13872 32852 13878 32904
rect 14016 32892 14044 33000
rect 14090 32988 14096 33000
rect 14148 32988 14154 33040
rect 14200 33028 14228 33068
rect 14274 33056 14280 33108
rect 14332 33096 14338 33108
rect 14550 33096 14556 33108
rect 14332 33068 14556 33096
rect 14332 33056 14338 33068
rect 14550 33056 14556 33068
rect 14608 33056 14614 33108
rect 14645 33099 14703 33105
rect 14645 33065 14657 33099
rect 14691 33096 14703 33099
rect 14826 33096 14832 33108
rect 14691 33068 14832 33096
rect 14691 33065 14703 33068
rect 14645 33059 14703 33065
rect 14826 33056 14832 33068
rect 14884 33056 14890 33108
rect 14921 33099 14979 33105
rect 14921 33065 14933 33099
rect 14967 33096 14979 33099
rect 15102 33096 15108 33108
rect 14967 33068 15108 33096
rect 14967 33065 14979 33068
rect 14921 33059 14979 33065
rect 15102 33056 15108 33068
rect 15160 33056 15166 33108
rect 15470 33096 15476 33108
rect 15212 33068 15476 33096
rect 14734 33028 14740 33040
rect 14200 33000 14740 33028
rect 14734 32988 14740 33000
rect 14792 33028 14798 33040
rect 15212 33028 15240 33068
rect 15470 33056 15476 33068
rect 15528 33056 15534 33108
rect 16206 33056 16212 33108
rect 16264 33096 16270 33108
rect 16301 33099 16359 33105
rect 16301 33096 16313 33099
rect 16264 33068 16313 33096
rect 16264 33056 16270 33068
rect 16301 33065 16313 33068
rect 16347 33065 16359 33099
rect 16301 33059 16359 33065
rect 16574 33056 16580 33108
rect 16632 33096 16638 33108
rect 17037 33099 17095 33105
rect 17037 33096 17049 33099
rect 16632 33068 17049 33096
rect 16632 33056 16638 33068
rect 17037 33065 17049 33068
rect 17083 33065 17095 33099
rect 17494 33096 17500 33108
rect 17037 33059 17095 33065
rect 17328 33068 17500 33096
rect 14792 33000 15240 33028
rect 14792 32988 14798 33000
rect 15378 32988 15384 33040
rect 15436 33028 15442 33040
rect 15657 33031 15715 33037
rect 15657 33028 15669 33031
rect 15436 33000 15669 33028
rect 15436 32988 15442 33000
rect 15657 32997 15669 33000
rect 15703 32997 15715 33031
rect 16022 33028 16028 33040
rect 15983 33000 16028 33028
rect 15657 32991 15715 32997
rect 14182 32960 14188 32972
rect 14095 32932 14188 32960
rect 14182 32920 14188 32932
rect 14240 32960 14246 32972
rect 14645 32963 14703 32969
rect 14645 32960 14657 32963
rect 14240 32932 14657 32960
rect 14240 32920 14246 32932
rect 14645 32929 14657 32932
rect 14691 32929 14703 32963
rect 15562 32960 15568 32972
rect 15523 32932 15568 32960
rect 14645 32923 14703 32929
rect 15562 32920 15568 32932
rect 15620 32920 15626 32972
rect 15672 32960 15700 32991
rect 16022 32988 16028 33000
rect 16080 32988 16086 33040
rect 17328 33028 17356 33068
rect 17494 33056 17500 33068
rect 17552 33056 17558 33108
rect 18598 33096 18604 33108
rect 18559 33068 18604 33096
rect 18598 33056 18604 33068
rect 18656 33056 18662 33108
rect 19610 33096 19616 33108
rect 19571 33068 19616 33096
rect 19610 33056 19616 33068
rect 19668 33056 19674 33108
rect 20717 33099 20775 33105
rect 20717 33065 20729 33099
rect 20763 33096 20775 33099
rect 20806 33096 20812 33108
rect 20763 33068 20812 33096
rect 20763 33065 20775 33068
rect 20717 33059 20775 33065
rect 20806 33056 20812 33068
rect 20864 33056 20870 33108
rect 22925 33099 22983 33105
rect 22925 33065 22937 33099
rect 22971 33096 22983 33099
rect 23382 33096 23388 33108
rect 22971 33068 23388 33096
rect 22971 33065 22983 33068
rect 22925 33059 22983 33065
rect 23382 33056 23388 33068
rect 23440 33056 23446 33108
rect 23661 33099 23719 33105
rect 23661 33065 23673 33099
rect 23707 33096 23719 33099
rect 23750 33096 23756 33108
rect 23707 33068 23756 33096
rect 23707 33065 23719 33068
rect 23661 33059 23719 33065
rect 23750 33056 23756 33068
rect 23808 33056 23814 33108
rect 25130 33096 25136 33108
rect 25091 33068 25136 33096
rect 25130 33056 25136 33068
rect 25188 33056 25194 33108
rect 23290 33028 23296 33040
rect 16316 33000 17356 33028
rect 23251 33000 23296 33028
rect 15930 32960 15936 32972
rect 15672 32932 15936 32960
rect 15930 32920 15936 32932
rect 15988 32920 15994 32972
rect 14366 32892 14372 32904
rect 14016 32864 14372 32892
rect 14366 32852 14372 32864
rect 14424 32852 14430 32904
rect 14550 32852 14556 32904
rect 14608 32892 14614 32904
rect 14826 32892 14832 32904
rect 14608 32864 14832 32892
rect 14608 32852 14614 32864
rect 14826 32852 14832 32864
rect 14884 32852 14890 32904
rect 14918 32852 14924 32904
rect 14976 32892 14982 32904
rect 15289 32895 15347 32901
rect 15289 32892 15301 32895
rect 14976 32864 15301 32892
rect 14976 32852 14982 32864
rect 15289 32861 15301 32864
rect 15335 32861 15347 32895
rect 15289 32855 15347 32861
rect 16316 32836 16344 33000
rect 23290 32988 23296 33000
rect 23348 32988 23354 33040
rect 17221 32963 17279 32969
rect 17221 32929 17233 32963
rect 17267 32960 17279 32963
rect 18230 32960 18236 32972
rect 17267 32932 18236 32960
rect 17267 32929 17279 32932
rect 17221 32923 17279 32929
rect 18230 32920 18236 32932
rect 18288 32960 18294 32972
rect 19150 32960 19156 32972
rect 18288 32932 19156 32960
rect 18288 32920 18294 32932
rect 19150 32920 19156 32932
rect 19208 32920 19214 32972
rect 19705 32963 19763 32969
rect 19705 32929 19717 32963
rect 19751 32960 19763 32963
rect 20901 32963 20959 32969
rect 19751 32932 20300 32960
rect 19751 32929 19763 32932
rect 19705 32923 19763 32929
rect 16482 32852 16488 32904
rect 16540 32892 16546 32904
rect 16850 32892 16856 32904
rect 16540 32864 16856 32892
rect 16540 32852 16546 32864
rect 16850 32852 16856 32864
rect 16908 32852 16914 32904
rect 17494 32892 17500 32904
rect 17455 32864 17500 32892
rect 17494 32852 17500 32864
rect 17552 32852 17558 32904
rect 14090 32824 14096 32836
rect 13556 32796 14096 32824
rect 9447 32793 9459 32796
rect 9401 32787 9459 32793
rect 6972 32728 8064 32756
rect 6972 32716 6978 32728
rect 10134 32716 10140 32768
rect 10192 32756 10198 32768
rect 11149 32759 11207 32765
rect 11149 32756 11161 32759
rect 10192 32728 11161 32756
rect 10192 32716 10198 32728
rect 11149 32725 11161 32728
rect 11195 32725 11207 32759
rect 11149 32719 11207 32725
rect 11422 32716 11428 32768
rect 11480 32756 11486 32768
rect 11885 32759 11943 32765
rect 11885 32756 11897 32759
rect 11480 32728 11897 32756
rect 11480 32716 11486 32728
rect 11885 32725 11897 32728
rect 11931 32725 11943 32759
rect 11885 32719 11943 32725
rect 12158 32716 12164 32768
rect 12216 32756 12222 32768
rect 13556 32756 13584 32796
rect 14090 32784 14096 32796
rect 14148 32784 14154 32836
rect 16298 32784 16304 32836
rect 16356 32784 16362 32836
rect 12216 32728 13584 32756
rect 12216 32716 12222 32728
rect 16574 32716 16580 32768
rect 16632 32756 16638 32768
rect 16669 32759 16727 32765
rect 16669 32756 16681 32759
rect 16632 32728 16681 32756
rect 16632 32716 16638 32728
rect 16669 32725 16681 32728
rect 16715 32725 16727 32759
rect 16669 32719 16727 32725
rect 17954 32716 17960 32768
rect 18012 32756 18018 32768
rect 19153 32759 19211 32765
rect 19153 32756 19165 32759
rect 18012 32728 19165 32756
rect 18012 32716 18018 32728
rect 19153 32725 19165 32728
rect 19199 32725 19211 32759
rect 19153 32719 19211 32725
rect 19889 32759 19947 32765
rect 19889 32725 19901 32759
rect 19935 32756 19947 32759
rect 19978 32756 19984 32768
rect 19935 32728 19984 32756
rect 19935 32725 19947 32728
rect 19889 32719 19947 32725
rect 19978 32716 19984 32728
rect 20036 32716 20042 32768
rect 20272 32765 20300 32932
rect 20901 32929 20913 32963
rect 20947 32960 20959 32963
rect 24302 32960 24308 32972
rect 20947 32932 24308 32960
rect 20947 32929 20959 32932
rect 20901 32923 20959 32929
rect 23768 32904 23796 32932
rect 24302 32920 24308 32932
rect 24360 32920 24366 32972
rect 21174 32892 21180 32904
rect 21087 32864 21180 32892
rect 21174 32852 21180 32864
rect 21232 32892 21238 32904
rect 21634 32892 21640 32904
rect 21232 32864 21640 32892
rect 21232 32852 21238 32864
rect 21634 32852 21640 32864
rect 21692 32852 21698 32904
rect 22278 32892 22284 32904
rect 22239 32864 22284 32892
rect 22278 32852 22284 32864
rect 22336 32852 22342 32904
rect 23750 32892 23756 32904
rect 23711 32864 23756 32892
rect 23750 32852 23756 32864
rect 23808 32852 23814 32904
rect 24026 32892 24032 32904
rect 23987 32864 24032 32892
rect 24026 32852 24032 32864
rect 24084 32852 24090 32904
rect 20257 32759 20315 32765
rect 20257 32725 20269 32759
rect 20303 32756 20315 32759
rect 20530 32756 20536 32768
rect 20303 32728 20536 32756
rect 20303 32725 20315 32728
rect 20257 32719 20315 32725
rect 20530 32716 20536 32728
rect 20588 32716 20594 32768
rect 21358 32716 21364 32768
rect 21416 32756 21422 32768
rect 22002 32756 22008 32768
rect 21416 32728 22008 32756
rect 21416 32716 21422 32728
rect 22002 32716 22008 32728
rect 22060 32716 22066 32768
rect 26237 32759 26295 32765
rect 26237 32725 26249 32759
rect 26283 32756 26295 32759
rect 26326 32756 26332 32768
rect 26283 32728 26332 32756
rect 26283 32725 26295 32728
rect 26237 32719 26295 32725
rect 26326 32716 26332 32728
rect 26384 32716 26390 32768
rect 1104 32666 28888 32688
rect 1104 32614 5982 32666
rect 6034 32614 6046 32666
rect 6098 32614 6110 32666
rect 6162 32614 6174 32666
rect 6226 32614 15982 32666
rect 16034 32614 16046 32666
rect 16098 32614 16110 32666
rect 16162 32614 16174 32666
rect 16226 32614 25982 32666
rect 26034 32614 26046 32666
rect 26098 32614 26110 32666
rect 26162 32614 26174 32666
rect 26226 32614 28888 32666
rect 1104 32592 28888 32614
rect 3418 32552 3424 32564
rect 3379 32524 3424 32552
rect 3418 32512 3424 32524
rect 3476 32512 3482 32564
rect 4890 32552 4896 32564
rect 4851 32524 4896 32552
rect 4890 32512 4896 32524
rect 4948 32512 4954 32564
rect 5166 32552 5172 32564
rect 5127 32524 5172 32552
rect 5166 32512 5172 32524
rect 5224 32512 5230 32564
rect 5810 32512 5816 32564
rect 5868 32552 5874 32564
rect 6181 32555 6239 32561
rect 6181 32552 6193 32555
rect 5868 32524 6193 32552
rect 5868 32512 5874 32524
rect 6181 32521 6193 32524
rect 6227 32521 6239 32555
rect 7926 32552 7932 32564
rect 7887 32524 7932 32552
rect 6181 32515 6239 32521
rect 7926 32512 7932 32524
rect 7984 32552 7990 32564
rect 7984 32524 8524 32552
rect 7984 32512 7990 32524
rect 4249 32487 4307 32493
rect 4249 32453 4261 32487
rect 4295 32484 4307 32487
rect 5258 32484 5264 32496
rect 4295 32456 5264 32484
rect 4295 32453 4307 32456
rect 4249 32447 4307 32453
rect 5258 32444 5264 32456
rect 5316 32444 5322 32496
rect 7377 32487 7435 32493
rect 7377 32453 7389 32487
rect 7423 32484 7435 32487
rect 8110 32484 8116 32496
rect 7423 32456 8116 32484
rect 7423 32453 7435 32456
rect 7377 32447 7435 32453
rect 8110 32444 8116 32456
rect 8168 32444 8174 32496
rect 4617 32419 4675 32425
rect 4617 32385 4629 32419
rect 4663 32416 4675 32419
rect 8294 32416 8300 32428
rect 4663 32388 8300 32416
rect 4663 32385 4675 32388
rect 4617 32379 4675 32385
rect 8294 32376 8300 32388
rect 8352 32376 8358 32428
rect 8496 32425 8524 32524
rect 9398 32512 9404 32564
rect 9456 32552 9462 32564
rect 9677 32555 9735 32561
rect 9677 32552 9689 32555
rect 9456 32524 9689 32552
rect 9456 32512 9462 32524
rect 9677 32521 9689 32524
rect 9723 32552 9735 32555
rect 10226 32552 10232 32564
rect 9723 32524 10232 32552
rect 9723 32521 9735 32524
rect 9677 32515 9735 32521
rect 10226 32512 10232 32524
rect 10284 32512 10290 32564
rect 11885 32555 11943 32561
rect 11885 32521 11897 32555
rect 11931 32552 11943 32555
rect 12158 32552 12164 32564
rect 11931 32524 12164 32552
rect 11931 32521 11943 32524
rect 11885 32515 11943 32521
rect 12158 32512 12164 32524
rect 12216 32512 12222 32564
rect 12897 32555 12955 32561
rect 12897 32552 12909 32555
rect 12544 32524 12909 32552
rect 8662 32484 8668 32496
rect 8588 32456 8668 32484
rect 8481 32419 8539 32425
rect 8481 32385 8493 32419
rect 8527 32385 8539 32419
rect 8481 32379 8539 32385
rect 4709 32351 4767 32357
rect 4709 32317 4721 32351
rect 4755 32317 4767 32351
rect 4709 32311 4767 32317
rect 5721 32351 5779 32357
rect 5721 32317 5733 32351
rect 5767 32348 5779 32351
rect 7561 32351 7619 32357
rect 5767 32320 6500 32348
rect 5767 32317 5779 32320
rect 5721 32311 5779 32317
rect 4724 32280 4752 32311
rect 5626 32280 5632 32292
rect 4724 32252 5632 32280
rect 5626 32240 5632 32252
rect 5684 32240 5690 32292
rect 6472 32224 6500 32320
rect 7561 32317 7573 32351
rect 7607 32348 7619 32351
rect 7650 32348 7656 32360
rect 7607 32320 7656 32348
rect 7607 32317 7619 32320
rect 7561 32311 7619 32317
rect 7650 32308 7656 32320
rect 7708 32308 7714 32360
rect 8389 32351 8447 32357
rect 8389 32317 8401 32351
rect 8435 32348 8447 32351
rect 8588 32348 8616 32456
rect 8662 32444 8668 32456
rect 8720 32484 8726 32496
rect 12544 32484 12572 32524
rect 12897 32521 12909 32524
rect 12943 32521 12955 32555
rect 12897 32515 12955 32521
rect 13078 32512 13084 32564
rect 13136 32552 13142 32564
rect 13817 32555 13875 32561
rect 13817 32552 13829 32555
rect 13136 32524 13829 32552
rect 13136 32512 13142 32524
rect 13817 32521 13829 32524
rect 13863 32552 13875 32555
rect 15562 32552 15568 32564
rect 13863 32524 14044 32552
rect 13863 32521 13875 32524
rect 13817 32515 13875 32521
rect 8720 32456 8984 32484
rect 8720 32444 8726 32456
rect 8846 32416 8852 32428
rect 8435 32320 8616 32348
rect 8680 32388 8852 32416
rect 8435 32317 8447 32320
rect 8389 32311 8447 32317
rect 8680 32280 8708 32388
rect 8846 32376 8852 32388
rect 8904 32376 8910 32428
rect 8757 32351 8815 32357
rect 8757 32317 8769 32351
rect 8803 32348 8815 32351
rect 8956 32348 8984 32456
rect 12452 32456 12572 32484
rect 12713 32487 12771 32493
rect 8803 32320 8984 32348
rect 9217 32351 9275 32357
rect 8803 32317 8815 32320
rect 8757 32311 8815 32317
rect 9217 32317 9229 32351
rect 9263 32348 9275 32351
rect 10134 32348 10140 32360
rect 9263 32320 10140 32348
rect 9263 32317 9275 32320
rect 9217 32311 9275 32317
rect 10134 32308 10140 32320
rect 10192 32308 10198 32360
rect 10226 32308 10232 32360
rect 10284 32348 10290 32360
rect 10505 32351 10563 32357
rect 10505 32348 10517 32351
rect 10284 32320 10517 32348
rect 10284 32308 10290 32320
rect 10505 32317 10517 32320
rect 10551 32317 10563 32351
rect 10505 32311 10563 32317
rect 10594 32308 10600 32360
rect 10652 32348 10658 32360
rect 10873 32351 10931 32357
rect 10873 32348 10885 32351
rect 10652 32320 10885 32348
rect 10652 32308 10658 32320
rect 10873 32317 10885 32320
rect 10919 32317 10931 32351
rect 11238 32348 11244 32360
rect 11199 32320 11244 32348
rect 10873 32311 10931 32317
rect 11238 32308 11244 32320
rect 11296 32348 11302 32360
rect 12452 32348 12480 32456
rect 12713 32453 12725 32487
rect 12759 32484 12771 32487
rect 12759 32456 13768 32484
rect 12759 32453 12771 32456
rect 12713 32447 12771 32453
rect 12584 32419 12642 32425
rect 12584 32385 12596 32419
rect 12630 32416 12642 32419
rect 13262 32416 13268 32428
rect 12630 32388 13268 32416
rect 12630 32385 12642 32388
rect 12584 32379 12642 32385
rect 13262 32376 13268 32388
rect 13320 32376 13326 32428
rect 12776 32351 12834 32357
rect 12776 32348 12788 32351
rect 11296 32320 12480 32348
rect 12636 32320 12788 32348
rect 11296 32308 11302 32320
rect 8846 32280 8852 32292
rect 8404 32252 8708 32280
rect 8807 32252 8852 32280
rect 8404 32224 8432 32252
rect 8846 32240 8852 32252
rect 8904 32240 8910 32292
rect 12437 32283 12495 32289
rect 12437 32249 12449 32283
rect 12483 32280 12495 32283
rect 12526 32280 12532 32292
rect 12483 32252 12532 32280
rect 12483 32249 12495 32252
rect 12437 32243 12495 32249
rect 12526 32240 12532 32252
rect 12584 32240 12590 32292
rect 3878 32212 3884 32224
rect 3839 32184 3884 32212
rect 3878 32172 3884 32184
rect 3936 32172 3942 32224
rect 5442 32172 5448 32224
rect 5500 32212 5506 32224
rect 5902 32212 5908 32224
rect 5500 32184 5908 32212
rect 5500 32172 5506 32184
rect 5902 32172 5908 32184
rect 5960 32172 5966 32224
rect 6454 32172 6460 32224
rect 6512 32212 6518 32224
rect 6549 32215 6607 32221
rect 6549 32212 6561 32215
rect 6512 32184 6561 32212
rect 6512 32172 6518 32184
rect 6549 32181 6561 32184
rect 6595 32181 6607 32215
rect 6549 32175 6607 32181
rect 8386 32172 8392 32224
rect 8444 32172 8450 32224
rect 8665 32215 8723 32221
rect 8665 32181 8677 32215
rect 8711 32212 8723 32215
rect 8754 32212 8760 32224
rect 8711 32184 8760 32212
rect 8711 32181 8723 32184
rect 8665 32175 8723 32181
rect 8754 32172 8760 32184
rect 8812 32212 8818 32224
rect 9950 32212 9956 32224
rect 8812 32184 9956 32212
rect 8812 32172 8818 32184
rect 9950 32172 9956 32184
rect 10008 32172 10014 32224
rect 10134 32212 10140 32224
rect 10095 32184 10140 32212
rect 10134 32172 10140 32184
rect 10192 32172 10198 32224
rect 12250 32212 12256 32224
rect 12211 32184 12256 32212
rect 12250 32172 12256 32184
rect 12308 32212 12314 32224
rect 12636 32212 12664 32320
rect 12776 32317 12788 32320
rect 12822 32317 12834 32351
rect 13740 32348 13768 32456
rect 14016 32425 14044 32524
rect 15488 32524 15568 32552
rect 14001 32419 14059 32425
rect 14001 32385 14013 32419
rect 14047 32385 14059 32419
rect 14001 32379 14059 32385
rect 13740 32320 14780 32348
rect 12776 32311 12834 32317
rect 14752 32292 14780 32320
rect 14274 32280 14280 32292
rect 14235 32252 14280 32280
rect 14274 32240 14280 32252
rect 14332 32240 14338 32292
rect 14369 32283 14427 32289
rect 14369 32249 14381 32283
rect 14415 32249 14427 32283
rect 14734 32280 14740 32292
rect 14695 32252 14740 32280
rect 14369 32243 14427 32249
rect 12308 32184 12664 32212
rect 12308 32172 12314 32184
rect 12986 32172 12992 32224
rect 13044 32212 13050 32224
rect 13449 32215 13507 32221
rect 13449 32212 13461 32215
rect 13044 32184 13461 32212
rect 13044 32172 13050 32184
rect 13449 32181 13461 32184
rect 13495 32181 13507 32215
rect 13449 32175 13507 32181
rect 13998 32172 14004 32224
rect 14056 32212 14062 32224
rect 14185 32215 14243 32221
rect 14185 32212 14197 32215
rect 14056 32184 14197 32212
rect 14056 32172 14062 32184
rect 14185 32181 14197 32184
rect 14231 32181 14243 32215
rect 14384 32212 14412 32243
rect 14734 32240 14740 32252
rect 14792 32240 14798 32292
rect 15102 32212 15108 32224
rect 14384 32184 15108 32212
rect 14185 32175 14243 32181
rect 15102 32172 15108 32184
rect 15160 32172 15166 32224
rect 15381 32215 15439 32221
rect 15381 32181 15393 32215
rect 15427 32212 15439 32215
rect 15488 32212 15516 32524
rect 15562 32512 15568 32524
rect 15620 32512 15626 32564
rect 16666 32512 16672 32564
rect 16724 32552 16730 32564
rect 17773 32555 17831 32561
rect 17773 32552 17785 32555
rect 16724 32524 17785 32552
rect 16724 32512 16730 32524
rect 17773 32521 17785 32524
rect 17819 32521 17831 32555
rect 21174 32552 21180 32564
rect 21135 32524 21180 32552
rect 17773 32515 17831 32521
rect 21174 32512 21180 32524
rect 21232 32512 21238 32564
rect 23474 32552 23480 32564
rect 23435 32524 23480 32552
rect 23474 32512 23480 32524
rect 23532 32512 23538 32564
rect 18233 32487 18291 32493
rect 18233 32453 18245 32487
rect 18279 32484 18291 32487
rect 18690 32484 18696 32496
rect 18279 32456 18696 32484
rect 18279 32453 18291 32456
rect 18233 32447 18291 32453
rect 18690 32444 18696 32456
rect 18748 32444 18754 32496
rect 22278 32444 22284 32496
rect 22336 32484 22342 32496
rect 22465 32487 22523 32493
rect 22465 32484 22477 32487
rect 22336 32456 22477 32484
rect 22336 32444 22342 32456
rect 22465 32453 22477 32456
rect 22511 32453 22523 32487
rect 22465 32447 22523 32453
rect 22738 32444 22744 32496
rect 22796 32484 22802 32496
rect 23017 32487 23075 32493
rect 23017 32484 23029 32487
rect 22796 32456 23029 32484
rect 22796 32444 22802 32456
rect 23017 32453 23029 32456
rect 23063 32484 23075 32487
rect 27522 32484 27528 32496
rect 23063 32456 27528 32484
rect 23063 32453 23075 32456
rect 23017 32447 23075 32453
rect 27522 32444 27528 32456
rect 27580 32444 27586 32496
rect 15562 32376 15568 32428
rect 15620 32416 15626 32428
rect 15749 32419 15807 32425
rect 15749 32416 15761 32419
rect 15620 32388 15761 32416
rect 15620 32376 15626 32388
rect 15749 32385 15761 32388
rect 15795 32385 15807 32419
rect 15749 32379 15807 32385
rect 15764 32348 15792 32379
rect 15838 32376 15844 32428
rect 15896 32416 15902 32428
rect 15933 32419 15991 32425
rect 15933 32416 15945 32419
rect 15896 32388 15945 32416
rect 15896 32376 15902 32388
rect 15933 32385 15945 32388
rect 15979 32385 15991 32419
rect 15933 32379 15991 32385
rect 19061 32419 19119 32425
rect 19061 32385 19073 32419
rect 19107 32416 19119 32419
rect 19429 32419 19487 32425
rect 19429 32416 19441 32419
rect 19107 32388 19441 32416
rect 19107 32385 19119 32388
rect 19061 32379 19119 32385
rect 19429 32385 19441 32388
rect 19475 32416 19487 32419
rect 19794 32416 19800 32428
rect 19475 32388 19800 32416
rect 19475 32385 19487 32388
rect 19429 32379 19487 32385
rect 19794 32376 19800 32388
rect 19852 32376 19858 32428
rect 23106 32416 23112 32428
rect 21652 32388 23112 32416
rect 16393 32351 16451 32357
rect 16393 32348 16405 32351
rect 15764 32320 16405 32348
rect 16393 32317 16405 32320
rect 16439 32317 16451 32351
rect 16393 32311 16451 32317
rect 16577 32351 16635 32357
rect 16577 32317 16589 32351
rect 16623 32348 16635 32351
rect 16850 32348 16856 32360
rect 16623 32320 16856 32348
rect 16623 32317 16635 32320
rect 16577 32311 16635 32317
rect 16850 32308 16856 32320
rect 16908 32308 16914 32360
rect 16945 32351 17003 32357
rect 16945 32317 16957 32351
rect 16991 32317 17003 32351
rect 16945 32311 17003 32317
rect 17129 32351 17187 32357
rect 17129 32317 17141 32351
rect 17175 32348 17187 32351
rect 17770 32348 17776 32360
rect 17175 32320 17776 32348
rect 17175 32317 17187 32320
rect 17129 32311 17187 32317
rect 16960 32280 16988 32311
rect 17770 32308 17776 32320
rect 17828 32308 17834 32360
rect 18049 32351 18107 32357
rect 18049 32317 18061 32351
rect 18095 32317 18107 32351
rect 19150 32348 19156 32360
rect 19111 32320 19156 32348
rect 18049 32311 18107 32317
rect 17954 32280 17960 32292
rect 16960 32252 17960 32280
rect 17954 32240 17960 32252
rect 18012 32240 18018 32292
rect 18064 32280 18092 32311
rect 19150 32308 19156 32320
rect 19208 32308 19214 32360
rect 21652 32357 21680 32388
rect 23106 32376 23112 32388
rect 23164 32376 23170 32428
rect 21545 32351 21603 32357
rect 21545 32317 21557 32351
rect 21591 32348 21603 32351
rect 21637 32351 21695 32357
rect 21637 32348 21649 32351
rect 21591 32320 21649 32348
rect 21591 32317 21603 32320
rect 21545 32311 21603 32317
rect 21637 32317 21649 32320
rect 21683 32317 21695 32351
rect 21637 32311 21695 32317
rect 21726 32308 21732 32360
rect 21784 32348 21790 32360
rect 22005 32351 22063 32357
rect 22005 32348 22017 32351
rect 21784 32320 22017 32348
rect 21784 32308 21790 32320
rect 22005 32317 22017 32320
rect 22051 32317 22063 32351
rect 22554 32348 22560 32360
rect 22467 32320 22560 32348
rect 22005 32311 22063 32317
rect 22554 32308 22560 32320
rect 22612 32348 22618 32360
rect 23014 32348 23020 32360
rect 22612 32320 23020 32348
rect 22612 32308 22618 32320
rect 23014 32308 23020 32320
rect 23072 32308 23078 32360
rect 18138 32280 18144 32292
rect 18051 32252 18144 32280
rect 18138 32240 18144 32252
rect 18196 32280 18202 32292
rect 18509 32283 18567 32289
rect 18509 32280 18521 32283
rect 18196 32252 18521 32280
rect 18196 32240 18202 32252
rect 18509 32249 18521 32252
rect 18555 32249 18567 32283
rect 18509 32243 18567 32249
rect 20809 32283 20867 32289
rect 20809 32249 20821 32283
rect 20855 32280 20867 32283
rect 20855 32252 21680 32280
rect 20855 32249 20867 32252
rect 20809 32243 20867 32249
rect 21652 32224 21680 32252
rect 15562 32212 15568 32224
rect 15427 32184 15568 32212
rect 15427 32181 15439 32184
rect 15381 32175 15439 32181
rect 15562 32172 15568 32184
rect 15620 32172 15626 32224
rect 16942 32172 16948 32224
rect 17000 32212 17006 32224
rect 17405 32215 17463 32221
rect 17405 32212 17417 32215
rect 17000 32184 17417 32212
rect 17000 32172 17006 32184
rect 17405 32181 17417 32184
rect 17451 32212 17463 32215
rect 17494 32212 17500 32224
rect 17451 32184 17500 32212
rect 17451 32181 17463 32184
rect 17405 32175 17463 32181
rect 17494 32172 17500 32184
rect 17552 32172 17558 32224
rect 18230 32172 18236 32224
rect 18288 32212 18294 32224
rect 18598 32212 18604 32224
rect 18288 32184 18604 32212
rect 18288 32172 18294 32184
rect 18598 32172 18604 32184
rect 18656 32172 18662 32224
rect 21634 32172 21640 32224
rect 21692 32172 21698 32224
rect 23937 32215 23995 32221
rect 23937 32181 23949 32215
rect 23983 32212 23995 32215
rect 24026 32212 24032 32224
rect 23983 32184 24032 32212
rect 23983 32181 23995 32184
rect 23937 32175 23995 32181
rect 24026 32172 24032 32184
rect 24084 32172 24090 32224
rect 24305 32215 24363 32221
rect 24305 32181 24317 32215
rect 24351 32212 24363 32215
rect 24581 32215 24639 32221
rect 24581 32212 24593 32215
rect 24351 32184 24593 32212
rect 24351 32181 24363 32184
rect 24305 32175 24363 32181
rect 24581 32181 24593 32184
rect 24627 32212 24639 32215
rect 24670 32212 24676 32224
rect 24627 32184 24676 32212
rect 24627 32181 24639 32184
rect 24581 32175 24639 32181
rect 24670 32172 24676 32184
rect 24728 32172 24734 32224
rect 1104 32122 28888 32144
rect 1104 32070 10982 32122
rect 11034 32070 11046 32122
rect 11098 32070 11110 32122
rect 11162 32070 11174 32122
rect 11226 32070 20982 32122
rect 21034 32070 21046 32122
rect 21098 32070 21110 32122
rect 21162 32070 21174 32122
rect 21226 32070 28888 32122
rect 1104 32048 28888 32070
rect 2866 32008 2872 32020
rect 2827 31980 2872 32008
rect 2866 31968 2872 31980
rect 2924 31968 2930 32020
rect 4985 32011 5043 32017
rect 4985 31977 4997 32011
rect 5031 32008 5043 32011
rect 5074 32008 5080 32020
rect 5031 31980 5080 32008
rect 5031 31977 5043 31980
rect 4985 31971 5043 31977
rect 5074 31968 5080 31980
rect 5132 31968 5138 32020
rect 5258 32008 5264 32020
rect 5219 31980 5264 32008
rect 5258 31968 5264 31980
rect 5316 31968 5322 32020
rect 8294 32008 8300 32020
rect 5460 31980 7512 32008
rect 8255 31980 8300 32008
rect 3878 31900 3884 31952
rect 3936 31940 3942 31952
rect 4617 31943 4675 31949
rect 4617 31940 4629 31943
rect 3936 31912 4629 31940
rect 3936 31900 3942 31912
rect 4617 31909 4629 31912
rect 4663 31940 4675 31943
rect 5460 31940 5488 31980
rect 5718 31940 5724 31952
rect 4663 31912 5488 31940
rect 5679 31912 5724 31940
rect 4663 31909 4675 31912
rect 4617 31903 4675 31909
rect 5718 31900 5724 31912
rect 5776 31900 5782 31952
rect 7484 31949 7512 31980
rect 8294 31968 8300 31980
rect 8352 31968 8358 32020
rect 8481 32011 8539 32017
rect 8481 31977 8493 32011
rect 8527 32008 8539 32011
rect 8570 32008 8576 32020
rect 8527 31980 8576 32008
rect 8527 31977 8539 31980
rect 8481 31971 8539 31977
rect 8570 31968 8576 31980
rect 8628 31968 8634 32020
rect 9122 32008 9128 32020
rect 9083 31980 9128 32008
rect 9122 31968 9128 31980
rect 9180 31968 9186 32020
rect 9398 32008 9404 32020
rect 9359 31980 9404 32008
rect 9398 31968 9404 31980
rect 9456 32008 9462 32020
rect 9677 32011 9735 32017
rect 9677 32008 9689 32011
rect 9456 31980 9689 32008
rect 9456 31968 9462 31980
rect 9677 31977 9689 31980
rect 9723 31977 9735 32011
rect 10042 32008 10048 32020
rect 10003 31980 10048 32008
rect 9677 31971 9735 31977
rect 10042 31968 10048 31980
rect 10100 31968 10106 32020
rect 10318 31968 10324 32020
rect 10376 32008 10382 32020
rect 10781 32011 10839 32017
rect 10781 32008 10793 32011
rect 10376 31980 10793 32008
rect 10376 31968 10382 31980
rect 10781 31977 10793 31980
rect 10827 31977 10839 32011
rect 10781 31971 10839 31977
rect 11241 32011 11299 32017
rect 11241 31977 11253 32011
rect 11287 32008 11299 32011
rect 11287 31980 12296 32008
rect 11287 31977 11299 31980
rect 11241 31971 11299 31977
rect 7469 31943 7527 31949
rect 7469 31909 7481 31943
rect 7515 31940 7527 31943
rect 7650 31940 7656 31952
rect 7515 31912 7656 31940
rect 7515 31909 7527 31912
rect 7469 31903 7527 31909
rect 7650 31900 7656 31912
rect 7708 31900 7714 31952
rect 8312 31940 8340 31968
rect 9030 31940 9036 31952
rect 8312 31912 9036 31940
rect 9030 31900 9036 31912
rect 9088 31900 9094 31952
rect 1394 31832 1400 31884
rect 1452 31872 1458 31884
rect 1489 31875 1547 31881
rect 1489 31872 1501 31875
rect 1452 31844 1501 31872
rect 1452 31832 1458 31844
rect 1489 31841 1501 31844
rect 1535 31872 1547 31875
rect 1535 31844 1992 31872
rect 1535 31841 1547 31844
rect 1489 31835 1547 31841
rect 1964 31816 1992 31844
rect 5902 31832 5908 31884
rect 5960 31872 5966 31884
rect 6089 31875 6147 31881
rect 6089 31872 6101 31875
rect 5960 31844 6101 31872
rect 5960 31832 5966 31844
rect 6089 31841 6101 31844
rect 6135 31841 6147 31875
rect 6089 31835 6147 31841
rect 7926 31832 7932 31884
rect 7984 31872 7990 31884
rect 8573 31875 8631 31881
rect 8573 31872 8585 31875
rect 7984 31844 8585 31872
rect 7984 31832 7990 31844
rect 8573 31841 8585 31844
rect 8619 31872 8631 31875
rect 9306 31872 9312 31884
rect 8619 31844 9312 31872
rect 8619 31841 8631 31844
rect 8573 31835 8631 31841
rect 9306 31832 9312 31844
rect 9364 31832 9370 31884
rect 9677 31875 9735 31881
rect 9677 31841 9689 31875
rect 9723 31872 9735 31875
rect 9769 31875 9827 31881
rect 9769 31872 9781 31875
rect 9723 31844 9781 31872
rect 9723 31841 9735 31844
rect 9677 31835 9735 31841
rect 9769 31841 9781 31844
rect 9815 31841 9827 31875
rect 9950 31872 9956 31884
rect 9911 31844 9956 31872
rect 9769 31835 9827 31841
rect 9950 31832 9956 31844
rect 10008 31832 10014 31884
rect 10060 31872 10088 31968
rect 10137 31943 10195 31949
rect 10137 31909 10149 31943
rect 10183 31940 10195 31943
rect 10962 31940 10968 31952
rect 10183 31912 10968 31940
rect 10183 31909 10195 31912
rect 10137 31903 10195 31909
rect 10962 31900 10968 31912
rect 11020 31900 11026 31952
rect 12268 31940 12296 31980
rect 12618 31968 12624 32020
rect 12676 32008 12682 32020
rect 13633 32011 13691 32017
rect 13633 32008 13645 32011
rect 12676 31980 13645 32008
rect 12676 31968 12682 31980
rect 13633 31977 13645 31980
rect 13679 31977 13691 32011
rect 13633 31971 13691 31977
rect 13998 31968 14004 32020
rect 14056 32008 14062 32020
rect 14185 32011 14243 32017
rect 14185 32008 14197 32011
rect 14056 31980 14197 32008
rect 14056 31968 14062 31980
rect 14185 31977 14197 31980
rect 14231 31977 14243 32011
rect 14185 31971 14243 31977
rect 14921 32011 14979 32017
rect 14921 31977 14933 32011
rect 14967 32008 14979 32011
rect 15010 32008 15016 32020
rect 14967 31980 15016 32008
rect 14967 31977 14979 31980
rect 14921 31971 14979 31977
rect 15010 31968 15016 31980
rect 15068 31968 15074 32020
rect 15105 32011 15163 32017
rect 15105 31977 15117 32011
rect 15151 32008 15163 32011
rect 15473 32011 15531 32017
rect 15473 32008 15485 32011
rect 15151 31980 15485 32008
rect 15151 31977 15163 31980
rect 15105 31971 15163 31977
rect 15473 31977 15485 31980
rect 15519 31977 15531 32011
rect 15473 31971 15531 31977
rect 17770 31968 17776 32020
rect 17828 32008 17834 32020
rect 18233 32011 18291 32017
rect 18233 32008 18245 32011
rect 17828 31980 18245 32008
rect 17828 31968 17834 31980
rect 18233 31977 18245 31980
rect 18279 32008 18291 32011
rect 19518 32008 19524 32020
rect 18279 31980 19524 32008
rect 18279 31977 18291 31980
rect 18233 31971 18291 31977
rect 19518 31968 19524 31980
rect 19576 31968 19582 32020
rect 20438 31968 20444 32020
rect 20496 32008 20502 32020
rect 20625 32011 20683 32017
rect 20625 32008 20637 32011
rect 20496 31980 20637 32008
rect 20496 31968 20502 31980
rect 20625 31977 20637 31980
rect 20671 31977 20683 32011
rect 21726 32008 21732 32020
rect 21687 31980 21732 32008
rect 20625 31971 20683 31977
rect 21726 31968 21732 31980
rect 21784 31968 21790 32020
rect 22189 32011 22247 32017
rect 22189 31977 22201 32011
rect 22235 32008 22247 32011
rect 22554 32008 22560 32020
rect 22235 31980 22560 32008
rect 22235 31977 22247 31980
rect 22189 31971 22247 31977
rect 22554 31968 22560 31980
rect 22612 31968 22618 32020
rect 23474 32008 23480 32020
rect 23435 31980 23480 32008
rect 23474 31968 23480 31980
rect 23532 31968 23538 32020
rect 12342 31940 12348 31952
rect 12268 31912 12348 31940
rect 10318 31872 10324 31884
rect 10060 31844 10324 31872
rect 10318 31832 10324 31844
rect 10376 31832 10382 31884
rect 10502 31872 10508 31884
rect 10463 31844 10508 31872
rect 10502 31832 10508 31844
rect 10560 31832 10566 31884
rect 11790 31872 11796 31884
rect 11751 31844 11796 31872
rect 11790 31832 11796 31844
rect 11848 31832 11854 31884
rect 12158 31872 12164 31884
rect 12119 31844 12164 31872
rect 12158 31832 12164 31844
rect 12216 31832 12222 31884
rect 12268 31881 12296 31912
rect 12342 31900 12348 31912
rect 12400 31900 12406 31952
rect 12894 31900 12900 31952
rect 12952 31940 12958 31952
rect 13354 31940 13360 31952
rect 12952 31912 13360 31940
rect 12952 31900 12958 31912
rect 13354 31900 13360 31912
rect 13412 31900 13418 31952
rect 13538 31900 13544 31952
rect 13596 31940 13602 31952
rect 14274 31940 14280 31952
rect 13596 31912 14280 31940
rect 13596 31900 13602 31912
rect 14274 31900 14280 31912
rect 14332 31900 14338 31952
rect 17954 31940 17960 31952
rect 17915 31912 17960 31940
rect 17954 31900 17960 31912
rect 18012 31900 18018 31952
rect 19886 31900 19892 31952
rect 19944 31940 19950 31952
rect 20714 31940 20720 31952
rect 19944 31912 20720 31940
rect 19944 31900 19950 31912
rect 20714 31900 20720 31912
rect 20772 31900 20778 31952
rect 23106 31940 23112 31952
rect 23067 31912 23112 31940
rect 23106 31900 23112 31912
rect 23164 31900 23170 31952
rect 12253 31875 12311 31881
rect 12253 31841 12265 31875
rect 12299 31841 12311 31875
rect 12710 31872 12716 31884
rect 12253 31835 12311 31841
rect 12360 31844 12716 31872
rect 1670 31764 1676 31816
rect 1728 31804 1734 31816
rect 1765 31807 1823 31813
rect 1765 31804 1777 31807
rect 1728 31776 1777 31804
rect 1728 31764 1734 31776
rect 1765 31773 1777 31776
rect 1811 31773 1823 31807
rect 1765 31767 1823 31773
rect 1946 31764 1952 31816
rect 2004 31764 2010 31816
rect 5718 31764 5724 31816
rect 5776 31804 5782 31816
rect 5813 31807 5871 31813
rect 5813 31804 5825 31807
rect 5776 31776 5825 31804
rect 5776 31764 5782 31776
rect 5813 31773 5825 31776
rect 5859 31773 5871 31807
rect 5813 31767 5871 31773
rect 11238 31764 11244 31816
rect 11296 31804 11302 31816
rect 11333 31807 11391 31813
rect 11333 31804 11345 31807
rect 11296 31776 11345 31804
rect 11296 31764 11302 31776
rect 11333 31773 11345 31776
rect 11379 31773 11391 31807
rect 11333 31767 11391 31773
rect 8481 31739 8539 31745
rect 8481 31705 8493 31739
rect 8527 31736 8539 31739
rect 8754 31736 8760 31748
rect 8527 31708 8760 31736
rect 8527 31705 8539 31708
rect 8481 31699 8539 31705
rect 8754 31696 8760 31708
rect 8812 31696 8818 31748
rect 12158 31696 12164 31748
rect 12216 31736 12222 31748
rect 12268 31736 12296 31835
rect 12360 31816 12388 31844
rect 12710 31832 12716 31844
rect 12768 31832 12774 31884
rect 13170 31872 13176 31884
rect 13131 31844 13176 31872
rect 13170 31832 13176 31844
rect 13228 31832 13234 31884
rect 13449 31875 13507 31881
rect 13449 31841 13461 31875
rect 13495 31872 13507 31875
rect 13906 31872 13912 31884
rect 13495 31844 13912 31872
rect 13495 31841 13507 31844
rect 13449 31835 13507 31841
rect 13906 31832 13912 31844
rect 13964 31832 13970 31884
rect 13998 31832 14004 31884
rect 14056 31872 14062 31884
rect 14642 31872 14648 31884
rect 14056 31844 14648 31872
rect 14056 31832 14062 31844
rect 14642 31832 14648 31844
rect 14700 31832 14706 31884
rect 15286 31872 15292 31884
rect 15247 31844 15292 31872
rect 15286 31832 15292 31844
rect 15344 31832 15350 31884
rect 15838 31832 15844 31884
rect 15896 31872 15902 31884
rect 15896 31844 16620 31872
rect 15896 31832 15902 31844
rect 12342 31764 12348 31816
rect 12400 31764 12406 31816
rect 12802 31804 12808 31816
rect 12763 31776 12808 31804
rect 12802 31764 12808 31776
rect 12860 31764 12866 31816
rect 13265 31807 13323 31813
rect 13265 31773 13277 31807
rect 13311 31804 13323 31807
rect 13354 31804 13360 31816
rect 13311 31776 13360 31804
rect 13311 31773 13323 31776
rect 13265 31767 13323 31773
rect 13354 31764 13360 31776
rect 13412 31804 13418 31816
rect 13722 31804 13728 31816
rect 13412 31776 13728 31804
rect 13412 31764 13418 31776
rect 13722 31764 13728 31776
rect 13780 31764 13786 31816
rect 14366 31764 14372 31816
rect 14424 31804 14430 31816
rect 15105 31807 15163 31813
rect 15105 31804 15117 31807
rect 14424 31776 15117 31804
rect 14424 31764 14430 31776
rect 15105 31773 15117 31776
rect 15151 31773 15163 31807
rect 15105 31767 15163 31773
rect 15470 31764 15476 31816
rect 15528 31804 15534 31816
rect 16592 31813 16620 31844
rect 16850 31832 16856 31884
rect 16908 31872 16914 31884
rect 18601 31875 18659 31881
rect 18601 31872 18613 31875
rect 16908 31844 18613 31872
rect 16908 31832 16914 31844
rect 18601 31841 18613 31844
rect 18647 31872 18659 31875
rect 18874 31872 18880 31884
rect 18647 31844 18880 31872
rect 18647 31841 18659 31844
rect 18601 31835 18659 31841
rect 18874 31832 18880 31844
rect 18932 31872 18938 31884
rect 19429 31875 19487 31881
rect 19429 31872 19441 31875
rect 18932 31844 19441 31872
rect 18932 31832 18938 31844
rect 19429 31841 19441 31844
rect 19475 31841 19487 31875
rect 19429 31835 19487 31841
rect 19610 31832 19616 31884
rect 19668 31872 19674 31884
rect 19797 31875 19855 31881
rect 19797 31872 19809 31875
rect 19668 31844 19809 31872
rect 19668 31832 19674 31844
rect 19797 31841 19809 31844
rect 19843 31872 19855 31875
rect 20257 31875 20315 31881
rect 20257 31872 20269 31875
rect 19843 31844 20269 31872
rect 19843 31841 19855 31844
rect 19797 31835 19855 31841
rect 20257 31841 20269 31844
rect 20303 31841 20315 31875
rect 20993 31875 21051 31881
rect 20993 31872 21005 31875
rect 20257 31835 20315 31841
rect 20364 31844 21005 31872
rect 16117 31807 16175 31813
rect 16117 31804 16129 31807
rect 15528 31776 16129 31804
rect 15528 31764 15534 31776
rect 16117 31773 16129 31776
rect 16163 31773 16175 31807
rect 16117 31767 16175 31773
rect 16301 31807 16359 31813
rect 16301 31773 16313 31807
rect 16347 31773 16359 31807
rect 16301 31767 16359 31773
rect 16577 31807 16635 31813
rect 16577 31773 16589 31807
rect 16623 31804 16635 31807
rect 17494 31804 17500 31816
rect 16623 31776 17500 31804
rect 16623 31773 16635 31776
rect 16577 31767 16635 31773
rect 12216 31708 12296 31736
rect 12216 31696 12222 31708
rect 13078 31696 13084 31748
rect 13136 31736 13142 31748
rect 13630 31736 13636 31748
rect 13136 31708 13636 31736
rect 13136 31696 13142 31708
rect 13630 31696 13636 31708
rect 13688 31736 13694 31748
rect 14918 31736 14924 31748
rect 13688 31708 14924 31736
rect 13688 31696 13694 31708
rect 14918 31696 14924 31708
rect 14976 31736 14982 31748
rect 15749 31739 15807 31745
rect 15749 31736 15761 31739
rect 14976 31708 15761 31736
rect 14976 31696 14982 31708
rect 15749 31705 15761 31708
rect 15795 31705 15807 31739
rect 15749 31699 15807 31705
rect 15838 31696 15844 31748
rect 15896 31696 15902 31748
rect 7190 31628 7196 31680
rect 7248 31668 7254 31680
rect 7837 31671 7895 31677
rect 7837 31668 7849 31671
rect 7248 31640 7849 31668
rect 7248 31628 7254 31640
rect 7837 31637 7849 31640
rect 7883 31637 7895 31671
rect 7837 31631 7895 31637
rect 8938 31628 8944 31680
rect 8996 31668 9002 31680
rect 12710 31668 12716 31680
rect 8996 31640 12716 31668
rect 8996 31628 9002 31640
rect 12710 31628 12716 31640
rect 12768 31628 12774 31680
rect 15562 31628 15568 31680
rect 15620 31668 15626 31680
rect 15856 31668 15884 31696
rect 15620 31640 15884 31668
rect 16316 31668 16344 31767
rect 17494 31764 17500 31776
rect 17552 31764 17558 31816
rect 18966 31804 18972 31816
rect 18927 31776 18972 31804
rect 18966 31764 18972 31776
rect 19024 31764 19030 31816
rect 19337 31807 19395 31813
rect 19337 31773 19349 31807
rect 19383 31773 19395 31807
rect 19337 31767 19395 31773
rect 19058 31696 19064 31748
rect 19116 31736 19122 31748
rect 19352 31736 19380 31767
rect 19518 31764 19524 31816
rect 19576 31804 19582 31816
rect 19705 31807 19763 31813
rect 19705 31804 19717 31807
rect 19576 31776 19717 31804
rect 19576 31764 19582 31776
rect 19705 31773 19717 31776
rect 19751 31773 19763 31807
rect 19705 31767 19763 31773
rect 19978 31764 19984 31816
rect 20036 31804 20042 31816
rect 20364 31804 20392 31844
rect 20993 31841 21005 31844
rect 21039 31872 21051 31875
rect 21726 31872 21732 31884
rect 21039 31844 21732 31872
rect 21039 31841 21051 31844
rect 20993 31835 21051 31841
rect 21726 31832 21732 31844
rect 21784 31832 21790 31884
rect 22922 31872 22928 31884
rect 22883 31844 22928 31872
rect 22922 31832 22928 31844
rect 22980 31832 22986 31884
rect 23474 31832 23480 31884
rect 23532 31872 23538 31884
rect 23658 31872 23664 31884
rect 23532 31844 23664 31872
rect 23532 31832 23538 31844
rect 23658 31832 23664 31844
rect 23716 31832 23722 31884
rect 20036 31776 20392 31804
rect 20036 31764 20042 31776
rect 20806 31764 20812 31816
rect 20864 31804 20870 31816
rect 20901 31807 20959 31813
rect 20901 31804 20913 31807
rect 20864 31776 20913 31804
rect 20864 31764 20870 31776
rect 20901 31773 20913 31776
rect 20947 31773 20959 31807
rect 20901 31767 20959 31773
rect 19116 31708 19380 31736
rect 19116 31696 19122 31708
rect 17954 31668 17960 31680
rect 16316 31640 17960 31668
rect 15620 31628 15626 31640
rect 17954 31628 17960 31640
rect 18012 31628 18018 31680
rect 21174 31668 21180 31680
rect 21135 31640 21180 31668
rect 21174 31628 21180 31640
rect 21232 31628 21238 31680
rect 1104 31578 28888 31600
rect 1104 31526 5982 31578
rect 6034 31526 6046 31578
rect 6098 31526 6110 31578
rect 6162 31526 6174 31578
rect 6226 31526 15982 31578
rect 16034 31526 16046 31578
rect 16098 31526 16110 31578
rect 16162 31526 16174 31578
rect 16226 31526 25982 31578
rect 26034 31526 26046 31578
rect 26098 31526 26110 31578
rect 26162 31526 26174 31578
rect 26226 31526 28888 31578
rect 1104 31504 28888 31526
rect 6638 31464 6644 31476
rect 6599 31436 6644 31464
rect 6638 31424 6644 31436
rect 6696 31424 6702 31476
rect 7190 31424 7196 31476
rect 7248 31464 7254 31476
rect 7745 31467 7803 31473
rect 7745 31464 7757 31467
rect 7248 31436 7757 31464
rect 7248 31424 7254 31436
rect 7745 31433 7757 31436
rect 7791 31433 7803 31467
rect 7926 31464 7932 31476
rect 7887 31436 7932 31464
rect 7745 31427 7803 31433
rect 7926 31424 7932 31436
rect 7984 31424 7990 31476
rect 8202 31424 8208 31476
rect 8260 31464 8266 31476
rect 8478 31464 8484 31476
rect 8260 31436 8484 31464
rect 8260 31424 8266 31436
rect 8478 31424 8484 31436
rect 8536 31424 8542 31476
rect 8846 31464 8852 31476
rect 8807 31436 8852 31464
rect 8846 31424 8852 31436
rect 8904 31424 8910 31476
rect 11425 31467 11483 31473
rect 11425 31433 11437 31467
rect 11471 31464 11483 31467
rect 11514 31464 11520 31476
rect 11471 31436 11520 31464
rect 11471 31433 11483 31436
rect 11425 31427 11483 31433
rect 11514 31424 11520 31436
rect 11572 31464 11578 31476
rect 11790 31464 11796 31476
rect 11572 31436 11796 31464
rect 11572 31424 11578 31436
rect 11790 31424 11796 31436
rect 11848 31424 11854 31476
rect 11885 31467 11943 31473
rect 11885 31433 11897 31467
rect 11931 31464 11943 31467
rect 12713 31467 12771 31473
rect 11931 31436 12664 31464
rect 11931 31433 11943 31436
rect 11885 31427 11943 31433
rect 5534 31396 5540 31408
rect 5495 31368 5540 31396
rect 5534 31356 5540 31368
rect 5592 31356 5598 31408
rect 6273 31399 6331 31405
rect 6273 31365 6285 31399
rect 6319 31396 6331 31399
rect 6914 31396 6920 31408
rect 6319 31368 6920 31396
rect 6319 31365 6331 31368
rect 6273 31359 6331 31365
rect 6914 31356 6920 31368
rect 6972 31356 6978 31408
rect 7561 31399 7619 31405
rect 7561 31365 7573 31399
rect 7607 31396 7619 31399
rect 12434 31396 12440 31408
rect 7607 31368 12440 31396
rect 7607 31365 7619 31368
rect 7561 31359 7619 31365
rect 7009 31263 7067 31269
rect 7009 31229 7021 31263
rect 7055 31260 7067 31263
rect 7576 31260 7604 31359
rect 12434 31356 12440 31368
rect 12492 31356 12498 31408
rect 12636 31396 12664 31436
rect 12713 31433 12725 31467
rect 12759 31464 12771 31467
rect 13354 31464 13360 31476
rect 12759 31436 13360 31464
rect 12759 31433 12771 31436
rect 12713 31427 12771 31433
rect 13354 31424 13360 31436
rect 13412 31424 13418 31476
rect 13906 31464 13912 31476
rect 13867 31436 13912 31464
rect 13906 31424 13912 31436
rect 13964 31424 13970 31476
rect 14090 31424 14096 31476
rect 14148 31464 14154 31476
rect 14277 31467 14335 31473
rect 14277 31464 14289 31467
rect 14148 31436 14289 31464
rect 14148 31424 14154 31436
rect 14277 31433 14289 31436
rect 14323 31464 14335 31467
rect 14366 31464 14372 31476
rect 14323 31436 14372 31464
rect 14323 31433 14335 31436
rect 14277 31427 14335 31433
rect 14366 31424 14372 31436
rect 14424 31424 14430 31476
rect 15286 31424 15292 31476
rect 15344 31464 15350 31476
rect 15381 31467 15439 31473
rect 15381 31464 15393 31467
rect 15344 31436 15393 31464
rect 15344 31424 15350 31436
rect 15381 31433 15393 31436
rect 15427 31433 15439 31467
rect 16390 31464 16396 31476
rect 16351 31436 16396 31464
rect 15381 31427 15439 31433
rect 16390 31424 16396 31436
rect 16448 31424 16454 31476
rect 16758 31424 16764 31476
rect 16816 31464 16822 31476
rect 17313 31467 17371 31473
rect 17313 31464 17325 31467
rect 16816 31436 17325 31464
rect 16816 31424 16822 31436
rect 17313 31433 17325 31436
rect 17359 31433 17371 31467
rect 19610 31464 19616 31476
rect 19571 31436 19616 31464
rect 17313 31427 17371 31433
rect 19610 31424 19616 31436
rect 19668 31424 19674 31476
rect 21726 31464 21732 31476
rect 21687 31436 21732 31464
rect 21726 31424 21732 31436
rect 21784 31424 21790 31476
rect 14182 31396 14188 31408
rect 12636 31368 14188 31396
rect 14182 31356 14188 31368
rect 14240 31356 14246 31408
rect 16574 31396 16580 31408
rect 14292 31368 16580 31396
rect 7745 31331 7803 31337
rect 7745 31297 7757 31331
rect 7791 31328 7803 31331
rect 8021 31331 8079 31337
rect 8021 31328 8033 31331
rect 7791 31300 8033 31328
rect 7791 31297 7803 31300
rect 7745 31291 7803 31297
rect 8021 31297 8033 31300
rect 8067 31328 8079 31331
rect 8294 31328 8300 31340
rect 8067 31300 8300 31328
rect 8067 31297 8079 31300
rect 8021 31291 8079 31297
rect 8294 31288 8300 31300
rect 8352 31288 8358 31340
rect 8662 31288 8668 31340
rect 8720 31328 8726 31340
rect 8938 31328 8944 31340
rect 8720 31300 8944 31328
rect 8720 31288 8726 31300
rect 8938 31288 8944 31300
rect 8996 31288 9002 31340
rect 9309 31331 9367 31337
rect 9309 31297 9321 31331
rect 9355 31328 9367 31331
rect 10594 31328 10600 31340
rect 9355 31300 10600 31328
rect 9355 31297 9367 31300
rect 9309 31291 9367 31297
rect 10594 31288 10600 31300
rect 10652 31328 10658 31340
rect 10689 31331 10747 31337
rect 10689 31328 10701 31331
rect 10652 31300 10701 31328
rect 10652 31288 10658 31300
rect 10689 31297 10701 31300
rect 10735 31328 10747 31331
rect 11146 31328 11152 31340
rect 10735 31300 11152 31328
rect 10735 31297 10747 31300
rect 10689 31291 10747 31297
rect 11146 31288 11152 31300
rect 11204 31288 11210 31340
rect 11882 31288 11888 31340
rect 11940 31328 11946 31340
rect 12066 31328 12072 31340
rect 11940 31300 12072 31328
rect 11940 31288 11946 31300
rect 12066 31288 12072 31300
rect 12124 31288 12130 31340
rect 12618 31288 12624 31340
rect 12676 31328 12682 31340
rect 12805 31331 12863 31337
rect 12805 31328 12817 31331
rect 12676 31300 12817 31328
rect 12676 31288 12682 31300
rect 12805 31297 12817 31300
rect 12851 31328 12863 31331
rect 14292 31328 14320 31368
rect 16574 31356 16580 31368
rect 16632 31396 16638 31408
rect 16945 31399 17003 31405
rect 16945 31396 16957 31399
rect 16632 31368 16957 31396
rect 16632 31356 16638 31368
rect 16945 31365 16957 31368
rect 16991 31365 17003 31399
rect 16945 31359 17003 31365
rect 12851 31300 14320 31328
rect 12851 31297 12863 31300
rect 12805 31291 12863 31297
rect 7055 31232 7604 31260
rect 8113 31263 8171 31269
rect 7055 31229 7067 31232
rect 7009 31223 7067 31229
rect 8113 31229 8125 31263
rect 8159 31260 8171 31263
rect 8846 31260 8852 31272
rect 8159 31232 8852 31260
rect 8159 31229 8171 31232
rect 8113 31223 8171 31229
rect 8846 31220 8852 31232
rect 8904 31220 8910 31272
rect 9861 31263 9919 31269
rect 9861 31229 9873 31263
rect 9907 31229 9919 31263
rect 10042 31260 10048 31272
rect 10003 31232 10048 31260
rect 9861 31223 9919 31229
rect 1946 31192 1952 31204
rect 1907 31164 1952 31192
rect 1946 31152 1952 31164
rect 2004 31152 2010 31204
rect 8570 31192 8576 31204
rect 8531 31164 8576 31192
rect 8570 31152 8576 31164
rect 8628 31152 8634 31204
rect 9398 31192 9404 31204
rect 9359 31164 9404 31192
rect 9398 31152 9404 31164
rect 9456 31152 9462 31204
rect 9876 31192 9904 31223
rect 10042 31220 10048 31232
rect 10100 31220 10106 31272
rect 10321 31263 10379 31269
rect 10321 31229 10333 31263
rect 10367 31260 10379 31263
rect 10502 31260 10508 31272
rect 10367 31232 10508 31260
rect 10367 31229 10379 31232
rect 10321 31223 10379 31229
rect 10502 31220 10508 31232
rect 10560 31220 10566 31272
rect 10781 31263 10839 31269
rect 10781 31229 10793 31263
rect 10827 31229 10839 31263
rect 10781 31223 10839 31229
rect 9950 31192 9956 31204
rect 9876 31164 9956 31192
rect 9950 31152 9956 31164
rect 10008 31152 10014 31204
rect 1670 31124 1676 31136
rect 1583 31096 1676 31124
rect 1670 31084 1676 31096
rect 1728 31124 1734 31136
rect 2958 31124 2964 31136
rect 1728 31096 2964 31124
rect 1728 31084 1734 31096
rect 2958 31084 2964 31096
rect 3016 31084 3022 31136
rect 4798 31124 4804 31136
rect 4759 31096 4804 31124
rect 4798 31084 4804 31096
rect 4856 31084 4862 31136
rect 5169 31127 5227 31133
rect 5169 31093 5181 31127
rect 5215 31124 5227 31127
rect 5442 31124 5448 31136
rect 5215 31096 5448 31124
rect 5215 31093 5227 31096
rect 5169 31087 5227 31093
rect 5442 31084 5448 31096
rect 5500 31084 5506 31136
rect 5810 31124 5816 31136
rect 5771 31096 5816 31124
rect 5810 31084 5816 31096
rect 5868 31084 5874 31136
rect 7193 31127 7251 31133
rect 7193 31093 7205 31127
rect 7239 31124 7251 31127
rect 8662 31124 8668 31136
rect 7239 31096 8668 31124
rect 7239 31093 7251 31096
rect 7193 31087 7251 31093
rect 8662 31084 8668 31096
rect 8720 31084 8726 31136
rect 9122 31084 9128 31136
rect 9180 31124 9186 31136
rect 10796 31124 10824 31223
rect 10962 31220 10968 31272
rect 11020 31260 11026 31272
rect 11790 31260 11796 31272
rect 11020 31232 11796 31260
rect 11020 31220 11026 31232
rect 11790 31220 11796 31232
rect 11848 31220 11854 31272
rect 12710 31220 12716 31272
rect 12768 31260 12774 31272
rect 13354 31260 13360 31272
rect 12768 31232 13360 31260
rect 12768 31220 12774 31232
rect 13188 31201 13216 31232
rect 13354 31220 13360 31232
rect 13412 31260 13418 31272
rect 14182 31260 14188 31272
rect 13412 31232 14188 31260
rect 13412 31220 13418 31232
rect 14182 31220 14188 31232
rect 14240 31220 14246 31272
rect 14292 31204 14320 31300
rect 14366 31288 14372 31340
rect 14424 31328 14430 31340
rect 14826 31328 14832 31340
rect 14424 31300 14504 31328
rect 14424 31288 14430 31300
rect 13173 31195 13231 31201
rect 13173 31161 13185 31195
rect 13219 31161 13231 31195
rect 13173 31155 13231 31161
rect 13541 31195 13599 31201
rect 13541 31161 13553 31195
rect 13587 31192 13599 31195
rect 13722 31192 13728 31204
rect 13587 31164 13728 31192
rect 13587 31161 13599 31164
rect 13541 31155 13599 31161
rect 13722 31152 13728 31164
rect 13780 31152 13786 31204
rect 14274 31152 14280 31204
rect 14332 31192 14338 31204
rect 14369 31195 14427 31201
rect 14369 31192 14381 31195
rect 14332 31164 14381 31192
rect 14332 31152 14338 31164
rect 14369 31161 14381 31164
rect 14415 31161 14427 31195
rect 14476 31192 14504 31300
rect 14568 31300 14832 31328
rect 14568 31269 14596 31300
rect 14826 31288 14832 31300
rect 14884 31328 14890 31340
rect 15749 31331 15807 31337
rect 15749 31328 15761 31331
rect 14884 31300 15761 31328
rect 14884 31288 14890 31300
rect 15749 31297 15761 31300
rect 15795 31297 15807 31331
rect 15749 31291 15807 31297
rect 15838 31288 15844 31340
rect 15896 31328 15902 31340
rect 16298 31328 16304 31340
rect 15896 31300 16304 31328
rect 15896 31288 15902 31300
rect 16298 31288 16304 31300
rect 16356 31288 16362 31340
rect 17954 31288 17960 31340
rect 18012 31328 18018 31340
rect 18049 31331 18107 31337
rect 18049 31328 18061 31331
rect 18012 31300 18061 31328
rect 18012 31288 18018 31300
rect 18049 31297 18061 31300
rect 18095 31297 18107 31331
rect 21361 31331 21419 31337
rect 21361 31328 21373 31331
rect 18049 31291 18107 31297
rect 20548 31300 21373 31328
rect 20548 31272 20576 31300
rect 21361 31297 21373 31300
rect 21407 31297 21419 31331
rect 21361 31291 21419 31297
rect 23477 31331 23535 31337
rect 23477 31297 23489 31331
rect 23523 31328 23535 31331
rect 23934 31328 23940 31340
rect 23523 31300 23940 31328
rect 23523 31297 23535 31300
rect 23477 31291 23535 31297
rect 23934 31288 23940 31300
rect 23992 31288 23998 31340
rect 26053 31331 26111 31337
rect 26053 31297 26065 31331
rect 26099 31328 26111 31331
rect 27614 31328 27620 31340
rect 26099 31300 26464 31328
rect 27575 31300 27620 31328
rect 26099 31297 26111 31300
rect 26053 31291 26111 31297
rect 26436 31272 26464 31300
rect 27614 31288 27620 31300
rect 27672 31288 27678 31340
rect 14553 31263 14611 31269
rect 14553 31229 14565 31263
rect 14599 31229 14611 31263
rect 16482 31260 16488 31272
rect 16443 31232 16488 31260
rect 14553 31223 14611 31229
rect 16482 31220 16488 31232
rect 16540 31220 16546 31272
rect 16574 31220 16580 31272
rect 16632 31260 16638 31272
rect 17681 31263 17739 31269
rect 17681 31260 17693 31263
rect 16632 31232 17693 31260
rect 16632 31220 16638 31232
rect 17681 31229 17693 31232
rect 17727 31229 17739 31263
rect 18325 31263 18383 31269
rect 18325 31260 18337 31263
rect 17681 31223 17739 31229
rect 17972 31232 18337 31260
rect 14645 31195 14703 31201
rect 14645 31192 14657 31195
rect 14476 31164 14657 31192
rect 14369 31155 14427 31161
rect 14645 31161 14657 31164
rect 14691 31161 14703 31195
rect 14645 31155 14703 31161
rect 14737 31195 14795 31201
rect 14737 31161 14749 31195
rect 14783 31161 14795 31195
rect 15102 31192 15108 31204
rect 15063 31164 15108 31192
rect 14737 31155 14795 31161
rect 12250 31124 12256 31136
rect 9180 31096 10824 31124
rect 12211 31096 12256 31124
rect 9180 31084 9186 31096
rect 12250 31084 12256 31096
rect 12308 31084 12314 31136
rect 12526 31084 12532 31136
rect 12584 31124 12590 31136
rect 12989 31127 13047 31133
rect 12989 31124 13001 31127
rect 12584 31096 13001 31124
rect 12584 31084 12590 31096
rect 12989 31093 13001 31096
rect 13035 31093 13047 31127
rect 12989 31087 13047 31093
rect 13081 31127 13139 31133
rect 13081 31093 13093 31127
rect 13127 31124 13139 31127
rect 13814 31124 13820 31136
rect 13127 31096 13820 31124
rect 13127 31093 13139 31096
rect 13081 31087 13139 31093
rect 13814 31084 13820 31096
rect 13872 31084 13878 31136
rect 14752 31124 14780 31155
rect 15102 31152 15108 31164
rect 15160 31152 15166 31204
rect 16850 31152 16856 31204
rect 16908 31192 16914 31204
rect 17972 31192 18000 31232
rect 18325 31229 18337 31232
rect 18371 31260 18383 31263
rect 19058 31260 19064 31272
rect 18371 31232 19064 31260
rect 18371 31229 18383 31232
rect 18325 31223 18383 31229
rect 19058 31220 19064 31232
rect 19116 31220 19122 31272
rect 20530 31260 20536 31272
rect 20491 31232 20536 31260
rect 20530 31220 20536 31232
rect 20588 31220 20594 31272
rect 20717 31263 20775 31269
rect 20717 31229 20729 31263
rect 20763 31260 20775 31263
rect 20806 31260 20812 31272
rect 20763 31232 20812 31260
rect 20763 31229 20775 31232
rect 20717 31223 20775 31229
rect 20732 31192 20760 31223
rect 20806 31220 20812 31232
rect 20864 31220 20870 31272
rect 20898 31220 20904 31272
rect 20956 31260 20962 31272
rect 21913 31263 21971 31269
rect 21913 31260 21925 31263
rect 20956 31232 21925 31260
rect 20956 31220 20962 31232
rect 21913 31229 21925 31232
rect 21959 31260 21971 31263
rect 22373 31263 22431 31269
rect 22373 31260 22385 31263
rect 21959 31232 22385 31260
rect 21959 31229 21971 31232
rect 21913 31223 21971 31229
rect 22373 31229 22385 31232
rect 22419 31229 22431 31263
rect 22373 31223 22431 31229
rect 22833 31263 22891 31269
rect 22833 31229 22845 31263
rect 22879 31260 22891 31263
rect 22922 31260 22928 31272
rect 22879 31232 22928 31260
rect 22879 31229 22891 31232
rect 22833 31223 22891 31229
rect 22922 31220 22928 31232
rect 22980 31220 22986 31272
rect 23661 31263 23719 31269
rect 23661 31229 23673 31263
rect 23707 31260 23719 31263
rect 23750 31260 23756 31272
rect 23707 31232 23756 31260
rect 23707 31229 23719 31232
rect 23661 31223 23719 31229
rect 23750 31220 23756 31232
rect 23808 31260 23814 31272
rect 24670 31260 24676 31272
rect 23808 31232 24676 31260
rect 23808 31220 23814 31232
rect 24670 31220 24676 31232
rect 24728 31260 24734 31272
rect 25774 31260 25780 31272
rect 24728 31232 25780 31260
rect 24728 31220 24734 31232
rect 25774 31220 25780 31232
rect 25832 31260 25838 31272
rect 26145 31263 26203 31269
rect 26145 31260 26157 31263
rect 25832 31232 26157 31260
rect 25832 31220 25838 31232
rect 26145 31229 26157 31232
rect 26191 31260 26203 31263
rect 26234 31260 26240 31272
rect 26191 31232 26240 31260
rect 26191 31229 26203 31232
rect 26145 31223 26203 31229
rect 26234 31220 26240 31232
rect 26292 31220 26298 31272
rect 26418 31260 26424 31272
rect 26379 31232 26424 31260
rect 26418 31220 26424 31232
rect 26476 31220 26482 31272
rect 16908 31164 18000 31192
rect 20364 31164 20760 31192
rect 16908 31152 16914 31164
rect 15562 31124 15568 31136
rect 14752 31096 15568 31124
rect 15562 31084 15568 31096
rect 15620 31084 15626 31136
rect 19978 31124 19984 31136
rect 19939 31096 19984 31124
rect 19978 31084 19984 31096
rect 20036 31124 20042 31136
rect 20364 31133 20392 31164
rect 20349 31127 20407 31133
rect 20349 31124 20361 31127
rect 20036 31096 20361 31124
rect 20036 31084 20042 31096
rect 20349 31093 20361 31096
rect 20395 31093 20407 31127
rect 20732 31124 20760 31164
rect 21085 31195 21143 31201
rect 21085 31161 21097 31195
rect 21131 31192 21143 31195
rect 21726 31192 21732 31204
rect 21131 31164 21732 31192
rect 21131 31161 21143 31164
rect 21085 31155 21143 31161
rect 21726 31152 21732 31164
rect 21784 31152 21790 31204
rect 22097 31127 22155 31133
rect 22097 31124 22109 31127
rect 20732 31096 22109 31124
rect 20349 31087 20407 31093
rect 22097 31093 22109 31096
rect 22143 31093 22155 31127
rect 25038 31124 25044 31136
rect 24999 31096 25044 31124
rect 22097 31087 22155 31093
rect 25038 31084 25044 31096
rect 25096 31084 25102 31136
rect 1104 31034 28888 31056
rect 1104 30982 10982 31034
rect 11034 30982 11046 31034
rect 11098 30982 11110 31034
rect 11162 30982 11174 31034
rect 11226 30982 20982 31034
rect 21034 30982 21046 31034
rect 21098 30982 21110 31034
rect 21162 30982 21174 31034
rect 21226 30982 28888 31034
rect 1104 30960 28888 30982
rect 5997 30923 6055 30929
rect 5997 30889 6009 30923
rect 6043 30920 6055 30923
rect 6362 30920 6368 30932
rect 6043 30892 6368 30920
rect 6043 30889 6055 30892
rect 5997 30883 6055 30889
rect 6362 30880 6368 30892
rect 6420 30880 6426 30932
rect 7190 30880 7196 30932
rect 7248 30920 7254 30932
rect 7466 30920 7472 30932
rect 7248 30892 7472 30920
rect 7248 30880 7254 30892
rect 7466 30880 7472 30892
rect 7524 30880 7530 30932
rect 9953 30923 10011 30929
rect 9953 30889 9965 30923
rect 9999 30920 10011 30923
rect 10410 30920 10416 30932
rect 9999 30892 10416 30920
rect 9999 30889 10011 30892
rect 9953 30883 10011 30889
rect 10410 30880 10416 30892
rect 10468 30880 10474 30932
rect 10505 30923 10563 30929
rect 10505 30889 10517 30923
rect 10551 30920 10563 30923
rect 10870 30920 10876 30932
rect 10551 30892 10876 30920
rect 10551 30889 10563 30892
rect 10505 30883 10563 30889
rect 10870 30880 10876 30892
rect 10928 30880 10934 30932
rect 11701 30923 11759 30929
rect 11701 30889 11713 30923
rect 11747 30920 11759 30923
rect 12618 30920 12624 30932
rect 11747 30892 12624 30920
rect 11747 30889 11759 30892
rect 11701 30883 11759 30889
rect 12618 30880 12624 30892
rect 12676 30880 12682 30932
rect 13170 30880 13176 30932
rect 13228 30920 13234 30932
rect 13449 30923 13507 30929
rect 13449 30920 13461 30923
rect 13228 30892 13461 30920
rect 13228 30880 13234 30892
rect 13449 30889 13461 30892
rect 13495 30889 13507 30923
rect 13814 30920 13820 30932
rect 13775 30892 13820 30920
rect 13449 30883 13507 30889
rect 13814 30880 13820 30892
rect 13872 30880 13878 30932
rect 16666 30920 16672 30932
rect 16627 30892 16672 30920
rect 16666 30880 16672 30892
rect 16724 30880 16730 30932
rect 17954 30920 17960 30932
rect 17788 30892 17960 30920
rect 8754 30812 8760 30864
rect 8812 30852 8818 30864
rect 9401 30855 9459 30861
rect 9401 30852 9413 30855
rect 8812 30824 9413 30852
rect 8812 30812 8818 30824
rect 9401 30821 9413 30824
rect 9447 30852 9459 30855
rect 9582 30852 9588 30864
rect 9447 30824 9588 30852
rect 9447 30821 9459 30824
rect 9401 30815 9459 30821
rect 9582 30812 9588 30824
rect 9640 30852 9646 30864
rect 10321 30855 10379 30861
rect 10321 30852 10333 30855
rect 9640 30824 10333 30852
rect 9640 30812 9646 30824
rect 10321 30821 10333 30824
rect 10367 30821 10379 30855
rect 10689 30855 10747 30861
rect 10689 30852 10701 30855
rect 10321 30815 10379 30821
rect 10520 30824 10701 30852
rect 4798 30744 4804 30796
rect 4856 30784 4862 30796
rect 5718 30784 5724 30796
rect 4856 30756 5724 30784
rect 4856 30744 4862 30756
rect 5718 30744 5724 30756
rect 5776 30784 5782 30796
rect 6089 30787 6147 30793
rect 6089 30784 6101 30787
rect 5776 30756 6101 30784
rect 5776 30744 5782 30756
rect 6089 30753 6101 30756
rect 6135 30784 6147 30787
rect 6638 30784 6644 30796
rect 6135 30756 6644 30784
rect 6135 30753 6147 30756
rect 6089 30747 6147 30753
rect 6638 30744 6644 30756
rect 6696 30744 6702 30796
rect 8573 30787 8631 30793
rect 8573 30753 8585 30787
rect 8619 30784 8631 30787
rect 8662 30784 8668 30796
rect 8619 30756 8668 30784
rect 8619 30753 8631 30756
rect 8573 30747 8631 30753
rect 8662 30744 8668 30756
rect 8720 30744 8726 30796
rect 9122 30784 9128 30796
rect 9083 30756 9128 30784
rect 9122 30744 9128 30756
rect 9180 30744 9186 30796
rect 9306 30744 9312 30796
rect 9364 30784 9370 30796
rect 10042 30784 10048 30796
rect 9364 30756 10048 30784
rect 9364 30744 9370 30756
rect 10042 30744 10048 30756
rect 10100 30744 10106 30796
rect 6365 30719 6423 30725
rect 6365 30685 6377 30719
rect 6411 30716 6423 30719
rect 6822 30716 6828 30728
rect 6411 30688 6828 30716
rect 6411 30685 6423 30688
rect 6365 30679 6423 30685
rect 6822 30676 6828 30688
rect 6880 30676 6886 30728
rect 8113 30719 8171 30725
rect 8113 30685 8125 30719
rect 8159 30716 8171 30719
rect 9950 30716 9956 30728
rect 8159 30688 9956 30716
rect 8159 30685 8171 30688
rect 8113 30679 8171 30685
rect 9950 30676 9956 30688
rect 10008 30716 10014 30728
rect 10520 30716 10548 30824
rect 10689 30821 10701 30824
rect 10735 30821 10747 30855
rect 10689 30815 10747 30821
rect 10962 30812 10968 30864
rect 11020 30852 11026 30864
rect 11057 30855 11115 30861
rect 11057 30852 11069 30855
rect 11020 30824 11069 30852
rect 11020 30812 11026 30824
rect 11057 30821 11069 30824
rect 11103 30821 11115 30855
rect 11057 30815 11115 30821
rect 12250 30812 12256 30864
rect 12308 30852 12314 30864
rect 12713 30855 12771 30861
rect 12713 30852 12725 30855
rect 12308 30824 12725 30852
rect 12308 30812 12314 30824
rect 12713 30821 12725 30824
rect 12759 30821 12771 30855
rect 12713 30815 12771 30821
rect 12805 30855 12863 30861
rect 12805 30821 12817 30855
rect 12851 30852 12863 30855
rect 13078 30852 13084 30864
rect 12851 30824 13084 30852
rect 12851 30821 12863 30824
rect 12805 30815 12863 30821
rect 13078 30812 13084 30824
rect 13136 30812 13142 30864
rect 15010 30812 15016 30864
rect 15068 30852 15074 30864
rect 16301 30855 16359 30861
rect 16301 30852 16313 30855
rect 15068 30824 16313 30852
rect 15068 30812 15074 30824
rect 16301 30821 16313 30824
rect 16347 30821 16359 30855
rect 16301 30815 16359 30821
rect 10597 30787 10655 30793
rect 10597 30753 10609 30787
rect 10643 30753 10655 30787
rect 10597 30747 10655 30753
rect 10008 30688 10548 30716
rect 10612 30716 10640 30747
rect 11514 30744 11520 30796
rect 11572 30784 11578 30796
rect 12345 30787 12403 30793
rect 12345 30784 12357 30787
rect 11572 30756 12357 30784
rect 11572 30744 11578 30756
rect 12345 30753 12357 30756
rect 12391 30753 12403 30787
rect 12345 30747 12403 30753
rect 12434 30744 12440 30796
rect 12492 30784 12498 30796
rect 12621 30787 12679 30793
rect 12492 30756 12572 30784
rect 12492 30744 12498 30756
rect 10962 30716 10968 30728
rect 10612 30688 10968 30716
rect 10008 30676 10014 30688
rect 5626 30608 5632 30660
rect 5684 30608 5690 30660
rect 8757 30651 8815 30657
rect 8757 30617 8769 30651
rect 8803 30648 8815 30651
rect 8938 30648 8944 30660
rect 8803 30620 8944 30648
rect 8803 30617 8815 30620
rect 8757 30611 8815 30617
rect 8938 30608 8944 30620
rect 8996 30648 9002 30660
rect 10612 30648 10640 30688
rect 10962 30676 10968 30688
rect 11020 30676 11026 30728
rect 12069 30719 12127 30725
rect 12069 30685 12081 30719
rect 12115 30716 12127 30719
rect 12158 30716 12164 30728
rect 12115 30688 12164 30716
rect 12115 30685 12127 30688
rect 12069 30679 12127 30685
rect 12158 30676 12164 30688
rect 12216 30676 12222 30728
rect 12544 30716 12572 30756
rect 12621 30753 12633 30787
rect 12667 30784 12679 30787
rect 13170 30784 13176 30796
rect 12667 30756 12848 30784
rect 13131 30756 13176 30784
rect 12667 30753 12679 30756
rect 12621 30747 12679 30753
rect 12710 30716 12716 30728
rect 12544 30688 12716 30716
rect 12710 30676 12716 30688
rect 12768 30676 12774 30728
rect 12820 30716 12848 30756
rect 13170 30744 13176 30756
rect 13228 30744 13234 30796
rect 14185 30787 14243 30793
rect 14185 30753 14197 30787
rect 14231 30784 14243 30787
rect 14274 30784 14280 30796
rect 14231 30756 14280 30784
rect 14231 30753 14243 30756
rect 14185 30747 14243 30753
rect 14274 30744 14280 30756
rect 14332 30744 14338 30796
rect 14458 30744 14464 30796
rect 14516 30744 14522 30796
rect 15286 30784 15292 30796
rect 15247 30756 15292 30784
rect 15286 30744 15292 30756
rect 15344 30744 15350 30796
rect 15378 30744 15384 30796
rect 15436 30784 15442 30796
rect 15565 30787 15623 30793
rect 15565 30784 15577 30787
rect 15436 30756 15577 30784
rect 15436 30744 15442 30756
rect 15565 30753 15577 30756
rect 15611 30753 15623 30787
rect 15565 30747 15623 30753
rect 17681 30787 17739 30793
rect 17681 30753 17693 30787
rect 17727 30784 17739 30787
rect 17788 30784 17816 30892
rect 17954 30880 17960 30892
rect 18012 30880 18018 30932
rect 21910 30880 21916 30932
rect 21968 30920 21974 30932
rect 23750 30920 23756 30932
rect 21968 30892 23756 30920
rect 21968 30880 21974 30892
rect 23750 30880 23756 30892
rect 23808 30880 23814 30932
rect 21453 30855 21511 30861
rect 21453 30821 21465 30855
rect 21499 30852 21511 30855
rect 22186 30852 22192 30864
rect 21499 30824 22192 30852
rect 21499 30821 21511 30824
rect 21453 30815 21511 30821
rect 22186 30812 22192 30824
rect 22244 30812 22250 30864
rect 19150 30784 19156 30796
rect 17727 30756 19156 30784
rect 17727 30753 17739 30756
rect 17681 30747 17739 30753
rect 19150 30744 19156 30756
rect 19208 30744 19214 30796
rect 20898 30784 20904 30796
rect 20859 30756 20904 30784
rect 20898 30744 20904 30756
rect 20956 30744 20962 30796
rect 13262 30716 13268 30728
rect 12820 30688 13268 30716
rect 13262 30676 13268 30688
rect 13320 30676 13326 30728
rect 14476 30716 14504 30744
rect 13556 30688 14504 30716
rect 14737 30719 14795 30725
rect 8996 30620 10640 30648
rect 8996 30608 9002 30620
rect 11790 30608 11796 30660
rect 11848 30648 11854 30660
rect 12618 30648 12624 30660
rect 11848 30620 12624 30648
rect 11848 30608 11854 30620
rect 12618 30608 12624 30620
rect 12676 30648 12682 30660
rect 13446 30648 13452 30660
rect 12676 30620 13452 30648
rect 12676 30608 12682 30620
rect 13446 30608 13452 30620
rect 13504 30608 13510 30660
rect 5534 30580 5540 30592
rect 5495 30552 5540 30580
rect 5534 30540 5540 30552
rect 5592 30540 5598 30592
rect 5644 30580 5672 30608
rect 6362 30580 6368 30592
rect 5644 30552 6368 30580
rect 6362 30540 6368 30552
rect 6420 30540 6426 30592
rect 7466 30580 7472 30592
rect 7427 30552 7472 30580
rect 7466 30540 7472 30552
rect 7524 30540 7530 30592
rect 8481 30583 8539 30589
rect 8481 30549 8493 30583
rect 8527 30580 8539 30583
rect 9306 30580 9312 30592
rect 8527 30552 9312 30580
rect 8527 30549 8539 30552
rect 8481 30543 8539 30549
rect 9306 30540 9312 30552
rect 9364 30540 9370 30592
rect 9858 30540 9864 30592
rect 9916 30580 9922 30592
rect 10226 30580 10232 30592
rect 9916 30552 10232 30580
rect 9916 30540 9922 30552
rect 10226 30540 10232 30552
rect 10284 30540 10290 30592
rect 11514 30540 11520 30592
rect 11572 30580 11578 30592
rect 12161 30583 12219 30589
rect 12161 30580 12173 30583
rect 11572 30552 12173 30580
rect 11572 30540 11578 30552
rect 12161 30549 12173 30552
rect 12207 30549 12219 30583
rect 12161 30543 12219 30549
rect 13354 30540 13360 30592
rect 13412 30580 13418 30592
rect 13556 30580 13584 30688
rect 14737 30685 14749 30719
rect 14783 30716 14795 30719
rect 14918 30716 14924 30728
rect 14783 30688 14924 30716
rect 14783 30685 14795 30688
rect 14737 30679 14795 30685
rect 14918 30676 14924 30688
rect 14976 30676 14982 30728
rect 16025 30719 16083 30725
rect 16025 30685 16037 30719
rect 16071 30716 16083 30719
rect 16574 30716 16580 30728
rect 16071 30688 16580 30716
rect 16071 30685 16083 30688
rect 16025 30679 16083 30685
rect 16574 30676 16580 30688
rect 16632 30676 16638 30728
rect 16666 30676 16672 30728
rect 16724 30716 16730 30728
rect 17037 30719 17095 30725
rect 17037 30716 17049 30719
rect 16724 30688 17049 30716
rect 16724 30676 16730 30688
rect 17037 30685 17049 30688
rect 17083 30685 17095 30719
rect 17037 30679 17095 30685
rect 17957 30719 18015 30725
rect 17957 30685 17969 30719
rect 18003 30716 18015 30719
rect 18138 30716 18144 30728
rect 18003 30688 18144 30716
rect 18003 30685 18015 30688
rect 17957 30679 18015 30685
rect 18138 30676 18144 30688
rect 18196 30676 18202 30728
rect 19058 30676 19064 30728
rect 19116 30716 19122 30728
rect 19886 30716 19892 30728
rect 19116 30688 19892 30716
rect 19116 30676 19122 30688
rect 19886 30676 19892 30688
rect 19944 30716 19950 30728
rect 20349 30719 20407 30725
rect 20349 30716 20361 30719
rect 19944 30688 20361 30716
rect 19944 30676 19950 30688
rect 20349 30685 20361 30688
rect 20395 30685 20407 30719
rect 20349 30679 20407 30685
rect 21821 30719 21879 30725
rect 21821 30685 21833 30719
rect 21867 30716 21879 30719
rect 22186 30716 22192 30728
rect 21867 30688 22192 30716
rect 21867 30685 21879 30688
rect 21821 30679 21879 30685
rect 22186 30676 22192 30688
rect 22244 30716 22250 30728
rect 23382 30716 23388 30728
rect 22244 30688 23388 30716
rect 22244 30676 22250 30688
rect 23382 30676 23388 30688
rect 23440 30676 23446 30728
rect 13630 30608 13636 30660
rect 13688 30648 13694 30660
rect 14369 30651 14427 30657
rect 14369 30648 14381 30651
rect 13688 30620 14381 30648
rect 13688 30608 13694 30620
rect 14369 30617 14381 30620
rect 14415 30648 14427 30651
rect 14458 30648 14464 30660
rect 14415 30620 14464 30648
rect 14415 30617 14427 30620
rect 14369 30611 14427 30617
rect 14458 30608 14464 30620
rect 14516 30608 14522 30660
rect 15381 30651 15439 30657
rect 15381 30617 15393 30651
rect 15427 30648 15439 30651
rect 16298 30648 16304 30660
rect 15427 30620 16304 30648
rect 15427 30617 15439 30620
rect 15381 30611 15439 30617
rect 16298 30608 16304 30620
rect 16356 30608 16362 30660
rect 19334 30608 19340 30660
rect 19392 30648 19398 30660
rect 19981 30651 20039 30657
rect 19981 30648 19993 30651
rect 19392 30620 19993 30648
rect 19392 30608 19398 30620
rect 19981 30617 19993 30620
rect 20027 30617 20039 30651
rect 21082 30648 21088 30660
rect 21043 30620 21088 30648
rect 19981 30611 20039 30617
rect 21082 30608 21088 30620
rect 21140 30648 21146 30660
rect 22094 30648 22100 30660
rect 21140 30620 22100 30648
rect 21140 30608 21146 30620
rect 22094 30608 22100 30620
rect 22152 30608 22158 30660
rect 13412 30552 13584 30580
rect 13412 30540 13418 30552
rect 14734 30540 14740 30592
rect 14792 30580 14798 30592
rect 15013 30583 15071 30589
rect 15013 30580 15025 30583
rect 14792 30552 15025 30580
rect 14792 30540 14798 30552
rect 15013 30549 15025 30552
rect 15059 30549 15071 30583
rect 15013 30543 15071 30549
rect 17589 30583 17647 30589
rect 17589 30549 17601 30583
rect 17635 30580 17647 30583
rect 17954 30580 17960 30592
rect 17635 30552 17960 30580
rect 17635 30549 17647 30552
rect 17589 30543 17647 30549
rect 17954 30540 17960 30552
rect 18012 30540 18018 30592
rect 19058 30580 19064 30592
rect 19019 30552 19064 30580
rect 19058 30540 19064 30552
rect 19116 30540 19122 30592
rect 19610 30580 19616 30592
rect 19571 30552 19616 30580
rect 19610 30540 19616 30552
rect 19668 30540 19674 30592
rect 25774 30540 25780 30592
rect 25832 30580 25838 30592
rect 26145 30583 26203 30589
rect 26145 30580 26157 30583
rect 25832 30552 26157 30580
rect 25832 30540 25838 30552
rect 26145 30549 26157 30552
rect 26191 30549 26203 30583
rect 26145 30543 26203 30549
rect 1104 30490 28888 30512
rect 1104 30438 5982 30490
rect 6034 30438 6046 30490
rect 6098 30438 6110 30490
rect 6162 30438 6174 30490
rect 6226 30438 15982 30490
rect 16034 30438 16046 30490
rect 16098 30438 16110 30490
rect 16162 30438 16174 30490
rect 16226 30438 25982 30490
rect 26034 30438 26046 30490
rect 26098 30438 26110 30490
rect 26162 30438 26174 30490
rect 26226 30438 28888 30490
rect 1104 30416 28888 30438
rect 8662 30376 8668 30388
rect 8623 30348 8668 30376
rect 8662 30336 8668 30348
rect 8720 30336 8726 30388
rect 9766 30336 9772 30388
rect 9824 30376 9830 30388
rect 10597 30379 10655 30385
rect 9824 30348 9996 30376
rect 9824 30336 9830 30348
rect 9968 30320 9996 30348
rect 10597 30345 10609 30379
rect 10643 30376 10655 30379
rect 10870 30376 10876 30388
rect 10643 30348 10876 30376
rect 10643 30345 10655 30348
rect 10597 30339 10655 30345
rect 10870 30336 10876 30348
rect 10928 30376 10934 30388
rect 11517 30379 11575 30385
rect 11517 30376 11529 30379
rect 10928 30348 11529 30376
rect 10928 30336 10934 30348
rect 11517 30345 11529 30348
rect 11563 30345 11575 30379
rect 11517 30339 11575 30345
rect 11885 30379 11943 30385
rect 11885 30345 11897 30379
rect 11931 30376 11943 30379
rect 12342 30376 12348 30388
rect 11931 30348 12348 30376
rect 11931 30345 11943 30348
rect 11885 30339 11943 30345
rect 5258 30308 5264 30320
rect 5219 30280 5264 30308
rect 5258 30268 5264 30280
rect 5316 30268 5322 30320
rect 5997 30311 6055 30317
rect 5997 30277 6009 30311
rect 6043 30308 6055 30311
rect 7466 30308 7472 30320
rect 6043 30280 7472 30308
rect 6043 30277 6055 30280
rect 5997 30271 6055 30277
rect 7466 30268 7472 30280
rect 7524 30268 7530 30320
rect 9950 30268 9956 30320
rect 10008 30268 10014 30320
rect 5626 30240 5632 30252
rect 5539 30212 5632 30240
rect 5626 30200 5632 30212
rect 5684 30240 5690 30252
rect 7101 30243 7159 30249
rect 5684 30212 6868 30240
rect 5684 30200 5690 30212
rect 6840 30184 6868 30212
rect 7101 30209 7113 30243
rect 7147 30240 7159 30243
rect 7190 30240 7196 30252
rect 7147 30212 7196 30240
rect 7147 30209 7159 30212
rect 7101 30203 7159 30209
rect 7190 30200 7196 30212
rect 7248 30200 7254 30252
rect 7484 30240 7512 30268
rect 7484 30212 7880 30240
rect 4433 30175 4491 30181
rect 4433 30141 4445 30175
rect 4479 30172 4491 30175
rect 4801 30175 4859 30181
rect 4801 30172 4813 30175
rect 4479 30144 4813 30172
rect 4479 30141 4491 30144
rect 4433 30135 4491 30141
rect 4801 30141 4813 30144
rect 4847 30172 4859 30175
rect 5534 30172 5540 30184
rect 4847 30144 5540 30172
rect 4847 30141 4859 30144
rect 4801 30135 4859 30141
rect 5534 30132 5540 30144
rect 5592 30172 5598 30184
rect 6641 30175 6699 30181
rect 6641 30172 6653 30175
rect 5592 30144 6653 30172
rect 5592 30132 5598 30144
rect 6641 30141 6653 30144
rect 6687 30141 6699 30175
rect 6641 30135 6699 30141
rect 6822 30132 6828 30184
rect 6880 30172 6886 30184
rect 7285 30175 7343 30181
rect 7285 30172 7297 30175
rect 6880 30144 7297 30172
rect 6880 30132 6886 30144
rect 7285 30141 7297 30144
rect 7331 30141 7343 30175
rect 7466 30172 7472 30184
rect 7427 30144 7472 30172
rect 7285 30135 7343 30141
rect 7466 30132 7472 30144
rect 7524 30132 7530 30184
rect 7852 30181 7880 30212
rect 8570 30200 8576 30252
rect 8628 30240 8634 30252
rect 10229 30243 10287 30249
rect 10229 30240 10241 30243
rect 8628 30212 10241 30240
rect 8628 30200 8634 30212
rect 10229 30209 10241 30212
rect 10275 30209 10287 30243
rect 10229 30203 10287 30209
rect 10502 30200 10508 30252
rect 10560 30240 10566 30252
rect 10873 30243 10931 30249
rect 10873 30240 10885 30243
rect 10560 30212 10885 30240
rect 10560 30200 10566 30212
rect 10873 30209 10885 30212
rect 10919 30209 10931 30243
rect 11422 30240 11428 30252
rect 10873 30203 10931 30209
rect 11164 30212 11428 30240
rect 7837 30175 7895 30181
rect 7837 30141 7849 30175
rect 7883 30141 7895 30175
rect 7837 30135 7895 30141
rect 7926 30132 7932 30184
rect 7984 30172 7990 30184
rect 9125 30175 9183 30181
rect 7984 30144 8077 30172
rect 7984 30132 7990 30144
rect 9125 30141 9137 30175
rect 9171 30172 9183 30175
rect 9769 30175 9827 30181
rect 9769 30172 9781 30175
rect 9171 30144 9781 30172
rect 9171 30141 9183 30144
rect 9125 30135 9183 30141
rect 9769 30141 9781 30144
rect 9815 30141 9827 30175
rect 10042 30172 10048 30184
rect 10003 30144 10048 30172
rect 9769 30135 9827 30141
rect 6365 30107 6423 30113
rect 6365 30073 6377 30107
rect 6411 30104 6423 30107
rect 7484 30104 7512 30132
rect 6411 30076 7512 30104
rect 6411 30073 6423 30076
rect 6365 30067 6423 30073
rect 7650 30064 7656 30116
rect 7708 30104 7714 30116
rect 7944 30104 7972 30132
rect 7708 30076 7972 30104
rect 9217 30107 9275 30113
rect 7708 30064 7714 30076
rect 9217 30073 9229 30107
rect 9263 30104 9275 30107
rect 9582 30104 9588 30116
rect 9263 30076 9588 30104
rect 9263 30073 9275 30076
rect 9217 30067 9275 30073
rect 9582 30064 9588 30076
rect 9640 30064 9646 30116
rect 9784 30104 9812 30135
rect 10042 30132 10048 30144
rect 10100 30132 10106 30184
rect 11164 30172 11192 30212
rect 11422 30200 11428 30212
rect 11480 30200 11486 30252
rect 10152 30144 11192 30172
rect 11333 30175 11391 30181
rect 10152 30104 10180 30144
rect 11333 30141 11345 30175
rect 11379 30172 11391 30175
rect 11900 30172 11928 30339
rect 12342 30336 12348 30348
rect 12400 30336 12406 30388
rect 12894 30336 12900 30388
rect 12952 30376 12958 30388
rect 15378 30376 15384 30388
rect 12952 30348 15384 30376
rect 12952 30336 12958 30348
rect 15378 30336 15384 30348
rect 15436 30376 15442 30388
rect 16669 30379 16727 30385
rect 16669 30376 16681 30379
rect 15436 30348 16681 30376
rect 15436 30336 15442 30348
rect 16669 30345 16681 30348
rect 16715 30345 16727 30379
rect 16669 30339 16727 30345
rect 18138 30336 18144 30388
rect 18196 30376 18202 30388
rect 18506 30376 18512 30388
rect 18196 30348 18512 30376
rect 18196 30336 18202 30348
rect 18506 30336 18512 30348
rect 18564 30336 18570 30388
rect 20898 30376 20904 30388
rect 20859 30348 20904 30376
rect 20898 30336 20904 30348
rect 20956 30336 20962 30388
rect 14274 30308 14280 30320
rect 14235 30280 14280 30308
rect 14274 30268 14280 30280
rect 14332 30268 14338 30320
rect 14737 30311 14795 30317
rect 14737 30277 14749 30311
rect 14783 30308 14795 30311
rect 15286 30308 15292 30320
rect 14783 30280 15292 30308
rect 14783 30277 14795 30280
rect 14737 30271 14795 30277
rect 15286 30268 15292 30280
rect 15344 30268 15350 30320
rect 16298 30268 16304 30320
rect 16356 30308 16362 30320
rect 17037 30311 17095 30317
rect 17037 30308 17049 30311
rect 16356 30280 17049 30308
rect 16356 30268 16362 30280
rect 17037 30277 17049 30280
rect 17083 30308 17095 30311
rect 17494 30308 17500 30320
rect 17083 30280 17500 30308
rect 17083 30277 17095 30280
rect 17037 30271 17095 30277
rect 17494 30268 17500 30280
rect 17552 30268 17558 30320
rect 18325 30311 18383 30317
rect 18325 30277 18337 30311
rect 18371 30308 18383 30311
rect 19242 30308 19248 30320
rect 18371 30280 19248 30308
rect 18371 30277 18383 30280
rect 18325 30271 18383 30277
rect 19242 30268 19248 30280
rect 19300 30268 19306 30320
rect 20254 30308 20260 30320
rect 20215 30280 20260 30308
rect 20254 30268 20260 30280
rect 20312 30268 20318 30320
rect 12158 30200 12164 30252
rect 12216 30240 12222 30252
rect 12897 30243 12955 30249
rect 12897 30240 12909 30243
rect 12216 30212 12909 30240
rect 12216 30200 12222 30212
rect 12897 30209 12909 30212
rect 12943 30240 12955 30243
rect 13354 30240 13360 30252
rect 12943 30212 13360 30240
rect 12943 30209 12955 30212
rect 12897 30203 12955 30209
rect 13354 30200 13360 30212
rect 13412 30200 13418 30252
rect 13633 30243 13691 30249
rect 13633 30209 13645 30243
rect 13679 30240 13691 30243
rect 13814 30240 13820 30252
rect 13679 30212 13820 30240
rect 13679 30209 13691 30212
rect 13633 30203 13691 30209
rect 13814 30200 13820 30212
rect 13872 30200 13878 30252
rect 13998 30200 14004 30252
rect 14056 30240 14062 30252
rect 14056 30212 15148 30240
rect 14056 30200 14062 30212
rect 15120 30184 15148 30212
rect 17218 30200 17224 30252
rect 17276 30240 17282 30252
rect 17405 30243 17463 30249
rect 17405 30240 17417 30243
rect 17276 30212 17417 30240
rect 17276 30200 17282 30212
rect 17405 30209 17417 30212
rect 17451 30240 17463 30243
rect 17773 30243 17831 30249
rect 17773 30240 17785 30243
rect 17451 30212 17785 30240
rect 17451 30209 17463 30212
rect 17405 30203 17463 30209
rect 17773 30209 17785 30212
rect 17819 30240 17831 30243
rect 18506 30240 18512 30252
rect 17819 30212 18512 30240
rect 17819 30209 17831 30212
rect 17773 30203 17831 30209
rect 18506 30200 18512 30212
rect 18564 30200 18570 30252
rect 19889 30243 19947 30249
rect 19889 30240 19901 30243
rect 19076 30212 19901 30240
rect 19076 30184 19104 30212
rect 19889 30209 19901 30212
rect 19935 30209 19947 30243
rect 19889 30203 19947 30209
rect 14734 30172 14740 30184
rect 11379 30144 11928 30172
rect 14695 30144 14740 30172
rect 11379 30141 11391 30144
rect 11333 30135 11391 30141
rect 14734 30132 14740 30144
rect 14792 30132 14798 30184
rect 14918 30172 14924 30184
rect 14879 30144 14924 30172
rect 14918 30132 14924 30144
rect 14976 30132 14982 30184
rect 15102 30132 15108 30184
rect 15160 30172 15166 30184
rect 15289 30175 15347 30181
rect 15289 30172 15301 30175
rect 15160 30144 15301 30172
rect 15160 30132 15166 30144
rect 15289 30141 15301 30144
rect 15335 30141 15347 30175
rect 15930 30172 15936 30184
rect 15891 30144 15936 30172
rect 15289 30135 15347 30141
rect 15930 30132 15936 30144
rect 15988 30132 15994 30184
rect 16393 30175 16451 30181
rect 16393 30141 16405 30175
rect 16439 30172 16451 30175
rect 16482 30172 16488 30184
rect 16439 30144 16488 30172
rect 16439 30141 16451 30144
rect 16393 30135 16451 30141
rect 16482 30132 16488 30144
rect 16540 30132 16546 30184
rect 17954 30132 17960 30184
rect 18012 30172 18018 30184
rect 18598 30172 18604 30184
rect 18012 30144 18604 30172
rect 18012 30132 18018 30144
rect 18598 30132 18604 30144
rect 18656 30172 18662 30184
rect 18693 30175 18751 30181
rect 18693 30172 18705 30175
rect 18656 30144 18705 30172
rect 18656 30132 18662 30144
rect 18693 30141 18705 30144
rect 18739 30141 18751 30175
rect 19058 30172 19064 30184
rect 19019 30144 19064 30172
rect 18693 30135 18751 30141
rect 9784 30076 10180 30104
rect 11422 30064 11428 30116
rect 11480 30104 11486 30116
rect 13081 30107 13139 30113
rect 13081 30104 13093 30107
rect 11480 30076 13093 30104
rect 11480 30064 11486 30076
rect 13081 30073 13093 30076
rect 13127 30073 13139 30107
rect 13081 30067 13139 30073
rect 13265 30107 13323 30113
rect 13265 30073 13277 30107
rect 13311 30104 13323 30107
rect 13538 30104 13544 30116
rect 13311 30076 13544 30104
rect 13311 30073 13323 30076
rect 13265 30067 13323 30073
rect 13538 30064 13544 30076
rect 13596 30064 13602 30116
rect 13998 30064 14004 30116
rect 14056 30104 14062 30116
rect 14182 30104 14188 30116
rect 14056 30076 14188 30104
rect 14056 30064 14062 30076
rect 14182 30064 14188 30076
rect 14240 30064 14246 30116
rect 14274 30064 14280 30116
rect 14332 30104 14338 30116
rect 16666 30104 16672 30116
rect 14332 30076 16672 30104
rect 14332 30064 14338 30076
rect 16666 30064 16672 30076
rect 16724 30104 16730 30116
rect 18708 30104 18736 30135
rect 19058 30132 19064 30144
rect 19116 30132 19122 30184
rect 19153 30175 19211 30181
rect 19153 30141 19165 30175
rect 19199 30172 19211 30175
rect 20070 30172 20076 30184
rect 19199 30144 19380 30172
rect 20031 30144 20076 30172
rect 19199 30141 19211 30144
rect 19153 30135 19211 30141
rect 18874 30104 18880 30116
rect 16724 30076 18000 30104
rect 18708 30076 18880 30104
rect 16724 30064 16730 30076
rect 17972 30048 18000 30076
rect 18874 30064 18880 30076
rect 18932 30104 18938 30116
rect 19242 30104 19248 30116
rect 18932 30076 19248 30104
rect 18932 30064 18938 30076
rect 19242 30064 19248 30076
rect 19300 30064 19306 30116
rect 19352 30048 19380 30144
rect 20070 30132 20076 30144
rect 20128 30172 20134 30184
rect 20533 30175 20591 30181
rect 20533 30172 20545 30175
rect 20128 30144 20545 30172
rect 20128 30132 20134 30144
rect 20533 30141 20545 30144
rect 20579 30141 20591 30175
rect 20533 30135 20591 30141
rect 19426 30064 19432 30116
rect 19484 30104 19490 30116
rect 21269 30107 21327 30113
rect 21269 30104 21281 30107
rect 19484 30076 21281 30104
rect 19484 30064 19490 30076
rect 21269 30073 21281 30076
rect 21315 30104 21327 30107
rect 21634 30104 21640 30116
rect 21315 30076 21640 30104
rect 21315 30073 21327 30076
rect 21269 30067 21327 30073
rect 21634 30064 21640 30076
rect 21692 30064 21698 30116
rect 4249 30039 4307 30045
rect 4249 30005 4261 30039
rect 4295 30036 4307 30039
rect 4614 30036 4620 30048
rect 4295 30008 4620 30036
rect 4295 30005 4307 30008
rect 4249 29999 4307 30005
rect 4614 29996 4620 30008
rect 4672 29996 4678 30048
rect 6457 30039 6515 30045
rect 6457 30005 6469 30039
rect 6503 30036 6515 30039
rect 6638 30036 6644 30048
rect 6503 30008 6644 30036
rect 6503 30005 6515 30008
rect 6457 29999 6515 30005
rect 6638 29996 6644 30008
rect 6696 30036 6702 30048
rect 6914 30036 6920 30048
rect 6696 30008 6920 30036
rect 6696 29996 6702 30008
rect 6914 29996 6920 30008
rect 6972 29996 6978 30048
rect 8294 29996 8300 30048
rect 8352 30036 8358 30048
rect 8846 30036 8852 30048
rect 8352 30008 8852 30036
rect 8352 29996 8358 30008
rect 8846 29996 8852 30008
rect 8904 29996 8910 30048
rect 10134 29996 10140 30048
rect 10192 30036 10198 30048
rect 12161 30039 12219 30045
rect 12161 30036 12173 30039
rect 10192 30008 12173 30036
rect 10192 29996 10198 30008
rect 12161 30005 12173 30008
rect 12207 30036 12219 30039
rect 12250 30036 12256 30048
rect 12207 30008 12256 30036
rect 12207 30005 12219 30008
rect 12161 29999 12219 30005
rect 12250 29996 12256 30008
rect 12308 29996 12314 30048
rect 12434 29996 12440 30048
rect 12492 30036 12498 30048
rect 12805 30039 12863 30045
rect 12805 30036 12817 30039
rect 12492 30008 12817 30036
rect 12492 29996 12498 30008
rect 12805 30005 12817 30008
rect 12851 30036 12863 30039
rect 13173 30039 13231 30045
rect 13173 30036 13185 30039
rect 12851 30008 13185 30036
rect 12851 30005 12863 30008
rect 12805 29999 12863 30005
rect 13173 30005 13185 30008
rect 13219 30036 13231 30039
rect 15010 30036 15016 30048
rect 13219 30008 15016 30036
rect 13219 30005 13231 30008
rect 13173 29999 13231 30005
rect 15010 29996 15016 30008
rect 15068 29996 15074 30048
rect 15378 29996 15384 30048
rect 15436 30036 15442 30048
rect 17494 30036 17500 30048
rect 15436 30008 17500 30036
rect 15436 29996 15442 30008
rect 17494 29996 17500 30008
rect 17552 29996 17558 30048
rect 17954 29996 17960 30048
rect 18012 29996 18018 30048
rect 19334 29996 19340 30048
rect 19392 30036 19398 30048
rect 19521 30039 19579 30045
rect 19521 30036 19533 30039
rect 19392 30008 19533 30036
rect 19392 29996 19398 30008
rect 19521 30005 19533 30008
rect 19567 30036 19579 30039
rect 19610 30036 19616 30048
rect 19567 30008 19616 30036
rect 19567 30005 19579 30008
rect 19521 29999 19579 30005
rect 19610 29996 19616 30008
rect 19668 29996 19674 30048
rect 1104 29946 28888 29968
rect 1104 29894 10982 29946
rect 11034 29894 11046 29946
rect 11098 29894 11110 29946
rect 11162 29894 11174 29946
rect 11226 29894 20982 29946
rect 21034 29894 21046 29946
rect 21098 29894 21110 29946
rect 21162 29894 21174 29946
rect 21226 29894 28888 29946
rect 1104 29872 28888 29894
rect 6546 29832 6552 29844
rect 6507 29804 6552 29832
rect 6546 29792 6552 29804
rect 6604 29792 6610 29844
rect 8294 29832 8300 29844
rect 8255 29804 8300 29832
rect 8294 29792 8300 29804
rect 8352 29792 8358 29844
rect 8570 29792 8576 29844
rect 8628 29832 8634 29844
rect 9033 29835 9091 29841
rect 9033 29832 9045 29835
rect 8628 29804 9045 29832
rect 8628 29792 8634 29804
rect 9033 29801 9045 29804
rect 9079 29801 9091 29835
rect 9033 29795 9091 29801
rect 9306 29792 9312 29844
rect 9364 29832 9370 29844
rect 9401 29835 9459 29841
rect 9401 29832 9413 29835
rect 9364 29804 9413 29832
rect 9364 29792 9370 29804
rect 9401 29801 9413 29804
rect 9447 29801 9459 29835
rect 9401 29795 9459 29801
rect 11790 29792 11796 29844
rect 11848 29832 11854 29844
rect 11848 29804 13124 29832
rect 11848 29792 11854 29804
rect 6181 29767 6239 29773
rect 6181 29733 6193 29767
rect 6227 29764 6239 29767
rect 6822 29764 6828 29776
rect 6227 29736 6828 29764
rect 6227 29733 6239 29736
rect 6181 29727 6239 29733
rect 6822 29724 6828 29736
rect 6880 29724 6886 29776
rect 6917 29767 6975 29773
rect 6917 29733 6929 29767
rect 6963 29764 6975 29767
rect 7650 29764 7656 29776
rect 6963 29736 7656 29764
rect 6963 29733 6975 29736
rect 6917 29727 6975 29733
rect 7650 29724 7656 29736
rect 7708 29724 7714 29776
rect 7929 29767 7987 29773
rect 7929 29733 7941 29767
rect 7975 29764 7987 29767
rect 10042 29764 10048 29776
rect 7975 29736 10048 29764
rect 7975 29733 7987 29736
rect 7929 29727 7987 29733
rect 10042 29724 10048 29736
rect 10100 29724 10106 29776
rect 12342 29764 12348 29776
rect 12303 29736 12348 29764
rect 12342 29724 12348 29736
rect 12400 29724 12406 29776
rect 12437 29767 12495 29773
rect 12437 29733 12449 29767
rect 12483 29764 12495 29767
rect 12894 29764 12900 29776
rect 12483 29736 12900 29764
rect 12483 29733 12495 29736
rect 12437 29727 12495 29733
rect 12894 29724 12900 29736
rect 12952 29724 12958 29776
rect 13096 29764 13124 29804
rect 13170 29792 13176 29844
rect 13228 29832 13234 29844
rect 13354 29832 13360 29844
rect 13228 29804 13360 29832
rect 13228 29792 13234 29804
rect 13354 29792 13360 29804
rect 13412 29832 13418 29844
rect 13449 29835 13507 29841
rect 13449 29832 13461 29835
rect 13412 29804 13461 29832
rect 13412 29792 13418 29804
rect 13449 29801 13461 29804
rect 13495 29801 13507 29835
rect 13449 29795 13507 29801
rect 15010 29792 15016 29844
rect 15068 29832 15074 29844
rect 15746 29832 15752 29844
rect 15068 29804 15752 29832
rect 15068 29792 15074 29804
rect 15746 29792 15752 29804
rect 15804 29792 15810 29844
rect 16393 29835 16451 29841
rect 16393 29801 16405 29835
rect 16439 29832 16451 29835
rect 16439 29804 17264 29832
rect 16439 29801 16451 29804
rect 16393 29795 16451 29801
rect 14642 29764 14648 29776
rect 13096 29736 14648 29764
rect 14642 29724 14648 29736
rect 14700 29724 14706 29776
rect 15102 29764 15108 29776
rect 15063 29736 15108 29764
rect 15102 29724 15108 29736
rect 15160 29724 15166 29776
rect 15378 29764 15384 29776
rect 15212 29736 15384 29764
rect 7009 29699 7067 29705
rect 7009 29665 7021 29699
rect 7055 29696 7067 29699
rect 7098 29696 7104 29708
rect 7055 29668 7104 29696
rect 7055 29665 7067 29668
rect 7009 29659 7067 29665
rect 7098 29656 7104 29668
rect 7156 29656 7162 29708
rect 8110 29696 8116 29708
rect 8071 29668 8116 29696
rect 8110 29656 8116 29668
rect 8168 29656 8174 29708
rect 9214 29696 9220 29708
rect 8220 29668 9220 29696
rect 5445 29631 5503 29637
rect 5445 29597 5457 29631
rect 5491 29628 5503 29631
rect 6914 29628 6920 29640
rect 5491 29600 6920 29628
rect 5491 29597 5503 29600
rect 5445 29591 5503 29597
rect 6914 29588 6920 29600
rect 6972 29588 6978 29640
rect 7561 29631 7619 29637
rect 7561 29597 7573 29631
rect 7607 29628 7619 29631
rect 8220 29628 8248 29668
rect 9214 29656 9220 29668
rect 9272 29696 9278 29708
rect 10505 29699 10563 29705
rect 10505 29696 10517 29699
rect 9272 29668 10517 29696
rect 9272 29656 9278 29668
rect 10505 29665 10517 29668
rect 10551 29665 10563 29699
rect 12253 29699 12311 29705
rect 12253 29696 12265 29699
rect 10505 29659 10563 29665
rect 11532 29668 12265 29696
rect 7607 29600 8248 29628
rect 9677 29631 9735 29637
rect 7607 29597 7619 29600
rect 7561 29591 7619 29597
rect 9677 29597 9689 29631
rect 9723 29628 9735 29631
rect 9858 29628 9864 29640
rect 9723 29600 9864 29628
rect 9723 29597 9735 29600
rect 9677 29591 9735 29597
rect 9858 29588 9864 29600
rect 9916 29588 9922 29640
rect 10134 29588 10140 29640
rect 10192 29628 10198 29640
rect 10229 29631 10287 29637
rect 10229 29628 10241 29631
rect 10192 29600 10241 29628
rect 10192 29588 10198 29600
rect 10229 29597 10241 29600
rect 10275 29597 10287 29631
rect 10229 29591 10287 29597
rect 10410 29588 10416 29640
rect 10468 29628 10474 29640
rect 10689 29631 10747 29637
rect 10689 29628 10701 29631
rect 10468 29600 10701 29628
rect 10468 29588 10474 29600
rect 10689 29597 10701 29600
rect 10735 29597 10747 29631
rect 10689 29591 10747 29597
rect 7193 29563 7251 29569
rect 7193 29529 7205 29563
rect 7239 29560 7251 29563
rect 11422 29560 11428 29572
rect 7239 29532 11428 29560
rect 7239 29529 7251 29532
rect 7193 29523 7251 29529
rect 11422 29520 11428 29532
rect 11480 29560 11486 29572
rect 11532 29569 11560 29668
rect 12253 29665 12265 29668
rect 12299 29696 12311 29699
rect 13262 29696 13268 29708
rect 12299 29668 13268 29696
rect 12299 29665 12311 29668
rect 12253 29659 12311 29665
rect 13262 29656 13268 29668
rect 13320 29656 13326 29708
rect 13630 29696 13636 29708
rect 13591 29668 13636 29696
rect 13630 29656 13636 29668
rect 13688 29656 13694 29708
rect 13814 29705 13820 29708
rect 13780 29699 13820 29705
rect 13780 29665 13792 29699
rect 13780 29659 13820 29665
rect 13814 29656 13820 29659
rect 13872 29656 13878 29708
rect 15212 29696 15240 29736
rect 15378 29724 15384 29736
rect 15436 29724 15442 29776
rect 16206 29724 16212 29776
rect 16264 29764 16270 29776
rect 17037 29767 17095 29773
rect 17037 29764 17049 29767
rect 16264 29736 17049 29764
rect 16264 29724 16270 29736
rect 17037 29733 17049 29736
rect 17083 29733 17095 29767
rect 17037 29727 17095 29733
rect 14016 29668 15240 29696
rect 15289 29699 15347 29705
rect 12069 29631 12127 29637
rect 12069 29597 12081 29631
rect 12115 29628 12127 29631
rect 12710 29628 12716 29640
rect 12115 29600 12716 29628
rect 12115 29597 12127 29600
rect 12069 29591 12127 29597
rect 12710 29588 12716 29600
rect 12768 29588 12774 29640
rect 14016 29637 14044 29668
rect 15289 29665 15301 29699
rect 15335 29696 15347 29699
rect 16482 29696 16488 29708
rect 15335 29668 16488 29696
rect 15335 29665 15347 29668
rect 15289 29659 15347 29665
rect 16482 29656 16488 29668
rect 16540 29656 16546 29708
rect 16574 29656 16580 29708
rect 16632 29696 16638 29708
rect 16850 29696 16856 29708
rect 16632 29668 16856 29696
rect 16632 29656 16638 29668
rect 16850 29656 16856 29668
rect 16908 29656 16914 29708
rect 17129 29699 17187 29705
rect 17129 29665 17141 29699
rect 17175 29665 17187 29699
rect 17236 29696 17264 29804
rect 17494 29792 17500 29844
rect 17552 29832 17558 29844
rect 17865 29835 17923 29841
rect 17865 29832 17877 29835
rect 17552 29804 17877 29832
rect 17552 29792 17558 29804
rect 17865 29801 17877 29804
rect 17911 29801 17923 29835
rect 17865 29795 17923 29801
rect 18046 29792 18052 29844
rect 18104 29832 18110 29844
rect 19889 29835 19947 29841
rect 18104 29804 19196 29832
rect 18104 29792 18110 29804
rect 17589 29767 17647 29773
rect 17589 29733 17601 29767
rect 17635 29764 17647 29767
rect 17770 29764 17776 29776
rect 17635 29736 17776 29764
rect 17635 29733 17647 29736
rect 17589 29727 17647 29733
rect 17770 29724 17776 29736
rect 17828 29724 17834 29776
rect 18693 29767 18751 29773
rect 18693 29733 18705 29767
rect 18739 29764 18751 29767
rect 18874 29764 18880 29776
rect 18739 29736 18880 29764
rect 18739 29733 18751 29736
rect 18693 29727 18751 29733
rect 18874 29724 18880 29736
rect 18932 29724 18938 29776
rect 19168 29773 19196 29804
rect 19889 29801 19901 29835
rect 19935 29832 19947 29835
rect 20070 29832 20076 29844
rect 19935 29804 20076 29832
rect 19935 29801 19947 29804
rect 19889 29795 19947 29801
rect 20070 29792 20076 29804
rect 20128 29832 20134 29844
rect 20441 29835 20499 29841
rect 20441 29832 20453 29835
rect 20128 29804 20453 29832
rect 20128 29792 20134 29804
rect 20441 29801 20453 29804
rect 20487 29801 20499 29835
rect 20441 29795 20499 29801
rect 21637 29835 21695 29841
rect 21637 29801 21649 29835
rect 21683 29832 21695 29835
rect 21910 29832 21916 29844
rect 21683 29804 21916 29832
rect 21683 29801 21695 29804
rect 21637 29795 21695 29801
rect 21910 29792 21916 29804
rect 21968 29792 21974 29844
rect 19153 29767 19211 29773
rect 19153 29733 19165 29767
rect 19199 29733 19211 29767
rect 21177 29767 21235 29773
rect 21177 29764 21189 29767
rect 19153 29727 19211 29733
rect 20088 29736 21189 29764
rect 18601 29699 18659 29705
rect 17236 29668 17816 29696
rect 17129 29659 17187 29665
rect 12805 29631 12863 29637
rect 12805 29597 12817 29631
rect 12851 29628 12863 29631
rect 14001 29631 14059 29637
rect 14001 29628 14013 29631
rect 12851 29600 14013 29628
rect 12851 29597 12863 29600
rect 12805 29591 12863 29597
rect 14001 29597 14013 29600
rect 14047 29597 14059 29631
rect 14001 29591 14059 29597
rect 14182 29588 14188 29640
rect 14240 29628 14246 29640
rect 14645 29631 14703 29637
rect 14645 29628 14657 29631
rect 14240 29600 14657 29628
rect 14240 29588 14246 29600
rect 14645 29597 14657 29600
rect 14691 29628 14703 29631
rect 14918 29628 14924 29640
rect 14691 29600 14924 29628
rect 14691 29597 14703 29600
rect 14645 29591 14703 29597
rect 14918 29588 14924 29600
rect 14976 29588 14982 29640
rect 15657 29631 15715 29637
rect 15657 29597 15669 29631
rect 15703 29628 15715 29631
rect 16298 29628 16304 29640
rect 15703 29600 16304 29628
rect 15703 29597 15715 29600
rect 15657 29591 15715 29597
rect 16298 29588 16304 29600
rect 16356 29588 16362 29640
rect 16666 29588 16672 29640
rect 16724 29628 16730 29640
rect 17144 29628 17172 29659
rect 17788 29640 17816 29668
rect 18601 29665 18613 29699
rect 18647 29665 18659 29699
rect 18601 29659 18659 29665
rect 18769 29699 18827 29705
rect 18769 29665 18781 29699
rect 18815 29696 18827 29699
rect 19058 29696 19064 29708
rect 18815 29668 19064 29696
rect 18815 29665 18827 29668
rect 18769 29659 18827 29665
rect 16724 29600 17172 29628
rect 16724 29588 16730 29600
rect 17770 29588 17776 29640
rect 17828 29588 17834 29640
rect 18417 29631 18475 29637
rect 18417 29597 18429 29631
rect 18463 29597 18475 29631
rect 18417 29591 18475 29597
rect 11517 29563 11575 29569
rect 11517 29560 11529 29563
rect 11480 29532 11529 29560
rect 11480 29520 11486 29532
rect 11517 29529 11529 29532
rect 11563 29529 11575 29563
rect 12728 29560 12756 29588
rect 13081 29563 13139 29569
rect 13081 29560 13093 29563
rect 12728 29532 13093 29560
rect 11517 29523 11575 29529
rect 13081 29529 13093 29532
rect 13127 29560 13139 29563
rect 13354 29560 13360 29572
rect 13127 29532 13360 29560
rect 13127 29529 13139 29532
rect 13081 29523 13139 29529
rect 13354 29520 13360 29532
rect 13412 29520 13418 29572
rect 13538 29520 13544 29572
rect 13596 29560 13602 29572
rect 15565 29563 15623 29569
rect 15565 29560 15577 29563
rect 13596 29532 15577 29560
rect 13596 29520 13602 29532
rect 15565 29529 15577 29532
rect 15611 29560 15623 29563
rect 15611 29532 16712 29560
rect 15611 29529 15623 29532
rect 15565 29523 15623 29529
rect 5813 29495 5871 29501
rect 5813 29461 5825 29495
rect 5859 29492 5871 29495
rect 6546 29492 6552 29504
rect 5859 29464 6552 29492
rect 5859 29461 5871 29464
rect 5813 29455 5871 29461
rect 6546 29452 6552 29464
rect 6604 29452 6610 29504
rect 9306 29452 9312 29504
rect 9364 29492 9370 29504
rect 9674 29492 9680 29504
rect 9364 29464 9680 29492
rect 9364 29452 9370 29464
rect 9674 29452 9680 29464
rect 9732 29452 9738 29504
rect 11054 29492 11060 29504
rect 11015 29464 11060 29492
rect 11054 29452 11060 29464
rect 11112 29452 11118 29504
rect 11977 29495 12035 29501
rect 11977 29461 11989 29495
rect 12023 29492 12035 29495
rect 12250 29492 12256 29504
rect 12023 29464 12256 29492
rect 12023 29461 12035 29464
rect 11977 29455 12035 29461
rect 12250 29452 12256 29464
rect 12308 29492 12314 29504
rect 12526 29492 12532 29504
rect 12308 29464 12532 29492
rect 12308 29452 12314 29464
rect 12526 29452 12532 29464
rect 12584 29452 12590 29504
rect 13906 29492 13912 29504
rect 13867 29464 13912 29492
rect 13906 29452 13912 29464
rect 13964 29452 13970 29504
rect 14274 29492 14280 29504
rect 14235 29464 14280 29492
rect 14274 29452 14280 29464
rect 14332 29452 14338 29504
rect 15378 29452 15384 29504
rect 15436 29501 15442 29504
rect 15436 29495 15485 29501
rect 15436 29461 15439 29495
rect 15473 29461 15485 29495
rect 15746 29492 15752 29504
rect 15707 29464 15752 29492
rect 15436 29455 15485 29461
rect 15436 29452 15442 29455
rect 15746 29452 15752 29464
rect 15804 29452 15810 29504
rect 16684 29501 16712 29532
rect 16758 29520 16764 29572
rect 16816 29560 16822 29572
rect 18233 29563 18291 29569
rect 18233 29560 18245 29563
rect 16816 29532 18245 29560
rect 16816 29520 16822 29532
rect 18233 29529 18245 29532
rect 18279 29529 18291 29563
rect 18233 29523 18291 29529
rect 16669 29495 16727 29501
rect 16669 29461 16681 29495
rect 16715 29461 16727 29495
rect 18432 29492 18460 29591
rect 18616 29560 18644 29659
rect 19058 29656 19064 29668
rect 19116 29656 19122 29708
rect 19521 29699 19579 29705
rect 19521 29665 19533 29699
rect 19567 29696 19579 29699
rect 19886 29696 19892 29708
rect 19567 29668 19892 29696
rect 19567 29665 19579 29668
rect 19521 29659 19579 29665
rect 19886 29656 19892 29668
rect 19944 29656 19950 29708
rect 19150 29588 19156 29640
rect 19208 29628 19214 29640
rect 20088 29628 20116 29736
rect 21177 29733 21189 29736
rect 21223 29764 21235 29767
rect 22186 29764 22192 29776
rect 21223 29736 22192 29764
rect 21223 29733 21235 29736
rect 21177 29727 21235 29733
rect 22186 29724 22192 29736
rect 22244 29724 22250 29776
rect 20165 29699 20223 29705
rect 20165 29665 20177 29699
rect 20211 29696 20223 29699
rect 20346 29696 20352 29708
rect 20211 29668 20352 29696
rect 20211 29665 20223 29668
rect 20165 29659 20223 29665
rect 20346 29656 20352 29668
rect 20404 29696 20410 29708
rect 21818 29696 21824 29708
rect 20404 29668 21824 29696
rect 20404 29656 20410 29668
rect 21818 29656 21824 29668
rect 21876 29656 21882 29708
rect 19208 29600 20116 29628
rect 19208 29588 19214 29600
rect 19981 29563 20039 29569
rect 18616 29532 19932 29560
rect 19352 29504 19380 29532
rect 18874 29492 18880 29504
rect 18432 29464 18880 29492
rect 16669 29455 16727 29461
rect 18874 29452 18880 29464
rect 18932 29452 18938 29504
rect 19334 29452 19340 29504
rect 19392 29452 19398 29504
rect 19904 29492 19932 29532
rect 19981 29529 19993 29563
rect 20027 29560 20039 29563
rect 20088 29560 20116 29600
rect 20027 29532 20116 29560
rect 20027 29529 20039 29532
rect 19981 29523 20039 29529
rect 22370 29492 22376 29504
rect 19904 29464 22376 29492
rect 22370 29452 22376 29464
rect 22428 29452 22434 29504
rect 1104 29402 28888 29424
rect 1104 29350 5982 29402
rect 6034 29350 6046 29402
rect 6098 29350 6110 29402
rect 6162 29350 6174 29402
rect 6226 29350 15982 29402
rect 16034 29350 16046 29402
rect 16098 29350 16110 29402
rect 16162 29350 16174 29402
rect 16226 29350 25982 29402
rect 26034 29350 26046 29402
rect 26098 29350 26110 29402
rect 26162 29350 26174 29402
rect 26226 29350 28888 29402
rect 1104 29328 28888 29350
rect 6638 29288 6644 29300
rect 6599 29260 6644 29288
rect 6638 29248 6644 29260
rect 6696 29248 6702 29300
rect 7098 29288 7104 29300
rect 7059 29260 7104 29288
rect 7098 29248 7104 29260
rect 7156 29248 7162 29300
rect 9122 29288 9128 29300
rect 9083 29260 9128 29288
rect 9122 29248 9128 29260
rect 9180 29248 9186 29300
rect 11422 29288 11428 29300
rect 11383 29260 11428 29288
rect 11422 29248 11428 29260
rect 11480 29288 11486 29300
rect 11701 29291 11759 29297
rect 11701 29288 11713 29291
rect 11480 29260 11713 29288
rect 11480 29248 11486 29260
rect 11701 29257 11713 29260
rect 11747 29257 11759 29291
rect 11701 29251 11759 29257
rect 12342 29248 12348 29300
rect 12400 29288 12406 29300
rect 12621 29291 12679 29297
rect 12621 29288 12633 29291
rect 12400 29260 12633 29288
rect 12400 29248 12406 29260
rect 12621 29257 12633 29260
rect 12667 29257 12679 29291
rect 14645 29291 14703 29297
rect 12621 29251 12679 29257
rect 13004 29260 13584 29288
rect 9306 29180 9312 29232
rect 9364 29220 9370 29232
rect 9401 29223 9459 29229
rect 9401 29220 9413 29223
rect 9364 29192 9413 29220
rect 9364 29180 9370 29192
rect 9401 29189 9413 29192
rect 9447 29189 9459 29223
rect 9401 29183 9459 29189
rect 9677 29223 9735 29229
rect 9677 29189 9689 29223
rect 9723 29220 9735 29223
rect 10502 29220 10508 29232
rect 9723 29192 10508 29220
rect 9723 29189 9735 29192
rect 9677 29183 9735 29189
rect 10502 29180 10508 29192
rect 10560 29180 10566 29232
rect 12161 29223 12219 29229
rect 12161 29189 12173 29223
rect 12207 29220 12219 29223
rect 12710 29220 12716 29232
rect 12207 29192 12716 29220
rect 12207 29189 12219 29192
rect 12161 29183 12219 29189
rect 12452 29164 12480 29192
rect 12710 29180 12716 29192
rect 12768 29180 12774 29232
rect 7745 29155 7803 29161
rect 7745 29121 7757 29155
rect 7791 29152 7803 29155
rect 8757 29155 8815 29161
rect 8757 29152 8769 29155
rect 7791 29124 8769 29152
rect 7791 29121 7803 29124
rect 7745 29115 7803 29121
rect 8757 29121 8769 29124
rect 8803 29152 8815 29155
rect 10410 29152 10416 29164
rect 8803 29124 10416 29152
rect 8803 29121 8815 29124
rect 8757 29115 8815 29121
rect 10410 29112 10416 29124
rect 10468 29112 10474 29164
rect 11054 29112 11060 29164
rect 11112 29152 11118 29164
rect 11422 29152 11428 29164
rect 11112 29124 11428 29152
rect 11112 29112 11118 29124
rect 11422 29112 11428 29124
rect 11480 29112 11486 29164
rect 12434 29112 12440 29164
rect 12492 29112 12498 29164
rect 13004 29152 13032 29260
rect 12636 29124 13032 29152
rect 13081 29155 13139 29161
rect 5537 29087 5595 29093
rect 5537 29053 5549 29087
rect 5583 29084 5595 29087
rect 6178 29084 6184 29096
rect 5583 29056 6184 29084
rect 5583 29053 5595 29056
rect 5537 29047 5595 29053
rect 6178 29044 6184 29056
rect 6236 29044 6242 29096
rect 6273 29087 6331 29093
rect 6273 29053 6285 29087
rect 6319 29084 6331 29087
rect 6822 29084 6828 29096
rect 6319 29056 6828 29084
rect 6319 29053 6331 29056
rect 6273 29047 6331 29053
rect 6822 29044 6828 29056
rect 6880 29084 6886 29096
rect 8202 29084 8208 29096
rect 6880 29056 8208 29084
rect 6880 29044 6886 29056
rect 8202 29044 8208 29056
rect 8260 29044 8266 29096
rect 8297 29087 8355 29093
rect 8297 29053 8309 29087
rect 8343 29084 8355 29087
rect 9122 29084 9128 29096
rect 8343 29056 9128 29084
rect 8343 29053 8355 29056
rect 8297 29047 8355 29053
rect 8680 29028 8708 29056
rect 9122 29044 9128 29056
rect 9180 29044 9186 29096
rect 9398 29044 9404 29096
rect 9456 29084 9462 29096
rect 10229 29087 10287 29093
rect 10229 29084 10241 29087
rect 9456 29056 10241 29084
rect 9456 29044 9462 29056
rect 10229 29053 10241 29056
rect 10275 29053 10287 29087
rect 10229 29047 10287 29053
rect 10321 29087 10379 29093
rect 10321 29053 10333 29087
rect 10367 29053 10379 29087
rect 10321 29047 10379 29053
rect 10597 29087 10655 29093
rect 10597 29053 10609 29087
rect 10643 29084 10655 29087
rect 10686 29084 10692 29096
rect 10643 29056 10692 29084
rect 10643 29053 10655 29056
rect 10597 29047 10655 29053
rect 1394 28976 1400 29028
rect 1452 29016 1458 29028
rect 1946 29016 1952 29028
rect 1452 28988 1952 29016
rect 1452 28976 1458 28988
rect 1946 28976 1952 28988
rect 2004 29016 2010 29028
rect 4614 29016 4620 29028
rect 2004 28988 4620 29016
rect 2004 28976 2010 28988
rect 4614 28976 4620 28988
rect 4672 28976 4678 29028
rect 5442 28976 5448 29028
rect 5500 29016 5506 29028
rect 5810 29016 5816 29028
rect 5500 28988 5816 29016
rect 5500 28976 5506 28988
rect 5810 28976 5816 28988
rect 5868 28976 5874 29028
rect 8110 29016 8116 29028
rect 8071 28988 8116 29016
rect 8110 28976 8116 28988
rect 8168 28976 8174 29028
rect 8662 28976 8668 29028
rect 8720 28976 8726 29028
rect 9306 28976 9312 29028
rect 9364 29016 9370 29028
rect 10336 29016 10364 29047
rect 9364 28988 10364 29016
rect 9364 28976 9370 28988
rect 8938 28908 8944 28960
rect 8996 28948 9002 28960
rect 9490 28948 9496 28960
rect 8996 28920 9496 28948
rect 8996 28908 9002 28920
rect 9490 28908 9496 28920
rect 9548 28908 9554 28960
rect 9766 28908 9772 28960
rect 9824 28948 9830 28960
rect 10612 28948 10640 29047
rect 10686 29044 10692 29056
rect 10744 29044 10750 29096
rect 10781 29087 10839 29093
rect 10781 29053 10793 29087
rect 10827 29084 10839 29087
rect 10870 29084 10876 29096
rect 10827 29056 10876 29084
rect 10827 29053 10839 29056
rect 10781 29047 10839 29053
rect 10870 29044 10876 29056
rect 10928 29044 10934 29096
rect 12636 29028 12664 29124
rect 13081 29121 13093 29155
rect 13127 29152 13139 29155
rect 13127 29124 13492 29152
rect 13127 29121 13139 29124
rect 13081 29115 13139 29121
rect 13170 29084 13176 29096
rect 13131 29056 13176 29084
rect 13170 29044 13176 29056
rect 13228 29044 13234 29096
rect 12618 29016 12624 29028
rect 12268 28988 12624 29016
rect 9824 28920 10640 28948
rect 9824 28908 9830 28920
rect 10870 28908 10876 28960
rect 10928 28948 10934 28960
rect 12268 28948 12296 28988
rect 12618 28976 12624 28988
rect 12676 28976 12682 29028
rect 13372 29016 13400 29124
rect 13464 29093 13492 29124
rect 13449 29087 13507 29093
rect 13449 29053 13461 29087
rect 13495 29053 13507 29087
rect 13556 29084 13584 29260
rect 14645 29257 14657 29291
rect 14691 29288 14703 29291
rect 15102 29288 15108 29300
rect 14691 29260 15108 29288
rect 14691 29257 14703 29260
rect 14645 29251 14703 29257
rect 15102 29248 15108 29260
rect 15160 29248 15166 29300
rect 15286 29248 15292 29300
rect 15344 29288 15350 29300
rect 15749 29291 15807 29297
rect 15749 29288 15761 29291
rect 15344 29260 15761 29288
rect 15344 29248 15350 29260
rect 15749 29257 15761 29260
rect 15795 29257 15807 29291
rect 15749 29251 15807 29257
rect 16390 29248 16396 29300
rect 16448 29297 16454 29300
rect 16448 29291 16497 29297
rect 16448 29257 16451 29291
rect 16485 29257 16497 29291
rect 16448 29251 16497 29257
rect 16577 29291 16635 29297
rect 16577 29257 16589 29291
rect 16623 29288 16635 29291
rect 16758 29288 16764 29300
rect 16623 29260 16764 29288
rect 16623 29257 16635 29260
rect 16577 29251 16635 29257
rect 16448 29248 16454 29251
rect 16758 29248 16764 29260
rect 16816 29248 16822 29300
rect 16850 29248 16856 29300
rect 16908 29288 16914 29300
rect 17313 29291 17371 29297
rect 17313 29288 17325 29291
rect 16908 29260 17325 29288
rect 16908 29248 16914 29260
rect 17313 29257 17325 29260
rect 17359 29257 17371 29291
rect 17313 29251 17371 29257
rect 18046 29248 18052 29300
rect 18104 29288 18110 29300
rect 18325 29291 18383 29297
rect 18325 29288 18337 29291
rect 18104 29260 18337 29288
rect 18104 29248 18110 29260
rect 18325 29257 18337 29260
rect 18371 29257 18383 29291
rect 18325 29251 18383 29257
rect 18506 29248 18512 29300
rect 18564 29288 18570 29300
rect 19613 29291 19671 29297
rect 19613 29288 19625 29291
rect 18564 29260 19625 29288
rect 18564 29248 18570 29260
rect 19613 29257 19625 29260
rect 19659 29257 19671 29291
rect 19886 29288 19892 29300
rect 19847 29260 19892 29288
rect 19613 29251 19671 29257
rect 19886 29248 19892 29260
rect 19944 29248 19950 29300
rect 20990 29288 20996 29300
rect 20951 29260 20996 29288
rect 20990 29248 20996 29260
rect 21048 29248 21054 29300
rect 21729 29291 21787 29297
rect 21729 29257 21741 29291
rect 21775 29288 21787 29291
rect 21818 29288 21824 29300
rect 21775 29260 21824 29288
rect 21775 29257 21787 29260
rect 21729 29251 21787 29257
rect 21818 29248 21824 29260
rect 21876 29248 21882 29300
rect 13906 29180 13912 29232
rect 13964 29220 13970 29232
rect 17218 29220 17224 29232
rect 13964 29192 15516 29220
rect 13964 29180 13970 29192
rect 14844 29164 14872 29192
rect 13630 29112 13636 29164
rect 13688 29152 13694 29164
rect 13688 29124 13768 29152
rect 13688 29112 13694 29124
rect 13556 29056 13676 29084
rect 13449 29047 13507 29053
rect 13533 29019 13591 29025
rect 13372 28988 13492 29016
rect 10928 28920 12296 28948
rect 10928 28908 10934 28920
rect 13262 28908 13268 28960
rect 13320 28948 13326 28960
rect 13357 28951 13415 28957
rect 13357 28948 13369 28951
rect 13320 28920 13369 28948
rect 13320 28908 13326 28920
rect 13357 28917 13369 28920
rect 13403 28917 13415 28951
rect 13464 28948 13492 28988
rect 13533 28985 13545 29019
rect 13579 29016 13591 29019
rect 13648 29016 13676 29056
rect 13579 28988 13676 29016
rect 13740 29016 13768 29124
rect 14826 29112 14832 29164
rect 14884 29112 14890 29164
rect 15102 29112 15108 29164
rect 15160 29112 15166 29164
rect 15488 29161 15516 29192
rect 15672 29192 17224 29220
rect 15473 29155 15531 29161
rect 15473 29121 15485 29155
rect 15519 29121 15531 29155
rect 15473 29115 15531 29121
rect 13814 29044 13820 29096
rect 13872 29084 13878 29096
rect 14277 29087 14335 29093
rect 13872 29056 14228 29084
rect 13872 29044 13878 29056
rect 13909 29019 13967 29025
rect 13909 29016 13921 29019
rect 13740 28988 13921 29016
rect 13579 28985 13591 28988
rect 13533 28979 13591 28985
rect 13909 28985 13921 28988
rect 13955 28985 13967 29019
rect 13909 28979 13967 28985
rect 13814 28948 13820 28960
rect 13464 28920 13820 28948
rect 13357 28911 13415 28917
rect 13814 28908 13820 28920
rect 13872 28908 13878 28960
rect 14200 28948 14228 29056
rect 14277 29053 14289 29087
rect 14323 29084 14335 29087
rect 14642 29084 14648 29096
rect 14323 29056 14648 29084
rect 14323 29053 14335 29056
rect 14277 29047 14335 29053
rect 14642 29044 14648 29056
rect 14700 29084 14706 29096
rect 14918 29084 14924 29096
rect 14700 29056 14924 29084
rect 14700 29044 14706 29056
rect 14918 29044 14924 29056
rect 14976 29044 14982 29096
rect 15120 29084 15148 29112
rect 15028 29056 15148 29084
rect 14737 29019 14795 29025
rect 14737 28985 14749 29019
rect 14783 29016 14795 29019
rect 15028 29016 15056 29056
rect 14783 28988 15056 29016
rect 15105 29019 15163 29025
rect 14783 28985 14795 28988
rect 14737 28979 14795 28985
rect 15105 28985 15117 29019
rect 15151 29016 15163 29019
rect 15672 29016 15700 29192
rect 17218 29180 17224 29192
rect 17276 29180 17282 29232
rect 17865 29223 17923 29229
rect 17865 29189 17877 29223
rect 17911 29220 17923 29223
rect 18690 29220 18696 29232
rect 17911 29192 18696 29220
rect 17911 29189 17923 29192
rect 17865 29183 17923 29189
rect 16669 29155 16727 29161
rect 16669 29121 16681 29155
rect 16715 29152 16727 29155
rect 16715 29124 16804 29152
rect 16715 29121 16727 29124
rect 16669 29115 16727 29121
rect 15746 29044 15752 29096
rect 15804 29084 15810 29096
rect 16301 29087 16359 29093
rect 16301 29084 16313 29087
rect 15804 29056 16313 29084
rect 15804 29044 15810 29056
rect 16301 29053 16313 29056
rect 16347 29084 16359 29087
rect 16574 29084 16580 29096
rect 16347 29056 16580 29084
rect 16347 29053 16359 29056
rect 16301 29047 16359 29053
rect 16574 29044 16580 29056
rect 16632 29044 16638 29096
rect 15151 28988 15700 29016
rect 15151 28985 15163 28988
rect 15105 28979 15163 28985
rect 14918 28948 14924 28960
rect 14200 28920 14924 28948
rect 14918 28908 14924 28920
rect 14976 28948 14982 28960
rect 15013 28951 15071 28957
rect 15013 28948 15025 28951
rect 14976 28920 15025 28948
rect 14976 28908 14982 28920
rect 15013 28917 15025 28920
rect 15059 28948 15071 28951
rect 15746 28948 15752 28960
rect 15059 28920 15752 28948
rect 15059 28917 15071 28920
rect 15013 28911 15071 28917
rect 15746 28908 15752 28920
rect 15804 28908 15810 28960
rect 16114 28948 16120 28960
rect 16075 28920 16120 28948
rect 16114 28908 16120 28920
rect 16172 28908 16178 28960
rect 16776 28948 16804 29124
rect 17034 29112 17040 29164
rect 17092 29152 17098 29164
rect 17402 29152 17408 29164
rect 17092 29124 17408 29152
rect 17092 29112 17098 29124
rect 17402 29112 17408 29124
rect 17460 29112 17466 29164
rect 17880 29152 17908 29183
rect 18690 29180 18696 29192
rect 18748 29180 18754 29232
rect 18874 29220 18880 29232
rect 18835 29192 18880 29220
rect 18874 29180 18880 29192
rect 18932 29180 18938 29232
rect 19058 29180 19064 29232
rect 19116 29220 19122 29232
rect 19334 29220 19340 29232
rect 19116 29192 19340 29220
rect 19116 29180 19122 29192
rect 19334 29180 19340 29192
rect 19392 29220 19398 29232
rect 19392 29192 19437 29220
rect 19392 29180 19398 29192
rect 17512 29124 17908 29152
rect 18049 29155 18107 29161
rect 17218 29044 17224 29096
rect 17276 29084 17282 29096
rect 17512 29084 17540 29124
rect 18049 29121 18061 29155
rect 18095 29152 18107 29155
rect 18414 29152 18420 29164
rect 18095 29124 18420 29152
rect 18095 29121 18107 29124
rect 18049 29115 18107 29121
rect 18414 29112 18420 29124
rect 18472 29152 18478 29164
rect 20257 29155 20315 29161
rect 20257 29152 20269 29155
rect 18472 29124 20269 29152
rect 18472 29112 18478 29124
rect 20257 29121 20269 29124
rect 20303 29121 20315 29155
rect 20257 29115 20315 29121
rect 17276 29056 17540 29084
rect 17276 29044 17282 29056
rect 17770 29044 17776 29096
rect 17828 29044 17834 29096
rect 18141 29087 18199 29093
rect 18141 29053 18153 29087
rect 18187 29084 18199 29087
rect 18690 29084 18696 29096
rect 18187 29056 18696 29084
rect 18187 29053 18199 29056
rect 18141 29047 18199 29053
rect 18690 29044 18696 29056
rect 18748 29044 18754 29096
rect 19426 29084 19432 29096
rect 19387 29056 19432 29084
rect 19426 29044 19432 29056
rect 19484 29084 19490 29096
rect 20625 29087 20683 29093
rect 20625 29084 20637 29087
rect 19484 29056 20637 29084
rect 19484 29044 19490 29056
rect 20625 29053 20637 29056
rect 20671 29053 20683 29087
rect 20625 29047 20683 29053
rect 17034 29016 17040 29028
rect 16995 28988 17040 29016
rect 17034 28976 17040 28988
rect 17092 28976 17098 29028
rect 17788 29016 17816 29044
rect 17144 28988 17816 29016
rect 17144 28948 17172 28988
rect 18874 28976 18880 29028
rect 18932 29016 18938 29028
rect 18932 28988 19380 29016
rect 18932 28976 18938 28988
rect 16776 28920 17172 28948
rect 19352 28948 19380 28988
rect 19426 28948 19432 28960
rect 19352 28920 19432 28948
rect 19426 28908 19432 28920
rect 19484 28908 19490 28960
rect 1104 28858 28888 28880
rect 1104 28806 10982 28858
rect 11034 28806 11046 28858
rect 11098 28806 11110 28858
rect 11162 28806 11174 28858
rect 11226 28806 20982 28858
rect 21034 28806 21046 28858
rect 21098 28806 21110 28858
rect 21162 28806 21174 28858
rect 21226 28806 28888 28858
rect 1104 28784 28888 28806
rect 5534 28744 5540 28756
rect 5495 28716 5540 28744
rect 5534 28704 5540 28716
rect 5592 28704 5598 28756
rect 6178 28744 6184 28756
rect 6139 28716 6184 28744
rect 6178 28704 6184 28716
rect 6236 28704 6242 28756
rect 6546 28744 6552 28756
rect 6507 28716 6552 28744
rect 6546 28704 6552 28716
rect 6604 28704 6610 28756
rect 9398 28744 9404 28756
rect 9359 28716 9404 28744
rect 9398 28704 9404 28716
rect 9456 28704 9462 28756
rect 9674 28744 9680 28756
rect 9635 28716 9680 28744
rect 9674 28704 9680 28716
rect 9732 28704 9738 28756
rect 11422 28704 11428 28756
rect 11480 28744 11486 28756
rect 11480 28716 11744 28744
rect 11480 28704 11486 28716
rect 9122 28676 9128 28688
rect 9083 28648 9128 28676
rect 9122 28636 9128 28648
rect 9180 28636 9186 28688
rect 11606 28676 11612 28688
rect 10796 28648 11612 28676
rect 1394 28608 1400 28620
rect 1355 28580 1400 28608
rect 1394 28568 1400 28580
rect 1452 28568 1458 28620
rect 5718 28608 5724 28620
rect 5679 28580 5724 28608
rect 5718 28568 5724 28580
rect 5776 28568 5782 28620
rect 8478 28568 8484 28620
rect 8536 28608 8542 28620
rect 8573 28611 8631 28617
rect 8573 28608 8585 28611
rect 8536 28580 8585 28608
rect 8536 28568 8542 28580
rect 8573 28577 8585 28580
rect 8619 28608 8631 28611
rect 9214 28608 9220 28620
rect 8619 28580 9220 28608
rect 8619 28577 8631 28580
rect 8573 28571 8631 28577
rect 9214 28568 9220 28580
rect 9272 28568 9278 28620
rect 9398 28568 9404 28620
rect 9456 28608 9462 28620
rect 10796 28617 10824 28648
rect 11606 28636 11612 28648
rect 11664 28636 11670 28688
rect 10781 28611 10839 28617
rect 10781 28608 10793 28611
rect 9456 28580 10793 28608
rect 9456 28568 9462 28580
rect 10781 28577 10793 28580
rect 10827 28577 10839 28611
rect 10781 28571 10839 28577
rect 11333 28611 11391 28617
rect 11333 28577 11345 28611
rect 11379 28608 11391 28611
rect 11514 28608 11520 28620
rect 11379 28580 11520 28608
rect 11379 28577 11391 28580
rect 11333 28571 11391 28577
rect 11514 28568 11520 28580
rect 11572 28568 11578 28620
rect 11716 28608 11744 28716
rect 12526 28704 12532 28756
rect 12584 28744 12590 28756
rect 13078 28744 13084 28756
rect 12584 28716 13084 28744
rect 12584 28704 12590 28716
rect 12342 28636 12348 28688
rect 12400 28676 12406 28688
rect 12912 28685 12940 28716
rect 13078 28704 13084 28716
rect 13136 28704 13142 28756
rect 13170 28704 13176 28756
rect 13228 28744 13234 28756
rect 14001 28747 14059 28753
rect 14001 28744 14013 28747
rect 13228 28716 14013 28744
rect 13228 28704 13234 28716
rect 14001 28713 14013 28716
rect 14047 28744 14059 28747
rect 15378 28744 15384 28756
rect 14047 28716 15384 28744
rect 14047 28713 14059 28716
rect 14001 28707 14059 28713
rect 15378 28704 15384 28716
rect 15436 28704 15442 28756
rect 15565 28747 15623 28753
rect 15565 28713 15577 28747
rect 15611 28744 15623 28747
rect 15746 28744 15752 28756
rect 15611 28716 15752 28744
rect 15611 28713 15623 28716
rect 15565 28707 15623 28713
rect 15746 28704 15752 28716
rect 15804 28704 15810 28756
rect 16298 28744 16304 28756
rect 16259 28716 16304 28744
rect 16298 28704 16304 28716
rect 16356 28704 16362 28756
rect 16574 28704 16580 28756
rect 16632 28744 16638 28756
rect 17497 28747 17555 28753
rect 17497 28744 17509 28747
rect 16632 28716 17509 28744
rect 16632 28704 16638 28716
rect 17497 28713 17509 28716
rect 17543 28713 17555 28747
rect 18141 28747 18199 28753
rect 18141 28744 18153 28747
rect 17497 28707 17555 28713
rect 17696 28716 18153 28744
rect 12805 28679 12863 28685
rect 12805 28676 12817 28679
rect 12400 28648 12817 28676
rect 12400 28636 12406 28648
rect 12805 28645 12817 28648
rect 12851 28645 12863 28679
rect 12805 28639 12863 28645
rect 12897 28679 12955 28685
rect 12897 28645 12909 28679
rect 12943 28645 12955 28679
rect 12897 28639 12955 28645
rect 13262 28636 13268 28688
rect 13320 28676 13326 28688
rect 13633 28679 13691 28685
rect 13633 28676 13645 28679
rect 13320 28648 13645 28676
rect 13320 28636 13326 28648
rect 13633 28645 13645 28648
rect 13679 28676 13691 28679
rect 15286 28676 15292 28688
rect 13679 28648 15292 28676
rect 13679 28645 13691 28648
rect 13633 28639 13691 28645
rect 15286 28636 15292 28648
rect 15344 28676 15350 28688
rect 15473 28679 15531 28685
rect 15473 28676 15485 28679
rect 15344 28648 15485 28676
rect 15344 28636 15350 28648
rect 15473 28645 15485 28648
rect 15519 28645 15531 28679
rect 15473 28639 15531 28645
rect 15657 28679 15715 28685
rect 15657 28645 15669 28679
rect 15703 28645 15715 28679
rect 15657 28639 15715 28645
rect 11624 28580 11744 28608
rect 12069 28611 12127 28617
rect 11624 28552 11652 28580
rect 12069 28577 12081 28611
rect 12115 28608 12127 28611
rect 12437 28611 12495 28617
rect 12437 28608 12449 28611
rect 12115 28580 12449 28608
rect 12115 28577 12127 28580
rect 12069 28571 12127 28577
rect 12437 28577 12449 28580
rect 12483 28608 12495 28611
rect 12710 28608 12716 28620
rect 12483 28580 12716 28608
rect 12483 28577 12495 28580
rect 12437 28571 12495 28577
rect 12710 28568 12716 28580
rect 12768 28568 12774 28620
rect 13722 28568 13728 28620
rect 13780 28608 13786 28620
rect 14093 28611 14151 28617
rect 14093 28608 14105 28611
rect 13780 28580 14105 28608
rect 13780 28568 13786 28580
rect 14093 28577 14105 28580
rect 14139 28608 14151 28611
rect 14550 28608 14556 28620
rect 14139 28580 14556 28608
rect 14139 28577 14151 28580
rect 14093 28571 14151 28577
rect 14550 28568 14556 28580
rect 14608 28568 14614 28620
rect 14918 28608 14924 28620
rect 14879 28580 14924 28608
rect 14918 28568 14924 28580
rect 14976 28568 14982 28620
rect 15672 28608 15700 28639
rect 15580 28580 15700 28608
rect 15764 28608 15792 28704
rect 16022 28636 16028 28688
rect 16080 28676 16086 28688
rect 16853 28679 16911 28685
rect 16080 28648 16528 28676
rect 16080 28636 16086 28648
rect 16390 28608 16396 28620
rect 15764 28580 16396 28608
rect 1578 28500 1584 28552
rect 1636 28540 1642 28552
rect 1673 28543 1731 28549
rect 1673 28540 1685 28543
rect 1636 28512 1685 28540
rect 1636 28500 1642 28512
rect 1673 28509 1685 28512
rect 1719 28509 1731 28543
rect 1673 28503 1731 28509
rect 6917 28543 6975 28549
rect 6917 28509 6929 28543
rect 6963 28540 6975 28543
rect 7745 28543 7803 28549
rect 7745 28540 7757 28543
rect 6963 28512 7757 28540
rect 6963 28509 6975 28512
rect 6917 28503 6975 28509
rect 7745 28509 7757 28512
rect 7791 28540 7803 28543
rect 7834 28540 7840 28552
rect 7791 28512 7840 28540
rect 7791 28509 7803 28512
rect 7745 28503 7803 28509
rect 7834 28500 7840 28512
rect 7892 28500 7898 28552
rect 8297 28543 8355 28549
rect 8297 28540 8309 28543
rect 8220 28512 8309 28540
rect 7285 28475 7343 28481
rect 7285 28441 7297 28475
rect 7331 28472 7343 28475
rect 7926 28472 7932 28484
rect 7331 28444 7932 28472
rect 7331 28441 7343 28444
rect 7285 28435 7343 28441
rect 7926 28432 7932 28444
rect 7984 28432 7990 28484
rect 8220 28416 8248 28512
rect 8297 28509 8309 28512
rect 8343 28509 8355 28543
rect 8297 28503 8355 28509
rect 8386 28500 8392 28552
rect 8444 28540 8450 28552
rect 8757 28543 8815 28549
rect 8757 28540 8769 28543
rect 8444 28512 8769 28540
rect 8444 28500 8450 28512
rect 8757 28509 8769 28512
rect 8803 28509 8815 28543
rect 11422 28540 11428 28552
rect 11383 28512 11428 28540
rect 8757 28503 8815 28509
rect 11422 28500 11428 28512
rect 11480 28500 11486 28552
rect 11606 28500 11612 28552
rect 11664 28500 11670 28552
rect 11698 28500 11704 28552
rect 11756 28540 11762 28552
rect 12529 28543 12587 28549
rect 12529 28540 12541 28543
rect 11756 28512 12541 28540
rect 11756 28500 11762 28512
rect 12529 28509 12541 28512
rect 12575 28509 12587 28543
rect 13262 28540 13268 28552
rect 13223 28512 13268 28540
rect 12529 28503 12587 28509
rect 13262 28500 13268 28512
rect 13320 28500 13326 28552
rect 13814 28500 13820 28552
rect 13872 28540 13878 28552
rect 15289 28543 15347 28549
rect 15289 28540 15301 28543
rect 13872 28512 15301 28540
rect 13872 28500 13878 28512
rect 15289 28509 15301 28512
rect 15335 28540 15347 28543
rect 15378 28540 15384 28552
rect 15335 28512 15384 28540
rect 15335 28509 15347 28512
rect 15289 28503 15347 28509
rect 15378 28500 15384 28512
rect 15436 28500 15442 28552
rect 9490 28432 9496 28484
rect 9548 28472 9554 28484
rect 9677 28475 9735 28481
rect 9677 28472 9689 28475
rect 9548 28444 9689 28472
rect 9548 28432 9554 28444
rect 9677 28441 9689 28444
rect 9723 28472 9735 28475
rect 10321 28475 10379 28481
rect 10321 28472 10333 28475
rect 9723 28444 10333 28472
rect 9723 28441 9735 28444
rect 9677 28435 9735 28441
rect 10321 28441 10333 28444
rect 10367 28441 10379 28475
rect 10321 28435 10379 28441
rect 10410 28432 10416 28484
rect 10468 28472 10474 28484
rect 10689 28475 10747 28481
rect 10689 28472 10701 28475
rect 10468 28444 10701 28472
rect 10468 28432 10474 28444
rect 10689 28441 10701 28444
rect 10735 28441 10747 28475
rect 10689 28435 10747 28441
rect 13354 28432 13360 28484
rect 13412 28472 13418 28484
rect 14277 28475 14335 28481
rect 14277 28472 14289 28475
rect 13412 28444 14289 28472
rect 13412 28432 13418 28444
rect 14277 28441 14289 28444
rect 14323 28441 14335 28475
rect 14277 28435 14335 28441
rect 14366 28432 14372 28484
rect 14424 28472 14430 28484
rect 14553 28475 14611 28481
rect 14553 28472 14565 28475
rect 14424 28444 14565 28472
rect 14424 28432 14430 28444
rect 14553 28441 14565 28444
rect 14599 28472 14611 28475
rect 14918 28472 14924 28484
rect 14599 28444 14924 28472
rect 14599 28441 14611 28444
rect 14553 28435 14611 28441
rect 14918 28432 14924 28444
rect 14976 28432 14982 28484
rect 15580 28472 15608 28580
rect 16390 28568 16396 28580
rect 16448 28568 16454 28620
rect 15654 28500 15660 28552
rect 15712 28540 15718 28552
rect 16025 28543 16083 28549
rect 16025 28540 16037 28543
rect 15712 28512 16037 28540
rect 15712 28500 15718 28512
rect 16025 28509 16037 28512
rect 16071 28509 16083 28543
rect 16025 28503 16083 28509
rect 15930 28472 15936 28484
rect 15580 28444 15936 28472
rect 15930 28432 15936 28444
rect 15988 28432 15994 28484
rect 16114 28432 16120 28484
rect 16172 28432 16178 28484
rect 16500 28472 16528 28648
rect 16853 28645 16865 28679
rect 16899 28676 16911 28679
rect 17034 28676 17040 28688
rect 16899 28648 17040 28676
rect 16899 28645 16911 28648
rect 16853 28639 16911 28645
rect 17034 28636 17040 28648
rect 17092 28636 17098 28688
rect 17218 28636 17224 28688
rect 17276 28676 17282 28688
rect 17276 28648 17632 28676
rect 17276 28636 17282 28648
rect 17604 28552 17632 28648
rect 16850 28500 16856 28552
rect 16908 28540 16914 28552
rect 17000 28543 17058 28549
rect 17000 28540 17012 28543
rect 16908 28512 17012 28540
rect 16908 28500 16914 28512
rect 17000 28509 17012 28512
rect 17046 28509 17058 28543
rect 17218 28540 17224 28552
rect 17179 28512 17224 28540
rect 17000 28503 17058 28509
rect 17218 28500 17224 28512
rect 17276 28500 17282 28552
rect 17586 28500 17592 28552
rect 17644 28500 17650 28552
rect 17696 28472 17724 28716
rect 18141 28713 18153 28716
rect 18187 28744 18199 28747
rect 18690 28744 18696 28756
rect 18187 28716 18696 28744
rect 18187 28713 18199 28716
rect 18141 28707 18199 28713
rect 18690 28704 18696 28716
rect 18748 28704 18754 28756
rect 18874 28744 18880 28756
rect 18835 28716 18880 28744
rect 18874 28704 18880 28716
rect 18932 28704 18938 28756
rect 19334 28744 19340 28756
rect 19295 28716 19340 28744
rect 19334 28704 19340 28716
rect 19392 28704 19398 28756
rect 19981 28747 20039 28753
rect 19981 28713 19993 28747
rect 20027 28744 20039 28747
rect 20070 28744 20076 28756
rect 20027 28716 20076 28744
rect 20027 28713 20039 28716
rect 19981 28707 20039 28713
rect 20070 28704 20076 28716
rect 20128 28704 20134 28756
rect 20346 28744 20352 28756
rect 20307 28716 20352 28744
rect 20346 28704 20352 28716
rect 20404 28704 20410 28756
rect 17954 28568 17960 28620
rect 18012 28608 18018 28620
rect 18417 28611 18475 28617
rect 18417 28608 18429 28611
rect 18012 28580 18429 28608
rect 18012 28568 18018 28580
rect 18417 28577 18429 28580
rect 18463 28608 18475 28611
rect 18506 28608 18512 28620
rect 18463 28580 18512 28608
rect 18463 28577 18475 28580
rect 18417 28571 18475 28577
rect 18506 28568 18512 28580
rect 18564 28568 18570 28620
rect 19426 28608 19432 28620
rect 19387 28580 19432 28608
rect 19426 28568 19432 28580
rect 19484 28568 19490 28620
rect 16500 28444 17724 28472
rect 2961 28407 3019 28413
rect 2961 28373 2973 28407
rect 3007 28404 3019 28407
rect 4062 28404 4068 28416
rect 3007 28376 4068 28404
rect 3007 28373 3019 28376
rect 2961 28367 3019 28373
rect 4062 28364 4068 28376
rect 4120 28364 4126 28416
rect 7653 28407 7711 28413
rect 7653 28373 7665 28407
rect 7699 28404 7711 28407
rect 8202 28404 8208 28416
rect 7699 28376 8208 28404
rect 7699 28373 7711 28376
rect 7653 28367 7711 28373
rect 8202 28364 8208 28376
rect 8260 28364 8266 28416
rect 9766 28364 9772 28416
rect 9824 28404 9830 28416
rect 9861 28407 9919 28413
rect 9861 28404 9873 28407
rect 9824 28376 9873 28404
rect 9824 28364 9830 28376
rect 9861 28373 9873 28376
rect 9907 28373 9919 28407
rect 9861 28367 9919 28373
rect 13906 28364 13912 28416
rect 13964 28404 13970 28416
rect 16132 28404 16160 28432
rect 13964 28376 16160 28404
rect 13964 28364 13970 28376
rect 16574 28364 16580 28416
rect 16632 28404 16638 28416
rect 16669 28407 16727 28413
rect 16669 28404 16681 28407
rect 16632 28376 16681 28404
rect 16632 28364 16638 28376
rect 16669 28373 16681 28376
rect 16715 28373 16727 28407
rect 16669 28367 16727 28373
rect 17034 28364 17040 28416
rect 17092 28404 17098 28416
rect 17129 28407 17187 28413
rect 17129 28404 17141 28407
rect 17092 28376 17141 28404
rect 17092 28364 17098 28376
rect 17129 28373 17141 28376
rect 17175 28373 17187 28407
rect 17129 28367 17187 28373
rect 18046 28364 18052 28416
rect 18104 28404 18110 28416
rect 18601 28407 18659 28413
rect 18601 28404 18613 28407
rect 18104 28376 18613 28404
rect 18104 28364 18110 28376
rect 18601 28373 18613 28376
rect 18647 28373 18659 28407
rect 19610 28404 19616 28416
rect 19571 28376 19616 28404
rect 18601 28367 18659 28373
rect 19610 28364 19616 28376
rect 19668 28364 19674 28416
rect 21729 28407 21787 28413
rect 21729 28373 21741 28407
rect 21775 28404 21787 28407
rect 22554 28404 22560 28416
rect 21775 28376 22560 28404
rect 21775 28373 21787 28376
rect 21729 28367 21787 28373
rect 22554 28364 22560 28376
rect 22612 28364 22618 28416
rect 1104 28314 28888 28336
rect 1104 28262 5982 28314
rect 6034 28262 6046 28314
rect 6098 28262 6110 28314
rect 6162 28262 6174 28314
rect 6226 28262 15982 28314
rect 16034 28262 16046 28314
rect 16098 28262 16110 28314
rect 16162 28262 16174 28314
rect 16226 28262 25982 28314
rect 26034 28262 26046 28314
rect 26098 28262 26110 28314
rect 26162 28262 26174 28314
rect 26226 28262 28888 28314
rect 1104 28240 28888 28262
rect 3142 28200 3148 28212
rect 3103 28172 3148 28200
rect 3142 28160 3148 28172
rect 3200 28160 3206 28212
rect 7282 28160 7288 28212
rect 7340 28200 7346 28212
rect 7834 28200 7840 28212
rect 7340 28172 7840 28200
rect 7340 28160 7346 28172
rect 7834 28160 7840 28172
rect 7892 28160 7898 28212
rect 8386 28160 8392 28212
rect 8444 28200 8450 28212
rect 8938 28200 8944 28212
rect 8444 28172 8800 28200
rect 8899 28172 8944 28200
rect 8444 28160 8450 28172
rect 7193 28135 7251 28141
rect 7193 28101 7205 28135
rect 7239 28132 7251 28135
rect 8662 28132 8668 28144
rect 7239 28104 8668 28132
rect 7239 28101 7251 28104
rect 7193 28095 7251 28101
rect 8662 28092 8668 28104
rect 8720 28092 8726 28144
rect 8772 28132 8800 28172
rect 8938 28160 8944 28172
rect 8996 28160 9002 28212
rect 11241 28203 11299 28209
rect 9416 28172 9996 28200
rect 9309 28135 9367 28141
rect 9309 28132 9321 28135
rect 8772 28104 9321 28132
rect 9309 28101 9321 28104
rect 9355 28101 9367 28135
rect 9309 28095 9367 28101
rect 1394 28024 1400 28076
rect 1452 28064 1458 28076
rect 1581 28067 1639 28073
rect 1581 28064 1593 28067
rect 1452 28036 1593 28064
rect 1452 28024 1458 28036
rect 1581 28033 1593 28036
rect 1627 28033 1639 28067
rect 1581 28027 1639 28033
rect 6822 28024 6828 28076
rect 6880 28064 6886 28076
rect 9416 28064 9444 28172
rect 9858 28132 9864 28144
rect 6880 28036 9444 28064
rect 9600 28104 9864 28132
rect 6880 28024 6886 28036
rect 1854 27996 1860 28008
rect 1815 27968 1860 27996
rect 1854 27956 1860 27968
rect 1912 27956 1918 28008
rect 6641 27999 6699 28005
rect 6641 27965 6653 27999
rect 6687 27996 6699 27999
rect 7009 27999 7067 28005
rect 7009 27996 7021 27999
rect 6687 27968 7021 27996
rect 6687 27965 6699 27968
rect 6641 27959 6699 27965
rect 7009 27965 7021 27968
rect 7055 27996 7067 27999
rect 7098 27996 7104 28008
rect 7055 27968 7104 27996
rect 7055 27965 7067 27968
rect 7009 27959 7067 27965
rect 7098 27956 7104 27968
rect 7156 27956 7162 28008
rect 8021 27999 8079 28005
rect 8021 27965 8033 27999
rect 8067 27996 8079 27999
rect 8573 27999 8631 28005
rect 8573 27996 8585 27999
rect 8067 27968 8585 27996
rect 8067 27965 8079 27968
rect 8021 27959 8079 27965
rect 8573 27965 8585 27968
rect 8619 27996 8631 27999
rect 9306 27996 9312 28008
rect 8619 27968 9312 27996
rect 8619 27965 8631 27968
rect 8573 27959 8631 27965
rect 9306 27956 9312 27968
rect 9364 27956 9370 28008
rect 9493 27999 9551 28005
rect 9493 27965 9505 27999
rect 9539 27996 9551 27999
rect 9600 27996 9628 28104
rect 9858 28092 9864 28104
rect 9916 28092 9922 28144
rect 9968 28073 9996 28172
rect 11241 28169 11253 28203
rect 11287 28200 11299 28203
rect 12526 28200 12532 28212
rect 11287 28172 12532 28200
rect 11287 28169 11299 28172
rect 11241 28163 11299 28169
rect 12526 28160 12532 28172
rect 12584 28160 12590 28212
rect 13722 28200 13728 28212
rect 13683 28172 13728 28200
rect 13722 28160 13728 28172
rect 13780 28160 13786 28212
rect 14090 28160 14096 28212
rect 14148 28200 14154 28212
rect 14366 28200 14372 28212
rect 14148 28172 14372 28200
rect 14148 28160 14154 28172
rect 14366 28160 14372 28172
rect 14424 28160 14430 28212
rect 16209 28203 16267 28209
rect 16209 28200 16221 28203
rect 14476 28172 16221 28200
rect 11609 28135 11667 28141
rect 11609 28101 11621 28135
rect 11655 28132 11667 28135
rect 11885 28135 11943 28141
rect 11885 28132 11897 28135
rect 11655 28104 11897 28132
rect 11655 28101 11667 28104
rect 11609 28095 11667 28101
rect 11885 28101 11897 28104
rect 11931 28132 11943 28135
rect 12434 28132 12440 28144
rect 11931 28104 12440 28132
rect 11931 28101 11943 28104
rect 11885 28095 11943 28101
rect 12434 28092 12440 28104
rect 12492 28092 12498 28144
rect 12710 28132 12716 28144
rect 12623 28104 12716 28132
rect 9953 28067 10011 28073
rect 9953 28033 9965 28067
rect 9999 28033 10011 28067
rect 9953 28027 10011 28033
rect 10318 28024 10324 28076
rect 10376 28064 10382 28076
rect 12161 28067 12219 28073
rect 12161 28064 12173 28067
rect 10376 28036 12173 28064
rect 10376 28024 10382 28036
rect 12161 28033 12173 28036
rect 12207 28064 12219 28067
rect 12207 28036 12480 28064
rect 12207 28033 12219 28036
rect 12161 28027 12219 28033
rect 12452 28008 12480 28036
rect 9539 27968 9628 27996
rect 9539 27965 9551 27968
rect 9493 27959 9551 27965
rect 5629 27931 5687 27937
rect 5629 27897 5641 27931
rect 5675 27928 5687 27931
rect 5718 27928 5724 27940
rect 5675 27900 5724 27928
rect 5675 27897 5687 27900
rect 5629 27891 5687 27897
rect 5718 27888 5724 27900
rect 5776 27928 5782 27940
rect 6454 27928 6460 27940
rect 5776 27900 6460 27928
rect 5776 27888 5782 27900
rect 6454 27888 6460 27900
rect 6512 27888 6518 27940
rect 7837 27931 7895 27937
rect 7837 27897 7849 27931
rect 7883 27928 7895 27931
rect 9214 27928 9220 27940
rect 7883 27900 9220 27928
rect 7883 27897 7895 27900
rect 7837 27891 7895 27897
rect 9214 27888 9220 27900
rect 9272 27888 9278 27940
rect 9508 27928 9536 27959
rect 9674 27956 9680 28008
rect 9732 27996 9738 28008
rect 10042 27996 10048 28008
rect 9732 27968 9777 27996
rect 10003 27968 10048 27996
rect 9732 27956 9738 27968
rect 10042 27956 10048 27968
rect 10100 27956 10106 28008
rect 10686 27956 10692 28008
rect 10744 27996 10750 28008
rect 11333 27999 11391 28005
rect 11333 27996 11345 27999
rect 10744 27968 11345 27996
rect 10744 27956 10750 27968
rect 11333 27965 11345 27968
rect 11379 27996 11391 27999
rect 11609 27999 11667 28005
rect 11609 27996 11621 27999
rect 11379 27968 11621 27996
rect 11379 27965 11391 27968
rect 11333 27959 11391 27965
rect 11609 27965 11621 27968
rect 11655 27965 11667 27999
rect 12434 27996 12440 28008
rect 12347 27968 12440 27996
rect 11609 27959 11667 27965
rect 12434 27956 12440 27968
rect 12492 27956 12498 28008
rect 12636 28005 12664 28104
rect 12710 28092 12716 28104
rect 12768 28132 12774 28144
rect 14476 28132 14504 28172
rect 16209 28169 16221 28172
rect 16255 28169 16267 28203
rect 16390 28200 16396 28212
rect 16351 28172 16396 28200
rect 16209 28163 16267 28169
rect 16390 28160 16396 28172
rect 16448 28160 16454 28212
rect 16758 28200 16764 28212
rect 16719 28172 16764 28200
rect 16758 28160 16764 28172
rect 16816 28160 16822 28212
rect 17218 28160 17224 28212
rect 17276 28200 17282 28212
rect 17681 28203 17739 28209
rect 17681 28200 17693 28203
rect 17276 28172 17693 28200
rect 17276 28160 17282 28172
rect 17681 28169 17693 28172
rect 17727 28169 17739 28203
rect 19426 28200 19432 28212
rect 19387 28172 19432 28200
rect 17681 28163 17739 28169
rect 19426 28160 19432 28172
rect 19484 28160 19490 28212
rect 20346 28160 20352 28212
rect 20404 28200 20410 28212
rect 20901 28203 20959 28209
rect 20901 28200 20913 28203
rect 20404 28172 20913 28200
rect 20404 28160 20410 28172
rect 20901 28169 20913 28172
rect 20947 28169 20959 28203
rect 21542 28200 21548 28212
rect 21503 28172 21548 28200
rect 20901 28163 20959 28169
rect 21542 28160 21548 28172
rect 21600 28200 21606 28212
rect 21600 28172 21772 28200
rect 21600 28160 21606 28172
rect 12768 28104 14504 28132
rect 12768 28092 12774 28104
rect 14918 28092 14924 28144
rect 14976 28132 14982 28144
rect 14976 28104 17724 28132
rect 14976 28092 14982 28104
rect 14090 28024 14096 28076
rect 14148 28064 14154 28076
rect 14277 28067 14335 28073
rect 14277 28064 14289 28067
rect 14148 28036 14289 28064
rect 14148 28024 14154 28036
rect 14277 28033 14289 28036
rect 14323 28033 14335 28067
rect 14277 28027 14335 28033
rect 15562 28024 15568 28076
rect 15620 28064 15626 28076
rect 16485 28067 16543 28073
rect 16485 28064 16497 28067
rect 15620 28036 16497 28064
rect 15620 28024 15626 28036
rect 16485 28033 16497 28036
rect 16531 28033 16543 28067
rect 17405 28067 17463 28073
rect 17405 28064 17417 28067
rect 16485 28027 16543 28033
rect 16592 28036 17417 28064
rect 12621 27999 12679 28005
rect 12621 27965 12633 27999
rect 12667 27965 12679 27999
rect 12621 27959 12679 27965
rect 12713 27999 12771 28005
rect 12713 27965 12725 27999
rect 12759 27965 12771 27999
rect 13170 27996 13176 28008
rect 13131 27968 13176 27996
rect 12713 27959 12771 27965
rect 9766 27928 9772 27940
rect 9324 27900 9536 27928
rect 9692 27900 9772 27928
rect 6273 27863 6331 27869
rect 6273 27829 6285 27863
rect 6319 27860 6331 27863
rect 6822 27860 6828 27872
rect 6319 27832 6828 27860
rect 6319 27829 6331 27832
rect 6273 27823 6331 27829
rect 6822 27820 6828 27832
rect 6880 27820 6886 27872
rect 8202 27860 8208 27872
rect 8163 27832 8208 27860
rect 8202 27820 8208 27832
rect 8260 27820 8266 27872
rect 8478 27820 8484 27872
rect 8536 27860 8542 27872
rect 9324 27860 9352 27900
rect 9692 27872 9720 27900
rect 9766 27888 9772 27900
rect 9824 27888 9830 27940
rect 9858 27888 9864 27940
rect 9916 27928 9922 27940
rect 10134 27928 10140 27940
rect 9916 27900 10140 27928
rect 9916 27888 9922 27900
rect 10134 27888 10140 27900
rect 10192 27888 10198 27940
rect 10873 27931 10931 27937
rect 10873 27897 10885 27931
rect 10919 27928 10931 27931
rect 12728 27928 12756 27959
rect 13170 27956 13176 27968
rect 13228 27956 13234 28008
rect 13998 27956 14004 28008
rect 14056 27996 14062 28008
rect 14185 27999 14243 28005
rect 14185 27996 14197 27999
rect 14056 27968 14197 27996
rect 14056 27956 14062 27968
rect 14185 27965 14197 27968
rect 14231 27965 14243 27999
rect 14185 27959 14243 27965
rect 13078 27928 13084 27940
rect 10919 27900 13084 27928
rect 10919 27897 10931 27900
rect 10873 27891 10931 27897
rect 13078 27888 13084 27900
rect 13136 27888 13142 27940
rect 14200 27928 14228 27959
rect 14366 27956 14372 28008
rect 14424 27996 14430 28008
rect 14553 27999 14611 28005
rect 14553 27996 14565 27999
rect 14424 27968 14565 27996
rect 14424 27956 14430 27968
rect 14553 27965 14565 27968
rect 14599 27965 14611 27999
rect 14918 27996 14924 28008
rect 14879 27968 14924 27996
rect 14553 27959 14611 27965
rect 14918 27956 14924 27968
rect 14976 27956 14982 28008
rect 15102 27956 15108 28008
rect 15160 27996 15166 28008
rect 15657 27999 15715 28005
rect 15657 27996 15669 27999
rect 15160 27968 15669 27996
rect 15160 27956 15166 27968
rect 15657 27965 15669 27968
rect 15703 27996 15715 27999
rect 15930 27996 15936 28008
rect 15703 27968 15936 27996
rect 15703 27965 15715 27968
rect 15657 27959 15715 27965
rect 15930 27956 15936 27968
rect 15988 27956 15994 28008
rect 16206 27996 16212 28008
rect 16167 27968 16212 27996
rect 16206 27956 16212 27968
rect 16264 27956 16270 28008
rect 16592 28005 16620 28036
rect 17405 28033 17417 28036
rect 17451 28064 17463 28067
rect 17586 28064 17592 28076
rect 17451 28036 17592 28064
rect 17451 28033 17463 28036
rect 17405 28027 17463 28033
rect 17586 28024 17592 28036
rect 17644 28024 17650 28076
rect 17696 28064 17724 28104
rect 18230 28092 18236 28144
rect 18288 28132 18294 28144
rect 18325 28135 18383 28141
rect 18325 28132 18337 28135
rect 18288 28104 18337 28132
rect 18288 28092 18294 28104
rect 18325 28101 18337 28104
rect 18371 28101 18383 28135
rect 20714 28132 20720 28144
rect 20675 28104 20720 28132
rect 18325 28095 18383 28101
rect 20714 28092 20720 28104
rect 20772 28092 20778 28144
rect 19978 28064 19984 28076
rect 17696 28036 19984 28064
rect 16577 27999 16635 28005
rect 16577 27965 16589 27999
rect 16623 27965 16635 27999
rect 16577 27959 16635 27965
rect 17954 27956 17960 28008
rect 18012 27996 18018 28008
rect 18509 27999 18567 28005
rect 18509 27996 18521 27999
rect 18012 27968 18521 27996
rect 18012 27956 18018 27968
rect 18509 27965 18521 27968
rect 18555 27965 18567 27999
rect 18690 27996 18696 28008
rect 18651 27968 18696 27996
rect 18509 27959 18567 27965
rect 15562 27928 15568 27940
rect 14200 27900 15568 27928
rect 15562 27888 15568 27900
rect 15620 27888 15626 27940
rect 16025 27931 16083 27937
rect 16025 27897 16037 27931
rect 16071 27928 16083 27931
rect 16666 27928 16672 27940
rect 16071 27900 16672 27928
rect 16071 27897 16083 27900
rect 16025 27891 16083 27897
rect 8536 27832 9352 27860
rect 8536 27820 8542 27832
rect 9674 27820 9680 27872
rect 9732 27820 9738 27872
rect 11517 27863 11575 27869
rect 11517 27829 11529 27863
rect 11563 27860 11575 27863
rect 11698 27860 11704 27872
rect 11563 27832 11704 27860
rect 11563 27829 11575 27832
rect 11517 27823 11575 27829
rect 11698 27820 11704 27832
rect 11756 27820 11762 27872
rect 14093 27863 14151 27869
rect 14093 27829 14105 27863
rect 14139 27860 14151 27863
rect 14366 27860 14372 27872
rect 14139 27832 14372 27860
rect 14139 27829 14151 27832
rect 14093 27823 14151 27829
rect 14366 27820 14372 27832
rect 14424 27820 14430 27872
rect 15378 27820 15384 27872
rect 15436 27860 15442 27872
rect 16040 27860 16068 27891
rect 16666 27888 16672 27900
rect 16724 27888 16730 27940
rect 18524 27928 18552 27959
rect 18690 27956 18696 27968
rect 18748 27956 18754 28008
rect 18782 27956 18788 28008
rect 18840 27996 18846 28008
rect 19904 28005 19932 28036
rect 19978 28024 19984 28036
rect 20036 28064 20042 28076
rect 21744 28073 21772 28172
rect 20349 28067 20407 28073
rect 20349 28064 20361 28067
rect 20036 28036 20361 28064
rect 20036 28024 20042 28036
rect 20349 28033 20361 28036
rect 20395 28033 20407 28067
rect 20349 28027 20407 28033
rect 21729 28067 21787 28073
rect 21729 28033 21741 28067
rect 21775 28033 21787 28067
rect 21729 28027 21787 28033
rect 21910 28024 21916 28076
rect 21968 28064 21974 28076
rect 22649 28067 22707 28073
rect 22649 28064 22661 28067
rect 21968 28036 22661 28064
rect 21968 28024 21974 28036
rect 22649 28033 22661 28036
rect 22695 28064 22707 28067
rect 23382 28064 23388 28076
rect 22695 28036 23388 28064
rect 22695 28033 22707 28036
rect 22649 28027 22707 28033
rect 23382 28024 23388 28036
rect 23440 28024 23446 28076
rect 18877 27999 18935 28005
rect 18877 27996 18889 27999
rect 18840 27968 18889 27996
rect 18840 27956 18846 27968
rect 18877 27965 18889 27968
rect 18923 27965 18935 27999
rect 18877 27959 18935 27965
rect 19889 27999 19947 28005
rect 19889 27965 19901 27999
rect 19935 27965 19947 27999
rect 19889 27959 19947 27965
rect 20714 27956 20720 28008
rect 20772 27996 20778 28008
rect 21085 27999 21143 28005
rect 21085 27996 21097 27999
rect 20772 27968 21097 27996
rect 20772 27956 20778 27968
rect 21085 27965 21097 27968
rect 21131 27965 21143 27999
rect 22554 27996 22560 28008
rect 22467 27968 22560 27996
rect 21085 27959 21143 27965
rect 22554 27956 22560 27968
rect 22612 27996 22618 28008
rect 23658 27996 23664 28008
rect 22612 27968 23664 27996
rect 22612 27956 22618 27968
rect 23658 27956 23664 27968
rect 23716 27956 23722 28008
rect 19242 27928 19248 27940
rect 18524 27900 19248 27928
rect 19242 27888 19248 27900
rect 19300 27888 19306 27940
rect 21818 27928 21824 27940
rect 21779 27900 21824 27928
rect 21818 27888 21824 27900
rect 21876 27888 21882 27940
rect 20070 27860 20076 27872
rect 15436 27832 16068 27860
rect 20031 27832 20076 27860
rect 15436 27820 15442 27832
rect 20070 27820 20076 27832
rect 20128 27820 20134 27872
rect 1104 27770 28888 27792
rect 1104 27718 10982 27770
rect 11034 27718 11046 27770
rect 11098 27718 11110 27770
rect 11162 27718 11174 27770
rect 11226 27718 20982 27770
rect 21034 27718 21046 27770
rect 21098 27718 21110 27770
rect 21162 27718 21174 27770
rect 21226 27718 28888 27770
rect 1104 27696 28888 27718
rect 1394 27616 1400 27668
rect 1452 27656 1458 27668
rect 2317 27659 2375 27665
rect 2317 27656 2329 27659
rect 1452 27628 2329 27656
rect 1452 27616 1458 27628
rect 2317 27625 2329 27628
rect 2363 27625 2375 27659
rect 7374 27656 7380 27668
rect 7335 27628 7380 27656
rect 2317 27619 2375 27625
rect 7374 27616 7380 27628
rect 7432 27616 7438 27668
rect 8202 27616 8208 27668
rect 8260 27656 8266 27668
rect 13354 27656 13360 27668
rect 8260 27628 10180 27656
rect 13315 27628 13360 27656
rect 8260 27616 8266 27628
rect 4614 27588 4620 27600
rect 4575 27560 4620 27588
rect 4614 27548 4620 27560
rect 4672 27588 4678 27600
rect 7193 27591 7251 27597
rect 4672 27560 4844 27588
rect 4672 27548 4678 27560
rect 4816 27529 4844 27560
rect 7193 27557 7205 27591
rect 7239 27588 7251 27591
rect 8478 27588 8484 27600
rect 7239 27560 8484 27588
rect 7239 27557 7251 27560
rect 7193 27551 7251 27557
rect 8478 27548 8484 27560
rect 8536 27548 8542 27600
rect 9582 27548 9588 27600
rect 9640 27588 9646 27600
rect 9861 27591 9919 27597
rect 9861 27588 9873 27591
rect 9640 27560 9873 27588
rect 9640 27548 9646 27560
rect 9861 27557 9873 27560
rect 9907 27588 9919 27591
rect 10152 27588 10180 27628
rect 13354 27616 13360 27628
rect 13412 27616 13418 27668
rect 13906 27616 13912 27668
rect 13964 27616 13970 27668
rect 14458 27656 14464 27668
rect 14371 27628 14464 27656
rect 14458 27616 14464 27628
rect 14516 27656 14522 27668
rect 15102 27656 15108 27668
rect 14516 27628 15108 27656
rect 14516 27616 14522 27628
rect 15102 27616 15108 27628
rect 15160 27616 15166 27668
rect 15286 27616 15292 27668
rect 15344 27656 15350 27668
rect 15841 27659 15899 27665
rect 15841 27656 15853 27659
rect 15344 27628 15853 27656
rect 15344 27616 15350 27628
rect 15841 27625 15853 27628
rect 15887 27625 15899 27659
rect 15841 27619 15899 27625
rect 16206 27616 16212 27668
rect 16264 27656 16270 27668
rect 17586 27656 17592 27668
rect 16264 27628 17592 27656
rect 16264 27616 16270 27628
rect 17586 27616 17592 27628
rect 17644 27616 17650 27668
rect 18506 27656 18512 27668
rect 18467 27628 18512 27656
rect 18506 27616 18512 27628
rect 18564 27616 18570 27668
rect 18782 27616 18788 27668
rect 18840 27656 18846 27668
rect 18840 27628 19288 27656
rect 18840 27616 18846 27628
rect 9907 27560 10088 27588
rect 10152 27560 10916 27588
rect 9907 27557 9919 27560
rect 9861 27551 9919 27557
rect 4801 27523 4859 27529
rect 4801 27489 4813 27523
rect 4847 27489 4859 27523
rect 4801 27483 4859 27489
rect 6825 27523 6883 27529
rect 6825 27489 6837 27523
rect 6871 27520 6883 27523
rect 7926 27520 7932 27532
rect 6871 27492 7932 27520
rect 6871 27489 6883 27492
rect 6825 27483 6883 27489
rect 7926 27480 7932 27492
rect 7984 27480 7990 27532
rect 8297 27523 8355 27529
rect 8297 27489 8309 27523
rect 8343 27520 8355 27523
rect 8386 27520 8392 27532
rect 8343 27492 8392 27520
rect 8343 27489 8355 27492
rect 8297 27483 8355 27489
rect 8386 27480 8392 27492
rect 8444 27480 8450 27532
rect 10060 27529 10088 27560
rect 10045 27523 10103 27529
rect 10045 27489 10057 27523
rect 10091 27489 10103 27523
rect 10410 27520 10416 27532
rect 10371 27492 10416 27520
rect 10045 27483 10103 27489
rect 10410 27480 10416 27492
rect 10468 27480 10474 27532
rect 10888 27529 10916 27560
rect 11054 27548 11060 27600
rect 11112 27588 11118 27600
rect 11517 27591 11575 27597
rect 11517 27588 11529 27591
rect 11112 27560 11529 27588
rect 11112 27548 11118 27560
rect 11517 27557 11529 27560
rect 11563 27588 11575 27591
rect 13924 27588 13952 27616
rect 14550 27588 14556 27600
rect 11563 27560 12572 27588
rect 13924 27560 14556 27588
rect 11563 27557 11575 27560
rect 11517 27551 11575 27557
rect 10873 27523 10931 27529
rect 10873 27489 10885 27523
rect 10919 27489 10931 27523
rect 12066 27520 12072 27532
rect 12027 27492 12072 27520
rect 10873 27483 10931 27489
rect 12066 27480 12072 27492
rect 12124 27480 12130 27532
rect 12544 27529 12572 27560
rect 14550 27548 14556 27560
rect 14608 27548 14614 27600
rect 14829 27591 14887 27597
rect 14829 27557 14841 27591
rect 14875 27588 14887 27591
rect 15470 27588 15476 27600
rect 14875 27560 15476 27588
rect 14875 27557 14887 27560
rect 14829 27551 14887 27557
rect 15470 27548 15476 27560
rect 15528 27588 15534 27600
rect 16298 27588 16304 27600
rect 15528 27560 16304 27588
rect 15528 27548 15534 27560
rect 16298 27548 16304 27560
rect 16356 27548 16362 27600
rect 16390 27548 16396 27600
rect 16448 27548 16454 27600
rect 19260 27588 19288 27628
rect 19337 27591 19395 27597
rect 19337 27588 19349 27591
rect 19260 27560 19349 27588
rect 19337 27557 19349 27560
rect 19383 27557 19395 27591
rect 19337 27551 19395 27557
rect 20714 27548 20720 27600
rect 20772 27548 20778 27600
rect 20806 27548 20812 27600
rect 20864 27548 20870 27600
rect 21729 27591 21787 27597
rect 21729 27557 21741 27591
rect 21775 27588 21787 27591
rect 21910 27588 21916 27600
rect 21775 27560 21916 27588
rect 21775 27557 21787 27560
rect 21729 27551 21787 27557
rect 21910 27548 21916 27560
rect 21968 27548 21974 27600
rect 12529 27523 12587 27529
rect 12529 27489 12541 27523
rect 12575 27489 12587 27523
rect 13906 27520 13912 27532
rect 13867 27492 13912 27520
rect 12529 27483 12587 27489
rect 13906 27480 13912 27492
rect 13964 27480 13970 27532
rect 14458 27480 14464 27532
rect 14516 27520 14522 27532
rect 14642 27520 14648 27532
rect 14516 27492 14648 27520
rect 14516 27480 14522 27492
rect 14642 27480 14648 27492
rect 14700 27480 14706 27532
rect 15381 27523 15439 27529
rect 15381 27489 15393 27523
rect 15427 27520 15439 27523
rect 16408 27520 16436 27548
rect 16666 27520 16672 27532
rect 15427 27492 16436 27520
rect 16627 27492 16672 27520
rect 15427 27489 15439 27492
rect 15381 27483 15439 27489
rect 16666 27480 16672 27492
rect 16724 27480 16730 27532
rect 17586 27480 17592 27532
rect 17644 27520 17650 27532
rect 17770 27520 17776 27532
rect 17644 27492 17776 27520
rect 17644 27480 17650 27492
rect 17770 27480 17776 27492
rect 17828 27520 17834 27532
rect 18874 27520 18880 27532
rect 17828 27492 18184 27520
rect 18835 27492 18880 27520
rect 17828 27480 17834 27492
rect 5074 27452 5080 27464
rect 5035 27424 5080 27452
rect 5074 27412 5080 27424
rect 5132 27412 5138 27464
rect 7282 27412 7288 27464
rect 7340 27452 7346 27464
rect 7745 27455 7803 27461
rect 7745 27452 7757 27455
rect 7340 27424 7757 27452
rect 7340 27412 7346 27424
rect 7745 27421 7757 27424
rect 7791 27421 7803 27455
rect 7745 27415 7803 27421
rect 7834 27412 7840 27464
rect 7892 27452 7898 27464
rect 8205 27455 8263 27461
rect 8205 27452 8217 27455
rect 7892 27424 8217 27452
rect 7892 27412 7898 27424
rect 8205 27421 8217 27424
rect 8251 27452 8263 27455
rect 9030 27452 9036 27464
rect 8251 27424 9036 27452
rect 8251 27421 8263 27424
rect 8205 27415 8263 27421
rect 9030 27412 9036 27424
rect 9088 27412 9094 27464
rect 9125 27455 9183 27461
rect 9125 27421 9137 27455
rect 9171 27452 9183 27455
rect 11422 27452 11428 27464
rect 9171 27424 11428 27452
rect 9171 27421 9183 27424
rect 9125 27415 9183 27421
rect 11422 27412 11428 27424
rect 11480 27452 11486 27464
rect 12989 27455 13047 27461
rect 11480 27424 12112 27452
rect 11480 27412 11486 27424
rect 10318 27344 10324 27396
rect 10376 27384 10382 27396
rect 12084 27393 12112 27424
rect 12989 27421 13001 27455
rect 13035 27452 13047 27455
rect 13170 27452 13176 27464
rect 13035 27424 13176 27452
rect 13035 27421 13047 27424
rect 12989 27415 13047 27421
rect 13170 27412 13176 27424
rect 13228 27412 13234 27464
rect 16393 27455 16451 27461
rect 16393 27421 16405 27455
rect 16439 27452 16451 27455
rect 18046 27452 18052 27464
rect 16439 27424 18052 27452
rect 16439 27421 16451 27424
rect 16393 27415 16451 27421
rect 18046 27412 18052 27424
rect 18104 27412 18110 27464
rect 10873 27387 10931 27393
rect 10873 27384 10885 27387
rect 10376 27356 10885 27384
rect 10376 27344 10382 27356
rect 10873 27353 10885 27356
rect 10919 27353 10931 27387
rect 10873 27347 10931 27353
rect 12069 27387 12127 27393
rect 12069 27353 12081 27387
rect 12115 27353 12127 27387
rect 12069 27347 12127 27353
rect 12434 27344 12440 27396
rect 12492 27384 12498 27396
rect 14093 27387 14151 27393
rect 14093 27384 14105 27387
rect 12492 27356 14105 27384
rect 12492 27344 12498 27356
rect 14093 27353 14105 27356
rect 14139 27353 14151 27387
rect 18156 27384 18184 27492
rect 18874 27480 18880 27492
rect 18932 27480 18938 27532
rect 20070 27520 20076 27532
rect 20031 27492 20076 27520
rect 20070 27480 20076 27492
rect 20128 27480 20134 27532
rect 19334 27412 19340 27464
rect 19392 27452 19398 27464
rect 19705 27455 19763 27461
rect 19705 27452 19717 27455
rect 19392 27424 19717 27452
rect 19392 27412 19398 27424
rect 19705 27421 19717 27424
rect 19751 27421 19763 27455
rect 19705 27415 19763 27421
rect 19061 27387 19119 27393
rect 19061 27384 19073 27387
rect 18156 27356 19073 27384
rect 14093 27347 14151 27353
rect 19061 27353 19073 27356
rect 19107 27353 19119 27387
rect 19061 27347 19119 27353
rect 1578 27316 1584 27328
rect 1539 27288 1584 27316
rect 1578 27276 1584 27288
rect 1636 27276 1642 27328
rect 1854 27276 1860 27328
rect 1912 27316 1918 27328
rect 1949 27319 2007 27325
rect 1949 27316 1961 27319
rect 1912 27288 1961 27316
rect 1912 27276 1918 27288
rect 1949 27285 1961 27288
rect 1995 27285 2007 27319
rect 1949 27279 2007 27285
rect 5718 27276 5724 27328
rect 5776 27316 5782 27328
rect 6181 27319 6239 27325
rect 6181 27316 6193 27319
rect 5776 27288 6193 27316
rect 5776 27276 5782 27288
rect 6181 27285 6193 27288
rect 6227 27285 6239 27319
rect 6181 27279 6239 27285
rect 9214 27276 9220 27328
rect 9272 27316 9278 27328
rect 9401 27319 9459 27325
rect 9401 27316 9413 27319
rect 9272 27288 9413 27316
rect 9272 27276 9278 27288
rect 9401 27285 9413 27288
rect 9447 27316 9459 27319
rect 9490 27316 9496 27328
rect 9447 27288 9496 27316
rect 9447 27285 9459 27288
rect 9401 27279 9459 27285
rect 9490 27276 9496 27288
rect 9548 27276 9554 27328
rect 10962 27276 10968 27328
rect 11020 27316 11026 27328
rect 11606 27316 11612 27328
rect 11020 27288 11612 27316
rect 11020 27276 11026 27288
rect 11606 27276 11612 27288
rect 11664 27316 11670 27328
rect 11793 27319 11851 27325
rect 11793 27316 11805 27319
rect 11664 27288 11805 27316
rect 11664 27276 11670 27288
rect 11793 27285 11805 27288
rect 11839 27316 11851 27319
rect 12342 27316 12348 27328
rect 11839 27288 12348 27316
rect 11839 27285 11851 27288
rect 11793 27279 11851 27285
rect 12342 27276 12348 27288
rect 12400 27276 12406 27328
rect 13722 27316 13728 27328
rect 13683 27288 13728 27316
rect 13722 27276 13728 27288
rect 13780 27276 13786 27328
rect 14918 27276 14924 27328
rect 14976 27316 14982 27328
rect 15102 27316 15108 27328
rect 14976 27288 15108 27316
rect 14976 27276 14982 27288
rect 15102 27276 15108 27288
rect 15160 27276 15166 27328
rect 15286 27276 15292 27328
rect 15344 27316 15350 27328
rect 15565 27319 15623 27325
rect 15565 27316 15577 27319
rect 15344 27288 15577 27316
rect 15344 27276 15350 27288
rect 15565 27285 15577 27288
rect 15611 27285 15623 27319
rect 16298 27316 16304 27328
rect 16259 27288 16304 27316
rect 15565 27279 15623 27285
rect 16298 27276 16304 27288
rect 16356 27316 16362 27328
rect 17034 27316 17040 27328
rect 16356 27288 17040 27316
rect 16356 27276 16362 27288
rect 17034 27276 17040 27288
rect 17092 27276 17098 27328
rect 17770 27316 17776 27328
rect 17731 27288 17776 27316
rect 17770 27276 17776 27288
rect 17828 27276 17834 27328
rect 19886 27276 19892 27328
rect 19944 27316 19950 27328
rect 20732 27316 20760 27548
rect 20824 27464 20852 27548
rect 20806 27412 20812 27464
rect 20864 27412 20870 27464
rect 21085 27319 21143 27325
rect 21085 27316 21097 27319
rect 19944 27288 21097 27316
rect 19944 27276 19950 27288
rect 21085 27285 21097 27288
rect 21131 27285 21143 27319
rect 21085 27279 21143 27285
rect 1104 27226 28888 27248
rect 1104 27174 5982 27226
rect 6034 27174 6046 27226
rect 6098 27174 6110 27226
rect 6162 27174 6174 27226
rect 6226 27174 15982 27226
rect 16034 27174 16046 27226
rect 16098 27174 16110 27226
rect 16162 27174 16174 27226
rect 16226 27174 25982 27226
rect 26034 27174 26046 27226
rect 26098 27174 26110 27226
rect 26162 27174 26174 27226
rect 26226 27174 28888 27226
rect 1104 27152 28888 27174
rect 1394 27072 1400 27124
rect 1452 27112 1458 27124
rect 1581 27115 1639 27121
rect 1581 27112 1593 27115
rect 1452 27084 1593 27112
rect 1452 27072 1458 27084
rect 1581 27081 1593 27084
rect 1627 27081 1639 27115
rect 1581 27075 1639 27081
rect 6641 27115 6699 27121
rect 6641 27081 6653 27115
rect 6687 27112 6699 27115
rect 7834 27112 7840 27124
rect 6687 27084 7840 27112
rect 6687 27081 6699 27084
rect 6641 27075 6699 27081
rect 7834 27072 7840 27084
rect 7892 27072 7898 27124
rect 7926 27072 7932 27124
rect 7984 27112 7990 27124
rect 8297 27115 8355 27121
rect 8297 27112 8309 27115
rect 7984 27084 8309 27112
rect 7984 27072 7990 27084
rect 8297 27081 8309 27084
rect 8343 27081 8355 27115
rect 8297 27075 8355 27081
rect 8846 27072 8852 27124
rect 8904 27112 8910 27124
rect 8941 27115 8999 27121
rect 8941 27112 8953 27115
rect 8904 27084 8953 27112
rect 8904 27072 8910 27084
rect 8941 27081 8953 27084
rect 8987 27112 8999 27115
rect 8987 27084 10640 27112
rect 8987 27081 8999 27084
rect 8941 27075 8999 27081
rect 8386 27004 8392 27056
rect 8444 27044 8450 27056
rect 10505 27047 10563 27053
rect 10505 27044 10517 27047
rect 8444 27016 10517 27044
rect 8444 27004 8450 27016
rect 10505 27013 10517 27016
rect 10551 27013 10563 27047
rect 10505 27007 10563 27013
rect 4249 26979 4307 26985
rect 4249 26945 4261 26979
rect 4295 26976 4307 26979
rect 6273 26979 6331 26985
rect 4295 26948 5764 26976
rect 4295 26945 4307 26948
rect 4249 26939 4307 26945
rect 5736 26920 5764 26948
rect 6273 26945 6285 26979
rect 6319 26976 6331 26979
rect 6638 26976 6644 26988
rect 6319 26948 6644 26976
rect 6319 26945 6331 26948
rect 6273 26939 6331 26945
rect 6638 26936 6644 26948
rect 6696 26976 6702 26988
rect 7193 26979 7251 26985
rect 7193 26976 7205 26979
rect 6696 26948 7205 26976
rect 6696 26936 6702 26948
rect 7193 26945 7205 26948
rect 7239 26976 7251 26979
rect 8404 26976 8432 27004
rect 7239 26948 8432 26976
rect 7239 26945 7251 26948
rect 7193 26939 7251 26945
rect 4706 26908 4712 26920
rect 4667 26880 4712 26908
rect 4706 26868 4712 26880
rect 4764 26868 4770 26920
rect 5074 26868 5080 26920
rect 5132 26908 5138 26920
rect 5169 26911 5227 26917
rect 5169 26908 5181 26911
rect 5132 26880 5181 26908
rect 5132 26868 5138 26880
rect 5169 26877 5181 26880
rect 5215 26877 5227 26911
rect 5350 26908 5356 26920
rect 5311 26880 5356 26908
rect 5169 26871 5227 26877
rect 5350 26868 5356 26880
rect 5408 26868 5414 26920
rect 5718 26908 5724 26920
rect 5679 26880 5724 26908
rect 5718 26868 5724 26880
rect 5776 26868 5782 26920
rect 5905 26911 5963 26917
rect 5905 26877 5917 26911
rect 5951 26908 5963 26911
rect 6362 26908 6368 26920
rect 5951 26880 6368 26908
rect 5951 26877 5963 26880
rect 5905 26871 5963 26877
rect 4617 26843 4675 26849
rect 4617 26809 4629 26843
rect 4663 26840 4675 26843
rect 5920 26840 5948 26871
rect 6362 26868 6368 26880
rect 6420 26868 6426 26920
rect 6914 26908 6920 26920
rect 6875 26880 6920 26908
rect 6914 26868 6920 26880
rect 6972 26868 6978 26920
rect 8846 26868 8852 26920
rect 8904 26908 8910 26920
rect 9214 26908 9220 26920
rect 8904 26880 9220 26908
rect 8904 26868 8910 26880
rect 9214 26868 9220 26880
rect 9272 26908 9278 26920
rect 9582 26917 9588 26920
rect 9401 26911 9459 26917
rect 9401 26908 9413 26911
rect 9272 26880 9413 26908
rect 9272 26868 9278 26880
rect 9401 26877 9413 26880
rect 9447 26877 9459 26911
rect 9401 26871 9459 26877
rect 9570 26911 9588 26917
rect 9570 26877 9582 26911
rect 9570 26871 9588 26877
rect 9582 26868 9588 26871
rect 9640 26868 9646 26920
rect 10225 26911 10283 26917
rect 10225 26877 10237 26911
rect 10271 26877 10283 26911
rect 10225 26871 10283 26877
rect 10321 26911 10379 26917
rect 10321 26877 10333 26911
rect 10367 26908 10379 26911
rect 10612 26908 10640 27084
rect 10870 27072 10876 27124
rect 10928 27112 10934 27124
rect 11057 27115 11115 27121
rect 11057 27112 11069 27115
rect 10928 27084 11069 27112
rect 10928 27072 10934 27084
rect 11057 27081 11069 27084
rect 11103 27081 11115 27115
rect 11057 27075 11115 27081
rect 11885 27115 11943 27121
rect 11885 27081 11897 27115
rect 11931 27112 11943 27115
rect 12066 27112 12072 27124
rect 11931 27084 12072 27112
rect 11931 27081 11943 27084
rect 11885 27075 11943 27081
rect 12066 27072 12072 27084
rect 12124 27072 12130 27124
rect 12802 27072 12808 27124
rect 12860 27112 12866 27124
rect 13354 27112 13360 27124
rect 12860 27084 13360 27112
rect 12860 27072 12866 27084
rect 13354 27072 13360 27084
rect 13412 27072 13418 27124
rect 15562 27072 15568 27124
rect 15620 27112 15626 27124
rect 15746 27112 15752 27124
rect 15620 27084 15752 27112
rect 15620 27072 15626 27084
rect 15746 27072 15752 27084
rect 15804 27072 15810 27124
rect 15933 27115 15991 27121
rect 15933 27081 15945 27115
rect 15979 27112 15991 27115
rect 16390 27112 16396 27124
rect 15979 27084 16396 27112
rect 15979 27081 15991 27084
rect 15933 27075 15991 27081
rect 16390 27072 16396 27084
rect 16448 27072 16454 27124
rect 19518 27072 19524 27124
rect 19576 27112 19582 27124
rect 19613 27115 19671 27121
rect 19613 27112 19625 27115
rect 19576 27084 19625 27112
rect 19576 27072 19582 27084
rect 19613 27081 19625 27084
rect 19659 27112 19671 27115
rect 19794 27112 19800 27124
rect 19659 27084 19800 27112
rect 19659 27081 19671 27084
rect 19613 27075 19671 27081
rect 19794 27072 19800 27084
rect 19852 27072 19858 27124
rect 20070 27112 20076 27124
rect 20031 27084 20076 27112
rect 20070 27072 20076 27084
rect 20128 27072 20134 27124
rect 13906 27044 13912 27056
rect 13867 27016 13912 27044
rect 13906 27004 13912 27016
rect 13964 27004 13970 27056
rect 15102 27004 15108 27056
rect 15160 27044 15166 27056
rect 16025 27047 16083 27053
rect 16025 27044 16037 27047
rect 15160 27016 16037 27044
rect 15160 27004 15166 27016
rect 16025 27013 16037 27016
rect 16071 27044 16083 27047
rect 16209 27047 16267 27053
rect 16209 27044 16221 27047
rect 16071 27016 16221 27044
rect 16071 27013 16083 27016
rect 16025 27007 16083 27013
rect 16209 27013 16221 27016
rect 16255 27013 16267 27047
rect 16209 27007 16267 27013
rect 13173 26979 13231 26985
rect 13173 26945 13185 26979
rect 13219 26976 13231 26979
rect 13538 26976 13544 26988
rect 13219 26948 13544 26976
rect 13219 26945 13231 26948
rect 13173 26939 13231 26945
rect 13538 26936 13544 26948
rect 13596 26936 13602 26988
rect 15565 26979 15623 26985
rect 15565 26945 15577 26979
rect 15611 26976 15623 26979
rect 16574 26976 16580 26988
rect 15611 26948 16580 26976
rect 15611 26945 15623 26948
rect 15565 26939 15623 26945
rect 16574 26936 16580 26948
rect 16632 26936 16638 26988
rect 17865 26979 17923 26985
rect 17865 26945 17877 26979
rect 17911 26976 17923 26979
rect 18325 26979 18383 26985
rect 18325 26976 18337 26979
rect 17911 26948 18337 26976
rect 17911 26945 17923 26948
rect 17865 26939 17923 26945
rect 18325 26945 18337 26948
rect 18371 26976 18383 26979
rect 18414 26976 18420 26988
rect 18371 26948 18420 26976
rect 18371 26945 18383 26948
rect 18325 26939 18383 26945
rect 18414 26936 18420 26948
rect 18472 26936 18478 26988
rect 11054 26908 11060 26920
rect 10367 26880 11060 26908
rect 10367 26877 10379 26880
rect 10321 26871 10379 26877
rect 4663 26812 5948 26840
rect 4663 26809 4675 26812
rect 4617 26803 4675 26809
rect 3326 26732 3332 26784
rect 3384 26772 3390 26784
rect 3789 26775 3847 26781
rect 3789 26772 3801 26775
rect 3384 26744 3801 26772
rect 3384 26732 3390 26744
rect 3789 26741 3801 26744
rect 3835 26741 3847 26775
rect 9214 26772 9220 26784
rect 9175 26744 9220 26772
rect 3789 26735 3847 26741
rect 9214 26732 9220 26744
rect 9272 26772 9278 26784
rect 9582 26772 9588 26784
rect 9272 26744 9588 26772
rect 9272 26732 9278 26744
rect 9582 26732 9588 26744
rect 9640 26772 9646 26784
rect 10244 26772 10272 26871
rect 11054 26868 11060 26880
rect 11112 26868 11118 26920
rect 12618 26908 12624 26920
rect 12531 26880 12624 26908
rect 12618 26868 12624 26880
rect 12676 26908 12682 26920
rect 13722 26908 13728 26920
rect 12676 26880 13728 26908
rect 12676 26868 12682 26880
rect 13722 26868 13728 26880
rect 13780 26868 13786 26920
rect 13998 26868 14004 26920
rect 14056 26908 14062 26920
rect 14093 26911 14151 26917
rect 14093 26908 14105 26911
rect 14056 26880 14105 26908
rect 14056 26868 14062 26880
rect 14093 26877 14105 26880
rect 14139 26877 14151 26911
rect 14093 26871 14151 26877
rect 14553 26911 14611 26917
rect 14553 26877 14565 26911
rect 14599 26877 14611 26911
rect 15010 26908 15016 26920
rect 14971 26880 15016 26908
rect 14553 26871 14611 26877
rect 12437 26843 12495 26849
rect 12437 26809 12449 26843
rect 12483 26809 12495 26843
rect 12802 26840 12808 26852
rect 12715 26812 12808 26840
rect 12437 26803 12495 26809
rect 11514 26772 11520 26784
rect 9640 26744 10272 26772
rect 11475 26744 11520 26772
rect 9640 26732 9646 26744
rect 11514 26732 11520 26744
rect 11572 26732 11578 26784
rect 11698 26732 11704 26784
rect 11756 26772 11762 26784
rect 12250 26772 12256 26784
rect 11756 26744 12256 26772
rect 11756 26732 11762 26744
rect 12250 26732 12256 26744
rect 12308 26772 12314 26784
rect 12452 26772 12480 26803
rect 12802 26800 12808 26812
rect 12860 26840 12866 26852
rect 13538 26840 13544 26852
rect 12860 26812 13544 26840
rect 12860 26800 12866 26812
rect 13538 26800 13544 26812
rect 13596 26800 13602 26852
rect 13633 26843 13691 26849
rect 13633 26809 13645 26843
rect 13679 26840 13691 26843
rect 14568 26840 14596 26871
rect 15010 26868 15016 26880
rect 15068 26868 15074 26920
rect 15470 26908 15476 26920
rect 15431 26880 15476 26908
rect 15470 26868 15476 26880
rect 15528 26868 15534 26920
rect 16025 26911 16083 26917
rect 16025 26877 16037 26911
rect 16071 26908 16083 26911
rect 16393 26911 16451 26917
rect 16393 26908 16405 26911
rect 16071 26880 16405 26908
rect 16071 26877 16083 26880
rect 16025 26871 16083 26877
rect 16393 26877 16405 26880
rect 16439 26877 16451 26911
rect 16393 26871 16451 26877
rect 16485 26911 16543 26917
rect 16485 26877 16497 26911
rect 16531 26908 16543 26911
rect 17218 26908 17224 26920
rect 16531 26880 17224 26908
rect 16531 26877 16543 26880
rect 16485 26871 16543 26877
rect 15102 26840 15108 26852
rect 13679 26812 15108 26840
rect 13679 26809 13691 26812
rect 13633 26803 13691 26809
rect 15102 26800 15108 26812
rect 15160 26800 15166 26852
rect 12710 26772 12716 26784
rect 12308 26744 12480 26772
rect 12671 26744 12716 26772
rect 12308 26732 12314 26744
rect 12710 26732 12716 26744
rect 12768 26732 12774 26784
rect 14274 26732 14280 26784
rect 14332 26772 14338 26784
rect 16500 26772 16528 26871
rect 17218 26868 17224 26880
rect 17276 26868 17282 26920
rect 18046 26908 18052 26920
rect 17959 26880 18052 26908
rect 18046 26868 18052 26880
rect 18104 26908 18110 26920
rect 18690 26908 18696 26920
rect 18104 26880 18696 26908
rect 18104 26868 18110 26880
rect 18690 26868 18696 26880
rect 18748 26908 18754 26920
rect 19150 26908 19156 26920
rect 18748 26880 19156 26908
rect 18748 26868 18754 26880
rect 19150 26868 19156 26880
rect 19208 26868 19214 26920
rect 16942 26840 16948 26852
rect 16903 26812 16948 26840
rect 16942 26800 16948 26812
rect 17000 26800 17006 26852
rect 14332 26744 16528 26772
rect 14332 26732 14338 26744
rect 1104 26682 28888 26704
rect 1104 26630 10982 26682
rect 11034 26630 11046 26682
rect 11098 26630 11110 26682
rect 11162 26630 11174 26682
rect 11226 26630 20982 26682
rect 21034 26630 21046 26682
rect 21098 26630 21110 26682
rect 21162 26630 21174 26682
rect 21226 26630 28888 26682
rect 1104 26608 28888 26630
rect 6914 26528 6920 26580
rect 6972 26568 6978 26580
rect 7098 26568 7104 26580
rect 6972 26540 7104 26568
rect 6972 26528 6978 26540
rect 7098 26528 7104 26540
rect 7156 26528 7162 26580
rect 8110 26568 8116 26580
rect 8071 26540 8116 26568
rect 8110 26528 8116 26540
rect 8168 26528 8174 26580
rect 8754 26568 8760 26580
rect 8715 26540 8760 26568
rect 8754 26528 8760 26540
rect 8812 26528 8818 26580
rect 9125 26571 9183 26577
rect 9125 26537 9137 26571
rect 9171 26568 9183 26571
rect 9398 26568 9404 26580
rect 9171 26540 9404 26568
rect 9171 26537 9183 26540
rect 9125 26531 9183 26537
rect 9398 26528 9404 26540
rect 9456 26528 9462 26580
rect 11514 26528 11520 26580
rect 11572 26568 11578 26580
rect 11885 26571 11943 26577
rect 11885 26568 11897 26571
rect 11572 26540 11897 26568
rect 11572 26528 11578 26540
rect 11885 26537 11897 26540
rect 11931 26537 11943 26571
rect 11885 26531 11943 26537
rect 12161 26571 12219 26577
rect 12161 26537 12173 26571
rect 12207 26568 12219 26571
rect 12710 26568 12716 26580
rect 12207 26540 12716 26568
rect 12207 26537 12219 26540
rect 12161 26531 12219 26537
rect 3050 26500 3056 26512
rect 3011 26472 3056 26500
rect 3050 26460 3056 26472
rect 3108 26460 3114 26512
rect 8662 26460 8668 26512
rect 8720 26460 8726 26512
rect 9950 26460 9956 26512
rect 10008 26500 10014 26512
rect 11900 26500 11928 26531
rect 12710 26528 12716 26540
rect 12768 26568 12774 26580
rect 13170 26568 13176 26580
rect 12768 26540 13176 26568
rect 12768 26528 12774 26540
rect 13170 26528 13176 26540
rect 13228 26528 13234 26580
rect 13998 26528 14004 26580
rect 14056 26568 14062 26580
rect 14093 26571 14151 26577
rect 14093 26568 14105 26571
rect 14056 26540 14105 26568
rect 14056 26528 14062 26540
rect 14093 26537 14105 26540
rect 14139 26537 14151 26571
rect 14826 26568 14832 26580
rect 14787 26540 14832 26568
rect 14093 26531 14151 26537
rect 14826 26528 14832 26540
rect 14884 26528 14890 26580
rect 16209 26571 16267 26577
rect 16209 26537 16221 26571
rect 16255 26568 16267 26571
rect 16482 26568 16488 26580
rect 16255 26540 16488 26568
rect 16255 26537 16267 26540
rect 16209 26531 16267 26537
rect 16482 26528 16488 26540
rect 16540 26528 16546 26580
rect 16850 26568 16856 26580
rect 16811 26540 16856 26568
rect 16850 26528 16856 26540
rect 16908 26528 16914 26580
rect 16942 26528 16948 26580
rect 17000 26568 17006 26580
rect 18874 26568 18880 26580
rect 17000 26540 18880 26568
rect 17000 26528 17006 26540
rect 18874 26528 18880 26540
rect 18932 26528 18938 26580
rect 12434 26500 12440 26512
rect 10008 26472 10732 26500
rect 11900 26472 12440 26500
rect 10008 26460 10014 26472
rect 1394 26432 1400 26444
rect 1355 26404 1400 26432
rect 1394 26392 1400 26404
rect 1452 26432 1458 26444
rect 2130 26432 2136 26444
rect 1452 26404 2136 26432
rect 1452 26392 1458 26404
rect 2130 26392 2136 26404
rect 2188 26392 2194 26444
rect 4614 26392 4620 26444
rect 4672 26432 4678 26444
rect 5261 26435 5319 26441
rect 5261 26432 5273 26435
rect 4672 26404 5273 26432
rect 4672 26392 4678 26404
rect 5261 26401 5273 26404
rect 5307 26432 5319 26435
rect 5626 26432 5632 26444
rect 5307 26404 5632 26432
rect 5307 26401 5319 26404
rect 5261 26395 5319 26401
rect 5626 26392 5632 26404
rect 5684 26392 5690 26444
rect 8573 26435 8631 26441
rect 8573 26401 8585 26435
rect 8619 26432 8631 26435
rect 8680 26432 8708 26460
rect 10318 26432 10324 26444
rect 8619 26404 8708 26432
rect 10279 26404 10324 26432
rect 8619 26401 8631 26404
rect 8573 26395 8631 26401
rect 10318 26392 10324 26404
rect 10376 26392 10382 26444
rect 10502 26432 10508 26444
rect 10463 26404 10508 26432
rect 10502 26392 10508 26404
rect 10560 26392 10566 26444
rect 10704 26441 10732 26472
rect 12434 26460 12440 26472
rect 12492 26500 12498 26512
rect 12492 26472 13216 26500
rect 12492 26460 12498 26472
rect 10689 26435 10747 26441
rect 10689 26401 10701 26435
rect 10735 26401 10747 26435
rect 10689 26395 10747 26401
rect 12342 26392 12348 26444
rect 12400 26432 12406 26444
rect 12400 26404 12572 26432
rect 12400 26392 12406 26404
rect 1670 26364 1676 26376
rect 1631 26336 1676 26364
rect 1670 26324 1676 26336
rect 1728 26324 1734 26376
rect 5166 26324 5172 26376
rect 5224 26364 5230 26376
rect 5537 26367 5595 26373
rect 5537 26364 5549 26367
rect 5224 26336 5549 26364
rect 5224 26324 5230 26336
rect 5537 26333 5549 26336
rect 5583 26364 5595 26367
rect 7006 26364 7012 26376
rect 5583 26336 7012 26364
rect 5583 26333 5595 26336
rect 5537 26327 5595 26333
rect 7006 26324 7012 26336
rect 7064 26324 7070 26376
rect 7745 26367 7803 26373
rect 7745 26333 7757 26367
rect 7791 26364 7803 26367
rect 8202 26364 8208 26376
rect 7791 26336 8208 26364
rect 7791 26333 7803 26336
rect 7745 26327 7803 26333
rect 8202 26324 8208 26336
rect 8260 26364 8266 26376
rect 8662 26364 8668 26376
rect 8260 26336 8668 26364
rect 8260 26324 8266 26336
rect 8662 26324 8668 26336
rect 8720 26324 8726 26376
rect 9122 26324 9128 26376
rect 9180 26364 9186 26376
rect 9398 26364 9404 26376
rect 9180 26336 9404 26364
rect 9180 26324 9186 26336
rect 9398 26324 9404 26336
rect 9456 26324 9462 26376
rect 9861 26367 9919 26373
rect 9861 26333 9873 26367
rect 9907 26364 9919 26367
rect 10410 26364 10416 26376
rect 9907 26336 10416 26364
rect 9907 26333 9919 26336
rect 9861 26327 9919 26333
rect 10410 26324 10416 26336
rect 10468 26324 10474 26376
rect 3326 26256 3332 26308
rect 3384 26296 3390 26308
rect 5074 26296 5080 26308
rect 3384 26268 5080 26296
rect 3384 26256 3390 26268
rect 5074 26256 5080 26268
rect 5132 26256 5138 26308
rect 7282 26296 7288 26308
rect 7243 26268 7288 26296
rect 7282 26256 7288 26268
rect 7340 26256 7346 26308
rect 10520 26296 10548 26392
rect 10594 26324 10600 26376
rect 10652 26364 10658 26376
rect 11057 26367 11115 26373
rect 11057 26364 11069 26367
rect 10652 26336 11069 26364
rect 10652 26324 10658 26336
rect 11057 26333 11069 26336
rect 11103 26333 11115 26367
rect 11238 26364 11244 26376
rect 11199 26336 11244 26364
rect 11057 26327 11115 26333
rect 11238 26324 11244 26336
rect 11296 26324 11302 26376
rect 11422 26324 11428 26376
rect 11480 26364 11486 26376
rect 12158 26364 12164 26376
rect 11480 26336 12164 26364
rect 11480 26324 11486 26336
rect 12158 26324 12164 26336
rect 12216 26324 12222 26376
rect 12250 26324 12256 26376
rect 12308 26364 12314 26376
rect 12308 26336 12480 26364
rect 12308 26324 12314 26336
rect 9600 26268 10548 26296
rect 9600 26240 9628 26268
rect 11606 26256 11612 26308
rect 11664 26296 11670 26308
rect 11882 26296 11888 26308
rect 11664 26268 11888 26296
rect 11664 26256 11670 26268
rect 11882 26256 11888 26268
rect 11940 26256 11946 26308
rect 4801 26231 4859 26237
rect 4801 26197 4813 26231
rect 4847 26228 4859 26231
rect 5258 26228 5264 26240
rect 4847 26200 5264 26228
rect 4847 26197 4859 26200
rect 4801 26191 4859 26197
rect 5258 26188 5264 26200
rect 5316 26188 5322 26240
rect 5718 26188 5724 26240
rect 5776 26228 5782 26240
rect 6641 26231 6699 26237
rect 6641 26228 6653 26231
rect 5776 26200 6653 26228
rect 5776 26188 5782 26200
rect 6641 26197 6653 26200
rect 6687 26197 6699 26231
rect 6641 26191 6699 26197
rect 8481 26231 8539 26237
rect 8481 26197 8493 26231
rect 8527 26228 8539 26231
rect 9214 26228 9220 26240
rect 8527 26200 9220 26228
rect 8527 26197 8539 26200
rect 8481 26191 8539 26197
rect 9214 26188 9220 26200
rect 9272 26228 9278 26240
rect 9401 26231 9459 26237
rect 9401 26228 9413 26231
rect 9272 26200 9413 26228
rect 9272 26188 9278 26200
rect 9401 26197 9413 26200
rect 9447 26197 9459 26231
rect 9401 26191 9459 26197
rect 9582 26188 9588 26240
rect 9640 26188 9646 26240
rect 10870 26188 10876 26240
rect 10928 26228 10934 26240
rect 12161 26231 12219 26237
rect 12161 26228 12173 26231
rect 10928 26200 12173 26228
rect 10928 26188 10934 26200
rect 12161 26197 12173 26200
rect 12207 26228 12219 26231
rect 12253 26231 12311 26237
rect 12253 26228 12265 26231
rect 12207 26200 12265 26228
rect 12207 26197 12219 26200
rect 12161 26191 12219 26197
rect 12253 26197 12265 26200
rect 12299 26197 12311 26231
rect 12452 26228 12480 26336
rect 12544 26305 12572 26404
rect 12618 26392 12624 26444
rect 12676 26432 12682 26444
rect 13188 26441 13216 26472
rect 13354 26460 13360 26512
rect 13412 26500 13418 26512
rect 13538 26500 13544 26512
rect 13412 26472 13544 26500
rect 13412 26460 13418 26472
rect 13538 26460 13544 26472
rect 13596 26460 13602 26512
rect 15470 26460 15476 26512
rect 15528 26500 15534 26512
rect 15841 26503 15899 26509
rect 15841 26500 15853 26503
rect 15528 26472 15853 26500
rect 15528 26460 15534 26472
rect 15841 26469 15853 26472
rect 15887 26469 15899 26503
rect 15841 26463 15899 26469
rect 17865 26503 17923 26509
rect 17865 26469 17877 26503
rect 17911 26500 17923 26503
rect 17954 26500 17960 26512
rect 17911 26472 17960 26500
rect 17911 26469 17923 26472
rect 17865 26463 17923 26469
rect 17954 26460 17960 26472
rect 18012 26460 18018 26512
rect 18138 26500 18144 26512
rect 18099 26472 18144 26500
rect 18138 26460 18144 26472
rect 18196 26460 18202 26512
rect 18230 26460 18236 26512
rect 18288 26500 18294 26512
rect 18509 26503 18567 26509
rect 18509 26500 18521 26503
rect 18288 26472 18521 26500
rect 18288 26460 18294 26472
rect 18509 26469 18521 26472
rect 18555 26469 18567 26503
rect 18509 26463 18567 26469
rect 13081 26435 13139 26441
rect 13081 26432 13093 26435
rect 12676 26404 13093 26432
rect 12676 26392 12682 26404
rect 13081 26401 13093 26404
rect 13127 26401 13139 26435
rect 13081 26395 13139 26401
rect 13173 26435 13231 26441
rect 13173 26401 13185 26435
rect 13219 26432 13231 26435
rect 13262 26432 13268 26444
rect 13219 26404 13268 26432
rect 13219 26401 13231 26404
rect 13173 26395 13231 26401
rect 13262 26392 13268 26404
rect 13320 26392 13326 26444
rect 13449 26435 13507 26441
rect 13449 26401 13461 26435
rect 13495 26432 13507 26435
rect 13556 26432 13584 26460
rect 13495 26404 13584 26432
rect 15381 26435 15439 26441
rect 13495 26401 13507 26404
rect 13449 26395 13507 26401
rect 15381 26401 15393 26435
rect 15427 26432 15439 26435
rect 15562 26432 15568 26444
rect 15427 26404 15568 26432
rect 15427 26401 15439 26404
rect 15381 26395 15439 26401
rect 15562 26392 15568 26404
rect 15620 26392 15626 26444
rect 16666 26432 16672 26444
rect 15764 26404 16672 26432
rect 13354 26324 13360 26376
rect 13412 26364 13418 26376
rect 13541 26367 13599 26373
rect 13541 26364 13553 26367
rect 13412 26336 13553 26364
rect 13412 26324 13418 26336
rect 13541 26333 13553 26336
rect 13587 26333 13599 26367
rect 13541 26327 13599 26333
rect 15289 26367 15347 26373
rect 15289 26333 15301 26367
rect 15335 26364 15347 26367
rect 15470 26364 15476 26376
rect 15335 26336 15476 26364
rect 15335 26333 15347 26336
rect 15289 26327 15347 26333
rect 15470 26324 15476 26336
rect 15528 26364 15534 26376
rect 15764 26364 15792 26404
rect 16666 26392 16672 26404
rect 16724 26392 16730 26444
rect 17405 26435 17463 26441
rect 17405 26401 17417 26435
rect 17451 26432 17463 26435
rect 17770 26432 17776 26444
rect 17451 26404 17776 26432
rect 17451 26401 17463 26404
rect 17405 26395 17463 26401
rect 17770 26392 17776 26404
rect 17828 26392 17834 26444
rect 15528 26336 15792 26364
rect 15528 26324 15534 26336
rect 15838 26324 15844 26376
rect 15896 26364 15902 26376
rect 16298 26364 16304 26376
rect 15896 26336 16304 26364
rect 15896 26324 15902 26336
rect 16298 26324 16304 26336
rect 16356 26324 16362 26376
rect 17313 26367 17371 26373
rect 17313 26333 17325 26367
rect 17359 26364 17371 26367
rect 17586 26364 17592 26376
rect 17359 26336 17592 26364
rect 17359 26333 17371 26336
rect 17313 26327 17371 26333
rect 17586 26324 17592 26336
rect 17644 26324 17650 26376
rect 12529 26299 12587 26305
rect 12529 26265 12541 26299
rect 12575 26265 12587 26299
rect 12529 26259 12587 26265
rect 16942 26256 16948 26308
rect 17000 26296 17006 26308
rect 17494 26296 17500 26308
rect 17000 26268 17500 26296
rect 17000 26256 17006 26268
rect 17494 26256 17500 26268
rect 17552 26256 17558 26308
rect 12710 26228 12716 26240
rect 12452 26200 12716 26228
rect 12253 26191 12311 26197
rect 12710 26188 12716 26200
rect 12768 26188 12774 26240
rect 14553 26231 14611 26237
rect 14553 26197 14565 26231
rect 14599 26228 14611 26231
rect 15010 26228 15016 26240
rect 14599 26200 15016 26228
rect 14599 26197 14611 26200
rect 14553 26191 14611 26197
rect 15010 26188 15016 26200
rect 15068 26188 15074 26240
rect 16577 26231 16635 26237
rect 16577 26197 16589 26231
rect 16623 26228 16635 26231
rect 16666 26228 16672 26240
rect 16623 26200 16672 26228
rect 16623 26197 16635 26200
rect 16577 26191 16635 26197
rect 16666 26188 16672 26200
rect 16724 26188 16730 26240
rect 25130 26188 25136 26240
rect 25188 26228 25194 26240
rect 25314 26228 25320 26240
rect 25188 26200 25320 26228
rect 25188 26188 25194 26200
rect 25314 26188 25320 26200
rect 25372 26188 25378 26240
rect 1104 26138 28888 26160
rect 1104 26086 5982 26138
rect 6034 26086 6046 26138
rect 6098 26086 6110 26138
rect 6162 26086 6174 26138
rect 6226 26086 15982 26138
rect 16034 26086 16046 26138
rect 16098 26086 16110 26138
rect 16162 26086 16174 26138
rect 16226 26086 25982 26138
rect 26034 26086 26046 26138
rect 26098 26086 26110 26138
rect 26162 26086 26174 26138
rect 26226 26086 28888 26138
rect 1104 26064 28888 26086
rect 1670 26024 1676 26036
rect 1631 25996 1676 26024
rect 1670 25984 1676 25996
rect 1728 25984 1734 26036
rect 2041 26027 2099 26033
rect 2041 25993 2053 26027
rect 2087 26024 2099 26027
rect 2130 26024 2136 26036
rect 2087 25996 2136 26024
rect 2087 25993 2099 25996
rect 2041 25987 2099 25993
rect 2130 25984 2136 25996
rect 2188 25984 2194 26036
rect 6638 26024 6644 26036
rect 6599 25996 6644 26024
rect 6638 25984 6644 25996
rect 6696 25984 6702 26036
rect 7190 26024 7196 26036
rect 7151 25996 7196 26024
rect 7190 25984 7196 25996
rect 7248 25984 7254 26036
rect 8297 26027 8355 26033
rect 8297 25993 8309 26027
rect 8343 26024 8355 26027
rect 8570 26024 8576 26036
rect 8343 25996 8576 26024
rect 8343 25993 8355 25996
rect 8297 25987 8355 25993
rect 8570 25984 8576 25996
rect 8628 25984 8634 26036
rect 10686 26024 10692 26036
rect 10647 25996 10692 26024
rect 10686 25984 10692 25996
rect 10744 26024 10750 26036
rect 10744 25996 10824 26024
rect 10744 25984 10750 25996
rect 9122 25956 9128 25968
rect 8496 25928 9128 25956
rect 8496 25897 8524 25928
rect 9122 25916 9128 25928
rect 9180 25916 9186 25968
rect 10134 25956 10140 25968
rect 10047 25928 10140 25956
rect 10134 25916 10140 25928
rect 10192 25956 10198 25968
rect 10594 25956 10600 25968
rect 10192 25928 10600 25956
rect 10192 25916 10198 25928
rect 10594 25916 10600 25928
rect 10652 25916 10658 25968
rect 10796 25897 10824 25996
rect 11238 25984 11244 26036
rect 11296 26024 11302 26036
rect 11793 26027 11851 26033
rect 11793 26024 11805 26027
rect 11296 25996 11805 26024
rect 11296 25984 11302 25996
rect 11793 25993 11805 25996
rect 11839 26024 11851 26027
rect 13538 26024 13544 26036
rect 11839 25996 13544 26024
rect 11839 25993 11851 25996
rect 11793 25987 11851 25993
rect 13538 25984 13544 25996
rect 13596 26024 13602 26036
rect 14458 26024 14464 26036
rect 13596 25996 14464 26024
rect 13596 25984 13602 25996
rect 14458 25984 14464 25996
rect 14516 26024 14522 26036
rect 15749 26027 15807 26033
rect 15749 26024 15761 26027
rect 14516 25996 15761 26024
rect 14516 25984 14522 25996
rect 15749 25993 15761 25996
rect 15795 25993 15807 26027
rect 17770 26024 17776 26036
rect 17731 25996 17776 26024
rect 15749 25987 15807 25993
rect 11698 25916 11704 25968
rect 11756 25956 11762 25968
rect 12529 25959 12587 25965
rect 12529 25956 12541 25959
rect 11756 25928 12541 25956
rect 11756 25916 11762 25928
rect 12529 25925 12541 25928
rect 12575 25925 12587 25959
rect 12529 25919 12587 25925
rect 14277 25959 14335 25965
rect 14277 25925 14289 25959
rect 14323 25956 14335 25959
rect 14734 25956 14740 25968
rect 14323 25928 14740 25956
rect 14323 25925 14335 25928
rect 14277 25919 14335 25925
rect 14734 25916 14740 25928
rect 14792 25916 14798 25968
rect 4249 25891 4307 25897
rect 4249 25857 4261 25891
rect 4295 25888 4307 25891
rect 8481 25891 8539 25897
rect 4295 25860 5764 25888
rect 4295 25857 4307 25860
rect 4249 25851 4307 25857
rect 5736 25832 5764 25860
rect 8481 25857 8493 25891
rect 8527 25857 8539 25891
rect 8481 25851 8539 25857
rect 10781 25891 10839 25897
rect 10781 25857 10793 25891
rect 10827 25857 10839 25891
rect 10781 25851 10839 25857
rect 11517 25891 11575 25897
rect 11517 25857 11529 25891
rect 11563 25888 11575 25891
rect 11882 25888 11888 25900
rect 11563 25860 11888 25888
rect 11563 25857 11575 25860
rect 11517 25851 11575 25857
rect 11882 25848 11888 25860
rect 11940 25888 11946 25900
rect 12618 25888 12624 25900
rect 11940 25860 12624 25888
rect 11940 25848 11946 25860
rect 12618 25848 12624 25860
rect 12676 25848 12682 25900
rect 13262 25888 13268 25900
rect 13223 25860 13268 25888
rect 13262 25848 13268 25860
rect 13320 25848 13326 25900
rect 13630 25848 13636 25900
rect 13688 25888 13694 25900
rect 13998 25888 14004 25900
rect 13688 25860 14004 25888
rect 13688 25848 13694 25860
rect 13998 25848 14004 25860
rect 14056 25888 14062 25900
rect 14369 25891 14427 25897
rect 14369 25888 14381 25891
rect 14056 25860 14381 25888
rect 14056 25848 14062 25860
rect 14369 25857 14381 25860
rect 14415 25857 14427 25891
rect 15102 25888 15108 25900
rect 15063 25860 15108 25888
rect 14369 25851 14427 25857
rect 15102 25848 15108 25860
rect 15160 25848 15166 25900
rect 15764 25888 15792 25987
rect 17770 25984 17776 25996
rect 17828 25984 17834 26036
rect 18325 26027 18383 26033
rect 18325 25993 18337 26027
rect 18371 26024 18383 26027
rect 18414 26024 18420 26036
rect 18371 25996 18420 26024
rect 18371 25993 18383 25996
rect 18325 25987 18383 25993
rect 18414 25984 18420 25996
rect 18472 25984 18478 26036
rect 18690 26024 18696 26036
rect 18651 25996 18696 26024
rect 18690 25984 18696 25996
rect 18748 25984 18754 26036
rect 16393 25891 16451 25897
rect 16393 25888 16405 25891
rect 15764 25860 16405 25888
rect 16393 25857 16405 25860
rect 16439 25857 16451 25891
rect 16393 25851 16451 25857
rect 4154 25780 4160 25832
rect 4212 25820 4218 25832
rect 4709 25823 4767 25829
rect 4709 25820 4721 25823
rect 4212 25792 4721 25820
rect 4212 25780 4218 25792
rect 4709 25789 4721 25792
rect 4755 25789 4767 25823
rect 5166 25820 5172 25832
rect 5127 25792 5172 25820
rect 4709 25783 4767 25789
rect 5166 25780 5172 25792
rect 5224 25780 5230 25832
rect 5350 25820 5356 25832
rect 5311 25792 5356 25820
rect 5350 25780 5356 25792
rect 5408 25780 5414 25832
rect 5718 25820 5724 25832
rect 5679 25792 5724 25820
rect 5718 25780 5724 25792
rect 5776 25780 5782 25832
rect 5905 25823 5963 25829
rect 5905 25789 5917 25823
rect 5951 25820 5963 25823
rect 6362 25820 6368 25832
rect 5951 25792 6368 25820
rect 5951 25789 5963 25792
rect 5905 25783 5963 25789
rect 3881 25755 3939 25761
rect 3881 25721 3893 25755
rect 3927 25752 3939 25755
rect 5184 25752 5212 25780
rect 3927 25724 5212 25752
rect 3927 25721 3939 25724
rect 3881 25715 3939 25721
rect 4617 25687 4675 25693
rect 4617 25653 4629 25687
rect 4663 25684 4675 25687
rect 5920 25684 5948 25783
rect 6362 25780 6368 25792
rect 6420 25780 6426 25832
rect 7929 25823 7987 25829
rect 7929 25789 7941 25823
rect 7975 25820 7987 25823
rect 8573 25823 8631 25829
rect 8573 25820 8585 25823
rect 7975 25792 8585 25820
rect 7975 25789 7987 25792
rect 7929 25783 7987 25789
rect 8573 25789 8585 25792
rect 8619 25820 8631 25823
rect 9125 25823 9183 25829
rect 9125 25820 9137 25823
rect 8619 25792 9137 25820
rect 8619 25789 8631 25792
rect 8573 25783 8631 25789
rect 9125 25789 9137 25792
rect 9171 25820 9183 25823
rect 9214 25820 9220 25832
rect 9171 25792 9220 25820
rect 9171 25789 9183 25792
rect 9125 25783 9183 25789
rect 9214 25780 9220 25792
rect 9272 25780 9278 25832
rect 9309 25823 9367 25829
rect 9309 25789 9321 25823
rect 9355 25820 9367 25823
rect 12161 25823 12219 25829
rect 12161 25820 12173 25823
rect 9355 25792 12173 25820
rect 9355 25789 9367 25792
rect 9309 25783 9367 25789
rect 12161 25789 12173 25792
rect 12207 25789 12219 25823
rect 12161 25783 12219 25789
rect 7561 25755 7619 25761
rect 7561 25721 7573 25755
rect 7607 25752 7619 25755
rect 9324 25752 9352 25783
rect 7607 25724 9352 25752
rect 7607 25721 7619 25724
rect 7561 25715 7619 25721
rect 10870 25712 10876 25764
rect 10928 25752 10934 25764
rect 11057 25755 11115 25761
rect 11057 25752 11069 25755
rect 10928 25724 11069 25752
rect 10928 25712 10934 25724
rect 11057 25721 11069 25724
rect 11103 25721 11115 25755
rect 11057 25715 11115 25721
rect 11146 25712 11152 25764
rect 11204 25752 11210 25764
rect 12176 25752 12204 25783
rect 12250 25780 12256 25832
rect 12308 25820 12314 25832
rect 12437 25823 12495 25829
rect 12437 25820 12449 25823
rect 12308 25792 12449 25820
rect 12308 25780 12314 25792
rect 12437 25789 12449 25792
rect 12483 25789 12495 25823
rect 12986 25820 12992 25832
rect 12947 25792 12992 25820
rect 12437 25783 12495 25789
rect 12986 25780 12992 25792
rect 13044 25780 13050 25832
rect 16577 25823 16635 25829
rect 16577 25789 16589 25823
rect 16623 25820 16635 25823
rect 16666 25820 16672 25832
rect 16623 25792 16672 25820
rect 16623 25789 16635 25792
rect 16577 25783 16635 25789
rect 16666 25780 16672 25792
rect 16724 25780 16730 25832
rect 16850 25780 16856 25832
rect 16908 25820 16914 25832
rect 16945 25823 17003 25829
rect 16945 25820 16957 25823
rect 16908 25792 16957 25820
rect 16908 25780 16914 25792
rect 16945 25789 16957 25792
rect 16991 25789 17003 25823
rect 16945 25783 17003 25789
rect 17037 25823 17095 25829
rect 17037 25789 17049 25823
rect 17083 25789 17095 25823
rect 17037 25783 17095 25789
rect 13004 25752 13032 25780
rect 11204 25724 11249 25752
rect 12176 25724 13032 25752
rect 13909 25755 13967 25761
rect 11204 25712 11210 25724
rect 13909 25721 13921 25755
rect 13955 25752 13967 25755
rect 14550 25752 14556 25764
rect 13955 25724 14556 25752
rect 13955 25721 13967 25724
rect 13909 25715 13967 25721
rect 14550 25712 14556 25724
rect 14608 25712 14614 25764
rect 14734 25752 14740 25764
rect 14695 25724 14740 25752
rect 14734 25712 14740 25724
rect 14792 25712 14798 25764
rect 16022 25712 16028 25764
rect 16080 25752 16086 25764
rect 17052 25752 17080 25783
rect 17770 25752 17776 25764
rect 16080 25724 17776 25752
rect 16080 25712 16086 25724
rect 17770 25712 17776 25724
rect 17828 25712 17834 25764
rect 4663 25656 5948 25684
rect 4663 25653 4675 25656
rect 4617 25647 4675 25653
rect 8386 25644 8392 25696
rect 8444 25684 8450 25696
rect 9585 25687 9643 25693
rect 9585 25684 9597 25687
rect 8444 25656 9597 25684
rect 8444 25644 8450 25656
rect 9585 25653 9597 25656
rect 9631 25653 9643 25687
rect 9585 25647 9643 25653
rect 10686 25644 10692 25696
rect 10744 25684 10750 25696
rect 10965 25687 11023 25693
rect 10965 25684 10977 25687
rect 10744 25656 10977 25684
rect 10744 25644 10750 25656
rect 10965 25653 10977 25656
rect 11011 25684 11023 25687
rect 11514 25684 11520 25696
rect 11011 25656 11520 25684
rect 11011 25653 11023 25656
rect 10965 25647 11023 25653
rect 11514 25644 11520 25656
rect 11572 25644 11578 25696
rect 14645 25687 14703 25693
rect 14645 25653 14657 25687
rect 14691 25684 14703 25687
rect 14826 25684 14832 25696
rect 14691 25656 14832 25684
rect 14691 25653 14703 25656
rect 14645 25647 14703 25653
rect 14826 25644 14832 25656
rect 14884 25644 14890 25696
rect 15470 25684 15476 25696
rect 15431 25656 15476 25684
rect 15470 25644 15476 25656
rect 15528 25644 15534 25696
rect 16206 25684 16212 25696
rect 16167 25656 16212 25684
rect 16206 25644 16212 25656
rect 16264 25644 16270 25696
rect 16298 25644 16304 25696
rect 16356 25684 16362 25696
rect 16758 25684 16764 25696
rect 16356 25656 16764 25684
rect 16356 25644 16362 25656
rect 16758 25644 16764 25656
rect 16816 25644 16822 25696
rect 17497 25687 17555 25693
rect 17497 25653 17509 25687
rect 17543 25684 17555 25687
rect 17586 25684 17592 25696
rect 17543 25656 17592 25684
rect 17543 25653 17555 25656
rect 17497 25647 17555 25653
rect 17586 25644 17592 25656
rect 17644 25684 17650 25696
rect 18230 25684 18236 25696
rect 17644 25656 18236 25684
rect 17644 25644 17650 25656
rect 18230 25644 18236 25656
rect 18288 25644 18294 25696
rect 1104 25594 28888 25616
rect 1104 25542 10982 25594
rect 11034 25542 11046 25594
rect 11098 25542 11110 25594
rect 11162 25542 11174 25594
rect 11226 25542 20982 25594
rect 21034 25542 21046 25594
rect 21098 25542 21110 25594
rect 21162 25542 21174 25594
rect 21226 25542 28888 25594
rect 1104 25520 28888 25542
rect 1670 25480 1676 25492
rect 1631 25452 1676 25480
rect 1670 25440 1676 25452
rect 1728 25440 1734 25492
rect 5626 25480 5632 25492
rect 5587 25452 5632 25480
rect 5626 25440 5632 25452
rect 5684 25440 5690 25492
rect 7009 25483 7067 25489
rect 7009 25449 7021 25483
rect 7055 25480 7067 25483
rect 7098 25480 7104 25492
rect 7055 25452 7104 25480
rect 7055 25449 7067 25452
rect 7009 25443 7067 25449
rect 7098 25440 7104 25452
rect 7156 25440 7162 25492
rect 9122 25480 9128 25492
rect 9083 25452 9128 25480
rect 9122 25440 9128 25452
rect 9180 25440 9186 25492
rect 9493 25483 9551 25489
rect 9493 25449 9505 25483
rect 9539 25480 9551 25483
rect 9582 25480 9588 25492
rect 9539 25452 9588 25480
rect 9539 25449 9551 25452
rect 9493 25443 9551 25449
rect 9582 25440 9588 25452
rect 9640 25440 9646 25492
rect 9950 25480 9956 25492
rect 9911 25452 9956 25480
rect 9950 25440 9956 25452
rect 10008 25480 10014 25492
rect 10686 25480 10692 25492
rect 10008 25452 10692 25480
rect 10008 25440 10014 25452
rect 10686 25440 10692 25452
rect 10744 25440 10750 25492
rect 10870 25480 10876 25492
rect 10831 25452 10876 25480
rect 10870 25440 10876 25452
rect 10928 25440 10934 25492
rect 11241 25483 11299 25489
rect 11241 25449 11253 25483
rect 11287 25480 11299 25483
rect 11330 25480 11336 25492
rect 11287 25452 11336 25480
rect 11287 25449 11299 25452
rect 11241 25443 11299 25449
rect 11330 25440 11336 25452
rect 11388 25440 11394 25492
rect 12250 25440 12256 25492
rect 12308 25480 12314 25492
rect 12897 25483 12955 25489
rect 12897 25480 12909 25483
rect 12308 25452 12909 25480
rect 12308 25440 12314 25452
rect 12897 25449 12909 25452
rect 12943 25449 12955 25483
rect 14918 25480 14924 25492
rect 12897 25443 12955 25449
rect 13464 25452 14924 25480
rect 1762 25412 1768 25424
rect 1412 25384 1768 25412
rect 1412 25356 1440 25384
rect 1762 25372 1768 25384
rect 1820 25372 1826 25424
rect 1394 25344 1400 25356
rect 1355 25316 1400 25344
rect 1394 25304 1400 25316
rect 1452 25304 1458 25356
rect 1581 25347 1639 25353
rect 1581 25313 1593 25347
rect 1627 25344 1639 25347
rect 1946 25344 1952 25356
rect 1627 25316 1952 25344
rect 1627 25313 1639 25316
rect 1581 25307 1639 25313
rect 1946 25304 1952 25316
rect 2004 25304 2010 25356
rect 7116 25353 7144 25440
rect 13464 25421 13492 25452
rect 14918 25440 14924 25452
rect 14976 25440 14982 25492
rect 15562 25480 15568 25492
rect 15523 25452 15568 25480
rect 15562 25440 15568 25452
rect 15620 25440 15626 25492
rect 16022 25480 16028 25492
rect 15983 25452 16028 25480
rect 16022 25440 16028 25452
rect 16080 25440 16086 25492
rect 13449 25415 13507 25421
rect 10888 25384 12848 25412
rect 10888 25356 10916 25384
rect 7101 25347 7159 25353
rect 7101 25313 7113 25347
rect 7147 25313 7159 25347
rect 7101 25307 7159 25313
rect 9306 25304 9312 25356
rect 9364 25344 9370 25356
rect 9582 25344 9588 25356
rect 9364 25316 9588 25344
rect 9364 25304 9370 25316
rect 9582 25304 9588 25316
rect 9640 25304 9646 25356
rect 10042 25344 10048 25356
rect 9876 25316 10048 25344
rect 9876 25288 9904 25316
rect 10042 25304 10048 25316
rect 10100 25304 10106 25356
rect 10137 25347 10195 25353
rect 10137 25313 10149 25347
rect 10183 25344 10195 25347
rect 10502 25344 10508 25356
rect 10183 25316 10508 25344
rect 10183 25313 10195 25316
rect 10137 25307 10195 25313
rect 10502 25304 10508 25316
rect 10560 25304 10566 25356
rect 10870 25304 10876 25356
rect 10928 25304 10934 25356
rect 11698 25344 11704 25356
rect 11659 25316 11704 25344
rect 11698 25304 11704 25316
rect 11756 25304 11762 25356
rect 11900 25353 11928 25384
rect 11885 25347 11943 25353
rect 11885 25313 11897 25347
rect 11931 25313 11943 25347
rect 12066 25344 12072 25356
rect 12027 25316 12072 25344
rect 11885 25307 11943 25313
rect 12066 25304 12072 25316
rect 12124 25304 12130 25356
rect 12250 25344 12256 25356
rect 12211 25316 12256 25344
rect 12250 25304 12256 25316
rect 12308 25304 12314 25356
rect 12621 25347 12679 25353
rect 12621 25313 12633 25347
rect 12667 25344 12679 25347
rect 12710 25344 12716 25356
rect 12667 25316 12716 25344
rect 12667 25313 12679 25316
rect 12621 25307 12679 25313
rect 12710 25304 12716 25316
rect 12768 25304 12774 25356
rect 12820 25344 12848 25384
rect 13449 25381 13461 25415
rect 13495 25381 13507 25415
rect 13449 25375 13507 25381
rect 13998 25372 14004 25424
rect 14056 25412 14062 25424
rect 14461 25415 14519 25421
rect 14461 25412 14473 25415
rect 14056 25384 14473 25412
rect 14056 25372 14062 25384
rect 14461 25381 14473 25384
rect 14507 25381 14519 25415
rect 14461 25375 14519 25381
rect 16117 25347 16175 25353
rect 12820 25316 13952 25344
rect 7377 25279 7435 25285
rect 7377 25245 7389 25279
rect 7423 25276 7435 25279
rect 8386 25276 8392 25288
rect 7423 25248 8392 25276
rect 7423 25245 7435 25248
rect 7377 25239 7435 25245
rect 8386 25236 8392 25248
rect 8444 25236 8450 25288
rect 9858 25236 9864 25288
rect 9916 25236 9922 25288
rect 13814 25276 13820 25288
rect 13775 25248 13820 25276
rect 13814 25236 13820 25248
rect 13872 25236 13878 25288
rect 13924 25285 13952 25316
rect 16117 25313 16129 25347
rect 16163 25344 16175 25347
rect 16758 25344 16764 25356
rect 16163 25316 16764 25344
rect 16163 25313 16175 25316
rect 16117 25307 16175 25313
rect 16758 25304 16764 25316
rect 16816 25304 16822 25356
rect 13909 25279 13967 25285
rect 13909 25245 13921 25279
rect 13955 25245 13967 25279
rect 16390 25276 16396 25288
rect 16351 25248 16396 25276
rect 13909 25239 13967 25245
rect 16390 25236 16396 25248
rect 16448 25236 16454 25288
rect 5166 25168 5172 25220
rect 5224 25208 5230 25220
rect 5261 25211 5319 25217
rect 5261 25208 5273 25211
rect 5224 25180 5273 25208
rect 5224 25168 5230 25180
rect 5261 25177 5273 25180
rect 5307 25177 5319 25211
rect 5261 25171 5319 25177
rect 8846 25168 8852 25220
rect 8904 25208 8910 25220
rect 13262 25208 13268 25220
rect 8904 25180 13268 25208
rect 8904 25168 8910 25180
rect 13262 25168 13268 25180
rect 13320 25168 13326 25220
rect 4801 25143 4859 25149
rect 4801 25109 4813 25143
rect 4847 25140 4859 25143
rect 5350 25140 5356 25152
rect 4847 25112 5356 25140
rect 4847 25109 4859 25112
rect 4801 25103 4859 25109
rect 5350 25100 5356 25112
rect 5408 25140 5414 25152
rect 6638 25140 6644 25152
rect 5408 25112 6644 25140
rect 5408 25100 5414 25112
rect 6638 25100 6644 25112
rect 6696 25100 6702 25152
rect 8294 25100 8300 25152
rect 8352 25140 8358 25152
rect 8481 25143 8539 25149
rect 8481 25140 8493 25143
rect 8352 25112 8493 25140
rect 8352 25100 8358 25112
rect 8481 25109 8493 25112
rect 8527 25109 8539 25143
rect 8481 25103 8539 25109
rect 10321 25143 10379 25149
rect 10321 25109 10333 25143
rect 10367 25140 10379 25143
rect 10594 25140 10600 25152
rect 10367 25112 10600 25140
rect 10367 25109 10379 25112
rect 10321 25103 10379 25109
rect 10594 25100 10600 25112
rect 10652 25100 10658 25152
rect 11514 25100 11520 25152
rect 11572 25140 11578 25152
rect 11974 25140 11980 25152
rect 11572 25112 11980 25140
rect 11572 25100 11578 25112
rect 11974 25100 11980 25112
rect 12032 25100 12038 25152
rect 13354 25140 13360 25152
rect 13315 25112 13360 25140
rect 13354 25100 13360 25112
rect 13412 25100 13418 25152
rect 13538 25100 13544 25152
rect 13596 25149 13602 25152
rect 13596 25143 13645 25149
rect 13596 25109 13599 25143
rect 13633 25109 13645 25143
rect 13722 25140 13728 25152
rect 13683 25112 13728 25140
rect 13596 25103 13645 25109
rect 13596 25100 13602 25103
rect 13722 25100 13728 25112
rect 13780 25100 13786 25152
rect 16574 25100 16580 25152
rect 16632 25140 16638 25152
rect 16850 25140 16856 25152
rect 16632 25112 16856 25140
rect 16632 25100 16638 25112
rect 16850 25100 16856 25112
rect 16908 25140 16914 25152
rect 17497 25143 17555 25149
rect 17497 25140 17509 25143
rect 16908 25112 17509 25140
rect 16908 25100 16914 25112
rect 17497 25109 17509 25112
rect 17543 25109 17555 25143
rect 17497 25103 17555 25109
rect 1104 25050 28888 25072
rect 1104 24998 5982 25050
rect 6034 24998 6046 25050
rect 6098 24998 6110 25050
rect 6162 24998 6174 25050
rect 6226 24998 15982 25050
rect 16034 24998 16046 25050
rect 16098 24998 16110 25050
rect 16162 24998 16174 25050
rect 16226 24998 25982 25050
rect 26034 24998 26046 25050
rect 26098 24998 26110 25050
rect 26162 24998 26174 25050
rect 26226 24998 28888 25050
rect 1104 24976 28888 24998
rect 10502 24896 10508 24948
rect 10560 24936 10566 24948
rect 10781 24939 10839 24945
rect 10781 24936 10793 24939
rect 10560 24908 10793 24936
rect 10560 24896 10566 24908
rect 10781 24905 10793 24908
rect 10827 24905 10839 24939
rect 11882 24936 11888 24948
rect 11843 24908 11888 24936
rect 10781 24899 10839 24905
rect 11882 24896 11888 24908
rect 11940 24896 11946 24948
rect 14458 24896 14464 24948
rect 14516 24936 14522 24948
rect 16209 24939 16267 24945
rect 16209 24936 16221 24939
rect 14516 24908 16221 24936
rect 14516 24896 14522 24908
rect 16209 24905 16221 24908
rect 16255 24905 16267 24939
rect 16574 24936 16580 24948
rect 16535 24908 16580 24936
rect 16209 24899 16267 24905
rect 16574 24896 16580 24908
rect 16632 24896 16638 24948
rect 16758 24896 16764 24948
rect 16816 24936 16822 24948
rect 17313 24939 17371 24945
rect 17313 24936 17325 24939
rect 16816 24908 17325 24936
rect 16816 24896 16822 24908
rect 17313 24905 17325 24908
rect 17359 24936 17371 24939
rect 17681 24939 17739 24945
rect 17681 24936 17693 24939
rect 17359 24908 17693 24936
rect 17359 24905 17371 24908
rect 17313 24899 17371 24905
rect 17681 24905 17693 24908
rect 17727 24936 17739 24939
rect 18138 24936 18144 24948
rect 17727 24908 18144 24936
rect 17727 24905 17739 24908
rect 17681 24899 17739 24905
rect 18138 24896 18144 24908
rect 18196 24936 18202 24948
rect 18690 24936 18696 24948
rect 18196 24908 18696 24936
rect 18196 24896 18202 24908
rect 18690 24896 18696 24908
rect 18748 24896 18754 24948
rect 9125 24871 9183 24877
rect 9125 24837 9137 24871
rect 9171 24868 9183 24871
rect 9214 24868 9220 24880
rect 9171 24840 9220 24868
rect 9171 24837 9183 24840
rect 9125 24831 9183 24837
rect 9214 24828 9220 24840
rect 9272 24868 9278 24880
rect 9272 24840 10640 24868
rect 9272 24828 9278 24840
rect 10612 24812 10640 24840
rect 11974 24828 11980 24880
rect 12032 24868 12038 24880
rect 14734 24868 14740 24880
rect 12032 24840 14740 24868
rect 12032 24828 12038 24840
rect 14734 24828 14740 24840
rect 14792 24828 14798 24880
rect 6641 24803 6699 24809
rect 6641 24769 6653 24803
rect 6687 24800 6699 24803
rect 6687 24772 8064 24800
rect 6687 24769 6699 24772
rect 6641 24763 6699 24769
rect 2682 24692 2688 24744
rect 2740 24732 2746 24744
rect 8036 24741 8064 24772
rect 8110 24760 8116 24812
rect 8168 24800 8174 24812
rect 9677 24803 9735 24809
rect 8168 24772 8213 24800
rect 8168 24760 8174 24772
rect 9677 24769 9689 24803
rect 9723 24800 9735 24803
rect 9766 24800 9772 24812
rect 9723 24772 9772 24800
rect 9723 24769 9735 24772
rect 9677 24763 9735 24769
rect 9766 24760 9772 24772
rect 9824 24760 9830 24812
rect 10594 24800 10600 24812
rect 10555 24772 10600 24800
rect 10594 24760 10600 24772
rect 10652 24760 10658 24812
rect 12253 24803 12311 24809
rect 12253 24769 12265 24803
rect 12299 24800 12311 24803
rect 13354 24800 13360 24812
rect 12299 24772 13360 24800
rect 12299 24769 12311 24772
rect 12253 24763 12311 24769
rect 13354 24760 13360 24772
rect 13412 24800 13418 24812
rect 14277 24803 14335 24809
rect 14277 24800 14289 24803
rect 13412 24772 14289 24800
rect 13412 24760 13418 24772
rect 14277 24769 14289 24772
rect 14323 24769 14335 24803
rect 14277 24763 14335 24769
rect 7377 24735 7435 24741
rect 7377 24732 7389 24735
rect 2740 24704 7389 24732
rect 2740 24692 2746 24704
rect 7377 24701 7389 24704
rect 7423 24701 7435 24735
rect 7377 24695 7435 24701
rect 8021 24735 8079 24741
rect 8021 24701 8033 24735
rect 8067 24732 8079 24735
rect 8202 24732 8208 24744
rect 8067 24704 8208 24732
rect 8067 24701 8079 24704
rect 8021 24695 8079 24701
rect 8202 24692 8208 24704
rect 8260 24692 8266 24744
rect 8386 24732 8392 24744
rect 8347 24704 8392 24732
rect 8386 24692 8392 24704
rect 8444 24692 8450 24744
rect 8573 24735 8631 24741
rect 8573 24701 8585 24735
rect 8619 24732 8631 24735
rect 9030 24732 9036 24744
rect 8619 24704 9036 24732
rect 8619 24701 8631 24704
rect 8573 24695 8631 24701
rect 9030 24692 9036 24704
rect 9088 24692 9094 24744
rect 9493 24735 9551 24741
rect 9493 24701 9505 24735
rect 9539 24732 9551 24735
rect 10134 24732 10140 24744
rect 9539 24704 10140 24732
rect 9539 24701 9551 24704
rect 9493 24695 9551 24701
rect 10134 24692 10140 24704
rect 10192 24732 10198 24744
rect 10505 24735 10563 24741
rect 10505 24732 10517 24735
rect 10192 24704 10517 24732
rect 10192 24692 10198 24704
rect 10505 24701 10517 24704
rect 10551 24701 10563 24735
rect 10505 24695 10563 24701
rect 11425 24735 11483 24741
rect 11425 24701 11437 24735
rect 11471 24732 11483 24735
rect 12710 24732 12716 24744
rect 11471 24704 12716 24732
rect 11471 24701 11483 24704
rect 11425 24695 11483 24701
rect 12710 24692 12716 24704
rect 12768 24692 12774 24744
rect 12894 24732 12900 24744
rect 12855 24704 12900 24732
rect 12894 24692 12900 24704
rect 12952 24692 12958 24744
rect 13262 24732 13268 24744
rect 13223 24704 13268 24732
rect 13262 24692 13268 24704
rect 13320 24692 13326 24744
rect 14185 24735 14243 24741
rect 14185 24701 14197 24735
rect 14231 24732 14243 24735
rect 14458 24732 14464 24744
rect 14231 24704 14464 24732
rect 14231 24701 14243 24704
rect 14185 24695 14243 24701
rect 14458 24692 14464 24704
rect 14516 24732 14522 24744
rect 14921 24735 14979 24741
rect 14921 24732 14933 24735
rect 14516 24704 14933 24732
rect 14516 24692 14522 24704
rect 14921 24701 14933 24704
rect 14967 24732 14979 24735
rect 15286 24732 15292 24744
rect 14967 24704 15292 24732
rect 14967 24701 14979 24704
rect 14921 24695 14979 24701
rect 15286 24692 15292 24704
rect 15344 24692 15350 24744
rect 16025 24735 16083 24741
rect 16025 24701 16037 24735
rect 16071 24732 16083 24735
rect 16390 24732 16396 24744
rect 16071 24704 16396 24732
rect 16071 24701 16083 24704
rect 16025 24695 16083 24701
rect 16390 24692 16396 24704
rect 16448 24732 16454 24744
rect 18046 24732 18052 24744
rect 16448 24704 16896 24732
rect 18007 24704 18052 24732
rect 16448 24692 16454 24704
rect 1394 24624 1400 24676
rect 1452 24664 1458 24676
rect 1673 24667 1731 24673
rect 1673 24664 1685 24667
rect 1452 24636 1685 24664
rect 1452 24624 1458 24636
rect 1673 24633 1685 24636
rect 1719 24664 1731 24667
rect 2958 24664 2964 24676
rect 1719 24636 2964 24664
rect 1719 24633 1731 24636
rect 1673 24627 1731 24633
rect 2958 24624 2964 24636
rect 3016 24624 3022 24676
rect 7282 24664 7288 24676
rect 7195 24636 7288 24664
rect 7282 24624 7288 24636
rect 7340 24664 7346 24676
rect 8110 24664 8116 24676
rect 7340 24636 8116 24664
rect 7340 24624 7346 24636
rect 8110 24624 8116 24636
rect 8168 24624 8174 24676
rect 9769 24667 9827 24673
rect 9769 24633 9781 24667
rect 9815 24664 9827 24667
rect 9815 24636 10548 24664
rect 9815 24633 9827 24636
rect 9769 24627 9827 24633
rect 10520 24608 10548 24636
rect 12434 24624 12440 24676
rect 12492 24664 12498 24676
rect 13280 24664 13308 24692
rect 15657 24667 15715 24673
rect 15657 24664 15669 24667
rect 12492 24636 12537 24664
rect 13280 24636 15669 24664
rect 12492 24624 12498 24636
rect 15657 24633 15669 24636
rect 15703 24633 15715 24667
rect 15657 24627 15715 24633
rect 16868 24608 16896 24704
rect 18046 24692 18052 24704
rect 18104 24732 18110 24744
rect 18509 24735 18567 24741
rect 18509 24732 18521 24735
rect 18104 24704 18521 24732
rect 18104 24692 18110 24704
rect 18509 24701 18521 24704
rect 18555 24701 18567 24735
rect 18509 24695 18567 24701
rect 1946 24596 1952 24608
rect 1907 24568 1952 24596
rect 1946 24556 1952 24568
rect 2004 24556 2010 24608
rect 6273 24599 6331 24605
rect 6273 24565 6285 24599
rect 6319 24596 6331 24599
rect 8386 24596 8392 24608
rect 6319 24568 8392 24596
rect 6319 24565 6331 24568
rect 6273 24559 6331 24565
rect 8386 24556 8392 24568
rect 8444 24556 8450 24608
rect 9950 24556 9956 24608
rect 10008 24596 10014 24608
rect 10134 24596 10140 24608
rect 10008 24568 10140 24596
rect 10008 24556 10014 24568
rect 10134 24556 10140 24568
rect 10192 24556 10198 24608
rect 10502 24556 10508 24608
rect 10560 24556 10566 24608
rect 10781 24599 10839 24605
rect 10781 24565 10793 24599
rect 10827 24596 10839 24599
rect 11057 24599 11115 24605
rect 11057 24596 11069 24599
rect 10827 24568 11069 24596
rect 10827 24565 10839 24568
rect 10781 24559 10839 24565
rect 11057 24565 11069 24568
rect 11103 24596 11115 24599
rect 11606 24596 11612 24608
rect 11103 24568 11612 24596
rect 11103 24565 11115 24568
rect 11057 24559 11115 24565
rect 11606 24556 11612 24568
rect 11664 24556 11670 24608
rect 12986 24556 12992 24608
rect 13044 24596 13050 24608
rect 13725 24599 13783 24605
rect 13725 24596 13737 24599
rect 13044 24568 13737 24596
rect 13044 24556 13050 24568
rect 13725 24565 13737 24568
rect 13771 24596 13783 24599
rect 13814 24596 13820 24608
rect 13771 24568 13820 24596
rect 13771 24565 13783 24568
rect 13725 24559 13783 24565
rect 13814 24556 13820 24568
rect 13872 24556 13878 24608
rect 15381 24599 15439 24605
rect 15381 24565 15393 24599
rect 15427 24596 15439 24599
rect 15562 24596 15568 24608
rect 15427 24568 15568 24596
rect 15427 24565 15439 24568
rect 15381 24559 15439 24565
rect 15562 24556 15568 24568
rect 15620 24556 15626 24608
rect 16850 24596 16856 24608
rect 16811 24568 16856 24596
rect 16850 24556 16856 24568
rect 16908 24556 16914 24608
rect 18230 24596 18236 24608
rect 18191 24568 18236 24596
rect 18230 24556 18236 24568
rect 18288 24556 18294 24608
rect 1104 24506 28888 24528
rect 1104 24454 10982 24506
rect 11034 24454 11046 24506
rect 11098 24454 11110 24506
rect 11162 24454 11174 24506
rect 11226 24454 20982 24506
rect 21034 24454 21046 24506
rect 21098 24454 21110 24506
rect 21162 24454 21174 24506
rect 21226 24454 28888 24506
rect 1104 24432 28888 24454
rect 7098 24392 7104 24404
rect 7059 24364 7104 24392
rect 7098 24352 7104 24364
rect 7156 24352 7162 24404
rect 7837 24395 7895 24401
rect 7837 24361 7849 24395
rect 7883 24392 7895 24395
rect 8386 24392 8392 24404
rect 7883 24364 8392 24392
rect 7883 24361 7895 24364
rect 7837 24355 7895 24361
rect 8386 24352 8392 24364
rect 8444 24352 8450 24404
rect 9766 24352 9772 24404
rect 9824 24392 9830 24404
rect 9861 24395 9919 24401
rect 9861 24392 9873 24395
rect 9824 24364 9873 24392
rect 9824 24352 9830 24364
rect 9861 24361 9873 24364
rect 9907 24361 9919 24395
rect 9861 24355 9919 24361
rect 10505 24395 10563 24401
rect 10505 24361 10517 24395
rect 10551 24392 10563 24395
rect 10870 24392 10876 24404
rect 10551 24364 10876 24392
rect 10551 24361 10563 24364
rect 10505 24355 10563 24361
rect 10870 24352 10876 24364
rect 10928 24352 10934 24404
rect 11241 24395 11299 24401
rect 11241 24361 11253 24395
rect 11287 24392 11299 24395
rect 12250 24392 12256 24404
rect 11287 24364 12256 24392
rect 11287 24361 11299 24364
rect 11241 24355 11299 24361
rect 12250 24352 12256 24364
rect 12308 24352 12314 24404
rect 12526 24392 12532 24404
rect 12487 24364 12532 24392
rect 12526 24352 12532 24364
rect 12584 24352 12590 24404
rect 12710 24352 12716 24404
rect 12768 24392 12774 24404
rect 12805 24395 12863 24401
rect 12805 24392 12817 24395
rect 12768 24364 12817 24392
rect 12768 24352 12774 24364
rect 12805 24361 12817 24364
rect 12851 24361 12863 24395
rect 12805 24355 12863 24361
rect 13814 24352 13820 24404
rect 13872 24392 13878 24404
rect 14366 24392 14372 24404
rect 13872 24364 14372 24392
rect 13872 24352 13878 24364
rect 14366 24352 14372 24364
rect 14424 24352 14430 24404
rect 14918 24392 14924 24404
rect 14879 24364 14924 24392
rect 14918 24352 14924 24364
rect 14976 24352 14982 24404
rect 15473 24395 15531 24401
rect 15473 24392 15485 24395
rect 15212 24364 15485 24392
rect 7469 24327 7527 24333
rect 7469 24293 7481 24327
rect 7515 24324 7527 24327
rect 9030 24324 9036 24336
rect 7515 24296 9036 24324
rect 7515 24293 7527 24296
rect 7469 24287 7527 24293
rect 9030 24284 9036 24296
rect 9088 24284 9094 24336
rect 10226 24284 10232 24336
rect 10284 24284 10290 24336
rect 10962 24284 10968 24336
rect 11020 24324 11026 24336
rect 11885 24327 11943 24333
rect 11885 24324 11897 24327
rect 11020 24296 11897 24324
rect 11020 24284 11026 24296
rect 11885 24293 11897 24296
rect 11931 24324 11943 24327
rect 12894 24324 12900 24336
rect 11931 24296 12900 24324
rect 11931 24293 11943 24296
rect 11885 24287 11943 24293
rect 12894 24284 12900 24296
rect 12952 24284 12958 24336
rect 13630 24324 13636 24336
rect 13004 24296 13636 24324
rect 10244 24256 10272 24284
rect 11422 24256 11428 24268
rect 10244 24228 11100 24256
rect 11383 24228 11428 24256
rect 11072 24188 11100 24228
rect 11422 24216 11428 24228
rect 11480 24216 11486 24268
rect 13004 24265 13032 24296
rect 13630 24284 13636 24296
rect 13688 24284 13694 24336
rect 14550 24284 14556 24336
rect 14608 24324 14614 24336
rect 15102 24324 15108 24336
rect 14608 24296 15108 24324
rect 14608 24284 14614 24296
rect 15102 24284 15108 24296
rect 15160 24324 15166 24336
rect 15212 24324 15240 24364
rect 15473 24361 15485 24364
rect 15519 24392 15531 24395
rect 17037 24395 17095 24401
rect 17037 24392 17049 24395
rect 15519 24364 17049 24392
rect 15519 24361 15531 24364
rect 15473 24355 15531 24361
rect 17037 24361 17049 24364
rect 17083 24361 17095 24395
rect 17037 24355 17095 24361
rect 17494 24352 17500 24404
rect 17552 24392 17558 24404
rect 18049 24395 18107 24401
rect 18049 24392 18061 24395
rect 17552 24364 18061 24392
rect 17552 24352 17558 24364
rect 18049 24361 18061 24364
rect 18095 24361 18107 24395
rect 18049 24355 18107 24361
rect 15160 24296 15240 24324
rect 15160 24284 15166 24296
rect 15286 24284 15292 24336
rect 15344 24324 15350 24336
rect 15565 24327 15623 24333
rect 15565 24324 15577 24327
rect 15344 24296 15577 24324
rect 15344 24284 15350 24296
rect 15565 24293 15577 24296
rect 15611 24293 15623 24327
rect 15565 24287 15623 24293
rect 15657 24327 15715 24333
rect 15657 24293 15669 24327
rect 15703 24324 15715 24327
rect 15703 24296 16436 24324
rect 15703 24293 15715 24296
rect 15657 24287 15715 24293
rect 12989 24259 13047 24265
rect 12989 24225 13001 24259
rect 13035 24225 13047 24259
rect 13170 24256 13176 24268
rect 13131 24228 13176 24256
rect 12989 24219 13047 24225
rect 13170 24216 13176 24228
rect 13228 24216 13234 24268
rect 13262 24216 13268 24268
rect 13320 24256 13326 24268
rect 13541 24259 13599 24265
rect 13541 24256 13553 24259
rect 13320 24228 13553 24256
rect 13320 24216 13326 24228
rect 13541 24225 13553 24228
rect 13587 24225 13599 24259
rect 16298 24256 16304 24268
rect 13541 24219 13599 24225
rect 15304 24228 16304 24256
rect 11330 24188 11336 24200
rect 11072 24160 11336 24188
rect 11330 24148 11336 24160
rect 11388 24148 11394 24200
rect 13722 24148 13728 24200
rect 13780 24188 13786 24200
rect 13998 24188 14004 24200
rect 13780 24160 14004 24188
rect 13780 24148 13786 24160
rect 13998 24148 14004 24160
rect 14056 24148 14062 24200
rect 15304 24197 15332 24228
rect 16298 24216 16304 24228
rect 16356 24216 16362 24268
rect 15289 24191 15347 24197
rect 15289 24157 15301 24191
rect 15335 24157 15347 24191
rect 15289 24151 15347 24157
rect 16025 24191 16083 24197
rect 16025 24157 16037 24191
rect 16071 24157 16083 24191
rect 16025 24151 16083 24157
rect 9493 24123 9551 24129
rect 9493 24089 9505 24123
rect 9539 24120 9551 24123
rect 11790 24120 11796 24132
rect 9539 24092 11796 24120
rect 9539 24089 9551 24092
rect 9493 24083 9551 24089
rect 11790 24080 11796 24092
rect 11848 24080 11854 24132
rect 14274 24080 14280 24132
rect 14332 24120 14338 24132
rect 16040 24120 16068 24151
rect 16408 24129 16436 24296
rect 16853 24259 16911 24265
rect 16853 24225 16865 24259
rect 16899 24256 16911 24259
rect 17865 24259 17923 24265
rect 17865 24256 17877 24259
rect 16899 24228 17877 24256
rect 16899 24225 16911 24228
rect 16853 24219 16911 24225
rect 17865 24225 17877 24228
rect 17911 24256 17923 24259
rect 19058 24256 19064 24268
rect 17911 24228 19064 24256
rect 17911 24225 17923 24228
rect 17865 24219 17923 24225
rect 19058 24216 19064 24228
rect 19116 24216 19122 24268
rect 14332 24092 16068 24120
rect 16393 24123 16451 24129
rect 14332 24080 14338 24092
rect 16393 24089 16405 24123
rect 16439 24120 16451 24123
rect 16761 24123 16819 24129
rect 16761 24120 16773 24123
rect 16439 24092 16773 24120
rect 16439 24089 16451 24092
rect 16393 24083 16451 24089
rect 16761 24089 16773 24092
rect 16807 24120 16819 24123
rect 16850 24120 16856 24132
rect 16807 24092 16856 24120
rect 16807 24089 16819 24092
rect 16761 24083 16819 24089
rect 16850 24080 16856 24092
rect 16908 24120 16914 24132
rect 17954 24120 17960 24132
rect 16908 24092 17960 24120
rect 16908 24080 16914 24092
rect 17954 24080 17960 24092
rect 18012 24080 18018 24132
rect 10870 24052 10876 24064
rect 10831 24024 10876 24052
rect 10870 24012 10876 24024
rect 10928 24012 10934 24064
rect 14185 24055 14243 24061
rect 14185 24021 14197 24055
rect 14231 24052 14243 24055
rect 14366 24052 14372 24064
rect 14231 24024 14372 24052
rect 14231 24021 14243 24024
rect 14185 24015 14243 24021
rect 14366 24012 14372 24024
rect 14424 24012 14430 24064
rect 14553 24055 14611 24061
rect 14553 24021 14565 24055
rect 14599 24052 14611 24055
rect 14918 24052 14924 24064
rect 14599 24024 14924 24052
rect 14599 24021 14611 24024
rect 14553 24015 14611 24021
rect 14918 24012 14924 24024
rect 14976 24012 14982 24064
rect 15470 24012 15476 24064
rect 15528 24052 15534 24064
rect 17494 24052 17500 24064
rect 15528 24024 17500 24052
rect 15528 24012 15534 24024
rect 17494 24012 17500 24024
rect 17552 24012 17558 24064
rect 1104 23962 28888 23984
rect 1104 23910 5982 23962
rect 6034 23910 6046 23962
rect 6098 23910 6110 23962
rect 6162 23910 6174 23962
rect 6226 23910 15982 23962
rect 16034 23910 16046 23962
rect 16098 23910 16110 23962
rect 16162 23910 16174 23962
rect 16226 23910 25982 23962
rect 26034 23910 26046 23962
rect 26098 23910 26110 23962
rect 26162 23910 26174 23962
rect 26226 23910 28888 23962
rect 1104 23888 28888 23910
rect 7098 23848 7104 23860
rect 7059 23820 7104 23848
rect 7098 23808 7104 23820
rect 7156 23808 7162 23860
rect 8570 23848 8576 23860
rect 8531 23820 8576 23848
rect 8570 23808 8576 23820
rect 8628 23808 8634 23860
rect 9674 23808 9680 23860
rect 9732 23848 9738 23860
rect 10318 23848 10324 23860
rect 9732 23820 10324 23848
rect 9732 23808 9738 23820
rect 10318 23808 10324 23820
rect 10376 23808 10382 23860
rect 10689 23851 10747 23857
rect 10689 23817 10701 23851
rect 10735 23848 10747 23851
rect 10962 23848 10968 23860
rect 10735 23820 10968 23848
rect 10735 23817 10747 23820
rect 10689 23811 10747 23817
rect 10962 23808 10968 23820
rect 11020 23808 11026 23860
rect 11422 23808 11428 23860
rect 11480 23848 11486 23860
rect 13357 23851 13415 23857
rect 11480 23820 11836 23848
rect 11480 23808 11486 23820
rect 8588 23644 8616 23808
rect 11057 23783 11115 23789
rect 11057 23749 11069 23783
rect 11103 23780 11115 23783
rect 11698 23780 11704 23792
rect 11103 23752 11704 23780
rect 11103 23749 11115 23752
rect 11057 23743 11115 23749
rect 11698 23740 11704 23752
rect 11756 23740 11762 23792
rect 8757 23647 8815 23653
rect 8757 23644 8769 23647
rect 8588 23616 8769 23644
rect 8757 23613 8769 23616
rect 8803 23613 8815 23647
rect 8757 23607 8815 23613
rect 11425 23647 11483 23653
rect 11425 23613 11437 23647
rect 11471 23644 11483 23647
rect 11808 23644 11836 23820
rect 13357 23817 13369 23851
rect 13403 23848 13415 23851
rect 13630 23848 13636 23860
rect 13403 23820 13636 23848
rect 13403 23817 13415 23820
rect 13357 23811 13415 23817
rect 13630 23808 13636 23820
rect 13688 23848 13694 23860
rect 13998 23848 14004 23860
rect 13688 23820 14004 23848
rect 13688 23808 13694 23820
rect 13998 23808 14004 23820
rect 14056 23808 14062 23860
rect 15841 23851 15899 23857
rect 15841 23848 15853 23851
rect 14108 23820 15853 23848
rect 12250 23740 12256 23792
rect 12308 23780 12314 23792
rect 13170 23780 13176 23792
rect 12308 23752 13176 23780
rect 12308 23740 12314 23752
rect 13170 23740 13176 23752
rect 13228 23740 13234 23792
rect 13538 23740 13544 23792
rect 13596 23780 13602 23792
rect 14108 23780 14136 23820
rect 15841 23817 15853 23820
rect 15887 23848 15899 23851
rect 16298 23848 16304 23860
rect 15887 23820 16304 23848
rect 15887 23817 15899 23820
rect 15841 23811 15899 23817
rect 16298 23808 16304 23820
rect 16356 23808 16362 23860
rect 16390 23808 16396 23860
rect 16448 23848 16454 23860
rect 16945 23851 17003 23857
rect 16945 23848 16957 23851
rect 16448 23820 16957 23848
rect 16448 23808 16454 23820
rect 16945 23817 16957 23820
rect 16991 23848 17003 23851
rect 18325 23851 18383 23857
rect 18325 23848 18337 23851
rect 16991 23820 18337 23848
rect 16991 23817 17003 23820
rect 16945 23811 17003 23817
rect 18325 23817 18337 23820
rect 18371 23848 18383 23851
rect 19058 23848 19064 23860
rect 18371 23820 19064 23848
rect 18371 23817 18383 23820
rect 18325 23811 18383 23817
rect 19058 23808 19064 23820
rect 19116 23808 19122 23860
rect 16482 23780 16488 23792
rect 13596 23752 14136 23780
rect 16443 23752 16488 23780
rect 13596 23740 13602 23752
rect 16482 23740 16488 23752
rect 16540 23740 16546 23792
rect 12986 23712 12992 23724
rect 12947 23684 12992 23712
rect 12986 23672 12992 23684
rect 13044 23672 13050 23724
rect 15286 23672 15292 23724
rect 15344 23712 15350 23724
rect 15344 23684 15424 23712
rect 15344 23672 15350 23684
rect 12253 23647 12311 23653
rect 12253 23644 12265 23647
rect 11471 23616 12265 23644
rect 11471 23613 11483 23616
rect 11425 23607 11483 23613
rect 12253 23613 12265 23616
rect 12299 23613 12311 23647
rect 12253 23607 12311 23613
rect 8570 23536 8576 23588
rect 8628 23576 8634 23588
rect 8665 23579 8723 23585
rect 8665 23576 8677 23579
rect 8628 23548 8677 23576
rect 8628 23536 8634 23548
rect 8665 23545 8677 23548
rect 8711 23545 8723 23579
rect 12268 23576 12296 23607
rect 12342 23604 12348 23656
rect 12400 23644 12406 23656
rect 12437 23647 12495 23653
rect 12437 23644 12449 23647
rect 12400 23616 12449 23644
rect 12400 23604 12406 23616
rect 12437 23613 12449 23616
rect 12483 23613 12495 23647
rect 12437 23607 12495 23613
rect 12529 23647 12587 23653
rect 12529 23613 12541 23647
rect 12575 23644 12587 23647
rect 13909 23647 13967 23653
rect 12575 23613 12613 23644
rect 12529 23607 12613 23613
rect 13909 23613 13921 23647
rect 13955 23644 13967 23647
rect 14274 23644 14280 23656
rect 13955 23616 14280 23644
rect 13955 23613 13967 23616
rect 13909 23607 13967 23613
rect 12585 23576 12613 23607
rect 14274 23604 14280 23616
rect 14332 23604 14338 23656
rect 14366 23604 14372 23656
rect 14424 23644 14430 23656
rect 14645 23647 14703 23653
rect 14645 23644 14657 23647
rect 14424 23616 14657 23644
rect 14424 23604 14430 23616
rect 14645 23613 14657 23616
rect 14691 23613 14703 23647
rect 14826 23644 14832 23656
rect 14787 23616 14832 23644
rect 14645 23607 14703 23613
rect 13446 23576 13452 23588
rect 12268 23548 13452 23576
rect 8665 23539 8723 23545
rect 13446 23536 13452 23548
rect 13504 23536 13510 23588
rect 14660 23576 14688 23607
rect 14826 23604 14832 23616
rect 14884 23604 14890 23656
rect 14918 23604 14924 23656
rect 14976 23644 14982 23656
rect 15197 23647 15255 23653
rect 15197 23644 15209 23647
rect 14976 23616 15209 23644
rect 14976 23604 14982 23616
rect 15197 23613 15209 23616
rect 15243 23613 15255 23647
rect 15197 23607 15255 23613
rect 15286 23576 15292 23588
rect 14660 23548 15292 23576
rect 15286 23536 15292 23548
rect 15344 23536 15350 23588
rect 11698 23468 11704 23520
rect 11756 23508 11762 23520
rect 11793 23511 11851 23517
rect 11793 23508 11805 23511
rect 11756 23480 11805 23508
rect 11756 23468 11762 23480
rect 11793 23477 11805 23480
rect 11839 23508 11851 23511
rect 12250 23508 12256 23520
rect 11839 23480 12256 23508
rect 11839 23477 11851 23480
rect 11793 23471 11851 23477
rect 12250 23468 12256 23480
rect 12308 23468 12314 23520
rect 14277 23511 14335 23517
rect 14277 23477 14289 23511
rect 14323 23508 14335 23511
rect 14642 23508 14648 23520
rect 14323 23480 14648 23508
rect 14323 23477 14335 23480
rect 14277 23471 14335 23477
rect 14642 23468 14648 23480
rect 14700 23468 14706 23520
rect 15396 23508 15424 23684
rect 16298 23644 16304 23656
rect 16259 23616 16304 23644
rect 16298 23604 16304 23616
rect 16356 23644 16362 23656
rect 18230 23644 18236 23656
rect 16356 23616 18236 23644
rect 16356 23604 16362 23616
rect 18230 23604 18236 23616
rect 18288 23604 18294 23656
rect 16209 23511 16267 23517
rect 16209 23508 16221 23511
rect 15396 23480 16221 23508
rect 16209 23477 16221 23480
rect 16255 23508 16267 23511
rect 16850 23508 16856 23520
rect 16255 23480 16856 23508
rect 16255 23477 16267 23480
rect 16209 23471 16267 23477
rect 16850 23468 16856 23480
rect 16908 23508 16914 23520
rect 17218 23508 17224 23520
rect 16908 23480 17224 23508
rect 16908 23468 16914 23480
rect 17218 23468 17224 23480
rect 17276 23468 17282 23520
rect 1104 23418 28888 23440
rect 1104 23366 10982 23418
rect 11034 23366 11046 23418
rect 11098 23366 11110 23418
rect 11162 23366 11174 23418
rect 11226 23366 20982 23418
rect 21034 23366 21046 23418
rect 21098 23366 21110 23418
rect 21162 23366 21174 23418
rect 21226 23366 28888 23418
rect 1104 23344 28888 23366
rect 8478 23264 8484 23316
rect 8536 23304 8542 23316
rect 8757 23307 8815 23313
rect 8757 23304 8769 23307
rect 8536 23276 8769 23304
rect 8536 23264 8542 23276
rect 8757 23273 8769 23276
rect 8803 23273 8815 23307
rect 8757 23267 8815 23273
rect 11330 23264 11336 23316
rect 11388 23304 11394 23316
rect 11425 23307 11483 23313
rect 11425 23304 11437 23307
rect 11388 23276 11437 23304
rect 11388 23264 11394 23276
rect 11425 23273 11437 23276
rect 11471 23273 11483 23307
rect 11425 23267 11483 23273
rect 11514 23264 11520 23316
rect 11572 23304 11578 23316
rect 11885 23307 11943 23313
rect 11885 23304 11897 23307
rect 11572 23276 11897 23304
rect 11572 23264 11578 23276
rect 11885 23273 11897 23276
rect 11931 23273 11943 23307
rect 12066 23304 12072 23316
rect 12027 23276 12072 23304
rect 11885 23267 11943 23273
rect 10137 23239 10195 23245
rect 10137 23205 10149 23239
rect 10183 23236 10195 23239
rect 10778 23236 10784 23248
rect 10183 23208 10784 23236
rect 10183 23205 10195 23208
rect 10137 23199 10195 23205
rect 10778 23196 10784 23208
rect 10836 23196 10842 23248
rect 11900 23236 11928 23267
rect 12066 23264 12072 23276
rect 12124 23264 12130 23316
rect 13906 23264 13912 23316
rect 13964 23304 13970 23316
rect 14366 23304 14372 23316
rect 13964 23276 14372 23304
rect 13964 23264 13970 23276
rect 14366 23264 14372 23276
rect 14424 23264 14430 23316
rect 14461 23307 14519 23313
rect 14461 23273 14473 23307
rect 14507 23304 14519 23307
rect 14826 23304 14832 23316
rect 14507 23276 14832 23304
rect 14507 23273 14519 23276
rect 14461 23267 14519 23273
rect 14568 23248 14596 23276
rect 14826 23264 14832 23276
rect 14884 23264 14890 23316
rect 15102 23304 15108 23316
rect 15063 23276 15108 23304
rect 15102 23264 15108 23276
rect 15160 23264 15166 23316
rect 15286 23264 15292 23316
rect 15344 23304 15350 23316
rect 18138 23304 18144 23316
rect 15344 23276 16068 23304
rect 18099 23276 18144 23304
rect 15344 23264 15350 23276
rect 12342 23236 12348 23248
rect 11900 23208 12348 23236
rect 12084 23180 12112 23208
rect 12342 23196 12348 23208
rect 12400 23196 12406 23248
rect 14550 23196 14556 23248
rect 14608 23196 14614 23248
rect 15120 23236 15148 23264
rect 15473 23239 15531 23245
rect 15473 23236 15485 23239
rect 15120 23208 15485 23236
rect 15473 23205 15485 23208
rect 15519 23205 15531 23239
rect 15654 23236 15660 23248
rect 15615 23208 15660 23236
rect 15473 23199 15531 23205
rect 15654 23196 15660 23208
rect 15712 23196 15718 23248
rect 16040 23245 16068 23276
rect 18138 23264 18144 23276
rect 18196 23264 18202 23316
rect 16025 23239 16083 23245
rect 16025 23205 16037 23239
rect 16071 23205 16083 23239
rect 16025 23199 16083 23205
rect 6638 23128 6644 23180
rect 6696 23168 6702 23180
rect 6822 23168 6828 23180
rect 6696 23140 6828 23168
rect 6696 23128 6702 23140
rect 6822 23128 6828 23140
rect 6880 23128 6886 23180
rect 7190 23168 7196 23180
rect 7151 23140 7196 23168
rect 7190 23128 7196 23140
rect 7248 23128 7254 23180
rect 7377 23171 7435 23177
rect 7377 23137 7389 23171
rect 7423 23137 7435 23171
rect 8570 23168 8576 23180
rect 8531 23140 8576 23168
rect 7377 23131 7435 23137
rect 5534 23060 5540 23112
rect 5592 23100 5598 23112
rect 6181 23103 6239 23109
rect 6181 23100 6193 23103
rect 5592 23072 6193 23100
rect 5592 23060 5598 23072
rect 6181 23069 6193 23072
rect 6227 23069 6239 23103
rect 6914 23100 6920 23112
rect 6827 23072 6920 23100
rect 6181 23063 6239 23069
rect 6914 23060 6920 23072
rect 6972 23100 6978 23112
rect 7282 23100 7288 23112
rect 6972 23072 7288 23100
rect 6972 23060 6978 23072
rect 7282 23060 7288 23072
rect 7340 23060 7346 23112
rect 7392 23100 7420 23131
rect 8570 23128 8576 23140
rect 8628 23128 8634 23180
rect 10962 23168 10968 23180
rect 10923 23140 10968 23168
rect 10962 23128 10968 23140
rect 11020 23128 11026 23180
rect 11514 23168 11520 23180
rect 11072 23140 11520 23168
rect 9490 23100 9496 23112
rect 7392 23072 9496 23100
rect 6270 22992 6276 23044
rect 6328 23032 6334 23044
rect 7392 23032 7420 23072
rect 9490 23060 9496 23072
rect 9548 23060 9554 23112
rect 9950 23060 9956 23112
rect 10008 23100 10014 23112
rect 10689 23103 10747 23109
rect 10689 23100 10701 23103
rect 10008 23072 10701 23100
rect 10008 23060 10014 23072
rect 10689 23069 10701 23072
rect 10735 23100 10747 23103
rect 11072 23100 11100 23140
rect 11514 23128 11520 23140
rect 11572 23168 11578 23180
rect 11977 23171 12035 23177
rect 11977 23168 11989 23171
rect 11572 23140 11989 23168
rect 11572 23128 11578 23140
rect 11977 23137 11989 23140
rect 12023 23137 12035 23171
rect 11977 23131 12035 23137
rect 12066 23128 12072 23180
rect 12124 23128 12130 23180
rect 12526 23128 12532 23180
rect 12584 23168 12590 23180
rect 12805 23171 12863 23177
rect 12805 23168 12817 23171
rect 12584 23140 12817 23168
rect 12584 23128 12590 23140
rect 12805 23137 12817 23140
rect 12851 23137 12863 23171
rect 12805 23131 12863 23137
rect 12989 23171 13047 23177
rect 12989 23137 13001 23171
rect 13035 23168 13047 23171
rect 13170 23168 13176 23180
rect 13035 23140 13176 23168
rect 13035 23137 13047 23140
rect 12989 23131 13047 23137
rect 13170 23128 13176 23140
rect 13228 23128 13234 23180
rect 13538 23128 13544 23180
rect 13596 23168 13602 23180
rect 13909 23171 13967 23177
rect 13909 23168 13921 23171
rect 13596 23140 13921 23168
rect 13596 23128 13602 23140
rect 13909 23137 13921 23140
rect 13955 23137 13967 23171
rect 13909 23131 13967 23137
rect 15565 23171 15623 23177
rect 15565 23137 15577 23171
rect 15611 23168 15623 23171
rect 16482 23168 16488 23180
rect 15611 23140 16488 23168
rect 15611 23137 15623 23140
rect 15565 23131 15623 23137
rect 16482 23128 16488 23140
rect 16540 23128 16546 23180
rect 10735 23072 11100 23100
rect 10735 23069 10747 23072
rect 10689 23063 10747 23069
rect 11146 23060 11152 23112
rect 11204 23100 11210 23112
rect 14182 23100 14188 23112
rect 11204 23072 14188 23100
rect 11204 23060 11210 23072
rect 14182 23060 14188 23072
rect 14240 23060 14246 23112
rect 15286 23100 15292 23112
rect 15247 23072 15292 23100
rect 15286 23060 15292 23072
rect 15344 23060 15350 23112
rect 6328 23004 7420 23032
rect 6328 22992 6334 23004
rect 13722 22992 13728 23044
rect 13780 23032 13786 23044
rect 13817 23035 13875 23041
rect 13817 23032 13829 23035
rect 13780 23004 13829 23032
rect 13780 22992 13786 23004
rect 13817 23001 13829 23004
rect 13863 23032 13875 23035
rect 14642 23032 14648 23044
rect 13863 23004 14648 23032
rect 13863 23001 13875 23004
rect 13817 22995 13875 23001
rect 14642 22992 14648 23004
rect 14700 22992 14706 23044
rect 7745 22967 7803 22973
rect 7745 22933 7757 22967
rect 7791 22964 7803 22967
rect 7834 22964 7840 22976
rect 7791 22936 7840 22964
rect 7791 22933 7803 22936
rect 7745 22927 7803 22933
rect 7834 22924 7840 22936
rect 7892 22924 7898 22976
rect 13262 22924 13268 22976
rect 13320 22964 13326 22976
rect 13357 22967 13415 22973
rect 13357 22964 13369 22967
rect 13320 22936 13369 22964
rect 13320 22924 13326 22936
rect 13357 22933 13369 22936
rect 13403 22933 13415 22967
rect 13357 22927 13415 22933
rect 13998 22924 14004 22976
rect 14056 22964 14062 22976
rect 14093 22967 14151 22973
rect 14093 22964 14105 22967
rect 14056 22936 14105 22964
rect 14056 22924 14062 22936
rect 14093 22933 14105 22936
rect 14139 22933 14151 22967
rect 14093 22927 14151 22933
rect 14274 22924 14280 22976
rect 14332 22964 14338 22976
rect 15470 22964 15476 22976
rect 14332 22936 15476 22964
rect 14332 22924 14338 22936
rect 15470 22924 15476 22936
rect 15528 22924 15534 22976
rect 16298 22924 16304 22976
rect 16356 22964 16362 22976
rect 16393 22967 16451 22973
rect 16393 22964 16405 22967
rect 16356 22936 16405 22964
rect 16356 22924 16362 22936
rect 16393 22933 16405 22936
rect 16439 22964 16451 22967
rect 16758 22964 16764 22976
rect 16439 22936 16764 22964
rect 16439 22933 16451 22936
rect 16393 22927 16451 22933
rect 16758 22924 16764 22936
rect 16816 22924 16822 22976
rect 1104 22874 28888 22896
rect 1104 22822 5982 22874
rect 6034 22822 6046 22874
rect 6098 22822 6110 22874
rect 6162 22822 6174 22874
rect 6226 22822 15982 22874
rect 16034 22822 16046 22874
rect 16098 22822 16110 22874
rect 16162 22822 16174 22874
rect 16226 22822 25982 22874
rect 26034 22822 26046 22874
rect 26098 22822 26110 22874
rect 26162 22822 26174 22874
rect 26226 22822 28888 22874
rect 1104 22800 28888 22822
rect 5905 22763 5963 22769
rect 5905 22729 5917 22763
rect 5951 22760 5963 22763
rect 7190 22760 7196 22772
rect 5951 22732 7196 22760
rect 5951 22729 5963 22732
rect 5905 22723 5963 22729
rect 7190 22720 7196 22732
rect 7248 22760 7254 22772
rect 8205 22763 8263 22769
rect 8205 22760 8217 22763
rect 7248 22732 8217 22760
rect 7248 22720 7254 22732
rect 8205 22729 8217 22732
rect 8251 22729 8263 22763
rect 8205 22723 8263 22729
rect 9861 22763 9919 22769
rect 9861 22729 9873 22763
rect 9907 22760 9919 22763
rect 9950 22760 9956 22772
rect 9907 22732 9956 22760
rect 9907 22729 9919 22732
rect 9861 22723 9919 22729
rect 9950 22720 9956 22732
rect 10008 22720 10014 22772
rect 10229 22763 10287 22769
rect 10229 22729 10241 22763
rect 10275 22760 10287 22763
rect 11146 22760 11152 22772
rect 10275 22732 11152 22760
rect 10275 22729 10287 22732
rect 10229 22723 10287 22729
rect 11146 22720 11152 22732
rect 11204 22720 11210 22772
rect 11698 22760 11704 22772
rect 11659 22732 11704 22760
rect 11698 22720 11704 22732
rect 11756 22720 11762 22772
rect 13357 22763 13415 22769
rect 13357 22729 13369 22763
rect 13403 22760 13415 22763
rect 13814 22760 13820 22772
rect 13403 22732 13820 22760
rect 13403 22729 13415 22732
rect 13357 22723 13415 22729
rect 6270 22692 6276 22704
rect 6231 22664 6276 22692
rect 6270 22652 6276 22664
rect 6328 22652 6334 22704
rect 6638 22692 6644 22704
rect 6599 22664 6644 22692
rect 6638 22652 6644 22664
rect 6696 22652 6702 22704
rect 11514 22652 11520 22704
rect 11572 22692 11578 22704
rect 11977 22695 12035 22701
rect 11977 22692 11989 22695
rect 11572 22664 11989 22692
rect 11572 22652 11578 22664
rect 11977 22661 11989 22664
rect 12023 22692 12035 22695
rect 12618 22692 12624 22704
rect 12023 22664 12624 22692
rect 12023 22661 12035 22664
rect 11977 22655 12035 22661
rect 12618 22652 12624 22664
rect 12676 22652 12682 22704
rect 6822 22624 6828 22636
rect 6783 22596 6828 22624
rect 6822 22584 6828 22596
rect 6880 22584 6886 22636
rect 7098 22624 7104 22636
rect 7011 22596 7104 22624
rect 7098 22584 7104 22596
rect 7156 22624 7162 22636
rect 7282 22624 7288 22636
rect 7156 22596 7288 22624
rect 7156 22584 7162 22596
rect 7282 22584 7288 22596
rect 7340 22624 7346 22636
rect 7834 22624 7840 22636
rect 7340 22596 7840 22624
rect 7340 22584 7346 22596
rect 7834 22584 7840 22596
rect 7892 22584 7898 22636
rect 12434 22584 12440 22636
rect 12492 22624 12498 22636
rect 12894 22624 12900 22636
rect 12492 22596 12900 22624
rect 12492 22584 12498 22596
rect 12894 22584 12900 22596
rect 12952 22584 12958 22636
rect 8570 22516 8576 22568
rect 8628 22556 8634 22568
rect 8849 22559 8907 22565
rect 8849 22556 8861 22559
rect 8628 22528 8861 22556
rect 8628 22516 8634 22528
rect 8849 22525 8861 22528
rect 8895 22556 8907 22559
rect 9217 22559 9275 22565
rect 9217 22556 9229 22559
rect 8895 22528 9229 22556
rect 8895 22525 8907 22528
rect 8849 22519 8907 22525
rect 9217 22525 9229 22528
rect 9263 22556 9275 22559
rect 9309 22559 9367 22565
rect 9309 22556 9321 22559
rect 9263 22528 9321 22556
rect 9263 22525 9275 22528
rect 9217 22519 9275 22525
rect 9309 22525 9321 22528
rect 9355 22556 9367 22559
rect 10321 22559 10379 22565
rect 10321 22556 10333 22559
rect 9355 22528 10333 22556
rect 9355 22525 9367 22528
rect 9309 22519 9367 22525
rect 10321 22525 10333 22528
rect 10367 22556 10379 22559
rect 11149 22559 11207 22565
rect 11149 22556 11161 22559
rect 10367 22528 11161 22556
rect 10367 22525 10379 22528
rect 10321 22519 10379 22525
rect 11149 22525 11161 22528
rect 11195 22525 11207 22559
rect 11149 22519 11207 22525
rect 12529 22559 12587 22565
rect 12529 22525 12541 22559
rect 12575 22556 12587 22559
rect 13372 22556 13400 22723
rect 13814 22720 13820 22732
rect 13872 22760 13878 22772
rect 13998 22760 14004 22772
rect 13872 22732 14004 22760
rect 13872 22720 13878 22732
rect 13998 22720 14004 22732
rect 14056 22720 14062 22772
rect 15102 22720 15108 22772
rect 15160 22760 15166 22772
rect 15289 22763 15347 22769
rect 15289 22760 15301 22763
rect 15160 22732 15301 22760
rect 15160 22720 15166 22732
rect 15289 22729 15301 22732
rect 15335 22729 15347 22763
rect 15289 22723 15347 22729
rect 19610 22720 19616 22772
rect 19668 22760 19674 22772
rect 21266 22760 21272 22772
rect 19668 22732 21272 22760
rect 19668 22720 19674 22732
rect 21266 22720 21272 22732
rect 21324 22720 21330 22772
rect 13538 22652 13544 22704
rect 13596 22692 13602 22704
rect 13725 22695 13783 22701
rect 13725 22692 13737 22695
rect 13596 22664 13737 22692
rect 13596 22652 13602 22664
rect 13725 22661 13737 22664
rect 13771 22661 13783 22695
rect 13725 22655 13783 22661
rect 16117 22695 16175 22701
rect 16117 22661 16129 22695
rect 16163 22692 16175 22695
rect 16298 22692 16304 22704
rect 16163 22664 16304 22692
rect 16163 22661 16175 22664
rect 16117 22655 16175 22661
rect 13446 22584 13452 22636
rect 13504 22624 13510 22636
rect 13630 22624 13636 22636
rect 13504 22596 13636 22624
rect 13504 22584 13510 22596
rect 13630 22584 13636 22596
rect 13688 22584 13694 22636
rect 12575 22528 13400 22556
rect 12575 22525 12587 22528
rect 12529 22519 12587 22525
rect 8938 22448 8944 22500
rect 8996 22488 9002 22500
rect 9398 22488 9404 22500
rect 8996 22460 9404 22488
rect 8996 22448 9002 22460
rect 9398 22448 9404 22460
rect 9456 22448 9462 22500
rect 10873 22491 10931 22497
rect 10873 22457 10885 22491
rect 10919 22488 10931 22491
rect 10962 22488 10968 22500
rect 10919 22460 10968 22488
rect 10919 22457 10931 22460
rect 10873 22451 10931 22457
rect 10962 22448 10968 22460
rect 11020 22488 11026 22500
rect 11330 22488 11336 22500
rect 11020 22460 11336 22488
rect 11020 22448 11026 22460
rect 11330 22448 11336 22460
rect 11388 22448 11394 22500
rect 12986 22488 12992 22500
rect 12947 22460 12992 22488
rect 12986 22448 12992 22460
rect 13044 22448 13050 22500
rect 5537 22423 5595 22429
rect 5537 22389 5549 22423
rect 5583 22420 5595 22423
rect 7098 22420 7104 22432
rect 5583 22392 7104 22420
rect 5583 22389 5595 22392
rect 5537 22383 5595 22389
rect 7098 22380 7104 22392
rect 7156 22380 7162 22432
rect 9490 22420 9496 22432
rect 9451 22392 9496 22420
rect 9490 22380 9496 22392
rect 9548 22380 9554 22432
rect 10042 22380 10048 22432
rect 10100 22420 10106 22432
rect 10505 22423 10563 22429
rect 10505 22420 10517 22423
rect 10100 22392 10517 22420
rect 10100 22380 10106 22392
rect 10505 22389 10517 22392
rect 10551 22389 10563 22423
rect 13740 22420 13768 22655
rect 16298 22652 16304 22664
rect 16356 22692 16362 22704
rect 16482 22692 16488 22704
rect 16356 22664 16488 22692
rect 16356 22652 16362 22664
rect 16482 22652 16488 22664
rect 16540 22652 16546 22704
rect 14826 22584 14832 22636
rect 14884 22624 14890 22636
rect 14921 22627 14979 22633
rect 14921 22624 14933 22627
rect 14884 22596 14933 22624
rect 14884 22584 14890 22596
rect 14921 22593 14933 22596
rect 14967 22593 14979 22627
rect 14921 22587 14979 22593
rect 17865 22627 17923 22633
rect 17865 22593 17877 22627
rect 17911 22624 17923 22627
rect 18325 22627 18383 22633
rect 18325 22624 18337 22627
rect 17911 22596 18337 22624
rect 17911 22593 17923 22596
rect 17865 22587 17923 22593
rect 18325 22593 18337 22596
rect 18371 22624 18383 22627
rect 18414 22624 18420 22636
rect 18371 22596 18420 22624
rect 18371 22593 18383 22596
rect 18325 22587 18383 22593
rect 18414 22584 18420 22596
rect 18472 22584 18478 22636
rect 25866 22584 25872 22636
rect 25924 22624 25930 22636
rect 26053 22627 26111 22633
rect 26053 22624 26065 22627
rect 25924 22596 26065 22624
rect 25924 22584 25930 22596
rect 26053 22593 26065 22596
rect 26099 22624 26111 22627
rect 26421 22627 26479 22633
rect 26421 22624 26433 22627
rect 26099 22596 26433 22624
rect 26099 22593 26111 22596
rect 26053 22587 26111 22593
rect 26421 22593 26433 22596
rect 26467 22593 26479 22627
rect 26421 22587 26479 22593
rect 14093 22559 14151 22565
rect 14093 22525 14105 22559
rect 14139 22525 14151 22559
rect 14274 22556 14280 22568
rect 14235 22528 14280 22556
rect 14093 22519 14151 22525
rect 14108 22488 14136 22519
rect 14274 22516 14280 22528
rect 14332 22516 14338 22568
rect 14642 22556 14648 22568
rect 14603 22528 14648 22556
rect 14642 22516 14648 22528
rect 14700 22516 14706 22568
rect 15286 22516 15292 22568
rect 15344 22556 15350 22568
rect 15565 22559 15623 22565
rect 15565 22556 15577 22559
rect 15344 22528 15577 22556
rect 15344 22516 15350 22528
rect 15565 22525 15577 22528
rect 15611 22525 15623 22559
rect 15565 22519 15623 22525
rect 15654 22516 15660 22568
rect 15712 22556 15718 22568
rect 16393 22559 16451 22565
rect 16393 22556 16405 22559
rect 15712 22528 16405 22556
rect 15712 22516 15718 22528
rect 16393 22525 16405 22528
rect 16439 22525 16451 22559
rect 16393 22519 16451 22525
rect 18049 22559 18107 22565
rect 18049 22525 18061 22559
rect 18095 22556 18107 22559
rect 18138 22556 18144 22568
rect 18095 22528 18144 22556
rect 18095 22525 18107 22528
rect 18049 22519 18107 22525
rect 18138 22516 18144 22528
rect 18196 22516 18202 22568
rect 26142 22556 26148 22568
rect 26103 22528 26148 22556
rect 26142 22516 26148 22528
rect 26200 22516 26206 22568
rect 14918 22488 14924 22500
rect 14108 22460 14924 22488
rect 14918 22448 14924 22460
rect 14976 22448 14982 22500
rect 15470 22448 15476 22500
rect 15528 22488 15534 22500
rect 16666 22488 16672 22500
rect 15528 22460 16672 22488
rect 15528 22448 15534 22460
rect 16666 22448 16672 22460
rect 16724 22448 16730 22500
rect 15378 22420 15384 22432
rect 13740 22392 15384 22420
rect 10505 22383 10563 22389
rect 15378 22380 15384 22392
rect 15436 22380 15442 22432
rect 15565 22423 15623 22429
rect 15565 22389 15577 22423
rect 15611 22420 15623 22423
rect 15657 22423 15715 22429
rect 15657 22420 15669 22423
rect 15611 22392 15669 22420
rect 15611 22389 15623 22392
rect 15565 22383 15623 22389
rect 15657 22389 15669 22392
rect 15703 22389 15715 22423
rect 15657 22383 15715 22389
rect 15838 22380 15844 22432
rect 15896 22420 15902 22432
rect 16390 22420 16396 22432
rect 15896 22392 16396 22420
rect 15896 22380 15902 22392
rect 16390 22380 16396 22392
rect 16448 22380 16454 22432
rect 16574 22380 16580 22432
rect 16632 22420 16638 22432
rect 16761 22423 16819 22429
rect 16761 22420 16773 22423
rect 16632 22392 16773 22420
rect 16632 22380 16638 22392
rect 16761 22389 16773 22392
rect 16807 22389 16819 22423
rect 16761 22383 16819 22389
rect 19334 22380 19340 22432
rect 19392 22420 19398 22432
rect 19429 22423 19487 22429
rect 19429 22420 19441 22423
rect 19392 22392 19441 22420
rect 19392 22380 19398 22392
rect 19429 22389 19441 22392
rect 19475 22389 19487 22423
rect 27706 22420 27712 22432
rect 27667 22392 27712 22420
rect 19429 22383 19487 22389
rect 27706 22380 27712 22392
rect 27764 22380 27770 22432
rect 1104 22330 28888 22352
rect 1104 22278 10982 22330
rect 11034 22278 11046 22330
rect 11098 22278 11110 22330
rect 11162 22278 11174 22330
rect 11226 22278 20982 22330
rect 21034 22278 21046 22330
rect 21098 22278 21110 22330
rect 21162 22278 21174 22330
rect 21226 22278 28888 22330
rect 1104 22256 28888 22278
rect 9490 22176 9496 22228
rect 9548 22216 9554 22228
rect 9548 22188 10640 22216
rect 9548 22176 9554 22188
rect 10612 22148 10640 22188
rect 12894 22176 12900 22228
rect 12952 22216 12958 22228
rect 12989 22219 13047 22225
rect 12989 22216 13001 22219
rect 12952 22188 13001 22216
rect 12952 22176 12958 22188
rect 12989 22185 13001 22188
rect 13035 22185 13047 22219
rect 12989 22179 13047 22185
rect 14093 22219 14151 22225
rect 14093 22185 14105 22219
rect 14139 22216 14151 22219
rect 14274 22216 14280 22228
rect 14139 22188 14280 22216
rect 14139 22185 14151 22188
rect 14093 22179 14151 22185
rect 14274 22176 14280 22188
rect 14332 22176 14338 22228
rect 14461 22219 14519 22225
rect 14461 22185 14473 22219
rect 14507 22216 14519 22219
rect 14918 22216 14924 22228
rect 14507 22188 14924 22216
rect 14507 22185 14519 22188
rect 14461 22179 14519 22185
rect 14918 22176 14924 22188
rect 14976 22176 14982 22228
rect 16574 22176 16580 22228
rect 16632 22176 16638 22228
rect 17037 22219 17095 22225
rect 17037 22185 17049 22219
rect 17083 22185 17095 22219
rect 17037 22179 17095 22185
rect 14734 22148 14740 22160
rect 10612 22120 14740 22148
rect 14734 22108 14740 22120
rect 14792 22108 14798 22160
rect 16592 22148 16620 22176
rect 17052 22148 17080 22179
rect 18414 22176 18420 22228
rect 18472 22216 18478 22228
rect 18874 22216 18880 22228
rect 18472 22188 18880 22216
rect 18472 22176 18478 22188
rect 18874 22176 18880 22188
rect 18932 22176 18938 22228
rect 25774 22176 25780 22228
rect 25832 22216 25838 22228
rect 26142 22216 26148 22228
rect 25832 22188 26148 22216
rect 25832 22176 25838 22188
rect 26142 22176 26148 22188
rect 26200 22176 26206 22228
rect 16500 22120 16620 22148
rect 16684 22120 18644 22148
rect 6089 22083 6147 22089
rect 6089 22049 6101 22083
rect 6135 22080 6147 22083
rect 6822 22080 6828 22092
rect 6135 22052 6828 22080
rect 6135 22049 6147 22052
rect 6089 22043 6147 22049
rect 6288 22024 6316 22052
rect 6822 22040 6828 22052
rect 6880 22040 6886 22092
rect 8570 22080 8576 22092
rect 8531 22052 8576 22080
rect 8570 22040 8576 22052
rect 8628 22040 8634 22092
rect 12066 22040 12072 22092
rect 12124 22080 12130 22092
rect 12161 22083 12219 22089
rect 12161 22080 12173 22083
rect 12124 22052 12173 22080
rect 12124 22040 12130 22052
rect 12161 22049 12173 22052
rect 12207 22080 12219 22083
rect 12250 22080 12256 22092
rect 12207 22052 12256 22080
rect 12207 22049 12219 22052
rect 12161 22043 12219 22049
rect 12250 22040 12256 22052
rect 12308 22040 12314 22092
rect 13265 22083 13323 22089
rect 13265 22049 13277 22083
rect 13311 22049 13323 22083
rect 15381 22083 15439 22089
rect 15381 22080 15393 22083
rect 13265 22043 13323 22049
rect 15028 22052 15393 22080
rect 6270 21972 6276 22024
rect 6328 21972 6334 22024
rect 6362 21972 6368 22024
rect 6420 22012 6426 22024
rect 6420 21984 6465 22012
rect 6420 21972 6426 21984
rect 8294 21972 8300 22024
rect 8352 22012 8358 22024
rect 9493 22015 9551 22021
rect 9493 22012 9505 22015
rect 8352 21984 9505 22012
rect 8352 21972 8358 21984
rect 9493 21981 9505 21984
rect 9539 22012 9551 22015
rect 9677 22015 9735 22021
rect 9677 22012 9689 22015
rect 9539 21984 9689 22012
rect 9539 21981 9551 21984
rect 9493 21975 9551 21981
rect 9677 21981 9689 21984
rect 9723 21981 9735 22015
rect 9950 22012 9956 22024
rect 9911 21984 9956 22012
rect 9677 21975 9735 21981
rect 9950 21972 9956 21984
rect 10008 21972 10014 22024
rect 13170 22012 13176 22024
rect 13131 21984 13176 22012
rect 13170 21972 13176 21984
rect 13228 21972 13234 22024
rect 12345 21947 12403 21953
rect 12345 21913 12357 21947
rect 12391 21944 12403 21947
rect 13280 21944 13308 22043
rect 15028 22024 15056 22052
rect 15381 22049 15393 22052
rect 15427 22049 15439 22083
rect 15381 22043 15439 22049
rect 16500 22024 16528 22120
rect 16574 22040 16580 22092
rect 16632 22080 16638 22092
rect 16684 22080 16712 22120
rect 18616 22092 18644 22120
rect 16632 22052 16712 22080
rect 16632 22040 16638 22052
rect 16758 22040 16764 22092
rect 16816 22080 16822 22092
rect 16853 22083 16911 22089
rect 16853 22080 16865 22083
rect 16816 22052 16865 22080
rect 16816 22040 16822 22052
rect 16853 22049 16865 22052
rect 16899 22049 16911 22083
rect 16853 22043 16911 22049
rect 18598 22040 18604 22092
rect 18656 22080 18662 22092
rect 18969 22083 19027 22089
rect 18969 22080 18981 22083
rect 18656 22052 18981 22080
rect 18656 22040 18662 22052
rect 18969 22049 18981 22052
rect 19015 22049 19027 22083
rect 19334 22080 19340 22092
rect 19295 22052 19340 22080
rect 18969 22043 19027 22049
rect 19334 22040 19340 22052
rect 19392 22040 19398 22092
rect 15010 21972 15016 22024
rect 15068 21972 15074 22024
rect 15102 21972 15108 22024
rect 15160 22012 15166 22024
rect 15289 22015 15347 22021
rect 15289 22012 15301 22015
rect 15160 21984 15301 22012
rect 15160 21972 15166 21984
rect 15289 21981 15301 21984
rect 15335 22012 15347 22015
rect 16117 22015 16175 22021
rect 16117 22012 16129 22015
rect 15335 21984 16129 22012
rect 15335 21981 15347 21984
rect 15289 21975 15347 21981
rect 16117 21981 16129 21984
rect 16163 21981 16175 22015
rect 16117 21975 16175 21981
rect 16482 21972 16488 22024
rect 16540 21972 16546 22024
rect 17034 21972 17040 22024
rect 17092 22012 17098 22024
rect 17494 22012 17500 22024
rect 17092 21984 17500 22012
rect 17092 21972 17098 21984
rect 17494 21972 17500 21984
rect 17552 21972 17558 22024
rect 18414 22012 18420 22024
rect 18375 21984 18420 22012
rect 18414 21972 18420 21984
rect 18472 21972 18478 22024
rect 19058 22012 19064 22024
rect 18892 21984 19064 22012
rect 18892 21956 18920 21984
rect 19058 21972 19064 21984
rect 19116 21972 19122 22024
rect 19242 22012 19248 22024
rect 19203 21984 19248 22012
rect 19242 21972 19248 21984
rect 19300 21972 19306 22024
rect 13814 21944 13820 21956
rect 12391 21916 13820 21944
rect 12391 21913 12403 21916
rect 12345 21907 12403 21913
rect 13814 21904 13820 21916
rect 13872 21904 13878 21956
rect 18874 21904 18880 21956
rect 18932 21904 18938 21956
rect 7653 21879 7711 21885
rect 7653 21845 7665 21879
rect 7699 21876 7711 21879
rect 7926 21876 7932 21888
rect 7699 21848 7932 21876
rect 7699 21845 7711 21848
rect 7653 21839 7711 21845
rect 7926 21836 7932 21848
rect 7984 21836 7990 21888
rect 8754 21876 8760 21888
rect 8715 21848 8760 21876
rect 8754 21836 8760 21848
rect 8812 21836 8818 21888
rect 11241 21879 11299 21885
rect 11241 21845 11253 21879
rect 11287 21876 11299 21879
rect 11698 21876 11704 21888
rect 11287 21848 11704 21876
rect 11287 21845 11299 21848
rect 11241 21839 11299 21845
rect 11698 21836 11704 21848
rect 11756 21836 11762 21888
rect 12069 21879 12127 21885
rect 12069 21845 12081 21879
rect 12115 21876 12127 21879
rect 12250 21876 12256 21888
rect 12115 21848 12256 21876
rect 12115 21845 12127 21848
rect 12069 21839 12127 21845
rect 12250 21836 12256 21848
rect 12308 21876 12314 21888
rect 12434 21876 12440 21888
rect 12308 21848 12440 21876
rect 12308 21836 12314 21848
rect 12434 21836 12440 21848
rect 12492 21836 12498 21888
rect 12710 21876 12716 21888
rect 12671 21848 12716 21876
rect 12710 21836 12716 21848
rect 12768 21836 12774 21888
rect 13446 21876 13452 21888
rect 13407 21848 13452 21876
rect 13446 21836 13452 21848
rect 13504 21836 13510 21888
rect 14182 21836 14188 21888
rect 14240 21876 14246 21888
rect 15565 21879 15623 21885
rect 15565 21876 15577 21879
rect 14240 21848 15577 21876
rect 14240 21836 14246 21848
rect 15565 21845 15577 21848
rect 15611 21845 15623 21879
rect 16666 21876 16672 21888
rect 16627 21848 16672 21876
rect 15565 21839 15623 21845
rect 16666 21836 16672 21848
rect 16724 21836 16730 21888
rect 18138 21876 18144 21888
rect 18099 21848 18144 21876
rect 18138 21836 18144 21848
rect 18196 21836 18202 21888
rect 1104 21786 28888 21808
rect 1104 21734 5982 21786
rect 6034 21734 6046 21786
rect 6098 21734 6110 21786
rect 6162 21734 6174 21786
rect 6226 21734 15982 21786
rect 16034 21734 16046 21786
rect 16098 21734 16110 21786
rect 16162 21734 16174 21786
rect 16226 21734 25982 21786
rect 26034 21734 26046 21786
rect 26098 21734 26110 21786
rect 26162 21734 26174 21786
rect 26226 21734 28888 21786
rect 1104 21712 28888 21734
rect 8570 21672 8576 21684
rect 8531 21644 8576 21672
rect 8570 21632 8576 21644
rect 8628 21632 8634 21684
rect 9769 21675 9827 21681
rect 9769 21641 9781 21675
rect 9815 21672 9827 21675
rect 9950 21672 9956 21684
rect 9815 21644 9956 21672
rect 9815 21641 9827 21644
rect 9769 21635 9827 21641
rect 9950 21632 9956 21644
rect 10008 21632 10014 21684
rect 10778 21672 10784 21684
rect 10739 21644 10784 21672
rect 10778 21632 10784 21644
rect 10836 21632 10842 21684
rect 11885 21675 11943 21681
rect 11885 21641 11897 21675
rect 11931 21672 11943 21675
rect 12066 21672 12072 21684
rect 11931 21644 12072 21672
rect 11931 21641 11943 21644
rect 11885 21635 11943 21641
rect 12066 21632 12072 21644
rect 12124 21672 12130 21684
rect 12618 21672 12624 21684
rect 12124 21644 12624 21672
rect 12124 21632 12130 21644
rect 12618 21632 12624 21644
rect 12676 21632 12682 21684
rect 13814 21672 13820 21684
rect 13775 21644 13820 21672
rect 13814 21632 13820 21644
rect 13872 21672 13878 21684
rect 16298 21672 16304 21684
rect 13872 21644 16304 21672
rect 13872 21632 13878 21644
rect 16298 21632 16304 21644
rect 16356 21632 16362 21684
rect 16390 21632 16396 21684
rect 16448 21672 16454 21684
rect 16758 21672 16764 21684
rect 16448 21644 16764 21672
rect 16448 21632 16454 21644
rect 16758 21632 16764 21644
rect 16816 21672 16822 21684
rect 17405 21675 17463 21681
rect 17405 21672 17417 21675
rect 16816 21644 17417 21672
rect 16816 21632 16822 21644
rect 17405 21641 17417 21644
rect 17451 21641 17463 21675
rect 17678 21672 17684 21684
rect 17639 21644 17684 21672
rect 17405 21635 17463 21641
rect 17678 21632 17684 21644
rect 17736 21632 17742 21684
rect 19334 21672 19340 21684
rect 19295 21644 19340 21672
rect 19334 21632 19340 21644
rect 19392 21632 19398 21684
rect 5905 21607 5963 21613
rect 5905 21573 5917 21607
rect 5951 21604 5963 21607
rect 6362 21604 6368 21616
rect 5951 21576 6368 21604
rect 5951 21573 5963 21576
rect 5905 21567 5963 21573
rect 6362 21564 6368 21576
rect 6420 21564 6426 21616
rect 9125 21607 9183 21613
rect 9125 21573 9137 21607
rect 9171 21573 9183 21607
rect 9125 21567 9183 21573
rect 6641 21539 6699 21545
rect 6641 21505 6653 21539
rect 6687 21536 6699 21539
rect 7377 21539 7435 21545
rect 7377 21536 7389 21539
rect 6687 21508 7389 21536
rect 6687 21505 6699 21508
rect 6641 21499 6699 21505
rect 7377 21505 7389 21508
rect 7423 21536 7435 21539
rect 8846 21536 8852 21548
rect 7423 21508 8852 21536
rect 7423 21505 7435 21508
rect 7377 21499 7435 21505
rect 8846 21496 8852 21508
rect 8904 21536 8910 21548
rect 9140 21536 9168 21567
rect 8904 21508 9168 21536
rect 10796 21536 10824 21632
rect 13170 21564 13176 21616
rect 13228 21564 13234 21616
rect 17770 21604 17776 21616
rect 16592 21576 17776 21604
rect 12253 21539 12311 21545
rect 10796 21508 11100 21536
rect 8904 21496 8910 21508
rect 7561 21471 7619 21477
rect 7561 21468 7573 21471
rect 6656 21440 7573 21468
rect 6656 21412 6684 21440
rect 7561 21437 7573 21440
rect 7607 21437 7619 21471
rect 7926 21468 7932 21480
rect 7887 21440 7932 21468
rect 7561 21431 7619 21437
rect 7926 21428 7932 21440
rect 7984 21428 7990 21480
rect 8021 21471 8079 21477
rect 8021 21437 8033 21471
rect 8067 21468 8079 21471
rect 8754 21468 8760 21480
rect 8067 21440 8760 21468
rect 8067 21437 8079 21440
rect 8021 21431 8079 21437
rect 6638 21360 6644 21412
rect 6696 21360 6702 21412
rect 6914 21400 6920 21412
rect 6875 21372 6920 21400
rect 6914 21360 6920 21372
rect 6972 21360 6978 21412
rect 6273 21335 6331 21341
rect 6273 21301 6285 21335
rect 6319 21332 6331 21335
rect 7282 21332 7288 21344
rect 6319 21304 7288 21332
rect 6319 21301 6331 21304
rect 6273 21295 6331 21301
rect 7282 21292 7288 21304
rect 7340 21332 7346 21344
rect 8036 21332 8064 21431
rect 8754 21428 8760 21440
rect 8812 21428 8818 21480
rect 8938 21468 8944 21480
rect 8899 21440 8944 21468
rect 8938 21428 8944 21440
rect 8996 21428 9002 21480
rect 9490 21428 9496 21480
rect 9548 21468 9554 21480
rect 10137 21471 10195 21477
rect 10137 21468 10149 21471
rect 9548 21440 10149 21468
rect 9548 21428 9554 21440
rect 10137 21437 10149 21440
rect 10183 21468 10195 21471
rect 10594 21468 10600 21480
rect 10183 21440 10600 21468
rect 10183 21437 10195 21440
rect 10137 21431 10195 21437
rect 10594 21428 10600 21440
rect 10652 21428 10658 21480
rect 11072 21477 11100 21508
rect 12253 21505 12265 21539
rect 12299 21536 12311 21539
rect 13188 21536 13216 21564
rect 13814 21536 13820 21548
rect 12299 21508 12572 21536
rect 13188 21508 13820 21536
rect 12299 21505 12311 21508
rect 12253 21499 12311 21505
rect 10689 21471 10747 21477
rect 10689 21437 10701 21471
rect 10735 21468 10747 21471
rect 10965 21471 11023 21477
rect 10965 21468 10977 21471
rect 10735 21440 10977 21468
rect 10735 21437 10747 21440
rect 10689 21431 10747 21437
rect 10965 21437 10977 21440
rect 11011 21437 11023 21471
rect 10965 21431 11023 21437
rect 11057 21471 11115 21477
rect 11057 21437 11069 21471
rect 11103 21468 11115 21471
rect 12434 21468 12440 21480
rect 11103 21440 12440 21468
rect 11103 21437 11115 21440
rect 11057 21431 11115 21437
rect 12434 21428 12440 21440
rect 12492 21428 12498 21480
rect 12544 21477 12572 21508
rect 13814 21496 13820 21508
rect 13872 21496 13878 21548
rect 13998 21496 14004 21548
rect 14056 21536 14062 21548
rect 16592 21545 16620 21576
rect 17420 21548 17448 21576
rect 17770 21564 17776 21576
rect 17828 21564 17834 21616
rect 18782 21604 18788 21616
rect 17880 21576 18788 21604
rect 14553 21539 14611 21545
rect 14553 21536 14565 21539
rect 14056 21508 14565 21536
rect 14056 21496 14062 21508
rect 14553 21505 14565 21508
rect 14599 21505 14611 21539
rect 14553 21499 14611 21505
rect 16209 21539 16267 21545
rect 16209 21505 16221 21539
rect 16255 21536 16267 21539
rect 16577 21539 16635 21545
rect 16577 21536 16589 21539
rect 16255 21508 16589 21536
rect 16255 21505 16267 21508
rect 16209 21499 16267 21505
rect 16577 21505 16589 21508
rect 16623 21505 16635 21539
rect 16577 21499 16635 21505
rect 17402 21496 17408 21548
rect 17460 21496 17466 21548
rect 17678 21496 17684 21548
rect 17736 21536 17742 21548
rect 17880 21545 17908 21576
rect 18782 21564 18788 21576
rect 18840 21564 18846 21616
rect 17865 21539 17923 21545
rect 17865 21536 17877 21539
rect 17736 21508 17877 21536
rect 17736 21496 17742 21508
rect 17865 21505 17877 21508
rect 17911 21505 17923 21539
rect 18046 21536 18052 21548
rect 18007 21508 18052 21536
rect 17865 21499 17923 21505
rect 18046 21496 18052 21508
rect 18104 21496 18110 21548
rect 12529 21471 12587 21477
rect 12529 21437 12541 21471
rect 12575 21437 12587 21471
rect 12529 21431 12587 21437
rect 11514 21400 11520 21412
rect 11475 21372 11520 21400
rect 11514 21360 11520 21372
rect 11572 21360 11578 21412
rect 12544 21400 12572 21431
rect 12710 21428 12716 21480
rect 12768 21468 12774 21480
rect 13170 21468 13176 21480
rect 12768 21440 13176 21468
rect 12768 21428 12774 21440
rect 13170 21428 13176 21440
rect 13228 21468 13234 21480
rect 13265 21471 13323 21477
rect 13265 21468 13277 21471
rect 13228 21440 13277 21468
rect 13228 21428 13234 21440
rect 13265 21437 13277 21440
rect 13311 21437 13323 21471
rect 13446 21468 13452 21480
rect 13407 21440 13452 21468
rect 13265 21431 13323 21437
rect 13446 21428 13452 21440
rect 13504 21428 13510 21480
rect 14645 21471 14703 21477
rect 14645 21437 14657 21471
rect 14691 21468 14703 21471
rect 16482 21468 16488 21480
rect 14691 21440 14725 21468
rect 16443 21440 16488 21468
rect 14691 21437 14703 21440
rect 14645 21431 14703 21437
rect 14274 21400 14280 21412
rect 12544 21372 14280 21400
rect 14274 21360 14280 21372
rect 14332 21360 14338 21412
rect 14461 21403 14519 21409
rect 14461 21369 14473 21403
rect 14507 21400 14519 21403
rect 14660 21400 14688 21431
rect 16482 21428 16488 21440
rect 16540 21428 16546 21480
rect 16666 21428 16672 21480
rect 16724 21468 16730 21480
rect 17129 21471 17187 21477
rect 16724 21440 16769 21468
rect 16724 21428 16730 21440
rect 17129 21437 17141 21471
rect 17175 21468 17187 21471
rect 18138 21468 18144 21480
rect 17175 21440 18144 21468
rect 17175 21437 17187 21440
rect 17129 21431 17187 21437
rect 18138 21428 18144 21440
rect 18196 21468 18202 21480
rect 18509 21471 18567 21477
rect 18509 21468 18521 21471
rect 18196 21440 18521 21468
rect 18196 21428 18202 21440
rect 18509 21437 18521 21440
rect 18555 21437 18567 21471
rect 18509 21431 18567 21437
rect 18693 21471 18751 21477
rect 18693 21437 18705 21471
rect 18739 21437 18751 21471
rect 18800 21468 18828 21564
rect 18877 21471 18935 21477
rect 18877 21468 18889 21471
rect 18800 21440 18889 21468
rect 18693 21431 18751 21437
rect 18877 21437 18889 21440
rect 18923 21437 18935 21471
rect 18877 21431 18935 21437
rect 15654 21400 15660 21412
rect 14507 21372 15660 21400
rect 14507 21369 14519 21372
rect 14461 21363 14519 21369
rect 15654 21360 15660 21372
rect 15712 21360 15718 21412
rect 16758 21360 16764 21412
rect 16816 21400 16822 21412
rect 18708 21400 18736 21431
rect 19705 21403 19763 21409
rect 19705 21400 19717 21403
rect 16816 21372 19717 21400
rect 16816 21360 16822 21372
rect 19705 21369 19717 21372
rect 19751 21369 19763 21403
rect 19705 21363 19763 21369
rect 25038 21360 25044 21412
rect 25096 21400 25102 21412
rect 25314 21400 25320 21412
rect 25096 21372 25320 21400
rect 25096 21360 25102 21372
rect 25314 21360 25320 21372
rect 25372 21360 25378 21412
rect 7340 21304 8064 21332
rect 9953 21335 10011 21341
rect 7340 21292 7346 21304
rect 9953 21301 9965 21335
rect 9999 21332 10011 21335
rect 10318 21332 10324 21344
rect 9999 21304 10324 21332
rect 9999 21301 10011 21304
rect 9953 21295 10011 21301
rect 10318 21292 10324 21304
rect 10376 21292 10382 21344
rect 10505 21335 10563 21341
rect 10505 21301 10517 21335
rect 10551 21332 10563 21335
rect 10594 21332 10600 21344
rect 10551 21304 10600 21332
rect 10551 21301 10563 21304
rect 10505 21295 10563 21301
rect 10594 21292 10600 21304
rect 10652 21332 10658 21344
rect 10689 21335 10747 21341
rect 10689 21332 10701 21335
rect 10652 21304 10701 21332
rect 10652 21292 10658 21304
rect 10689 21301 10701 21304
rect 10735 21301 10747 21335
rect 10689 21295 10747 21301
rect 12250 21292 12256 21344
rect 12308 21332 12314 21344
rect 12529 21335 12587 21341
rect 12529 21332 12541 21335
rect 12308 21304 12541 21332
rect 12308 21292 12314 21304
rect 12529 21301 12541 21304
rect 12575 21301 12587 21335
rect 12529 21295 12587 21301
rect 15010 21292 15016 21344
rect 15068 21332 15074 21344
rect 15565 21335 15623 21341
rect 15565 21332 15577 21335
rect 15068 21304 15577 21332
rect 15068 21292 15074 21304
rect 15565 21301 15577 21304
rect 15611 21332 15623 21335
rect 15930 21332 15936 21344
rect 15611 21304 15936 21332
rect 15611 21301 15623 21304
rect 15565 21295 15623 21301
rect 15930 21292 15936 21304
rect 15988 21292 15994 21344
rect 16206 21292 16212 21344
rect 16264 21332 16270 21344
rect 16301 21335 16359 21341
rect 16301 21332 16313 21335
rect 16264 21304 16313 21332
rect 16264 21292 16270 21304
rect 16301 21301 16313 21304
rect 16347 21301 16359 21335
rect 16301 21295 16359 21301
rect 16482 21292 16488 21344
rect 16540 21332 16546 21344
rect 17681 21335 17739 21341
rect 17681 21332 17693 21335
rect 16540 21304 17693 21332
rect 16540 21292 16546 21304
rect 17681 21301 17693 21304
rect 17727 21301 17739 21335
rect 17681 21295 17739 21301
rect 1104 21242 28888 21264
rect 1104 21190 10982 21242
rect 11034 21190 11046 21242
rect 11098 21190 11110 21242
rect 11162 21190 11174 21242
rect 11226 21190 20982 21242
rect 21034 21190 21046 21242
rect 21098 21190 21110 21242
rect 21162 21190 21174 21242
rect 21226 21190 28888 21242
rect 1104 21168 28888 21190
rect 6181 21131 6239 21137
rect 6181 21097 6193 21131
rect 6227 21128 6239 21131
rect 6270 21128 6276 21140
rect 6227 21100 6276 21128
rect 6227 21097 6239 21100
rect 6181 21091 6239 21097
rect 6270 21088 6276 21100
rect 6328 21088 6334 21140
rect 6638 21088 6644 21140
rect 6696 21128 6702 21140
rect 6917 21131 6975 21137
rect 6917 21128 6929 21131
rect 6696 21100 6929 21128
rect 6696 21088 6702 21100
rect 6917 21097 6929 21100
rect 6963 21097 6975 21131
rect 6917 21091 6975 21097
rect 7377 21131 7435 21137
rect 7377 21097 7389 21131
rect 7423 21128 7435 21131
rect 7926 21128 7932 21140
rect 7423 21100 7932 21128
rect 7423 21097 7435 21100
rect 7377 21091 7435 21097
rect 7926 21088 7932 21100
rect 7984 21088 7990 21140
rect 8938 21128 8944 21140
rect 8899 21100 8944 21128
rect 8938 21088 8944 21100
rect 8996 21088 9002 21140
rect 9490 21128 9496 21140
rect 9451 21100 9496 21128
rect 9490 21088 9496 21100
rect 9548 21088 9554 21140
rect 9858 21128 9864 21140
rect 9819 21100 9864 21128
rect 9858 21088 9864 21100
rect 9916 21088 9922 21140
rect 10873 21131 10931 21137
rect 10873 21097 10885 21131
rect 10919 21128 10931 21131
rect 11422 21128 11428 21140
rect 10919 21100 11428 21128
rect 10919 21097 10931 21100
rect 10873 21091 10931 21097
rect 11422 21088 11428 21100
rect 11480 21088 11486 21140
rect 13078 21128 13084 21140
rect 13039 21100 13084 21128
rect 13078 21088 13084 21100
rect 13136 21088 13142 21140
rect 14274 21088 14280 21140
rect 14332 21128 14338 21140
rect 14369 21131 14427 21137
rect 14369 21128 14381 21131
rect 14332 21100 14381 21128
rect 14332 21088 14338 21100
rect 14369 21097 14381 21100
rect 14415 21097 14427 21131
rect 14369 21091 14427 21097
rect 14734 21088 14740 21140
rect 14792 21128 14798 21140
rect 15933 21131 15991 21137
rect 15933 21128 15945 21131
rect 14792 21100 15945 21128
rect 14792 21088 14798 21100
rect 15933 21097 15945 21100
rect 15979 21128 15991 21131
rect 16482 21128 16488 21140
rect 15979 21100 16488 21128
rect 15979 21097 15991 21100
rect 15933 21091 15991 21097
rect 16482 21088 16488 21100
rect 16540 21088 16546 21140
rect 16666 21088 16672 21140
rect 16724 21128 16730 21140
rect 17773 21131 17831 21137
rect 17773 21128 17785 21131
rect 16724 21100 17785 21128
rect 16724 21088 16730 21100
rect 17773 21097 17785 21100
rect 17819 21097 17831 21131
rect 17773 21091 17831 21097
rect 18417 21131 18475 21137
rect 18417 21097 18429 21131
rect 18463 21128 18475 21131
rect 19242 21128 19248 21140
rect 18463 21100 19248 21128
rect 18463 21097 18475 21100
rect 18417 21091 18475 21097
rect 19242 21088 19248 21100
rect 19300 21088 19306 21140
rect 3142 21060 3148 21072
rect 3103 21032 3148 21060
rect 3142 21020 3148 21032
rect 3200 21020 3206 21072
rect 12066 21060 12072 21072
rect 11072 21032 12072 21060
rect 11072 21004 11100 21032
rect 12066 21020 12072 21032
rect 12124 21020 12130 21072
rect 12529 21063 12587 21069
rect 12529 21029 12541 21063
rect 12575 21060 12587 21063
rect 13446 21060 13452 21072
rect 12575 21032 13452 21060
rect 12575 21029 12587 21032
rect 12529 21023 12587 21029
rect 13446 21020 13452 21032
rect 13504 21020 13510 21072
rect 13814 21020 13820 21072
rect 13872 21060 13878 21072
rect 14093 21063 14151 21069
rect 14093 21060 14105 21063
rect 13872 21032 14105 21060
rect 13872 21020 13878 21032
rect 14093 21029 14105 21032
rect 14139 21060 14151 21063
rect 14642 21060 14648 21072
rect 14139 21032 14648 21060
rect 14139 21029 14151 21032
rect 14093 21023 14151 21029
rect 14642 21020 14648 21032
rect 14700 21020 14706 21072
rect 18598 21020 18604 21072
rect 18656 21060 18662 21072
rect 18693 21063 18751 21069
rect 18693 21060 18705 21063
rect 18656 21032 18705 21060
rect 18656 21020 18662 21032
rect 18693 21029 18705 21032
rect 18739 21029 18751 21063
rect 18693 21023 18751 21029
rect 1578 20952 1584 21004
rect 1636 20992 1642 21004
rect 1765 20995 1823 21001
rect 1765 20992 1777 20995
rect 1636 20964 1777 20992
rect 1636 20952 1642 20964
rect 1765 20961 1777 20964
rect 1811 20961 1823 20995
rect 1765 20955 1823 20961
rect 9677 20995 9735 21001
rect 9677 20961 9689 20995
rect 9723 20992 9735 20995
rect 9858 20992 9864 21004
rect 9723 20964 9864 20992
rect 9723 20961 9735 20964
rect 9677 20955 9735 20961
rect 9858 20952 9864 20964
rect 9916 20992 9922 21004
rect 10042 20992 10048 21004
rect 9916 20964 10048 20992
rect 9916 20952 9922 20964
rect 10042 20952 10048 20964
rect 10100 20952 10106 21004
rect 11054 20992 11060 21004
rect 10967 20964 11060 20992
rect 11054 20952 11060 20964
rect 11112 20952 11118 21004
rect 11149 20995 11207 21001
rect 11149 20961 11161 20995
rect 11195 20961 11207 20995
rect 11149 20955 11207 20961
rect 1489 20927 1547 20933
rect 1489 20893 1501 20927
rect 1535 20924 1547 20927
rect 2130 20924 2136 20936
rect 1535 20896 2136 20924
rect 1535 20893 1547 20896
rect 1489 20887 1547 20893
rect 2130 20884 2136 20896
rect 2188 20884 2194 20936
rect 10870 20884 10876 20936
rect 10928 20924 10934 20936
rect 11164 20924 11192 20955
rect 11514 20952 11520 21004
rect 11572 20992 11578 21004
rect 12805 20995 12863 21001
rect 12805 20992 12817 20995
rect 11572 20964 12817 20992
rect 11572 20952 11578 20964
rect 12805 20961 12817 20964
rect 12851 20961 12863 20995
rect 12986 20992 12992 21004
rect 12947 20964 12992 20992
rect 12805 20955 12863 20961
rect 12986 20952 12992 20964
rect 13044 20952 13050 21004
rect 14182 20992 14188 21004
rect 14143 20964 14188 20992
rect 14182 20952 14188 20964
rect 14240 20952 14246 21004
rect 15381 20995 15439 21001
rect 15381 20961 15393 20995
rect 15427 20992 15439 20995
rect 15470 20992 15476 21004
rect 15427 20964 15476 20992
rect 15427 20961 15439 20964
rect 15381 20955 15439 20961
rect 15470 20952 15476 20964
rect 15528 20952 15534 21004
rect 15562 20952 15568 21004
rect 15620 20992 15626 21004
rect 15930 20992 15936 21004
rect 15620 20964 15936 20992
rect 15620 20952 15626 20964
rect 15930 20952 15936 20964
rect 15988 20992 15994 21004
rect 18966 20992 18972 21004
rect 15988 20964 18972 20992
rect 15988 20952 15994 20964
rect 18966 20952 18972 20964
rect 19024 20952 19030 21004
rect 22462 20952 22468 21004
rect 22520 20992 22526 21004
rect 22649 20995 22707 21001
rect 22649 20992 22661 20995
rect 22520 20964 22661 20992
rect 22520 20952 22526 20964
rect 22649 20961 22661 20964
rect 22695 20961 22707 20995
rect 22649 20955 22707 20961
rect 22922 20952 22928 21004
rect 22980 20952 22986 21004
rect 10928 20896 11192 20924
rect 10928 20884 10934 20896
rect 11698 20884 11704 20936
rect 11756 20924 11762 20936
rect 11974 20924 11980 20936
rect 11756 20896 11980 20924
rect 11756 20884 11762 20896
rect 11974 20884 11980 20896
rect 12032 20884 12038 20936
rect 16298 20884 16304 20936
rect 16356 20924 16362 20936
rect 16393 20927 16451 20933
rect 16393 20924 16405 20927
rect 16356 20896 16405 20924
rect 16356 20884 16362 20896
rect 16393 20893 16405 20896
rect 16439 20893 16451 20927
rect 16666 20924 16672 20936
rect 16627 20896 16672 20924
rect 16393 20887 16451 20893
rect 16666 20884 16672 20896
rect 16724 20884 16730 20936
rect 22373 20927 22431 20933
rect 22373 20893 22385 20927
rect 22419 20924 22431 20927
rect 22940 20924 22968 20952
rect 22419 20896 22968 20924
rect 22419 20893 22431 20896
rect 22373 20887 22431 20893
rect 10413 20859 10471 20865
rect 10413 20825 10425 20859
rect 10459 20856 10471 20859
rect 10962 20856 10968 20868
rect 10459 20828 10968 20856
rect 10459 20825 10471 20828
rect 10413 20819 10471 20825
rect 10962 20816 10968 20828
rect 11020 20816 11026 20868
rect 12069 20859 12127 20865
rect 12069 20856 12081 20859
rect 11072 20828 12081 20856
rect 10042 20748 10048 20800
rect 10100 20788 10106 20800
rect 10594 20788 10600 20800
rect 10100 20760 10600 20788
rect 10100 20748 10106 20760
rect 10594 20748 10600 20760
rect 10652 20788 10658 20800
rect 11072 20788 11100 20828
rect 12069 20825 12081 20828
rect 12115 20856 12127 20859
rect 12250 20856 12256 20868
rect 12115 20828 12256 20856
rect 12115 20825 12127 20828
rect 12069 20819 12127 20825
rect 12250 20816 12256 20828
rect 12308 20816 12314 20868
rect 14737 20859 14795 20865
rect 14737 20825 14749 20859
rect 14783 20856 14795 20859
rect 16316 20856 16344 20884
rect 14783 20828 16344 20856
rect 14783 20825 14795 20828
rect 14737 20819 14795 20825
rect 11330 20788 11336 20800
rect 10652 20760 11100 20788
rect 11291 20760 11336 20788
rect 10652 20748 10658 20760
rect 11330 20748 11336 20760
rect 11388 20788 11394 20800
rect 11974 20788 11980 20800
rect 11388 20760 11980 20788
rect 11388 20748 11394 20760
rect 11974 20748 11980 20760
rect 12032 20748 12038 20800
rect 13630 20788 13636 20800
rect 13591 20760 13636 20788
rect 13630 20748 13636 20760
rect 13688 20748 13694 20800
rect 15010 20788 15016 20800
rect 14971 20760 15016 20788
rect 15010 20748 15016 20760
rect 15068 20748 15074 20800
rect 15565 20791 15623 20797
rect 15565 20757 15577 20791
rect 15611 20788 15623 20791
rect 15654 20788 15660 20800
rect 15611 20760 15660 20788
rect 15611 20757 15623 20760
rect 15565 20751 15623 20757
rect 15654 20748 15660 20760
rect 15712 20748 15718 20800
rect 16301 20791 16359 20797
rect 16301 20757 16313 20791
rect 16347 20788 16359 20791
rect 16666 20788 16672 20800
rect 16347 20760 16672 20788
rect 16347 20757 16359 20760
rect 16301 20751 16359 20757
rect 16666 20748 16672 20760
rect 16724 20748 16730 20800
rect 19058 20748 19064 20800
rect 19116 20788 19122 20800
rect 19153 20791 19211 20797
rect 19153 20788 19165 20791
rect 19116 20760 19165 20788
rect 19116 20748 19122 20760
rect 19153 20757 19165 20760
rect 19199 20788 19211 20791
rect 19242 20788 19248 20800
rect 19199 20760 19248 20788
rect 19199 20757 19211 20760
rect 19153 20751 19211 20757
rect 19242 20748 19248 20760
rect 19300 20748 19306 20800
rect 23750 20788 23756 20800
rect 23711 20760 23756 20788
rect 23750 20748 23756 20760
rect 23808 20748 23814 20800
rect 1104 20698 28888 20720
rect 1104 20646 5982 20698
rect 6034 20646 6046 20698
rect 6098 20646 6110 20698
rect 6162 20646 6174 20698
rect 6226 20646 15982 20698
rect 16034 20646 16046 20698
rect 16098 20646 16110 20698
rect 16162 20646 16174 20698
rect 16226 20646 25982 20698
rect 26034 20646 26046 20698
rect 26098 20646 26110 20698
rect 26162 20646 26174 20698
rect 26226 20646 28888 20698
rect 1104 20624 28888 20646
rect 2041 20587 2099 20593
rect 2041 20553 2053 20587
rect 2087 20584 2099 20587
rect 2130 20584 2136 20596
rect 2087 20556 2136 20584
rect 2087 20553 2099 20556
rect 2041 20547 2099 20553
rect 2130 20544 2136 20556
rect 2188 20544 2194 20596
rect 9401 20587 9459 20593
rect 9401 20553 9413 20587
rect 9447 20584 9459 20587
rect 9490 20584 9496 20596
rect 9447 20556 9496 20584
rect 9447 20553 9459 20556
rect 9401 20547 9459 20553
rect 9490 20544 9496 20556
rect 9548 20544 9554 20596
rect 10134 20584 10140 20596
rect 10095 20556 10140 20584
rect 10134 20544 10140 20556
rect 10192 20544 10198 20596
rect 10226 20544 10232 20596
rect 10284 20584 10290 20596
rect 10870 20584 10876 20596
rect 10284 20556 10876 20584
rect 10284 20544 10290 20556
rect 10870 20544 10876 20556
rect 10928 20584 10934 20596
rect 11609 20587 11667 20593
rect 11609 20584 11621 20587
rect 10928 20556 11621 20584
rect 10928 20544 10934 20556
rect 11609 20553 11621 20556
rect 11655 20553 11667 20587
rect 11609 20547 11667 20553
rect 12253 20587 12311 20593
rect 12253 20553 12265 20587
rect 12299 20584 12311 20587
rect 12986 20584 12992 20596
rect 12299 20556 12992 20584
rect 12299 20553 12311 20556
rect 12253 20547 12311 20553
rect 12986 20544 12992 20556
rect 13044 20544 13050 20596
rect 15470 20584 15476 20596
rect 15431 20556 15476 20584
rect 15470 20544 15476 20556
rect 15528 20544 15534 20596
rect 16666 20584 16672 20596
rect 16408 20556 16672 20584
rect 10152 20448 10180 20544
rect 12618 20476 12624 20528
rect 12676 20516 12682 20528
rect 12805 20519 12863 20525
rect 12805 20516 12817 20519
rect 12676 20488 12817 20516
rect 12676 20476 12682 20488
rect 12805 20485 12817 20488
rect 12851 20485 12863 20519
rect 12805 20479 12863 20485
rect 13265 20519 13323 20525
rect 13265 20485 13277 20519
rect 13311 20516 13323 20519
rect 13722 20516 13728 20528
rect 13311 20488 13728 20516
rect 13311 20485 13323 20488
rect 13265 20479 13323 20485
rect 10686 20448 10692 20460
rect 10152 20420 10692 20448
rect 10686 20408 10692 20420
rect 10744 20448 10750 20460
rect 10873 20451 10931 20457
rect 10873 20448 10885 20451
rect 10744 20420 10885 20448
rect 10744 20408 10750 20420
rect 10873 20417 10885 20420
rect 10919 20417 10931 20451
rect 10873 20411 10931 20417
rect 10962 20340 10968 20392
rect 11020 20380 11026 20392
rect 11149 20383 11207 20389
rect 11149 20380 11161 20383
rect 11020 20352 11161 20380
rect 11020 20340 11026 20352
rect 11149 20349 11161 20352
rect 11195 20349 11207 20383
rect 11330 20380 11336 20392
rect 11291 20352 11336 20380
rect 11149 20343 11207 20349
rect 11330 20340 11336 20352
rect 11388 20340 11394 20392
rect 10318 20312 10324 20324
rect 10279 20284 10324 20312
rect 10318 20272 10324 20284
rect 10376 20272 10382 20324
rect 12820 20312 12848 20479
rect 13722 20476 13728 20488
rect 13780 20476 13786 20528
rect 12986 20408 12992 20460
rect 13044 20448 13050 20460
rect 13044 20420 13860 20448
rect 13044 20408 13050 20420
rect 13265 20383 13323 20389
rect 13265 20349 13277 20383
rect 13311 20380 13323 20383
rect 13446 20380 13452 20392
rect 13311 20352 13452 20380
rect 13311 20349 13323 20352
rect 13265 20343 13323 20349
rect 13446 20340 13452 20352
rect 13504 20340 13510 20392
rect 13630 20380 13636 20392
rect 13591 20352 13636 20380
rect 13630 20340 13636 20352
rect 13688 20340 13694 20392
rect 13832 20389 13860 20420
rect 16206 20408 16212 20460
rect 16264 20448 16270 20460
rect 16408 20457 16436 20556
rect 16666 20544 16672 20556
rect 16724 20584 16730 20596
rect 17402 20584 17408 20596
rect 16724 20556 17408 20584
rect 16724 20544 16730 20556
rect 17402 20544 17408 20556
rect 17460 20544 17466 20596
rect 17678 20544 17684 20596
rect 17736 20584 17742 20596
rect 17773 20587 17831 20593
rect 17773 20584 17785 20587
rect 17736 20556 17785 20584
rect 17736 20544 17742 20556
rect 17773 20553 17785 20556
rect 17819 20553 17831 20587
rect 17773 20547 17831 20553
rect 22833 20587 22891 20593
rect 22833 20553 22845 20587
rect 22879 20584 22891 20587
rect 22922 20584 22928 20596
rect 22879 20556 22928 20584
rect 22879 20553 22891 20556
rect 22833 20547 22891 20553
rect 16482 20476 16488 20528
rect 16540 20516 16546 20528
rect 16540 20488 16804 20516
rect 16540 20476 16546 20488
rect 16776 20457 16804 20488
rect 16393 20451 16451 20457
rect 16393 20448 16405 20451
rect 16264 20420 16405 20448
rect 16264 20408 16270 20420
rect 16393 20417 16405 20420
rect 16439 20417 16451 20451
rect 16393 20411 16451 20417
rect 16761 20451 16819 20457
rect 16761 20417 16773 20451
rect 16807 20417 16819 20451
rect 17788 20448 17816 20547
rect 22922 20544 22928 20556
rect 22980 20544 22986 20596
rect 18325 20519 18383 20525
rect 18325 20485 18337 20519
rect 18371 20516 18383 20519
rect 18506 20516 18512 20528
rect 18371 20488 18512 20516
rect 18371 20485 18383 20488
rect 18325 20479 18383 20485
rect 18506 20476 18512 20488
rect 18564 20476 18570 20528
rect 17788 20420 18920 20448
rect 16761 20411 16819 20417
rect 13817 20383 13875 20389
rect 13817 20349 13829 20383
rect 13863 20349 13875 20383
rect 14182 20380 14188 20392
rect 14143 20352 14188 20380
rect 13817 20343 13875 20349
rect 14182 20340 14188 20352
rect 14240 20340 14246 20392
rect 14553 20383 14611 20389
rect 14553 20349 14565 20383
rect 14599 20349 14611 20383
rect 14553 20343 14611 20349
rect 16485 20383 16543 20389
rect 16485 20349 16497 20383
rect 16531 20380 16543 20383
rect 16574 20380 16580 20392
rect 16531 20352 16580 20380
rect 16531 20349 16543 20352
rect 16485 20343 16543 20349
rect 14568 20312 14596 20343
rect 16574 20340 16580 20352
rect 16632 20340 16638 20392
rect 16850 20380 16856 20392
rect 16811 20352 16856 20380
rect 16850 20340 16856 20352
rect 16908 20340 16914 20392
rect 17497 20383 17555 20389
rect 17497 20349 17509 20383
rect 17543 20380 17555 20383
rect 18230 20380 18236 20392
rect 17543 20352 18236 20380
rect 17543 20349 17555 20352
rect 17497 20343 17555 20349
rect 18230 20340 18236 20352
rect 18288 20380 18294 20392
rect 18509 20383 18567 20389
rect 18509 20380 18521 20383
rect 18288 20352 18521 20380
rect 18288 20340 18294 20352
rect 18509 20349 18521 20352
rect 18555 20349 18567 20383
rect 18690 20380 18696 20392
rect 18651 20352 18696 20380
rect 18509 20343 18567 20349
rect 18690 20340 18696 20352
rect 18748 20340 18754 20392
rect 18892 20389 18920 20420
rect 18877 20383 18935 20389
rect 18877 20349 18889 20383
rect 18923 20349 18935 20383
rect 18877 20343 18935 20349
rect 12820 20284 14596 20312
rect 14826 20272 14832 20324
rect 14884 20312 14890 20324
rect 15841 20315 15899 20321
rect 15841 20312 15853 20315
rect 14884 20284 15853 20312
rect 14884 20272 14890 20284
rect 15841 20281 15853 20284
rect 15887 20281 15899 20315
rect 15841 20275 15899 20281
rect 1578 20244 1584 20256
rect 1539 20216 1584 20244
rect 1578 20204 1584 20216
rect 1636 20204 1642 20256
rect 9769 20247 9827 20253
rect 9769 20213 9781 20247
rect 9815 20244 9827 20247
rect 9858 20244 9864 20256
rect 9815 20216 9864 20244
rect 9815 20213 9827 20216
rect 9769 20207 9827 20213
rect 9858 20204 9864 20216
rect 9916 20204 9922 20256
rect 14642 20204 14648 20256
rect 14700 20244 14706 20256
rect 16758 20244 16764 20256
rect 14700 20216 16764 20244
rect 14700 20204 14706 20216
rect 16758 20204 16764 20216
rect 16816 20204 16822 20256
rect 22370 20244 22376 20256
rect 22331 20216 22376 20244
rect 22370 20204 22376 20216
rect 22428 20204 22434 20256
rect 1104 20154 28888 20176
rect 1104 20102 10982 20154
rect 11034 20102 11046 20154
rect 11098 20102 11110 20154
rect 11162 20102 11174 20154
rect 11226 20102 20982 20154
rect 21034 20102 21046 20154
rect 21098 20102 21110 20154
rect 21162 20102 21174 20154
rect 21226 20102 28888 20154
rect 1104 20080 28888 20102
rect 7466 20040 7472 20052
rect 7427 20012 7472 20040
rect 7466 20000 7472 20012
rect 7524 20000 7530 20052
rect 9953 20043 10011 20049
rect 9953 20009 9965 20043
rect 9999 20040 10011 20043
rect 10318 20040 10324 20052
rect 9999 20012 10324 20040
rect 9999 20009 10011 20012
rect 9953 20003 10011 20009
rect 10318 20000 10324 20012
rect 10376 20000 10382 20052
rect 10413 20043 10471 20049
rect 10413 20009 10425 20043
rect 10459 20040 10471 20043
rect 11330 20040 11336 20052
rect 10459 20012 11336 20040
rect 10459 20009 10471 20012
rect 10413 20003 10471 20009
rect 8757 19975 8815 19981
rect 8757 19941 8769 19975
rect 8803 19972 8815 19975
rect 10428 19972 10456 20003
rect 11330 20000 11336 20012
rect 11388 20000 11394 20052
rect 14185 20043 14243 20049
rect 14185 20040 14197 20043
rect 12728 20012 14197 20040
rect 8803 19944 10456 19972
rect 10781 19975 10839 19981
rect 8803 19941 8815 19944
rect 8757 19935 8815 19941
rect 10781 19941 10793 19975
rect 10827 19972 10839 19975
rect 10870 19972 10876 19984
rect 10827 19944 10876 19972
rect 10827 19941 10839 19944
rect 10781 19935 10839 19941
rect 10870 19932 10876 19944
rect 10928 19932 10934 19984
rect 12069 19975 12127 19981
rect 12069 19972 12081 19975
rect 11532 19944 12081 19972
rect 11532 19916 11560 19944
rect 12069 19941 12081 19944
rect 12115 19941 12127 19975
rect 12069 19935 12127 19941
rect 8202 19904 8208 19916
rect 8163 19876 8208 19904
rect 8202 19864 8208 19876
rect 8260 19864 8266 19916
rect 8297 19907 8355 19913
rect 8297 19873 8309 19907
rect 8343 19904 8355 19907
rect 8938 19904 8944 19916
rect 8343 19876 8944 19904
rect 8343 19873 8355 19876
rect 8297 19867 8355 19873
rect 8938 19864 8944 19876
rect 8996 19864 9002 19916
rect 11241 19907 11299 19913
rect 11241 19873 11253 19907
rect 11287 19904 11299 19907
rect 11514 19904 11520 19916
rect 11287 19876 11520 19904
rect 11287 19873 11299 19876
rect 11241 19867 11299 19873
rect 11514 19864 11520 19876
rect 11572 19864 11578 19916
rect 11609 19907 11667 19913
rect 11609 19873 11621 19907
rect 11655 19904 11667 19907
rect 12158 19904 12164 19916
rect 11655 19876 12164 19904
rect 11655 19873 11667 19876
rect 11609 19867 11667 19873
rect 12158 19864 12164 19876
rect 12216 19864 12222 19916
rect 12434 19864 12440 19916
rect 12492 19904 12498 19916
rect 12728 19913 12756 20012
rect 14185 20009 14197 20012
rect 14231 20009 14243 20043
rect 14185 20003 14243 20009
rect 14274 20000 14280 20052
rect 14332 20040 14338 20052
rect 14461 20043 14519 20049
rect 14461 20040 14473 20043
rect 14332 20012 14473 20040
rect 14332 20000 14338 20012
rect 14461 20009 14473 20012
rect 14507 20009 14519 20043
rect 14461 20003 14519 20009
rect 14734 20000 14740 20052
rect 14792 20040 14798 20052
rect 15473 20043 15531 20049
rect 15473 20040 15485 20043
rect 14792 20012 15485 20040
rect 14792 20000 14798 20012
rect 15473 20009 15485 20012
rect 15519 20009 15531 20043
rect 15473 20003 15531 20009
rect 15933 20043 15991 20049
rect 15933 20009 15945 20043
rect 15979 20040 15991 20043
rect 16482 20040 16488 20052
rect 15979 20012 16488 20040
rect 15979 20009 15991 20012
rect 15933 20003 15991 20009
rect 13170 19972 13176 19984
rect 13131 19944 13176 19972
rect 13170 19932 13176 19944
rect 13228 19932 13234 19984
rect 12713 19907 12771 19913
rect 12713 19904 12725 19907
rect 12492 19876 12725 19904
rect 12492 19864 12498 19876
rect 12713 19873 12725 19876
rect 12759 19873 12771 19907
rect 12713 19867 12771 19873
rect 12986 19864 12992 19916
rect 13044 19904 13050 19916
rect 13449 19907 13507 19913
rect 13449 19904 13461 19907
rect 13044 19876 13461 19904
rect 13044 19864 13050 19876
rect 13449 19873 13461 19876
rect 13495 19873 13507 19907
rect 13998 19904 14004 19916
rect 13911 19876 14004 19904
rect 13449 19867 13507 19873
rect 13998 19864 14004 19876
rect 14056 19904 14062 19916
rect 14752 19904 14780 20000
rect 15488 19972 15516 20003
rect 16482 20000 16488 20012
rect 16540 20000 16546 20052
rect 16574 19972 16580 19984
rect 15488 19944 16580 19972
rect 16574 19932 16580 19944
rect 16632 19932 16638 19984
rect 18966 19932 18972 19984
rect 19024 19972 19030 19984
rect 19518 19972 19524 19984
rect 19024 19944 19104 19972
rect 19479 19944 19524 19972
rect 19024 19932 19030 19944
rect 14056 19876 14780 19904
rect 15289 19907 15347 19913
rect 14056 19864 14062 19876
rect 15289 19873 15301 19907
rect 15335 19904 15347 19907
rect 15746 19904 15752 19916
rect 15335 19876 15752 19904
rect 15335 19873 15347 19876
rect 15289 19867 15347 19873
rect 15746 19864 15752 19876
rect 15804 19864 15810 19916
rect 16298 19864 16304 19916
rect 16356 19904 16362 19916
rect 16356 19876 16528 19904
rect 16356 19864 16362 19876
rect 16500 19848 16528 19876
rect 17402 19864 17408 19916
rect 17460 19904 17466 19916
rect 19076 19913 19104 19944
rect 19518 19932 19524 19944
rect 19576 19932 19582 19984
rect 19061 19907 19119 19913
rect 17460 19876 19012 19904
rect 17460 19864 17466 19876
rect 11422 19796 11428 19848
rect 11480 19836 11486 19848
rect 11701 19839 11759 19845
rect 11701 19836 11713 19839
rect 11480 19808 11713 19836
rect 11480 19796 11486 19808
rect 11701 19805 11713 19808
rect 11747 19805 11759 19839
rect 12618 19836 12624 19848
rect 12579 19808 12624 19836
rect 11701 19799 11759 19805
rect 12618 19796 12624 19808
rect 12676 19796 12682 19848
rect 16482 19836 16488 19848
rect 16443 19808 16488 19836
rect 16482 19796 16488 19808
rect 16540 19796 16546 19848
rect 16758 19836 16764 19848
rect 16719 19808 16764 19836
rect 16758 19796 16764 19808
rect 16816 19836 16822 19848
rect 18417 19839 18475 19845
rect 18417 19836 18429 19839
rect 16816 19808 18429 19836
rect 16816 19796 16822 19808
rect 18417 19805 18429 19808
rect 18463 19836 18475 19839
rect 18690 19836 18696 19848
rect 18463 19808 18696 19836
rect 18463 19805 18475 19808
rect 18417 19799 18475 19805
rect 18690 19796 18696 19808
rect 18748 19796 18754 19848
rect 18984 19845 19012 19876
rect 19061 19873 19073 19907
rect 19107 19873 19119 19907
rect 19061 19867 19119 19873
rect 18969 19839 19027 19845
rect 18969 19805 18981 19839
rect 19015 19836 19027 19839
rect 19242 19836 19248 19848
rect 19015 19808 19248 19836
rect 19015 19805 19027 19808
rect 18969 19799 19027 19805
rect 19242 19796 19248 19808
rect 19300 19796 19306 19848
rect 11238 19728 11244 19780
rect 11296 19768 11302 19780
rect 11606 19768 11612 19780
rect 11296 19740 11612 19768
rect 11296 19728 11302 19740
rect 11606 19728 11612 19740
rect 11664 19728 11670 19780
rect 12529 19771 12587 19777
rect 12529 19737 12541 19771
rect 12575 19768 12587 19771
rect 12894 19768 12900 19780
rect 12575 19740 12900 19768
rect 12575 19737 12587 19740
rect 12529 19731 12587 19737
rect 12894 19728 12900 19740
rect 12952 19768 12958 19780
rect 13170 19768 13176 19780
rect 12952 19740 13176 19768
rect 12952 19728 12958 19740
rect 13170 19728 13176 19740
rect 13228 19728 13234 19780
rect 7837 19703 7895 19709
rect 7837 19669 7849 19703
rect 7883 19700 7895 19703
rect 8110 19700 8116 19712
rect 7883 19672 8116 19700
rect 7883 19669 7895 19672
rect 7837 19663 7895 19669
rect 8110 19660 8116 19672
rect 8168 19660 8174 19712
rect 13446 19660 13452 19712
rect 13504 19700 13510 19712
rect 13817 19703 13875 19709
rect 13817 19700 13829 19703
rect 13504 19672 13829 19700
rect 13504 19660 13510 19672
rect 13817 19669 13829 19672
rect 13863 19669 13875 19703
rect 13817 19663 13875 19669
rect 14366 19660 14372 19712
rect 14424 19700 14430 19712
rect 14734 19700 14740 19712
rect 14424 19672 14740 19700
rect 14424 19660 14430 19672
rect 14734 19660 14740 19672
rect 14792 19700 14798 19712
rect 14829 19703 14887 19709
rect 14829 19700 14841 19703
rect 14792 19672 14841 19700
rect 14792 19660 14798 19672
rect 14829 19669 14841 19672
rect 14875 19669 14887 19703
rect 14829 19663 14887 19669
rect 16301 19703 16359 19709
rect 16301 19669 16313 19703
rect 16347 19700 16359 19703
rect 16850 19700 16856 19712
rect 16347 19672 16856 19700
rect 16347 19669 16359 19672
rect 16301 19663 16359 19669
rect 16850 19660 16856 19672
rect 16908 19660 16914 19712
rect 18049 19703 18107 19709
rect 18049 19669 18061 19703
rect 18095 19700 18107 19703
rect 18138 19700 18144 19712
rect 18095 19672 18144 19700
rect 18095 19669 18107 19672
rect 18049 19663 18107 19669
rect 18138 19660 18144 19672
rect 18196 19660 18202 19712
rect 1104 19610 28888 19632
rect 1104 19558 5982 19610
rect 6034 19558 6046 19610
rect 6098 19558 6110 19610
rect 6162 19558 6174 19610
rect 6226 19558 15982 19610
rect 16034 19558 16046 19610
rect 16098 19558 16110 19610
rect 16162 19558 16174 19610
rect 16226 19558 25982 19610
rect 26034 19558 26046 19610
rect 26098 19558 26110 19610
rect 26162 19558 26174 19610
rect 26226 19558 28888 19610
rect 1104 19536 28888 19558
rect 8938 19496 8944 19508
rect 8899 19468 8944 19496
rect 8938 19456 8944 19468
rect 8996 19456 9002 19508
rect 11425 19499 11483 19505
rect 11425 19465 11437 19499
rect 11471 19496 11483 19499
rect 11514 19496 11520 19508
rect 11471 19468 11520 19496
rect 11471 19465 11483 19468
rect 11425 19459 11483 19465
rect 11514 19456 11520 19468
rect 11572 19456 11578 19508
rect 11885 19499 11943 19505
rect 11885 19465 11897 19499
rect 11931 19496 11943 19499
rect 12158 19496 12164 19508
rect 11931 19468 12164 19496
rect 11931 19465 11943 19468
rect 11885 19459 11943 19465
rect 11057 19431 11115 19437
rect 11057 19397 11069 19431
rect 11103 19428 11115 19431
rect 11900 19428 11928 19459
rect 12158 19456 12164 19468
rect 12216 19456 12222 19508
rect 13998 19496 14004 19508
rect 13959 19468 14004 19496
rect 13998 19456 14004 19468
rect 14056 19456 14062 19508
rect 15381 19499 15439 19505
rect 15381 19465 15393 19499
rect 15427 19496 15439 19499
rect 15746 19496 15752 19508
rect 15427 19468 15752 19496
rect 15427 19465 15439 19468
rect 15381 19459 15439 19465
rect 15746 19456 15752 19468
rect 15804 19456 15810 19508
rect 16850 19496 16856 19508
rect 16811 19468 16856 19496
rect 16850 19456 16856 19468
rect 16908 19456 16914 19508
rect 17126 19456 17132 19508
rect 17184 19456 17190 19508
rect 18230 19456 18236 19508
rect 18288 19496 18294 19508
rect 18325 19499 18383 19505
rect 18325 19496 18337 19499
rect 18288 19468 18337 19496
rect 18288 19456 18294 19468
rect 18325 19465 18337 19468
rect 18371 19465 18383 19499
rect 18966 19496 18972 19508
rect 18927 19468 18972 19496
rect 18325 19459 18383 19465
rect 18966 19456 18972 19468
rect 19024 19456 19030 19508
rect 11103 19400 11928 19428
rect 11103 19397 11115 19400
rect 11057 19391 11115 19397
rect 7466 19320 7472 19372
rect 7524 19360 7530 19372
rect 7524 19332 8064 19360
rect 7524 19320 7530 19332
rect 7282 19292 7288 19304
rect 7243 19264 7288 19292
rect 7282 19252 7288 19264
rect 7340 19252 7346 19304
rect 8036 19301 8064 19332
rect 8110 19320 8116 19372
rect 8168 19360 8174 19372
rect 9490 19360 9496 19372
rect 8168 19332 9496 19360
rect 8168 19320 8174 19332
rect 9490 19320 9496 19332
rect 9548 19320 9554 19372
rect 10045 19363 10103 19369
rect 10045 19329 10057 19363
rect 10091 19360 10103 19363
rect 10318 19360 10324 19372
rect 10091 19332 10324 19360
rect 10091 19329 10103 19332
rect 10045 19323 10103 19329
rect 10318 19320 10324 19332
rect 10376 19320 10382 19372
rect 12434 19320 12440 19372
rect 12492 19360 12498 19372
rect 15473 19363 15531 19369
rect 12492 19332 12537 19360
rect 12492 19320 12498 19332
rect 15473 19329 15485 19363
rect 15519 19360 15531 19363
rect 16482 19360 16488 19372
rect 15519 19332 16488 19360
rect 15519 19329 15531 19332
rect 15473 19323 15531 19329
rect 16482 19320 16488 19332
rect 16540 19320 16546 19372
rect 16850 19320 16856 19372
rect 16908 19360 16914 19372
rect 17144 19360 17172 19456
rect 16908 19332 17172 19360
rect 16908 19320 16914 19332
rect 19242 19320 19248 19372
rect 19300 19320 19306 19372
rect 8021 19295 8079 19301
rect 8021 19261 8033 19295
rect 8067 19292 8079 19295
rect 8202 19292 8208 19304
rect 8067 19264 8208 19292
rect 8067 19261 8079 19264
rect 8021 19255 8079 19261
rect 8202 19252 8208 19264
rect 8260 19252 8266 19304
rect 8386 19252 8392 19304
rect 8444 19292 8450 19304
rect 8573 19295 8631 19301
rect 8444 19264 8489 19292
rect 8444 19252 8450 19264
rect 8573 19261 8585 19295
rect 8619 19261 8631 19295
rect 8573 19255 8631 19261
rect 7300 19224 7328 19252
rect 7300 19196 8386 19224
rect 6638 19156 6644 19168
rect 6599 19128 6644 19156
rect 6638 19116 6644 19128
rect 6696 19116 6702 19168
rect 7653 19159 7711 19165
rect 7653 19125 7665 19159
rect 7699 19156 7711 19159
rect 8018 19156 8024 19168
rect 7699 19128 8024 19156
rect 7699 19125 7711 19128
rect 7653 19119 7711 19125
rect 8018 19116 8024 19128
rect 8076 19116 8082 19168
rect 8358 19156 8386 19196
rect 8478 19156 8484 19168
rect 8358 19128 8484 19156
rect 8478 19116 8484 19128
rect 8536 19156 8542 19168
rect 8588 19156 8616 19255
rect 8938 19252 8944 19304
rect 8996 19292 9002 19304
rect 9306 19292 9312 19304
rect 8996 19264 9312 19292
rect 8996 19252 9002 19264
rect 9306 19252 9312 19264
rect 9364 19252 9370 19304
rect 10137 19295 10195 19301
rect 10137 19261 10149 19295
rect 10183 19292 10195 19295
rect 10226 19292 10232 19304
rect 10183 19264 10232 19292
rect 10183 19261 10195 19264
rect 10137 19255 10195 19261
rect 10226 19252 10232 19264
rect 10284 19252 10290 19304
rect 10505 19295 10563 19301
rect 10505 19261 10517 19295
rect 10551 19261 10563 19295
rect 10505 19255 10563 19261
rect 10597 19295 10655 19301
rect 10597 19261 10609 19295
rect 10643 19261 10655 19295
rect 10597 19255 10655 19261
rect 9490 19184 9496 19236
rect 9548 19224 9554 19236
rect 9548 19196 9904 19224
rect 9548 19184 9554 19196
rect 9766 19156 9772 19168
rect 8536 19128 8616 19156
rect 9727 19128 9772 19156
rect 8536 19116 8542 19128
rect 9766 19116 9772 19128
rect 9824 19116 9830 19168
rect 9876 19156 9904 19196
rect 9950 19184 9956 19236
rect 10008 19224 10014 19236
rect 10520 19224 10548 19255
rect 10008 19196 10548 19224
rect 10008 19184 10014 19196
rect 10042 19156 10048 19168
rect 9876 19128 10048 19156
rect 10042 19116 10048 19128
rect 10100 19156 10106 19168
rect 10612 19156 10640 19255
rect 12158 19252 12164 19304
rect 12216 19292 12222 19304
rect 12894 19292 12900 19304
rect 12216 19264 12664 19292
rect 12855 19264 12900 19292
rect 12216 19252 12222 19264
rect 11146 19184 11152 19236
rect 11204 19184 11210 19236
rect 12250 19224 12256 19236
rect 12211 19196 12256 19224
rect 12250 19184 12256 19196
rect 12308 19184 12314 19236
rect 12636 19224 12664 19264
rect 12894 19252 12900 19264
rect 12952 19252 12958 19304
rect 13078 19292 13084 19304
rect 13039 19264 13084 19292
rect 13078 19252 13084 19264
rect 13136 19252 13142 19304
rect 13265 19295 13323 19301
rect 13265 19261 13277 19295
rect 13311 19261 13323 19295
rect 13265 19255 13323 19261
rect 13280 19224 13308 19255
rect 14366 19252 14372 19304
rect 14424 19292 14430 19304
rect 14461 19295 14519 19301
rect 14461 19292 14473 19295
rect 14424 19264 14473 19292
rect 14424 19252 14430 19264
rect 14461 19261 14473 19264
rect 14507 19292 14519 19295
rect 14737 19295 14795 19301
rect 14737 19292 14749 19295
rect 14507 19264 14749 19292
rect 14507 19261 14519 19264
rect 14461 19255 14519 19261
rect 14737 19261 14749 19264
rect 14783 19261 14795 19295
rect 14737 19255 14795 19261
rect 15102 19252 15108 19304
rect 15160 19292 15166 19304
rect 15749 19295 15807 19301
rect 15749 19292 15761 19295
rect 15160 19264 15761 19292
rect 15160 19252 15166 19264
rect 15749 19261 15761 19264
rect 15795 19292 15807 19295
rect 16206 19292 16212 19304
rect 15795 19264 16212 19292
rect 15795 19261 15807 19264
rect 15749 19255 15807 19261
rect 16206 19252 16212 19264
rect 16264 19252 16270 19304
rect 16500 19292 16528 19320
rect 17402 19292 17408 19304
rect 16500 19264 17408 19292
rect 17402 19252 17408 19264
rect 17460 19252 17466 19304
rect 18049 19295 18107 19301
rect 18049 19292 18061 19295
rect 17788 19264 18061 19292
rect 12636 19196 13308 19224
rect 10100 19128 10640 19156
rect 11164 19156 11192 19184
rect 12636 19168 12664 19196
rect 17788 19168 17816 19264
rect 18049 19261 18061 19264
rect 18095 19261 18107 19295
rect 18049 19255 18107 19261
rect 18138 19252 18144 19304
rect 18196 19292 18202 19304
rect 19260 19292 19288 19320
rect 19337 19295 19395 19301
rect 19337 19292 19349 19295
rect 18196 19264 18241 19292
rect 19260 19264 19349 19292
rect 18196 19252 18202 19264
rect 19337 19261 19349 19264
rect 19383 19292 19395 19295
rect 19426 19292 19432 19304
rect 19383 19264 19432 19292
rect 19383 19261 19395 19264
rect 19337 19255 19395 19261
rect 19426 19252 19432 19264
rect 19484 19252 19490 19304
rect 12158 19156 12164 19168
rect 11164 19128 12164 19156
rect 10100 19116 10106 19128
rect 12158 19116 12164 19128
rect 12216 19116 12222 19168
rect 12618 19116 12624 19168
rect 12676 19116 12682 19168
rect 12894 19116 12900 19168
rect 12952 19156 12958 19168
rect 14642 19156 14648 19168
rect 12952 19128 14648 19156
rect 12952 19116 12958 19128
rect 14642 19116 14648 19128
rect 14700 19116 14706 19168
rect 14737 19159 14795 19165
rect 14737 19125 14749 19159
rect 14783 19156 14795 19159
rect 15013 19159 15071 19165
rect 15013 19156 15025 19159
rect 14783 19128 15025 19156
rect 14783 19125 14795 19128
rect 14737 19119 14795 19125
rect 15013 19125 15025 19128
rect 15059 19156 15071 19159
rect 15562 19156 15568 19168
rect 15059 19128 15568 19156
rect 15059 19125 15071 19128
rect 15013 19119 15071 19125
rect 15562 19116 15568 19128
rect 15620 19116 15626 19168
rect 16758 19116 16764 19168
rect 16816 19156 16822 19168
rect 17405 19159 17463 19165
rect 17405 19156 17417 19159
rect 16816 19128 17417 19156
rect 16816 19116 16822 19128
rect 17405 19125 17417 19128
rect 17451 19125 17463 19159
rect 17770 19156 17776 19168
rect 17731 19128 17776 19156
rect 17405 19119 17463 19125
rect 17770 19116 17776 19128
rect 17828 19116 17834 19168
rect 1104 19066 28888 19088
rect 1104 19014 10982 19066
rect 11034 19014 11046 19066
rect 11098 19014 11110 19066
rect 11162 19014 11174 19066
rect 11226 19014 20982 19066
rect 21034 19014 21046 19066
rect 21098 19014 21110 19066
rect 21162 19014 21174 19066
rect 21226 19014 28888 19066
rect 1104 18992 28888 19014
rect 6638 18912 6644 18964
rect 6696 18952 6702 18964
rect 8386 18952 8392 18964
rect 6696 18924 8392 18952
rect 6696 18912 6702 18924
rect 8386 18912 8392 18924
rect 8444 18952 8450 18964
rect 8481 18955 8539 18961
rect 8481 18952 8493 18955
rect 8444 18924 8493 18952
rect 8444 18912 8450 18924
rect 8481 18921 8493 18924
rect 8527 18921 8539 18955
rect 9950 18952 9956 18964
rect 9911 18924 9956 18952
rect 8481 18915 8539 18921
rect 9950 18912 9956 18924
rect 10008 18912 10014 18964
rect 10778 18952 10784 18964
rect 10739 18924 10784 18952
rect 10778 18912 10784 18924
rect 10836 18912 10842 18964
rect 12621 18955 12679 18961
rect 12621 18921 12633 18955
rect 12667 18952 12679 18955
rect 12710 18952 12716 18964
rect 12667 18924 12716 18952
rect 12667 18921 12679 18924
rect 12621 18915 12679 18921
rect 12710 18912 12716 18924
rect 12768 18912 12774 18964
rect 13078 18912 13084 18964
rect 13136 18952 13142 18964
rect 14001 18955 14059 18961
rect 14001 18952 14013 18955
rect 13136 18924 14013 18952
rect 13136 18912 13142 18924
rect 14001 18921 14013 18924
rect 14047 18921 14059 18955
rect 14001 18915 14059 18921
rect 14182 18912 14188 18964
rect 14240 18952 14246 18964
rect 14829 18955 14887 18961
rect 14829 18952 14841 18955
rect 14240 18924 14841 18952
rect 14240 18912 14246 18924
rect 14829 18921 14841 18924
rect 14875 18952 14887 18955
rect 15010 18952 15016 18964
rect 14875 18924 15016 18952
rect 14875 18921 14887 18924
rect 14829 18915 14887 18921
rect 15010 18912 15016 18924
rect 15068 18912 15074 18964
rect 15746 18952 15752 18964
rect 15707 18924 15752 18952
rect 15746 18912 15752 18924
rect 15804 18912 15810 18964
rect 16206 18912 16212 18964
rect 16264 18952 16270 18964
rect 16301 18955 16359 18961
rect 16301 18952 16313 18955
rect 16264 18924 16313 18952
rect 16264 18912 16270 18924
rect 16301 18921 16313 18924
rect 16347 18921 16359 18955
rect 18138 18952 18144 18964
rect 18099 18924 18144 18952
rect 16301 18915 16359 18921
rect 18138 18912 18144 18924
rect 18196 18912 18202 18964
rect 12529 18887 12587 18893
rect 12529 18853 12541 18887
rect 12575 18884 12587 18887
rect 13446 18884 13452 18896
rect 12575 18856 13452 18884
rect 12575 18853 12587 18856
rect 12529 18847 12587 18853
rect 13446 18844 13452 18856
rect 13504 18844 13510 18896
rect 7190 18776 7196 18828
rect 7248 18816 7254 18828
rect 7377 18819 7435 18825
rect 7377 18816 7389 18819
rect 7248 18788 7389 18816
rect 7248 18776 7254 18788
rect 7377 18785 7389 18788
rect 7423 18816 7435 18819
rect 8110 18816 8116 18828
rect 7423 18788 8116 18816
rect 7423 18785 7435 18788
rect 7377 18779 7435 18785
rect 8110 18776 8116 18788
rect 8168 18776 8174 18828
rect 10870 18776 10876 18828
rect 10928 18816 10934 18828
rect 11333 18819 11391 18825
rect 11333 18816 11345 18819
rect 10928 18788 11345 18816
rect 10928 18776 10934 18788
rect 11333 18785 11345 18788
rect 11379 18785 11391 18819
rect 11698 18816 11704 18828
rect 11659 18788 11704 18816
rect 11333 18779 11391 18785
rect 11698 18776 11704 18788
rect 11756 18776 11762 18828
rect 12434 18776 12440 18828
rect 12492 18816 12498 18828
rect 13541 18819 13599 18825
rect 13541 18816 13553 18819
rect 12492 18788 13553 18816
rect 12492 18776 12498 18788
rect 13541 18785 13553 18788
rect 13587 18785 13599 18819
rect 13541 18779 13599 18785
rect 15933 18819 15991 18825
rect 15933 18785 15945 18819
rect 15979 18816 15991 18819
rect 16298 18816 16304 18828
rect 15979 18788 16304 18816
rect 15979 18785 15991 18788
rect 15933 18779 15991 18785
rect 16298 18776 16304 18788
rect 16356 18776 16362 18828
rect 16574 18776 16580 18828
rect 16632 18816 16638 18828
rect 16945 18819 17003 18825
rect 16945 18816 16957 18819
rect 16632 18788 16957 18816
rect 16632 18776 16638 18788
rect 16945 18785 16957 18788
rect 16991 18816 17003 18819
rect 17678 18816 17684 18828
rect 16991 18788 17684 18816
rect 16991 18785 17003 18788
rect 16945 18779 17003 18785
rect 17678 18776 17684 18788
rect 17736 18776 17742 18828
rect 7098 18748 7104 18760
rect 7059 18720 7104 18748
rect 7098 18708 7104 18720
rect 7156 18708 7162 18760
rect 11422 18748 11428 18760
rect 11383 18720 11428 18748
rect 11422 18708 11428 18720
rect 11480 18708 11486 18760
rect 11609 18751 11667 18757
rect 11609 18717 11621 18751
rect 11655 18717 11667 18751
rect 12710 18748 12716 18760
rect 12671 18720 12716 18748
rect 11609 18711 11667 18717
rect 10502 18640 10508 18692
rect 10560 18680 10566 18692
rect 11624 18680 11652 18711
rect 12710 18708 12716 18720
rect 12768 18708 12774 18760
rect 13170 18708 13176 18760
rect 13228 18748 13234 18760
rect 13265 18751 13323 18757
rect 13265 18748 13277 18751
rect 13228 18720 13277 18748
rect 13228 18708 13234 18720
rect 13265 18717 13277 18720
rect 13311 18717 13323 18751
rect 13722 18748 13728 18760
rect 13683 18720 13728 18748
rect 13265 18711 13323 18717
rect 13722 18708 13728 18720
rect 13780 18708 13786 18760
rect 16853 18751 16911 18757
rect 16853 18748 16865 18751
rect 16500 18720 16865 18748
rect 10560 18652 11652 18680
rect 10560 18640 10566 18652
rect 3326 18572 3332 18624
rect 3384 18612 3390 18624
rect 9401 18615 9459 18621
rect 9401 18612 9413 18615
rect 3384 18584 9413 18612
rect 3384 18572 3390 18584
rect 9401 18581 9413 18584
rect 9447 18612 9459 18615
rect 9490 18612 9496 18624
rect 9447 18584 9496 18612
rect 9447 18581 9459 18584
rect 9401 18575 9459 18581
rect 9490 18572 9496 18584
rect 9548 18572 9554 18624
rect 10226 18612 10232 18624
rect 10187 18584 10232 18612
rect 10226 18572 10232 18584
rect 10284 18572 10290 18624
rect 11624 18612 11652 18652
rect 12434 18640 12440 18692
rect 12492 18680 12498 18692
rect 12621 18683 12679 18689
rect 12621 18680 12633 18683
rect 12492 18652 12633 18680
rect 12492 18640 12498 18652
rect 12621 18649 12633 18652
rect 12667 18680 12679 18683
rect 14369 18683 14427 18689
rect 14369 18680 14381 18683
rect 12667 18652 14381 18680
rect 12667 18649 12679 18652
rect 12621 18643 12679 18649
rect 14369 18649 14381 18652
rect 14415 18680 14427 18683
rect 15102 18680 15108 18692
rect 14415 18652 15108 18680
rect 14415 18649 14427 18652
rect 14369 18643 14427 18649
rect 15102 18640 15108 18652
rect 15160 18640 15166 18692
rect 16500 18624 16528 18720
rect 16853 18717 16865 18720
rect 16899 18717 16911 18751
rect 16853 18711 16911 18717
rect 16482 18612 16488 18624
rect 11624 18584 16488 18612
rect 16482 18572 16488 18584
rect 16540 18572 16546 18624
rect 16574 18572 16580 18624
rect 16632 18612 16638 18624
rect 16669 18615 16727 18621
rect 16669 18612 16681 18615
rect 16632 18584 16681 18612
rect 16632 18572 16638 18584
rect 16669 18581 16681 18584
rect 16715 18581 16727 18615
rect 17126 18612 17132 18624
rect 17087 18584 17132 18612
rect 16669 18575 16727 18581
rect 17126 18572 17132 18584
rect 17184 18572 17190 18624
rect 17402 18572 17408 18624
rect 17460 18612 17466 18624
rect 17681 18615 17739 18621
rect 17681 18612 17693 18615
rect 17460 18584 17693 18612
rect 17460 18572 17466 18584
rect 17681 18581 17693 18584
rect 17727 18581 17739 18615
rect 17681 18575 17739 18581
rect 1104 18522 28888 18544
rect 1104 18470 5982 18522
rect 6034 18470 6046 18522
rect 6098 18470 6110 18522
rect 6162 18470 6174 18522
rect 6226 18470 15982 18522
rect 16034 18470 16046 18522
rect 16098 18470 16110 18522
rect 16162 18470 16174 18522
rect 16226 18470 25982 18522
rect 26034 18470 26046 18522
rect 26098 18470 26110 18522
rect 26162 18470 26174 18522
rect 26226 18470 28888 18522
rect 1104 18448 28888 18470
rect 3237 18411 3295 18417
rect 3237 18377 3249 18411
rect 3283 18408 3295 18411
rect 3326 18408 3332 18420
rect 3283 18380 3332 18408
rect 3283 18377 3295 18380
rect 3237 18371 3295 18377
rect 3326 18368 3332 18380
rect 3384 18368 3390 18420
rect 7098 18368 7104 18420
rect 7156 18408 7162 18420
rect 7561 18411 7619 18417
rect 7561 18408 7573 18411
rect 7156 18380 7573 18408
rect 7156 18368 7162 18380
rect 7561 18377 7573 18380
rect 7607 18408 7619 18411
rect 7834 18408 7840 18420
rect 7607 18380 7840 18408
rect 7607 18377 7619 18380
rect 7561 18371 7619 18377
rect 7834 18368 7840 18380
rect 7892 18408 7898 18420
rect 8294 18408 8300 18420
rect 7892 18380 8300 18408
rect 7892 18368 7898 18380
rect 8294 18368 8300 18380
rect 8352 18368 8358 18420
rect 8662 18368 8668 18420
rect 8720 18408 8726 18420
rect 9217 18411 9275 18417
rect 9217 18408 9229 18411
rect 8720 18380 9229 18408
rect 8720 18368 8726 18380
rect 9217 18377 9229 18380
rect 9263 18377 9275 18411
rect 9217 18371 9275 18377
rect 7190 18340 7196 18352
rect 7151 18312 7196 18340
rect 7190 18300 7196 18312
rect 7248 18300 7254 18352
rect 9232 18340 9260 18371
rect 9950 18368 9956 18420
rect 10008 18408 10014 18420
rect 11057 18411 11115 18417
rect 11057 18408 11069 18411
rect 10008 18380 11069 18408
rect 10008 18368 10014 18380
rect 11057 18377 11069 18380
rect 11103 18408 11115 18411
rect 11698 18408 11704 18420
rect 11103 18380 11704 18408
rect 11103 18377 11115 18380
rect 11057 18371 11115 18377
rect 11698 18368 11704 18380
rect 11756 18368 11762 18420
rect 11974 18368 11980 18420
rect 12032 18408 12038 18420
rect 12161 18411 12219 18417
rect 12161 18408 12173 18411
rect 12032 18380 12173 18408
rect 12032 18368 12038 18380
rect 12161 18377 12173 18380
rect 12207 18408 12219 18411
rect 13722 18408 13728 18420
rect 12207 18380 13728 18408
rect 12207 18377 12219 18380
rect 12161 18371 12219 18377
rect 13722 18368 13728 18380
rect 13780 18368 13786 18420
rect 14366 18408 14372 18420
rect 14327 18380 14372 18408
rect 14366 18368 14372 18380
rect 14424 18368 14430 18420
rect 16298 18408 16304 18420
rect 16259 18380 16304 18408
rect 16298 18368 16304 18380
rect 16356 18408 16362 18420
rect 17037 18411 17095 18417
rect 17037 18408 17049 18411
rect 16356 18380 17049 18408
rect 16356 18368 16362 18380
rect 17037 18377 17049 18380
rect 17083 18377 17095 18411
rect 17310 18408 17316 18420
rect 17271 18380 17316 18408
rect 17037 18371 17095 18377
rect 17310 18368 17316 18380
rect 17368 18368 17374 18420
rect 17678 18408 17684 18420
rect 17639 18380 17684 18408
rect 17678 18368 17684 18380
rect 17736 18368 17742 18420
rect 9232 18312 10364 18340
rect 10336 18284 10364 18312
rect 10686 18300 10692 18352
rect 10744 18340 10750 18352
rect 11793 18343 11851 18349
rect 11793 18340 11805 18343
rect 10744 18312 11805 18340
rect 10744 18300 10750 18312
rect 11793 18309 11805 18312
rect 11839 18340 11851 18343
rect 13170 18340 13176 18352
rect 11839 18312 13176 18340
rect 11839 18309 11851 18312
rect 11793 18303 11851 18309
rect 13170 18300 13176 18312
rect 13228 18300 13234 18352
rect 15746 18340 15752 18352
rect 14844 18312 15752 18340
rect 9306 18232 9312 18284
rect 9364 18272 9370 18284
rect 9674 18272 9680 18284
rect 9364 18244 9680 18272
rect 9364 18232 9370 18244
rect 9674 18232 9680 18244
rect 9732 18232 9738 18284
rect 9769 18275 9827 18281
rect 9769 18241 9781 18275
rect 9815 18272 9827 18275
rect 10226 18272 10232 18284
rect 9815 18244 10232 18272
rect 9815 18241 9827 18244
rect 9769 18235 9827 18241
rect 10226 18232 10232 18244
rect 10284 18232 10290 18284
rect 10318 18232 10324 18284
rect 10376 18272 10382 18284
rect 10781 18275 10839 18281
rect 10781 18272 10793 18275
rect 10376 18244 10469 18272
rect 10520 18244 10793 18272
rect 10376 18232 10382 18244
rect 1854 18204 1860 18216
rect 1815 18176 1860 18204
rect 1854 18164 1860 18176
rect 1912 18164 1918 18216
rect 2133 18207 2191 18213
rect 2133 18204 2145 18207
rect 1964 18176 2145 18204
rect 1486 18028 1492 18080
rect 1544 18068 1550 18080
rect 1673 18071 1731 18077
rect 1673 18068 1685 18071
rect 1544 18040 1685 18068
rect 1544 18028 1550 18040
rect 1673 18037 1685 18040
rect 1719 18068 1731 18071
rect 1964 18068 1992 18176
rect 2133 18173 2145 18176
rect 2179 18173 2191 18207
rect 2133 18167 2191 18173
rect 8941 18207 8999 18213
rect 8941 18173 8953 18207
rect 8987 18204 8999 18207
rect 9582 18204 9588 18216
rect 8987 18176 9588 18204
rect 8987 18173 8999 18176
rect 8941 18167 8999 18173
rect 9582 18164 9588 18176
rect 9640 18164 9646 18216
rect 9692 18204 9720 18232
rect 10520 18204 10548 18244
rect 10781 18241 10793 18244
rect 10827 18241 10839 18275
rect 10781 18235 10839 18241
rect 12989 18275 13047 18281
rect 12989 18241 13001 18275
rect 13035 18272 13047 18275
rect 13188 18272 13216 18300
rect 13725 18275 13783 18281
rect 13725 18272 13737 18275
rect 13035 18244 13737 18272
rect 13035 18241 13047 18244
rect 12989 18235 13047 18241
rect 13725 18241 13737 18244
rect 13771 18241 13783 18275
rect 13725 18235 13783 18241
rect 9692 18176 10548 18204
rect 10597 18207 10655 18213
rect 10597 18173 10609 18207
rect 10643 18173 10655 18207
rect 10597 18167 10655 18173
rect 1719 18040 1992 18068
rect 9677 18071 9735 18077
rect 1719 18037 1731 18040
rect 1673 18031 1731 18037
rect 9677 18037 9689 18071
rect 9723 18068 9735 18071
rect 10612 18068 10640 18167
rect 11422 18164 11428 18216
rect 11480 18204 11486 18216
rect 12437 18207 12495 18213
rect 12437 18204 12449 18207
rect 11480 18176 12449 18204
rect 11480 18164 11486 18176
rect 12437 18173 12449 18176
rect 12483 18173 12495 18207
rect 12437 18167 12495 18173
rect 13265 18207 13323 18213
rect 13265 18173 13277 18207
rect 13311 18173 13323 18207
rect 13446 18204 13452 18216
rect 13407 18176 13452 18204
rect 13265 18167 13323 18173
rect 11238 18096 11244 18148
rect 11296 18096 11302 18148
rect 11517 18139 11575 18145
rect 11517 18105 11529 18139
rect 11563 18136 11575 18139
rect 13280 18136 13308 18167
rect 13446 18164 13452 18176
rect 13504 18164 13510 18216
rect 14642 18164 14648 18216
rect 14700 18204 14706 18216
rect 14844 18213 14872 18312
rect 15746 18300 15752 18312
rect 15804 18300 15810 18352
rect 16482 18300 16488 18352
rect 16540 18340 16546 18352
rect 16669 18343 16727 18349
rect 16669 18340 16681 18343
rect 16540 18312 16681 18340
rect 16540 18300 16546 18312
rect 16669 18309 16681 18312
rect 16715 18309 16727 18343
rect 16669 18303 16727 18309
rect 15010 18272 15016 18284
rect 14971 18244 15016 18272
rect 15010 18232 15016 18244
rect 15068 18232 15074 18284
rect 16574 18272 16580 18284
rect 15212 18244 16580 18272
rect 14829 18207 14887 18213
rect 14829 18204 14841 18207
rect 14700 18176 14841 18204
rect 14700 18164 14706 18176
rect 14829 18173 14841 18176
rect 14875 18173 14887 18207
rect 14829 18167 14887 18173
rect 15102 18164 15108 18216
rect 15160 18204 15166 18216
rect 15212 18213 15240 18244
rect 16574 18232 16580 18244
rect 16632 18232 16638 18284
rect 15197 18207 15255 18213
rect 15197 18204 15209 18207
rect 15160 18176 15209 18204
rect 15160 18164 15166 18176
rect 15197 18173 15209 18176
rect 15243 18173 15255 18207
rect 15197 18167 15255 18173
rect 15381 18207 15439 18213
rect 15381 18173 15393 18207
rect 15427 18173 15439 18207
rect 15381 18167 15439 18173
rect 13538 18136 13544 18148
rect 11563 18108 13544 18136
rect 11563 18105 11575 18108
rect 11517 18099 11575 18105
rect 13538 18096 13544 18108
rect 13596 18096 13602 18148
rect 11256 18068 11284 18096
rect 11698 18068 11704 18080
rect 9723 18040 11704 18068
rect 9723 18037 9735 18040
rect 9677 18031 9735 18037
rect 11698 18028 11704 18040
rect 11756 18028 11762 18080
rect 11974 18028 11980 18080
rect 12032 18068 12038 18080
rect 14734 18068 14740 18080
rect 12032 18040 14740 18068
rect 12032 18028 12038 18040
rect 14734 18028 14740 18040
rect 14792 18068 14798 18080
rect 15396 18068 15424 18167
rect 15562 18164 15568 18216
rect 15620 18204 15626 18216
rect 15749 18207 15807 18213
rect 15749 18204 15761 18207
rect 15620 18176 15761 18204
rect 15620 18164 15626 18176
rect 15749 18173 15761 18176
rect 15795 18173 15807 18207
rect 15749 18167 15807 18173
rect 16853 18207 16911 18213
rect 16853 18173 16865 18207
rect 16899 18204 16911 18207
rect 17310 18204 17316 18216
rect 16899 18176 17316 18204
rect 16899 18173 16911 18176
rect 16853 18167 16911 18173
rect 17310 18164 17316 18176
rect 17368 18164 17374 18216
rect 14792 18040 15424 18068
rect 14792 18028 14798 18040
rect 1104 17978 28888 18000
rect 1104 17926 10982 17978
rect 11034 17926 11046 17978
rect 11098 17926 11110 17978
rect 11162 17926 11174 17978
rect 11226 17926 20982 17978
rect 21034 17926 21046 17978
rect 21098 17926 21110 17978
rect 21162 17926 21174 17978
rect 21226 17926 28888 17978
rect 1104 17904 28888 17926
rect 8294 17864 8300 17876
rect 8255 17836 8300 17864
rect 8294 17824 8300 17836
rect 8352 17824 8358 17876
rect 9125 17867 9183 17873
rect 9125 17833 9137 17867
rect 9171 17864 9183 17867
rect 9306 17864 9312 17876
rect 9171 17836 9312 17864
rect 9171 17833 9183 17836
rect 9125 17827 9183 17833
rect 9306 17824 9312 17836
rect 9364 17824 9370 17876
rect 11422 17824 11428 17876
rect 11480 17864 11486 17876
rect 11609 17867 11667 17873
rect 11609 17864 11621 17867
rect 11480 17836 11621 17864
rect 11480 17824 11486 17836
rect 11609 17833 11621 17836
rect 11655 17833 11667 17867
rect 11609 17827 11667 17833
rect 12253 17867 12311 17873
rect 12253 17833 12265 17867
rect 12299 17864 12311 17867
rect 12342 17864 12348 17876
rect 12299 17836 12348 17864
rect 12299 17833 12311 17836
rect 12253 17827 12311 17833
rect 12342 17824 12348 17836
rect 12400 17824 12406 17876
rect 13538 17864 13544 17876
rect 13499 17836 13544 17864
rect 13538 17824 13544 17836
rect 13596 17824 13602 17876
rect 14642 17864 14648 17876
rect 14603 17836 14648 17864
rect 14642 17824 14648 17836
rect 14700 17824 14706 17876
rect 15562 17864 15568 17876
rect 15523 17836 15568 17864
rect 15562 17824 15568 17836
rect 15620 17824 15626 17876
rect 16298 17824 16304 17876
rect 16356 17824 16362 17876
rect 16482 17824 16488 17876
rect 16540 17864 16546 17876
rect 16761 17867 16819 17873
rect 16761 17864 16773 17867
rect 16540 17836 16773 17864
rect 16540 17824 16546 17836
rect 16761 17833 16773 17836
rect 16807 17833 16819 17867
rect 16761 17827 16819 17833
rect 17954 17824 17960 17876
rect 18012 17864 18018 17876
rect 18693 17867 18751 17873
rect 18693 17864 18705 17867
rect 18012 17836 18705 17864
rect 18012 17824 18018 17836
rect 18693 17833 18705 17836
rect 18739 17833 18751 17867
rect 18693 17827 18751 17833
rect 9674 17756 9680 17808
rect 9732 17796 9738 17808
rect 10321 17799 10379 17805
rect 10321 17796 10333 17799
rect 9732 17768 10333 17796
rect 9732 17756 9738 17768
rect 10321 17765 10333 17768
rect 10367 17796 10379 17799
rect 10870 17796 10876 17808
rect 10367 17768 10876 17796
rect 10367 17765 10379 17768
rect 10321 17759 10379 17765
rect 10870 17756 10876 17768
rect 10928 17756 10934 17808
rect 13722 17796 13728 17808
rect 12544 17768 13728 17796
rect 12544 17740 12572 17768
rect 13722 17756 13728 17768
rect 13780 17756 13786 17808
rect 16316 17796 16344 17824
rect 15948 17768 16344 17796
rect 11146 17728 11152 17740
rect 11107 17700 11152 17728
rect 11146 17688 11152 17700
rect 11204 17688 11210 17740
rect 12526 17728 12532 17740
rect 12439 17700 12532 17728
rect 12526 17688 12532 17700
rect 12584 17688 12590 17740
rect 12986 17688 12992 17740
rect 13044 17728 13050 17740
rect 13081 17731 13139 17737
rect 13081 17728 13093 17731
rect 13044 17700 13093 17728
rect 13044 17688 13050 17700
rect 13081 17697 13093 17700
rect 13127 17697 13139 17731
rect 13262 17728 13268 17740
rect 13175 17700 13268 17728
rect 13081 17691 13139 17697
rect 13262 17688 13268 17700
rect 13320 17728 13326 17740
rect 15948 17737 15976 17768
rect 15105 17731 15163 17737
rect 15105 17728 15117 17731
rect 13320 17700 15117 17728
rect 13320 17688 13326 17700
rect 15105 17697 15117 17700
rect 15151 17728 15163 17731
rect 15933 17731 15991 17737
rect 15151 17700 15884 17728
rect 15151 17697 15163 17700
rect 15105 17691 15163 17697
rect 5166 17620 5172 17672
rect 5224 17660 5230 17672
rect 9401 17663 9459 17669
rect 9401 17660 9413 17663
rect 5224 17632 9413 17660
rect 5224 17620 5230 17632
rect 9401 17629 9413 17632
rect 9447 17660 9459 17663
rect 9582 17660 9588 17672
rect 9447 17632 9588 17660
rect 9447 17629 9459 17632
rect 9401 17623 9459 17629
rect 9582 17620 9588 17632
rect 9640 17620 9646 17672
rect 10318 17620 10324 17672
rect 10376 17660 10382 17672
rect 10873 17663 10931 17669
rect 10873 17660 10885 17663
rect 10376 17632 10885 17660
rect 10376 17620 10382 17632
rect 10873 17629 10885 17632
rect 10919 17629 10931 17663
rect 11330 17660 11336 17672
rect 11291 17632 11336 17660
rect 10873 17623 10931 17629
rect 11330 17620 11336 17632
rect 11388 17620 11394 17672
rect 12158 17620 12164 17672
rect 12216 17660 12222 17672
rect 12345 17663 12403 17669
rect 12345 17660 12357 17663
rect 12216 17632 12357 17660
rect 12216 17620 12222 17632
rect 12345 17629 12357 17632
rect 12391 17660 12403 17663
rect 12618 17660 12624 17672
rect 12391 17632 12624 17660
rect 12391 17629 12403 17632
rect 12345 17623 12403 17629
rect 12618 17620 12624 17632
rect 12676 17620 12682 17672
rect 14185 17663 14243 17669
rect 14185 17629 14197 17663
rect 14231 17660 14243 17663
rect 15010 17660 15016 17672
rect 14231 17632 15016 17660
rect 14231 17629 14243 17632
rect 14185 17623 14243 17629
rect 15010 17620 15016 17632
rect 15068 17620 15074 17672
rect 15746 17660 15752 17672
rect 15707 17632 15752 17660
rect 15746 17620 15752 17632
rect 15804 17620 15810 17672
rect 15856 17660 15884 17700
rect 15933 17697 15945 17731
rect 15979 17697 15991 17731
rect 15933 17691 15991 17697
rect 16301 17731 16359 17737
rect 16301 17697 16313 17731
rect 16347 17728 16359 17731
rect 16482 17728 16488 17740
rect 16347 17700 16488 17728
rect 16347 17697 16359 17700
rect 16301 17691 16359 17697
rect 16482 17688 16488 17700
rect 16540 17688 16546 17740
rect 17402 17688 17408 17740
rect 17460 17728 17466 17740
rect 17589 17731 17647 17737
rect 17589 17728 17601 17731
rect 17460 17700 17601 17728
rect 17460 17688 17466 17700
rect 17589 17697 17601 17700
rect 17635 17697 17647 17731
rect 17589 17691 17647 17697
rect 16209 17663 16267 17669
rect 16209 17660 16221 17663
rect 15856 17632 16221 17660
rect 16209 17629 16221 17632
rect 16255 17629 16267 17663
rect 16209 17623 16267 17629
rect 17313 17663 17371 17669
rect 17313 17629 17325 17663
rect 17359 17629 17371 17663
rect 17313 17623 17371 17629
rect 10229 17595 10287 17601
rect 10229 17561 10241 17595
rect 10275 17592 10287 17595
rect 10778 17592 10784 17604
rect 10275 17564 10784 17592
rect 10275 17561 10287 17564
rect 10229 17555 10287 17561
rect 10778 17552 10784 17564
rect 10836 17552 10842 17604
rect 17328 17536 17356 17623
rect 1946 17524 1952 17536
rect 1907 17496 1952 17524
rect 1946 17484 1952 17496
rect 2004 17484 2010 17536
rect 17221 17527 17279 17533
rect 17221 17493 17233 17527
rect 17267 17524 17279 17527
rect 17310 17524 17316 17536
rect 17267 17496 17316 17524
rect 17267 17493 17279 17496
rect 17221 17487 17279 17493
rect 17310 17484 17316 17496
rect 17368 17484 17374 17536
rect 1104 17434 28888 17456
rect 1104 17382 5982 17434
rect 6034 17382 6046 17434
rect 6098 17382 6110 17434
rect 6162 17382 6174 17434
rect 6226 17382 15982 17434
rect 16034 17382 16046 17434
rect 16098 17382 16110 17434
rect 16162 17382 16174 17434
rect 16226 17382 25982 17434
rect 26034 17382 26046 17434
rect 26098 17382 26110 17434
rect 26162 17382 26174 17434
rect 26226 17382 28888 17434
rect 1104 17360 28888 17382
rect 2774 17280 2780 17332
rect 2832 17320 2838 17332
rect 8481 17323 8539 17329
rect 2832 17292 2877 17320
rect 2832 17280 2838 17292
rect 8481 17289 8493 17323
rect 8527 17320 8539 17323
rect 9398 17320 9404 17332
rect 8527 17292 9404 17320
rect 8527 17289 8539 17292
rect 8481 17283 8539 17289
rect 9398 17280 9404 17292
rect 9456 17280 9462 17332
rect 9861 17323 9919 17329
rect 9861 17289 9873 17323
rect 9907 17320 9919 17323
rect 9950 17320 9956 17332
rect 9907 17292 9956 17320
rect 9907 17289 9919 17292
rect 9861 17283 9919 17289
rect 9950 17280 9956 17292
rect 10008 17320 10014 17332
rect 10686 17320 10692 17332
rect 10008 17292 10692 17320
rect 10008 17280 10014 17292
rect 10686 17280 10692 17292
rect 10744 17320 10750 17332
rect 11885 17323 11943 17329
rect 10744 17292 11376 17320
rect 10744 17280 10750 17292
rect 8570 17212 8576 17264
rect 8628 17252 8634 17264
rect 8628 17224 9168 17252
rect 8628 17212 8634 17224
rect 1670 17184 1676 17196
rect 1631 17156 1676 17184
rect 1670 17144 1676 17156
rect 1728 17144 1734 17196
rect 8294 17144 8300 17196
rect 8352 17184 8358 17196
rect 8352 17156 8892 17184
rect 8352 17144 8358 17156
rect 1397 17119 1455 17125
rect 1397 17085 1409 17119
rect 1443 17116 1455 17119
rect 1946 17116 1952 17128
rect 1443 17088 1952 17116
rect 1443 17085 1455 17088
rect 1397 17079 1455 17085
rect 1946 17076 1952 17088
rect 2004 17076 2010 17128
rect 8864 17125 8892 17156
rect 8938 17144 8944 17196
rect 8996 17184 9002 17196
rect 9140 17193 9168 17224
rect 9674 17212 9680 17264
rect 9732 17252 9738 17264
rect 10137 17255 10195 17261
rect 10137 17252 10149 17255
rect 9732 17224 10149 17252
rect 9732 17212 9738 17224
rect 10137 17221 10149 17224
rect 10183 17252 10195 17255
rect 10226 17252 10232 17264
rect 10183 17224 10232 17252
rect 10183 17221 10195 17224
rect 10137 17215 10195 17221
rect 10226 17212 10232 17224
rect 10284 17252 10290 17264
rect 11146 17252 11152 17264
rect 10284 17224 11152 17252
rect 10284 17212 10290 17224
rect 11146 17212 11152 17224
rect 11204 17212 11210 17264
rect 9125 17187 9183 17193
rect 8996 17156 9041 17184
rect 8996 17144 9002 17156
rect 9125 17153 9137 17187
rect 9171 17153 9183 17187
rect 10778 17184 10784 17196
rect 10739 17156 10784 17184
rect 9125 17147 9183 17153
rect 10778 17144 10784 17156
rect 10836 17144 10842 17196
rect 11238 17184 11244 17196
rect 11199 17156 11244 17184
rect 11238 17144 11244 17156
rect 11296 17144 11302 17196
rect 8849 17119 8907 17125
rect 8849 17085 8861 17119
rect 8895 17085 8907 17119
rect 8849 17079 8907 17085
rect 9217 17119 9275 17125
rect 9217 17085 9229 17119
rect 9263 17085 9275 17119
rect 9217 17079 9275 17085
rect 7745 17051 7803 17057
rect 7745 17017 7757 17051
rect 7791 17048 7803 17051
rect 9232 17048 9260 17079
rect 10134 17076 10140 17128
rect 10192 17116 10198 17128
rect 10594 17116 10600 17128
rect 10192 17088 10600 17116
rect 10192 17076 10198 17088
rect 10594 17076 10600 17088
rect 10652 17076 10658 17128
rect 10870 17076 10876 17128
rect 10928 17116 10934 17128
rect 11348 17125 11376 17292
rect 11885 17289 11897 17323
rect 11931 17320 11943 17323
rect 12158 17320 12164 17332
rect 11931 17292 12164 17320
rect 11931 17289 11943 17292
rect 11885 17283 11943 17289
rect 12158 17280 12164 17292
rect 12216 17280 12222 17332
rect 12253 17323 12311 17329
rect 12253 17289 12265 17323
rect 12299 17320 12311 17323
rect 12986 17320 12992 17332
rect 12299 17292 12992 17320
rect 12299 17289 12311 17292
rect 12253 17283 12311 17289
rect 12986 17280 12992 17292
rect 13044 17280 13050 17332
rect 13814 17280 13820 17332
rect 13872 17320 13878 17332
rect 14001 17323 14059 17329
rect 14001 17320 14013 17323
rect 13872 17292 14013 17320
rect 13872 17280 13878 17292
rect 14001 17289 14013 17292
rect 14047 17320 14059 17323
rect 14458 17320 14464 17332
rect 14047 17292 14464 17320
rect 14047 17289 14059 17292
rect 14001 17283 14059 17289
rect 14458 17280 14464 17292
rect 14516 17280 14522 17332
rect 15289 17323 15347 17329
rect 15289 17289 15301 17323
rect 15335 17320 15347 17323
rect 15378 17320 15384 17332
rect 15335 17292 15384 17320
rect 15335 17289 15347 17292
rect 15289 17283 15347 17289
rect 15378 17280 15384 17292
rect 15436 17280 15442 17332
rect 15562 17280 15568 17332
rect 15620 17320 15626 17332
rect 15749 17323 15807 17329
rect 15749 17320 15761 17323
rect 15620 17292 15761 17320
rect 15620 17280 15626 17292
rect 15749 17289 15761 17292
rect 15795 17289 15807 17323
rect 15749 17283 15807 17289
rect 16209 17323 16267 17329
rect 16209 17289 16221 17323
rect 16255 17320 16267 17323
rect 16298 17320 16304 17332
rect 16255 17292 16304 17320
rect 16255 17289 16267 17292
rect 16209 17283 16267 17289
rect 15764 17252 15792 17283
rect 16298 17280 16304 17292
rect 16356 17280 16362 17332
rect 16482 17252 16488 17264
rect 15764 17224 16488 17252
rect 16482 17212 16488 17224
rect 16540 17212 16546 17264
rect 14182 17184 14188 17196
rect 14143 17156 14188 17184
rect 14182 17144 14188 17156
rect 14240 17144 14246 17196
rect 16301 17187 16359 17193
rect 16301 17153 16313 17187
rect 16347 17184 16359 17187
rect 16574 17184 16580 17196
rect 16347 17156 16580 17184
rect 16347 17153 16359 17156
rect 16301 17147 16359 17153
rect 16574 17144 16580 17156
rect 16632 17144 16638 17196
rect 16853 17187 16911 17193
rect 16853 17153 16865 17187
rect 16899 17184 16911 17187
rect 16942 17184 16948 17196
rect 16899 17156 16948 17184
rect 16899 17153 16911 17156
rect 16853 17147 16911 17153
rect 16942 17144 16948 17156
rect 17000 17144 17006 17196
rect 10965 17119 11023 17125
rect 10965 17116 10977 17119
rect 10928 17088 10977 17116
rect 10928 17076 10934 17088
rect 10965 17085 10977 17088
rect 11011 17085 11023 17119
rect 10965 17079 11023 17085
rect 11333 17119 11391 17125
rect 11333 17085 11345 17119
rect 11379 17085 11391 17119
rect 12710 17116 12716 17128
rect 12671 17088 12716 17116
rect 11333 17079 11391 17085
rect 12710 17076 12716 17088
rect 12768 17076 12774 17128
rect 13633 17119 13691 17125
rect 13633 17085 13645 17119
rect 13679 17116 13691 17119
rect 14274 17116 14280 17128
rect 13679 17088 14280 17116
rect 13679 17085 13691 17088
rect 13633 17079 13691 17085
rect 14274 17076 14280 17088
rect 14332 17076 14338 17128
rect 14458 17076 14464 17128
rect 14516 17116 14522 17128
rect 14829 17119 14887 17125
rect 14829 17116 14841 17119
rect 14516 17088 14841 17116
rect 14516 17076 14522 17088
rect 14829 17085 14841 17088
rect 14875 17085 14887 17119
rect 15010 17116 15016 17128
rect 14923 17088 15016 17116
rect 14829 17079 14887 17085
rect 15010 17076 15016 17088
rect 15068 17116 15074 17128
rect 15746 17116 15752 17128
rect 15068 17088 15752 17116
rect 15068 17076 15074 17088
rect 15746 17076 15752 17088
rect 15804 17076 15810 17128
rect 16393 17119 16451 17125
rect 16393 17085 16405 17119
rect 16439 17085 16451 17119
rect 17402 17116 17408 17128
rect 17363 17088 17408 17116
rect 16393 17079 16451 17085
rect 9674 17048 9680 17060
rect 7791 17020 9680 17048
rect 7791 17017 7803 17020
rect 7745 17011 7803 17017
rect 9674 17008 9680 17020
rect 9732 17008 9738 17060
rect 13265 17051 13323 17057
rect 13265 17017 13277 17051
rect 13311 17048 13323 17051
rect 15028 17048 15056 17076
rect 16408 17048 16436 17079
rect 17402 17076 17408 17088
rect 17460 17076 17466 17128
rect 16666 17048 16672 17060
rect 13311 17020 15056 17048
rect 15672 17020 16672 17048
rect 13311 17017 13323 17020
rect 13265 17011 13323 17017
rect 8113 16983 8171 16989
rect 8113 16949 8125 16983
rect 8159 16980 8171 16983
rect 8938 16980 8944 16992
rect 8159 16952 8944 16980
rect 8159 16949 8171 16952
rect 8113 16943 8171 16949
rect 8938 16940 8944 16952
rect 8996 16980 9002 16992
rect 9766 16980 9772 16992
rect 8996 16952 9772 16980
rect 8996 16940 9002 16952
rect 9766 16940 9772 16952
rect 9824 16940 9830 16992
rect 10594 16980 10600 16992
rect 10555 16952 10600 16980
rect 10594 16940 10600 16952
rect 10652 16940 10658 16992
rect 14274 16940 14280 16992
rect 14332 16980 14338 16992
rect 15672 16980 15700 17020
rect 16666 17008 16672 17020
rect 16724 17008 16730 17060
rect 14332 16952 15700 16980
rect 14332 16940 14338 16952
rect 17310 16940 17316 16992
rect 17368 16980 17374 16992
rect 17773 16983 17831 16989
rect 17773 16980 17785 16983
rect 17368 16952 17785 16980
rect 17368 16940 17374 16952
rect 17773 16949 17785 16952
rect 17819 16980 17831 16983
rect 18046 16980 18052 16992
rect 17819 16952 18052 16980
rect 17819 16949 17831 16952
rect 17773 16943 17831 16949
rect 18046 16940 18052 16952
rect 18104 16940 18110 16992
rect 1104 16890 28888 16912
rect 1104 16838 10982 16890
rect 11034 16838 11046 16890
rect 11098 16838 11110 16890
rect 11162 16838 11174 16890
rect 11226 16838 20982 16890
rect 21034 16838 21046 16890
rect 21098 16838 21110 16890
rect 21162 16838 21174 16890
rect 21226 16838 28888 16890
rect 1104 16816 28888 16838
rect 1670 16776 1676 16788
rect 1631 16748 1676 16776
rect 1670 16736 1676 16748
rect 1728 16736 1734 16788
rect 8297 16779 8355 16785
rect 8297 16745 8309 16779
rect 8343 16776 8355 16779
rect 8478 16776 8484 16788
rect 8343 16748 8484 16776
rect 8343 16745 8355 16748
rect 8297 16739 8355 16745
rect 8478 16736 8484 16748
rect 8536 16736 8542 16788
rect 9490 16776 9496 16788
rect 9451 16748 9496 16776
rect 9490 16736 9496 16748
rect 9548 16736 9554 16788
rect 10318 16776 10324 16788
rect 10279 16748 10324 16776
rect 10318 16736 10324 16748
rect 10376 16776 10382 16788
rect 10778 16776 10784 16788
rect 10376 16748 10784 16776
rect 10376 16736 10382 16748
rect 10778 16736 10784 16748
rect 10836 16776 10842 16788
rect 12437 16779 12495 16785
rect 10836 16748 11284 16776
rect 10836 16736 10842 16748
rect 7745 16711 7803 16717
rect 7745 16677 7757 16711
rect 7791 16708 7803 16711
rect 9306 16708 9312 16720
rect 7791 16680 9312 16708
rect 7791 16677 7803 16680
rect 7745 16671 7803 16677
rect 9306 16668 9312 16680
rect 9364 16668 9370 16720
rect 10045 16711 10103 16717
rect 10045 16677 10057 16711
rect 10091 16708 10103 16711
rect 10689 16711 10747 16717
rect 10689 16708 10701 16711
rect 10091 16680 10701 16708
rect 10091 16677 10103 16680
rect 10045 16671 10103 16677
rect 10689 16677 10701 16680
rect 10735 16708 10747 16711
rect 10870 16708 10876 16720
rect 10735 16680 10876 16708
rect 10735 16677 10747 16680
rect 10689 16671 10747 16677
rect 10870 16668 10876 16680
rect 10928 16668 10934 16720
rect 5810 16600 5816 16652
rect 5868 16640 5874 16652
rect 11256 16649 11284 16748
rect 12437 16745 12449 16779
rect 12483 16776 12495 16779
rect 13262 16776 13268 16788
rect 12483 16748 13268 16776
rect 12483 16745 12495 16748
rect 12437 16739 12495 16745
rect 13262 16736 13268 16748
rect 13320 16736 13326 16788
rect 14737 16779 14795 16785
rect 14737 16745 14749 16779
rect 14783 16776 14795 16779
rect 15562 16776 15568 16788
rect 14783 16748 15568 16776
rect 14783 16745 14795 16748
rect 14737 16739 14795 16745
rect 15562 16736 15568 16748
rect 15620 16736 15626 16788
rect 16666 16776 16672 16788
rect 16627 16748 16672 16776
rect 16666 16736 16672 16748
rect 16724 16736 16730 16788
rect 23658 16776 23664 16788
rect 23619 16748 23664 16776
rect 23658 16736 23664 16748
rect 23716 16736 23722 16788
rect 11698 16668 11704 16720
rect 11756 16668 11762 16720
rect 12066 16708 12072 16720
rect 11979 16680 12072 16708
rect 12066 16668 12072 16680
rect 12124 16708 12130 16720
rect 12710 16708 12716 16720
rect 12124 16680 12716 16708
rect 12124 16668 12130 16680
rect 12710 16668 12716 16680
rect 12768 16668 12774 16720
rect 13173 16711 13231 16717
rect 13173 16677 13185 16711
rect 13219 16708 13231 16711
rect 15010 16708 15016 16720
rect 13219 16680 14136 16708
rect 14971 16680 15016 16708
rect 13219 16677 13231 16680
rect 13173 16671 13231 16677
rect 6365 16643 6423 16649
rect 6365 16640 6377 16643
rect 5868 16612 6377 16640
rect 5868 16600 5874 16612
rect 6365 16609 6377 16612
rect 6411 16609 6423 16643
rect 6365 16603 6423 16609
rect 11241 16643 11299 16649
rect 11241 16609 11253 16643
rect 11287 16609 11299 16643
rect 11517 16643 11575 16649
rect 11517 16640 11529 16643
rect 11241 16603 11299 16609
rect 11348 16612 11529 16640
rect 11348 16584 11376 16612
rect 11517 16609 11529 16612
rect 11563 16640 11575 16643
rect 11716 16640 11744 16668
rect 14108 16652 14136 16680
rect 15010 16668 15016 16680
rect 15068 16668 15074 16720
rect 15102 16668 15108 16720
rect 15160 16708 15166 16720
rect 15160 16680 16160 16708
rect 15160 16668 15166 16680
rect 11563 16612 11744 16640
rect 11563 16609 11575 16612
rect 11517 16603 11575 16609
rect 12526 16600 12532 16652
rect 12584 16640 12590 16652
rect 12805 16643 12863 16649
rect 12805 16640 12817 16643
rect 12584 16612 12817 16640
rect 12584 16600 12590 16612
rect 12805 16609 12817 16612
rect 12851 16609 12863 16643
rect 13814 16640 13820 16652
rect 13775 16612 13820 16640
rect 12805 16603 12863 16609
rect 13814 16600 13820 16612
rect 13872 16600 13878 16652
rect 14090 16640 14096 16652
rect 14051 16612 14096 16640
rect 14090 16600 14096 16612
rect 14148 16600 14154 16652
rect 15470 16640 15476 16652
rect 15431 16612 15476 16640
rect 15470 16600 15476 16612
rect 15528 16600 15534 16652
rect 15838 16640 15844 16652
rect 15799 16612 15844 16640
rect 15838 16600 15844 16612
rect 15896 16600 15902 16652
rect 16132 16649 16160 16680
rect 16117 16643 16175 16649
rect 16117 16609 16129 16643
rect 16163 16640 16175 16643
rect 16574 16640 16580 16652
rect 16163 16612 16580 16640
rect 16163 16609 16175 16612
rect 16117 16603 16175 16609
rect 16574 16600 16580 16612
rect 16632 16600 16638 16652
rect 16758 16600 16764 16652
rect 16816 16640 16822 16652
rect 17221 16643 17279 16649
rect 17221 16640 17233 16643
rect 16816 16612 17233 16640
rect 16816 16600 16822 16612
rect 17221 16609 17233 16612
rect 17267 16640 17279 16643
rect 17310 16640 17316 16652
rect 17267 16612 17316 16640
rect 17267 16609 17279 16612
rect 17221 16603 17279 16609
rect 17310 16600 17316 16612
rect 17368 16600 17374 16652
rect 22281 16643 22339 16649
rect 22281 16609 22293 16643
rect 22327 16640 22339 16643
rect 22327 16612 22784 16640
rect 22327 16609 22339 16612
rect 22281 16603 22339 16609
rect 22756 16584 22784 16612
rect 6089 16575 6147 16581
rect 6089 16541 6101 16575
rect 6135 16572 6147 16575
rect 6546 16572 6552 16584
rect 6135 16544 6552 16572
rect 6135 16541 6147 16544
rect 6089 16535 6147 16541
rect 6546 16532 6552 16544
rect 6604 16532 6610 16584
rect 11330 16532 11336 16584
rect 11388 16532 11394 16584
rect 11701 16575 11759 16581
rect 11701 16541 11713 16575
rect 11747 16572 11759 16575
rect 11974 16572 11980 16584
rect 11747 16544 11980 16572
rect 11747 16541 11759 16544
rect 11701 16535 11759 16541
rect 11974 16532 11980 16544
rect 12032 16532 12038 16584
rect 13446 16572 13452 16584
rect 13407 16544 13452 16572
rect 13446 16532 13452 16544
rect 13504 16532 13510 16584
rect 14369 16575 14427 16581
rect 14369 16541 14381 16575
rect 14415 16572 14427 16575
rect 14642 16572 14648 16584
rect 14415 16544 14648 16572
rect 14415 16541 14427 16544
rect 14369 16535 14427 16541
rect 14642 16532 14648 16544
rect 14700 16532 14706 16584
rect 22462 16532 22468 16584
rect 22520 16572 22526 16584
rect 22557 16575 22615 16581
rect 22557 16572 22569 16575
rect 22520 16544 22569 16572
rect 22520 16532 22526 16544
rect 22557 16541 22569 16544
rect 22603 16541 22615 16575
rect 22557 16535 22615 16541
rect 22738 16532 22744 16584
rect 22796 16532 22802 16584
rect 1946 16396 1952 16448
rect 2004 16436 2010 16448
rect 2041 16439 2099 16445
rect 2041 16436 2053 16439
rect 2004 16408 2053 16436
rect 2004 16396 2010 16408
rect 2041 16405 2053 16408
rect 2087 16436 2099 16439
rect 3418 16436 3424 16448
rect 2087 16408 3424 16436
rect 2087 16405 2099 16408
rect 2041 16399 2099 16405
rect 3418 16396 3424 16408
rect 3476 16396 3482 16448
rect 17402 16436 17408 16448
rect 17363 16408 17408 16436
rect 17402 16396 17408 16408
rect 17460 16396 17466 16448
rect 1104 16346 28888 16368
rect 1104 16294 5982 16346
rect 6034 16294 6046 16346
rect 6098 16294 6110 16346
rect 6162 16294 6174 16346
rect 6226 16294 15982 16346
rect 16034 16294 16046 16346
rect 16098 16294 16110 16346
rect 16162 16294 16174 16346
rect 16226 16294 25982 16346
rect 26034 16294 26046 16346
rect 26098 16294 26110 16346
rect 26162 16294 26174 16346
rect 26226 16294 28888 16346
rect 1104 16272 28888 16294
rect 4985 16235 5043 16241
rect 4985 16201 4997 16235
rect 5031 16232 5043 16235
rect 5166 16232 5172 16244
rect 5031 16204 5172 16232
rect 5031 16201 5043 16204
rect 4985 16195 5043 16201
rect 5166 16192 5172 16204
rect 5224 16192 5230 16244
rect 6549 16235 6607 16241
rect 6549 16201 6561 16235
rect 6595 16232 6607 16235
rect 6638 16232 6644 16244
rect 6595 16204 6644 16232
rect 6595 16201 6607 16204
rect 6549 16195 6607 16201
rect 6638 16192 6644 16204
rect 6696 16232 6702 16244
rect 7834 16232 7840 16244
rect 6696 16204 7840 16232
rect 6696 16192 6702 16204
rect 7834 16192 7840 16204
rect 7892 16192 7898 16244
rect 9674 16232 9680 16244
rect 9635 16204 9680 16232
rect 9674 16192 9680 16204
rect 9732 16192 9738 16244
rect 10686 16192 10692 16244
rect 10744 16232 10750 16244
rect 10965 16235 11023 16241
rect 10965 16232 10977 16235
rect 10744 16204 10977 16232
rect 10744 16192 10750 16204
rect 10965 16201 10977 16204
rect 11011 16201 11023 16235
rect 10965 16195 11023 16201
rect 13814 16192 13820 16244
rect 13872 16232 13878 16244
rect 14001 16235 14059 16241
rect 14001 16232 14013 16235
rect 13872 16204 14013 16232
rect 13872 16192 13878 16204
rect 14001 16201 14013 16204
rect 14047 16201 14059 16235
rect 14001 16195 14059 16201
rect 15838 16192 15844 16244
rect 15896 16232 15902 16244
rect 16393 16235 16451 16241
rect 16393 16232 16405 16235
rect 15896 16204 16405 16232
rect 15896 16192 15902 16204
rect 16393 16201 16405 16204
rect 16439 16201 16451 16235
rect 16393 16195 16451 16201
rect 16574 16192 16580 16244
rect 16632 16232 16638 16244
rect 16761 16235 16819 16241
rect 16761 16232 16773 16235
rect 16632 16204 16773 16232
rect 16632 16192 16638 16204
rect 16761 16201 16773 16204
rect 16807 16201 16819 16235
rect 17310 16232 17316 16244
rect 17271 16204 17316 16232
rect 16761 16195 16819 16201
rect 17310 16192 17316 16204
rect 17368 16192 17374 16244
rect 19613 16235 19671 16241
rect 19613 16201 19625 16235
rect 19659 16232 19671 16235
rect 19702 16232 19708 16244
rect 19659 16204 19708 16232
rect 19659 16201 19671 16204
rect 19613 16195 19671 16201
rect 19702 16192 19708 16204
rect 19760 16192 19766 16244
rect 10597 16167 10655 16173
rect 10597 16133 10609 16167
rect 10643 16164 10655 16167
rect 10778 16164 10784 16176
rect 10643 16136 10784 16164
rect 10643 16133 10655 16136
rect 10597 16127 10655 16133
rect 10778 16124 10784 16136
rect 10836 16124 10842 16176
rect 15286 16124 15292 16176
rect 15344 16164 15350 16176
rect 16025 16167 16083 16173
rect 16025 16164 16037 16167
rect 15344 16136 16037 16164
rect 15344 16124 15350 16136
rect 16025 16133 16037 16136
rect 16071 16133 16083 16167
rect 16025 16127 16083 16133
rect 3329 16099 3387 16105
rect 3329 16065 3341 16099
rect 3375 16096 3387 16099
rect 8205 16099 8263 16105
rect 3375 16068 3740 16096
rect 3375 16065 3387 16068
rect 3329 16059 3387 16065
rect 3712 16040 3740 16068
rect 8205 16065 8217 16099
rect 8251 16096 8263 16099
rect 8251 16068 8616 16096
rect 8251 16065 8263 16068
rect 8205 16059 8263 16065
rect 3418 16028 3424 16040
rect 3379 16000 3424 16028
rect 3418 15988 3424 16000
rect 3476 15988 3482 16040
rect 3694 16028 3700 16040
rect 3655 16000 3700 16028
rect 3694 15988 3700 16000
rect 3752 15988 3758 16040
rect 7834 15988 7840 16040
rect 7892 16028 7898 16040
rect 8588 16037 8616 16068
rect 8297 16031 8355 16037
rect 8297 16028 8309 16031
rect 7892 16000 8309 16028
rect 7892 15988 7898 16000
rect 8297 15997 8309 16000
rect 8343 15997 8355 16031
rect 8297 15991 8355 15997
rect 8573 16031 8631 16037
rect 8573 15997 8585 16031
rect 8619 16028 8631 16031
rect 9582 16028 9588 16040
rect 8619 16000 9588 16028
rect 8619 15997 8631 16000
rect 8573 15991 8631 15997
rect 9582 15988 9588 16000
rect 9640 15988 9646 16040
rect 10134 15988 10140 16040
rect 10192 16028 10198 16040
rect 10778 16028 10784 16040
rect 10192 16000 10784 16028
rect 10192 15988 10198 16000
rect 10778 15988 10784 16000
rect 10836 16028 10842 16040
rect 11609 16031 11667 16037
rect 11609 16028 11621 16031
rect 10836 16000 11621 16028
rect 10836 15988 10842 16000
rect 11609 15997 11621 16000
rect 11655 15997 11667 16031
rect 11609 15991 11667 15997
rect 12253 16031 12311 16037
rect 12253 15997 12265 16031
rect 12299 16028 12311 16031
rect 12897 16031 12955 16037
rect 12897 16028 12909 16031
rect 12299 16000 12909 16028
rect 12299 15997 12311 16000
rect 12253 15991 12311 15997
rect 12897 15997 12909 16000
rect 12943 16028 12955 16031
rect 13078 16028 13084 16040
rect 12943 16000 13084 16028
rect 12943 15997 12955 16000
rect 12897 15991 12955 15997
rect 13078 15988 13084 16000
rect 13136 15988 13142 16040
rect 14645 16031 14703 16037
rect 14645 15997 14657 16031
rect 14691 15997 14703 16031
rect 14645 15991 14703 15997
rect 10321 15963 10379 15969
rect 10321 15929 10333 15963
rect 10367 15960 10379 15963
rect 11974 15960 11980 15972
rect 10367 15932 11980 15960
rect 10367 15929 10379 15932
rect 10321 15923 10379 15929
rect 11974 15920 11980 15932
rect 12032 15920 12038 15972
rect 13357 15963 13415 15969
rect 13357 15929 13369 15963
rect 13403 15960 13415 15963
rect 13446 15960 13452 15972
rect 13403 15932 13452 15960
rect 13403 15929 13415 15932
rect 13357 15923 13415 15929
rect 13446 15920 13452 15932
rect 13504 15960 13510 15972
rect 13633 15963 13691 15969
rect 13633 15960 13645 15963
rect 13504 15932 13645 15960
rect 13504 15920 13510 15932
rect 13633 15929 13645 15932
rect 13679 15929 13691 15963
rect 13633 15923 13691 15929
rect 13814 15920 13820 15972
rect 13872 15960 13878 15972
rect 14461 15963 14519 15969
rect 14461 15960 14473 15963
rect 13872 15932 14473 15960
rect 13872 15920 13878 15932
rect 14461 15929 14473 15932
rect 14507 15960 14519 15963
rect 14660 15960 14688 15991
rect 14734 15988 14740 16040
rect 14792 16028 14798 16040
rect 15105 16031 15163 16037
rect 15105 16028 15117 16031
rect 14792 16000 15117 16028
rect 14792 15988 14798 16000
rect 15105 15997 15117 16000
rect 15151 15997 15163 16031
rect 15562 16028 15568 16040
rect 15523 16000 15568 16028
rect 15105 15991 15163 15997
rect 15562 15988 15568 16000
rect 15620 15988 15626 16040
rect 15838 16028 15844 16040
rect 15799 16000 15844 16028
rect 15838 15988 15844 16000
rect 15896 15988 15902 16040
rect 18046 16028 18052 16040
rect 18007 16000 18052 16028
rect 18046 15988 18052 16000
rect 18104 15988 18110 16040
rect 18325 16031 18383 16037
rect 18325 16028 18337 16031
rect 18156 16000 18337 16028
rect 18156 15960 18184 16000
rect 18325 15997 18337 16000
rect 18371 15997 18383 16031
rect 18325 15991 18383 15997
rect 14507 15932 14688 15960
rect 17788 15932 18184 15960
rect 14507 15929 14519 15932
rect 14461 15923 14519 15929
rect 5810 15852 5816 15904
rect 5868 15892 5874 15904
rect 6089 15895 6147 15901
rect 6089 15892 6101 15895
rect 5868 15864 6101 15892
rect 5868 15852 5874 15864
rect 6089 15861 6101 15864
rect 6135 15861 6147 15895
rect 11330 15892 11336 15904
rect 11291 15864 11336 15892
rect 6089 15855 6147 15861
rect 11330 15852 11336 15864
rect 11388 15852 11394 15904
rect 17678 15852 17684 15904
rect 17736 15892 17742 15904
rect 17788 15901 17816 15932
rect 17773 15895 17831 15901
rect 17773 15892 17785 15895
rect 17736 15864 17785 15892
rect 17736 15852 17742 15864
rect 17773 15861 17785 15864
rect 17819 15861 17831 15895
rect 17773 15855 17831 15861
rect 22373 15895 22431 15901
rect 22373 15861 22385 15895
rect 22419 15892 22431 15895
rect 22462 15892 22468 15904
rect 22419 15864 22468 15892
rect 22419 15861 22431 15864
rect 22373 15855 22431 15861
rect 22462 15852 22468 15864
rect 22520 15852 22526 15904
rect 22738 15892 22744 15904
rect 22699 15864 22744 15892
rect 22738 15852 22744 15864
rect 22796 15852 22802 15904
rect 1104 15802 28888 15824
rect 1104 15750 10982 15802
rect 11034 15750 11046 15802
rect 11098 15750 11110 15802
rect 11162 15750 11174 15802
rect 11226 15750 20982 15802
rect 21034 15750 21046 15802
rect 21098 15750 21110 15802
rect 21162 15750 21174 15802
rect 21226 15750 28888 15802
rect 1104 15728 28888 15750
rect 3418 15648 3424 15700
rect 3476 15688 3482 15700
rect 3513 15691 3571 15697
rect 3513 15688 3525 15691
rect 3476 15660 3525 15688
rect 3476 15648 3482 15660
rect 3513 15657 3525 15660
rect 3559 15688 3571 15691
rect 6638 15688 6644 15700
rect 3559 15660 6644 15688
rect 3559 15657 3571 15660
rect 3513 15651 3571 15657
rect 6638 15648 6644 15660
rect 6696 15648 6702 15700
rect 10042 15688 10048 15700
rect 10003 15660 10048 15688
rect 10042 15648 10048 15660
rect 10100 15648 10106 15700
rect 10413 15691 10471 15697
rect 10413 15657 10425 15691
rect 10459 15688 10471 15691
rect 10870 15688 10876 15700
rect 10459 15660 10876 15688
rect 10459 15657 10471 15660
rect 10413 15651 10471 15657
rect 10870 15648 10876 15660
rect 10928 15648 10934 15700
rect 12529 15691 12587 15697
rect 12529 15657 12541 15691
rect 12575 15688 12587 15691
rect 14185 15691 14243 15697
rect 12575 15660 13768 15688
rect 12575 15657 12587 15660
rect 12529 15651 12587 15657
rect 7006 15620 7012 15632
rect 6840 15592 7012 15620
rect 6840 15561 6868 15592
rect 7006 15580 7012 15592
rect 7064 15580 7070 15632
rect 8662 15620 8668 15632
rect 8623 15592 8668 15620
rect 8662 15580 8668 15592
rect 8720 15580 8726 15632
rect 13354 15620 13360 15632
rect 13280 15592 13360 15620
rect 6825 15555 6883 15561
rect 6825 15521 6837 15555
rect 6871 15521 6883 15555
rect 7282 15552 7288 15564
rect 7243 15524 7288 15552
rect 6825 15515 6883 15521
rect 7282 15512 7288 15524
rect 7340 15512 7346 15564
rect 9861 15555 9919 15561
rect 9861 15521 9873 15555
rect 9907 15552 9919 15555
rect 10318 15552 10324 15564
rect 9907 15524 10324 15552
rect 9907 15521 9919 15524
rect 9861 15515 9919 15521
rect 10318 15512 10324 15524
rect 10376 15512 10382 15564
rect 12342 15512 12348 15564
rect 12400 15552 12406 15564
rect 12894 15552 12900 15564
rect 12400 15524 12900 15552
rect 12400 15512 12406 15524
rect 12894 15512 12900 15524
rect 12952 15552 12958 15564
rect 13280 15561 13308 15592
rect 13354 15580 13360 15592
rect 13412 15580 13418 15632
rect 13740 15561 13768 15660
rect 14185 15657 14197 15691
rect 14231 15688 14243 15691
rect 15105 15691 15163 15697
rect 15105 15688 15117 15691
rect 14231 15660 15117 15688
rect 14231 15657 14243 15660
rect 14185 15651 14243 15657
rect 15105 15657 15117 15660
rect 15151 15688 15163 15691
rect 15838 15688 15844 15700
rect 15151 15660 15844 15688
rect 15151 15657 15163 15660
rect 15105 15651 15163 15657
rect 15838 15648 15844 15660
rect 15896 15648 15902 15700
rect 14642 15620 14648 15632
rect 14603 15592 14648 15620
rect 14642 15580 14648 15592
rect 14700 15580 14706 15632
rect 15470 15620 15476 15632
rect 15431 15592 15476 15620
rect 15470 15580 15476 15592
rect 15528 15580 15534 15632
rect 13173 15555 13231 15561
rect 13173 15552 13185 15555
rect 12952 15524 13185 15552
rect 12952 15512 12958 15524
rect 13173 15521 13185 15524
rect 13219 15521 13231 15555
rect 13173 15515 13231 15521
rect 13265 15555 13323 15561
rect 13265 15521 13277 15555
rect 13311 15521 13323 15555
rect 13633 15555 13691 15561
rect 13633 15552 13645 15555
rect 13265 15515 13323 15521
rect 13372 15524 13645 15552
rect 6638 15444 6644 15496
rect 6696 15484 6702 15496
rect 7009 15487 7067 15493
rect 7009 15484 7021 15487
rect 6696 15456 7021 15484
rect 6696 15444 6702 15456
rect 7009 15453 7021 15456
rect 7055 15453 7067 15487
rect 7009 15447 7067 15453
rect 13372 15416 13400 15524
rect 13633 15521 13645 15524
rect 13679 15521 13691 15555
rect 13633 15515 13691 15521
rect 13725 15555 13783 15561
rect 13725 15521 13737 15555
rect 13771 15552 13783 15555
rect 13814 15552 13820 15564
rect 13771 15524 13820 15552
rect 13771 15521 13783 15524
rect 13725 15515 13783 15521
rect 13814 15512 13820 15524
rect 13872 15512 13878 15564
rect 16206 15552 16212 15564
rect 16167 15524 16212 15552
rect 16206 15512 16212 15524
rect 16264 15512 16270 15564
rect 15746 15444 15752 15496
rect 15804 15484 15810 15496
rect 15933 15487 15991 15493
rect 15933 15484 15945 15487
rect 15804 15456 15945 15484
rect 15804 15444 15810 15456
rect 15933 15453 15945 15456
rect 15979 15484 15991 15487
rect 18046 15484 18052 15496
rect 15979 15456 18052 15484
rect 15979 15453 15991 15456
rect 15933 15447 15991 15453
rect 18046 15444 18052 15456
rect 18104 15444 18110 15496
rect 13004 15388 13400 15416
rect 13004 15360 13032 15388
rect 12897 15351 12955 15357
rect 12897 15317 12909 15351
rect 12943 15348 12955 15351
rect 12986 15348 12992 15360
rect 12943 15320 12992 15348
rect 12943 15317 12955 15320
rect 12897 15311 12955 15317
rect 12986 15308 12992 15320
rect 13044 15308 13050 15360
rect 17310 15348 17316 15360
rect 17271 15320 17316 15348
rect 17310 15308 17316 15320
rect 17368 15308 17374 15360
rect 1104 15258 28888 15280
rect 1104 15206 5982 15258
rect 6034 15206 6046 15258
rect 6098 15206 6110 15258
rect 6162 15206 6174 15258
rect 6226 15206 15982 15258
rect 16034 15206 16046 15258
rect 16098 15206 16110 15258
rect 16162 15206 16174 15258
rect 16226 15206 25982 15258
rect 26034 15206 26046 15258
rect 26098 15206 26110 15258
rect 26162 15206 26174 15258
rect 26226 15206 28888 15258
rect 1104 15184 28888 15206
rect 6638 15144 6644 15156
rect 6599 15116 6644 15144
rect 6638 15104 6644 15116
rect 6696 15104 6702 15156
rect 7101 15147 7159 15153
rect 7101 15113 7113 15147
rect 7147 15144 7159 15147
rect 7282 15144 7288 15156
rect 7147 15116 7288 15144
rect 7147 15113 7159 15116
rect 7101 15107 7159 15113
rect 7282 15104 7288 15116
rect 7340 15104 7346 15156
rect 7834 15144 7840 15156
rect 7795 15116 7840 15144
rect 7834 15104 7840 15116
rect 7892 15104 7898 15156
rect 10318 15144 10324 15156
rect 10279 15116 10324 15144
rect 10318 15104 10324 15116
rect 10376 15104 10382 15156
rect 12253 15147 12311 15153
rect 12253 15113 12265 15147
rect 12299 15144 12311 15147
rect 12342 15144 12348 15156
rect 12299 15116 12348 15144
rect 12299 15113 12311 15116
rect 12253 15107 12311 15113
rect 12342 15104 12348 15116
rect 12400 15104 12406 15156
rect 13354 15104 13360 15156
rect 13412 15144 13418 15156
rect 13541 15147 13599 15153
rect 13541 15144 13553 15147
rect 13412 15116 13553 15144
rect 13412 15104 13418 15116
rect 13541 15113 13553 15116
rect 13587 15113 13599 15147
rect 13541 15107 13599 15113
rect 13630 15104 13636 15156
rect 13688 15144 13694 15156
rect 13817 15147 13875 15153
rect 13817 15144 13829 15147
rect 13688 15116 13829 15144
rect 13688 15104 13694 15116
rect 13817 15113 13829 15116
rect 13863 15144 13875 15147
rect 13909 15147 13967 15153
rect 13909 15144 13921 15147
rect 13863 15116 13921 15144
rect 13863 15113 13875 15116
rect 13817 15107 13875 15113
rect 13909 15113 13921 15116
rect 13955 15113 13967 15147
rect 13909 15107 13967 15113
rect 16025 15147 16083 15153
rect 16025 15113 16037 15147
rect 16071 15144 16083 15147
rect 16298 15144 16304 15156
rect 16071 15116 16304 15144
rect 16071 15113 16083 15116
rect 16025 15107 16083 15113
rect 16298 15104 16304 15116
rect 16356 15104 16362 15156
rect 8205 15011 8263 15017
rect 8205 14977 8217 15011
rect 8251 15008 8263 15011
rect 8573 15011 8631 15017
rect 8573 15008 8585 15011
rect 8251 14980 8585 15008
rect 8251 14977 8263 14980
rect 8205 14971 8263 14977
rect 8573 14977 8585 14980
rect 8619 15008 8631 15011
rect 10336 15008 10364 15104
rect 14918 15036 14924 15088
rect 14976 15076 14982 15088
rect 15197 15079 15255 15085
rect 15197 15076 15209 15079
rect 14976 15048 15209 15076
rect 14976 15036 14982 15048
rect 15197 15045 15209 15048
rect 15243 15045 15255 15079
rect 15197 15039 15255 15045
rect 13262 15008 13268 15020
rect 8619 14980 10364 15008
rect 13223 14980 13268 15008
rect 8619 14977 8631 14980
rect 8573 14971 8631 14977
rect 13262 14968 13268 14980
rect 13320 15008 13326 15020
rect 16485 15011 16543 15017
rect 13320 14980 14504 15008
rect 13320 14968 13326 14980
rect 14476 14952 14504 14980
rect 16485 14977 16497 15011
rect 16531 15008 16543 15011
rect 16531 14980 16712 15008
rect 16531 14977 16543 14980
rect 16485 14971 16543 14977
rect 7834 14900 7840 14952
rect 7892 14940 7898 14952
rect 8297 14943 8355 14949
rect 8297 14940 8309 14943
rect 7892 14912 8309 14940
rect 7892 14900 7898 14912
rect 8297 14909 8309 14912
rect 8343 14909 8355 14943
rect 8297 14903 8355 14909
rect 9858 14900 9864 14952
rect 9916 14940 9922 14952
rect 10781 14943 10839 14949
rect 10781 14940 10793 14943
rect 9916 14912 10793 14940
rect 9916 14900 9922 14912
rect 10781 14909 10793 14912
rect 10827 14940 10839 14943
rect 11241 14943 11299 14949
rect 11241 14940 11253 14943
rect 10827 14912 11253 14940
rect 10827 14909 10839 14912
rect 10781 14903 10839 14909
rect 11241 14909 11253 14912
rect 11287 14909 11299 14943
rect 11241 14903 11299 14909
rect 11885 14943 11943 14949
rect 11885 14909 11897 14943
rect 11931 14940 11943 14943
rect 12618 14940 12624 14952
rect 11931 14912 12624 14940
rect 11931 14909 11943 14912
rect 11885 14903 11943 14909
rect 12618 14900 12624 14912
rect 12676 14940 12682 14952
rect 13817 14943 13875 14949
rect 12676 14912 13308 14940
rect 12676 14900 12682 14912
rect 13280 14884 13308 14912
rect 13817 14909 13829 14943
rect 13863 14940 13875 14943
rect 14277 14943 14335 14949
rect 14277 14940 14289 14943
rect 13863 14912 14289 14940
rect 13863 14909 13875 14912
rect 13817 14903 13875 14909
rect 14277 14909 14289 14912
rect 14323 14909 14335 14943
rect 14277 14903 14335 14909
rect 14369 14943 14427 14949
rect 14369 14909 14381 14943
rect 14415 14909 14427 14943
rect 14369 14903 14427 14909
rect 13262 14832 13268 14884
rect 13320 14832 13326 14884
rect 14384 14872 14412 14903
rect 14458 14900 14464 14952
rect 14516 14940 14522 14952
rect 14737 14943 14795 14949
rect 14737 14940 14749 14943
rect 14516 14912 14749 14940
rect 14516 14900 14522 14912
rect 14737 14909 14749 14912
rect 14783 14909 14795 14943
rect 14737 14903 14795 14909
rect 14829 14943 14887 14949
rect 14829 14909 14841 14943
rect 14875 14940 14887 14943
rect 15010 14940 15016 14952
rect 14875 14912 15016 14940
rect 14875 14909 14887 14912
rect 14829 14903 14887 14909
rect 15010 14900 15016 14912
rect 15068 14900 15074 14952
rect 16684 14949 16712 14980
rect 16577 14943 16635 14949
rect 16577 14909 16589 14943
rect 16623 14909 16635 14943
rect 16577 14903 16635 14909
rect 16669 14943 16727 14949
rect 16669 14909 16681 14943
rect 16715 14940 16727 14943
rect 17310 14940 17316 14952
rect 16715 14912 17316 14940
rect 16715 14909 16727 14912
rect 16669 14903 16727 14909
rect 14918 14872 14924 14884
rect 14384 14844 14924 14872
rect 14918 14832 14924 14844
rect 14976 14832 14982 14884
rect 7006 14764 7012 14816
rect 7064 14804 7070 14816
rect 7377 14807 7435 14813
rect 7377 14804 7389 14807
rect 7064 14776 7389 14804
rect 7064 14764 7070 14776
rect 7377 14773 7389 14776
rect 7423 14773 7435 14807
rect 7377 14767 7435 14773
rect 8570 14764 8576 14816
rect 8628 14804 8634 14816
rect 9677 14807 9735 14813
rect 9677 14804 9689 14807
rect 8628 14776 9689 14804
rect 8628 14764 8634 14776
rect 9677 14773 9689 14776
rect 9723 14773 9735 14807
rect 9677 14767 9735 14773
rect 10318 14764 10324 14816
rect 10376 14804 10382 14816
rect 10965 14807 11023 14813
rect 10965 14804 10977 14807
rect 10376 14776 10977 14804
rect 10376 14764 10382 14776
rect 10965 14773 10977 14776
rect 11011 14773 11023 14807
rect 10965 14767 11023 14773
rect 11422 14764 11428 14816
rect 11480 14804 11486 14816
rect 11882 14804 11888 14816
rect 11480 14776 11888 14804
rect 11480 14764 11486 14776
rect 11882 14764 11888 14776
rect 11940 14764 11946 14816
rect 16592 14804 16620 14903
rect 17310 14900 17316 14912
rect 17368 14900 17374 14952
rect 17126 14872 17132 14884
rect 17087 14844 17132 14872
rect 17126 14832 17132 14844
rect 17184 14832 17190 14884
rect 17405 14807 17463 14813
rect 17405 14804 17417 14807
rect 16592 14776 17417 14804
rect 17405 14773 17417 14776
rect 17451 14804 17463 14807
rect 17770 14804 17776 14816
rect 17451 14776 17776 14804
rect 17451 14773 17463 14776
rect 17405 14767 17463 14773
rect 17770 14764 17776 14776
rect 17828 14764 17834 14816
rect 1104 14714 28888 14736
rect 1104 14662 10982 14714
rect 11034 14662 11046 14714
rect 11098 14662 11110 14714
rect 11162 14662 11174 14714
rect 11226 14662 20982 14714
rect 21034 14662 21046 14714
rect 21098 14662 21110 14714
rect 21162 14662 21174 14714
rect 21226 14662 28888 14714
rect 1104 14640 28888 14662
rect 7469 14603 7527 14609
rect 7469 14569 7481 14603
rect 7515 14600 7527 14603
rect 8570 14600 8576 14612
rect 7515 14572 8576 14600
rect 7515 14569 7527 14572
rect 7469 14563 7527 14569
rect 8570 14560 8576 14572
rect 8628 14560 8634 14612
rect 9766 14560 9772 14612
rect 9824 14600 9830 14612
rect 10137 14603 10195 14609
rect 10137 14600 10149 14603
rect 9824 14572 10149 14600
rect 9824 14560 9830 14572
rect 10137 14569 10149 14572
rect 10183 14569 10195 14603
rect 10137 14563 10195 14569
rect 11149 14603 11207 14609
rect 11149 14569 11161 14603
rect 11195 14600 11207 14603
rect 11790 14600 11796 14612
rect 11195 14572 11796 14600
rect 11195 14569 11207 14572
rect 11149 14563 11207 14569
rect 11790 14560 11796 14572
rect 11848 14560 11854 14612
rect 14458 14600 14464 14612
rect 14419 14572 14464 14600
rect 14458 14560 14464 14572
rect 14516 14560 14522 14612
rect 7558 14532 7564 14544
rect 7519 14504 7564 14532
rect 7558 14492 7564 14504
rect 7616 14492 7622 14544
rect 11514 14492 11520 14544
rect 11572 14532 11578 14544
rect 12253 14535 12311 14541
rect 12253 14532 12265 14535
rect 11572 14504 12265 14532
rect 11572 14492 11578 14504
rect 12253 14501 12265 14504
rect 12299 14501 12311 14535
rect 13722 14532 13728 14544
rect 13683 14504 13728 14532
rect 12253 14495 12311 14501
rect 8205 14467 8263 14473
rect 8205 14433 8217 14467
rect 8251 14464 8263 14467
rect 8294 14464 8300 14476
rect 8251 14436 8300 14464
rect 8251 14433 8263 14436
rect 8205 14427 8263 14433
rect 8294 14424 8300 14436
rect 8352 14424 8358 14476
rect 8570 14464 8576 14476
rect 8531 14436 8576 14464
rect 8570 14424 8576 14436
rect 8628 14424 8634 14476
rect 9582 14424 9588 14476
rect 9640 14464 9646 14476
rect 9950 14464 9956 14476
rect 9640 14436 9956 14464
rect 9640 14424 9646 14436
rect 9950 14424 9956 14436
rect 10008 14424 10014 14476
rect 10226 14424 10232 14476
rect 10284 14464 10290 14476
rect 10686 14464 10692 14476
rect 10284 14436 10692 14464
rect 10284 14424 10290 14436
rect 10686 14424 10692 14436
rect 10744 14464 10750 14476
rect 10965 14467 11023 14473
rect 10965 14464 10977 14467
rect 10744 14436 10977 14464
rect 10744 14424 10750 14436
rect 10965 14433 10977 14436
rect 11011 14433 11023 14467
rect 10965 14427 11023 14433
rect 8110 14396 8116 14408
rect 8071 14368 8116 14396
rect 8110 14356 8116 14368
rect 8168 14356 8174 14408
rect 8478 14396 8484 14408
rect 8439 14368 8484 14396
rect 8478 14356 8484 14368
rect 8536 14356 8542 14408
rect 12268 14396 12296 14495
rect 13722 14492 13728 14504
rect 13780 14492 13786 14544
rect 13814 14492 13820 14544
rect 13872 14532 13878 14544
rect 14185 14535 14243 14541
rect 14185 14532 14197 14535
rect 13872 14504 14197 14532
rect 13872 14492 13878 14504
rect 14185 14501 14197 14504
rect 14231 14532 14243 14535
rect 15010 14532 15016 14544
rect 14231 14504 15016 14532
rect 14231 14501 14243 14504
rect 14185 14495 14243 14501
rect 15010 14492 15016 14504
rect 15068 14492 15074 14544
rect 16298 14492 16304 14544
rect 16356 14532 16362 14544
rect 16356 14504 17356 14532
rect 16356 14492 16362 14504
rect 12621 14467 12679 14473
rect 12621 14433 12633 14467
rect 12667 14433 12679 14467
rect 13078 14464 13084 14476
rect 13039 14436 13084 14464
rect 12621 14427 12679 14433
rect 12342 14396 12348 14408
rect 12255 14368 12348 14396
rect 12342 14356 12348 14368
rect 12400 14396 12406 14408
rect 12437 14399 12495 14405
rect 12437 14396 12449 14399
rect 12400 14368 12449 14396
rect 12400 14356 12406 14368
rect 12437 14365 12449 14368
rect 12483 14365 12495 14399
rect 12437 14359 12495 14365
rect 8754 14288 8760 14340
rect 8812 14328 8818 14340
rect 9490 14328 9496 14340
rect 8812 14300 9496 14328
rect 8812 14288 8818 14300
rect 9490 14288 9496 14300
rect 9548 14328 9554 14340
rect 11606 14328 11612 14340
rect 9548 14300 11612 14328
rect 9548 14288 9554 14300
rect 11606 14288 11612 14300
rect 11664 14288 11670 14340
rect 12636 14328 12664 14427
rect 13078 14424 13084 14436
rect 13136 14424 13142 14476
rect 13173 14467 13231 14473
rect 13173 14433 13185 14467
rect 13219 14464 13231 14467
rect 14642 14464 14648 14476
rect 13219 14436 14648 14464
rect 13219 14433 13231 14436
rect 13173 14427 13231 14433
rect 14642 14424 14648 14436
rect 14700 14424 14706 14476
rect 17126 14464 17132 14476
rect 17087 14436 17132 14464
rect 17126 14424 17132 14436
rect 17184 14424 17190 14476
rect 17328 14473 17356 14504
rect 20438 14492 20444 14544
rect 20496 14532 20502 14544
rect 20622 14532 20628 14544
rect 20496 14504 20628 14532
rect 20496 14492 20502 14504
rect 20622 14492 20628 14504
rect 20680 14492 20686 14544
rect 17313 14467 17371 14473
rect 17313 14433 17325 14467
rect 17359 14464 17371 14467
rect 17402 14464 17408 14476
rect 17359 14436 17408 14464
rect 17359 14433 17371 14436
rect 17313 14427 17371 14433
rect 17402 14424 17408 14436
rect 17460 14424 17466 14476
rect 17497 14467 17555 14473
rect 17497 14433 17509 14467
rect 17543 14464 17555 14467
rect 17586 14464 17592 14476
rect 17543 14436 17592 14464
rect 17543 14433 17555 14436
rect 17497 14427 17555 14433
rect 17586 14424 17592 14436
rect 17644 14424 17650 14476
rect 14918 14396 14924 14408
rect 14879 14368 14924 14396
rect 14918 14356 14924 14368
rect 14976 14356 14982 14408
rect 13630 14328 13636 14340
rect 12636 14300 13636 14328
rect 13630 14288 13636 14300
rect 13688 14288 13694 14340
rect 16945 14331 17003 14337
rect 16945 14297 16957 14331
rect 16991 14328 17003 14331
rect 17770 14328 17776 14340
rect 16991 14300 17776 14328
rect 16991 14297 17003 14300
rect 16945 14291 17003 14297
rect 17770 14288 17776 14300
rect 17828 14288 17834 14340
rect 9122 14260 9128 14272
rect 9083 14232 9128 14260
rect 9122 14220 9128 14232
rect 9180 14220 9186 14272
rect 15746 14220 15752 14272
rect 15804 14260 15810 14272
rect 15933 14263 15991 14269
rect 15933 14260 15945 14263
rect 15804 14232 15945 14260
rect 15804 14220 15810 14232
rect 15933 14229 15945 14232
rect 15979 14229 15991 14263
rect 15933 14223 15991 14229
rect 1104 14170 28888 14192
rect 1104 14118 5982 14170
rect 6034 14118 6046 14170
rect 6098 14118 6110 14170
rect 6162 14118 6174 14170
rect 6226 14118 15982 14170
rect 16034 14118 16046 14170
rect 16098 14118 16110 14170
rect 16162 14118 16174 14170
rect 16226 14118 25982 14170
rect 26034 14118 26046 14170
rect 26098 14118 26110 14170
rect 26162 14118 26174 14170
rect 26226 14118 28888 14170
rect 1104 14096 28888 14118
rect 7285 14059 7343 14065
rect 7285 14025 7297 14059
rect 7331 14056 7343 14059
rect 8478 14056 8484 14068
rect 7331 14028 8484 14056
rect 7331 14025 7343 14028
rect 7285 14019 7343 14025
rect 8478 14016 8484 14028
rect 8536 14016 8542 14068
rect 9950 14056 9956 14068
rect 9911 14028 9956 14056
rect 9950 14016 9956 14028
rect 10008 14016 10014 14068
rect 10686 14056 10692 14068
rect 10647 14028 10692 14056
rect 10686 14016 10692 14028
rect 10744 14056 10750 14068
rect 11333 14059 11391 14065
rect 11333 14056 11345 14059
rect 10744 14028 11345 14056
rect 10744 14016 10750 14028
rect 11333 14025 11345 14028
rect 11379 14025 11391 14059
rect 11333 14019 11391 14025
rect 12158 14016 12164 14068
rect 12216 14056 12222 14068
rect 12897 14059 12955 14065
rect 12897 14056 12909 14059
rect 12216 14028 12909 14056
rect 12216 14016 12222 14028
rect 12897 14025 12909 14028
rect 12943 14056 12955 14059
rect 13078 14056 13084 14068
rect 12943 14028 13084 14056
rect 12943 14025 12955 14028
rect 12897 14019 12955 14025
rect 13078 14016 13084 14028
rect 13136 14016 13142 14068
rect 13541 14059 13599 14065
rect 13541 14025 13553 14059
rect 13587 14056 13599 14059
rect 13630 14056 13636 14068
rect 13587 14028 13636 14056
rect 13587 14025 13599 14028
rect 13541 14019 13599 14025
rect 13630 14016 13636 14028
rect 13688 14016 13694 14068
rect 14274 14056 14280 14068
rect 14235 14028 14280 14056
rect 14274 14016 14280 14028
rect 14332 14016 14338 14068
rect 15378 14056 15384 14068
rect 15339 14028 15384 14056
rect 15378 14016 15384 14028
rect 15436 14016 15442 14068
rect 17126 14056 17132 14068
rect 17087 14028 17132 14056
rect 17126 14016 17132 14028
rect 17184 14016 17190 14068
rect 17402 14056 17408 14068
rect 17363 14028 17408 14056
rect 17402 14016 17408 14028
rect 17460 14016 17466 14068
rect 7653 13991 7711 13997
rect 7653 13957 7665 13991
rect 7699 13988 7711 13991
rect 8110 13988 8116 14000
rect 7699 13960 8116 13988
rect 7699 13957 7711 13960
rect 7653 13951 7711 13957
rect 8110 13948 8116 13960
rect 8168 13948 8174 14000
rect 8496 13988 8524 14016
rect 16761 13991 16819 13997
rect 8496 13960 9352 13988
rect 8294 13880 8300 13932
rect 8352 13920 8358 13932
rect 9324 13929 9352 13960
rect 16761 13957 16773 13991
rect 16807 13988 16819 13991
rect 17586 13988 17592 14000
rect 16807 13960 17592 13988
rect 16807 13957 16819 13960
rect 16761 13951 16819 13957
rect 17586 13948 17592 13960
rect 17644 13948 17650 14000
rect 9309 13923 9367 13929
rect 8352 13892 9076 13920
rect 8352 13880 8358 13892
rect 8386 13852 8392 13864
rect 8347 13824 8392 13852
rect 8386 13812 8392 13824
rect 8444 13812 8450 13864
rect 8754 13852 8760 13864
rect 8496 13824 8760 13852
rect 8297 13787 8355 13793
rect 8297 13753 8309 13787
rect 8343 13784 8355 13787
rect 8496 13784 8524 13824
rect 8754 13812 8760 13824
rect 8812 13852 8818 13864
rect 9048 13861 9076 13892
rect 9309 13889 9321 13923
rect 9355 13889 9367 13923
rect 9309 13883 9367 13889
rect 11885 13923 11943 13929
rect 11885 13889 11897 13923
rect 11931 13920 11943 13923
rect 15562 13920 15568 13932
rect 11931 13892 13952 13920
rect 15523 13892 15568 13920
rect 11931 13889 11943 13892
rect 11885 13883 11943 13889
rect 8849 13855 8907 13861
rect 8849 13852 8861 13855
rect 8812 13824 8861 13852
rect 8812 13812 8818 13824
rect 8849 13821 8861 13824
rect 8895 13821 8907 13855
rect 8849 13815 8907 13821
rect 9033 13855 9091 13861
rect 9033 13821 9045 13855
rect 9079 13821 9091 13855
rect 9033 13815 9091 13821
rect 9122 13812 9128 13864
rect 9180 13852 9186 13864
rect 9401 13855 9459 13861
rect 9401 13852 9413 13855
rect 9180 13824 9413 13852
rect 9180 13812 9186 13824
rect 9401 13821 9413 13824
rect 9447 13821 9459 13855
rect 9401 13815 9459 13821
rect 10505 13855 10563 13861
rect 10505 13821 10517 13855
rect 10551 13852 10563 13855
rect 12158 13852 12164 13864
rect 10551 13824 10916 13852
rect 12119 13824 12164 13852
rect 10551 13821 10563 13824
rect 10505 13815 10563 13821
rect 8343 13756 8524 13784
rect 8343 13753 8355 13756
rect 8297 13747 8355 13753
rect 8938 13744 8944 13796
rect 8996 13784 9002 13796
rect 9214 13784 9220 13796
rect 8996 13756 9220 13784
rect 8996 13744 9002 13756
rect 9214 13744 9220 13756
rect 9272 13744 9278 13796
rect 9416 13784 9444 13815
rect 10042 13784 10048 13796
rect 9416 13756 10048 13784
rect 10042 13744 10048 13756
rect 10100 13744 10106 13796
rect 10888 13728 10916 13824
rect 12158 13812 12164 13824
rect 12216 13812 12222 13864
rect 12802 13852 12808 13864
rect 12763 13824 12808 13852
rect 12802 13812 12808 13824
rect 12860 13812 12866 13864
rect 13924 13861 13952 13892
rect 15562 13880 15568 13892
rect 15620 13880 15626 13932
rect 26053 13923 26111 13929
rect 26053 13889 26065 13923
rect 26099 13920 26111 13923
rect 27614 13920 27620 13932
rect 26099 13892 26464 13920
rect 27575 13892 27620 13920
rect 26099 13889 26111 13892
rect 26053 13883 26111 13889
rect 13909 13855 13967 13861
rect 13909 13821 13921 13855
rect 13955 13852 13967 13855
rect 14642 13852 14648 13864
rect 13955 13824 14648 13852
rect 13955 13821 13967 13824
rect 13909 13815 13967 13821
rect 14642 13812 14648 13824
rect 14700 13812 14706 13864
rect 15378 13812 15384 13864
rect 15436 13852 15442 13864
rect 26436 13861 26464 13892
rect 27614 13880 27620 13892
rect 27672 13880 27678 13932
rect 15657 13855 15715 13861
rect 15657 13852 15669 13855
rect 15436 13824 15669 13852
rect 15436 13812 15442 13824
rect 15657 13821 15669 13824
rect 15703 13821 15715 13855
rect 15657 13815 15715 13821
rect 26145 13855 26203 13861
rect 26145 13821 26157 13855
rect 26191 13821 26203 13855
rect 26145 13815 26203 13821
rect 26421 13855 26479 13861
rect 26421 13821 26433 13855
rect 26467 13852 26479 13855
rect 26510 13852 26516 13864
rect 26467 13824 26516 13852
rect 26467 13821 26479 13824
rect 26421 13815 26479 13821
rect 26160 13784 26188 13815
rect 26510 13812 26516 13824
rect 26568 13812 26574 13864
rect 26234 13784 26240 13796
rect 26160 13756 26240 13784
rect 26234 13744 26240 13756
rect 26292 13744 26298 13796
rect 10870 13676 10876 13728
rect 10928 13716 10934 13728
rect 10965 13719 11023 13725
rect 10965 13716 10977 13719
rect 10928 13688 10977 13716
rect 10928 13676 10934 13688
rect 10965 13685 10977 13688
rect 11011 13685 11023 13719
rect 10965 13679 11023 13685
rect 1104 13626 28888 13648
rect 1104 13574 10982 13626
rect 11034 13574 11046 13626
rect 11098 13574 11110 13626
rect 11162 13574 11174 13626
rect 11226 13574 20982 13626
rect 21034 13574 21046 13626
rect 21098 13574 21110 13626
rect 21162 13574 21174 13626
rect 21226 13574 28888 13626
rect 1104 13552 28888 13574
rect 7837 13515 7895 13521
rect 7837 13481 7849 13515
rect 7883 13512 7895 13515
rect 8294 13512 8300 13524
rect 7883 13484 8300 13512
rect 7883 13481 7895 13484
rect 7837 13475 7895 13481
rect 8294 13472 8300 13484
rect 8352 13512 8358 13524
rect 8757 13515 8815 13521
rect 8757 13512 8769 13515
rect 8352 13484 8769 13512
rect 8352 13472 8358 13484
rect 8757 13481 8769 13484
rect 8803 13481 8815 13515
rect 8757 13475 8815 13481
rect 12802 13472 12808 13524
rect 12860 13512 12866 13524
rect 12989 13515 13047 13521
rect 12989 13512 13001 13515
rect 12860 13484 13001 13512
rect 12860 13472 12866 13484
rect 12989 13481 13001 13484
rect 13035 13481 13047 13515
rect 22554 13512 22560 13524
rect 22515 13484 22560 13512
rect 12989 13475 13047 13481
rect 22554 13472 22560 13484
rect 22612 13472 22618 13524
rect 26234 13512 26240 13524
rect 26195 13484 26240 13512
rect 26234 13472 26240 13484
rect 26292 13472 26298 13524
rect 8478 13444 8484 13456
rect 8439 13416 8484 13444
rect 8478 13404 8484 13416
rect 8536 13404 8542 13456
rect 7374 13336 7380 13388
rect 7432 13376 7438 13388
rect 7469 13379 7527 13385
rect 7469 13376 7481 13379
rect 7432 13348 7481 13376
rect 7432 13336 7438 13348
rect 7469 13345 7481 13348
rect 7515 13345 7527 13379
rect 10686 13376 10692 13388
rect 10647 13348 10692 13376
rect 7469 13339 7527 13345
rect 10686 13336 10692 13348
rect 10744 13336 10750 13388
rect 12250 13376 12256 13388
rect 12211 13348 12256 13376
rect 12250 13336 12256 13348
rect 12308 13376 12314 13388
rect 13538 13376 13544 13388
rect 12308 13348 13544 13376
rect 12308 13336 12314 13348
rect 13538 13336 13544 13348
rect 13596 13336 13602 13388
rect 20530 13336 20536 13388
rect 20588 13376 20594 13388
rect 21177 13379 21235 13385
rect 21177 13376 21189 13379
rect 20588 13348 21189 13376
rect 20588 13336 20594 13348
rect 21177 13345 21189 13348
rect 21223 13376 21235 13379
rect 21542 13376 21548 13388
rect 21223 13348 21548 13376
rect 21223 13345 21235 13348
rect 21177 13339 21235 13345
rect 21542 13336 21548 13348
rect 21600 13336 21606 13388
rect 12161 13311 12219 13317
rect 12161 13277 12173 13311
rect 12207 13308 12219 13311
rect 12342 13308 12348 13320
rect 12207 13280 12348 13308
rect 12207 13277 12219 13280
rect 12161 13271 12219 13277
rect 12342 13268 12348 13280
rect 12400 13308 12406 13320
rect 13906 13308 13912 13320
rect 12400 13280 13912 13308
rect 12400 13268 12406 13280
rect 13906 13268 13912 13280
rect 13964 13268 13970 13320
rect 21450 13308 21456 13320
rect 21411 13280 21456 13308
rect 21450 13268 21456 13280
rect 21508 13268 21514 13320
rect 10778 13200 10784 13252
rect 10836 13240 10842 13252
rect 13725 13243 13783 13249
rect 13725 13240 13737 13243
rect 10836 13212 13737 13240
rect 10836 13200 10842 13212
rect 13725 13209 13737 13212
rect 13771 13209 13783 13243
rect 13725 13203 13783 13209
rect 7006 13132 7012 13184
rect 7064 13172 7070 13184
rect 7285 13175 7343 13181
rect 7285 13172 7297 13175
rect 7064 13144 7297 13172
rect 7064 13132 7070 13144
rect 7285 13141 7297 13144
rect 7331 13141 7343 13175
rect 11054 13172 11060 13184
rect 11015 13144 11060 13172
rect 7285 13135 7343 13141
rect 11054 13132 11060 13144
rect 11112 13132 11118 13184
rect 12342 13132 12348 13184
rect 12400 13172 12406 13184
rect 12437 13175 12495 13181
rect 12437 13172 12449 13175
rect 12400 13144 12449 13172
rect 12400 13132 12406 13144
rect 12437 13141 12449 13144
rect 12483 13141 12495 13175
rect 12437 13135 12495 13141
rect 25038 13132 25044 13184
rect 25096 13172 25102 13184
rect 26510 13172 26516 13184
rect 25096 13144 26516 13172
rect 25096 13132 25102 13144
rect 26510 13132 26516 13144
rect 26568 13132 26574 13184
rect 1104 13082 28888 13104
rect 1104 13030 5982 13082
rect 6034 13030 6046 13082
rect 6098 13030 6110 13082
rect 6162 13030 6174 13082
rect 6226 13030 15982 13082
rect 16034 13030 16046 13082
rect 16098 13030 16110 13082
rect 16162 13030 16174 13082
rect 16226 13030 25982 13082
rect 26034 13030 26046 13082
rect 26098 13030 26110 13082
rect 26162 13030 26174 13082
rect 26226 13030 28888 13082
rect 1104 13008 28888 13030
rect 7374 12968 7380 12980
rect 7335 12940 7380 12968
rect 7374 12928 7380 12940
rect 7432 12928 7438 12980
rect 10042 12968 10048 12980
rect 10003 12940 10048 12968
rect 10042 12928 10048 12940
rect 10100 12928 10106 12980
rect 10686 12968 10692 12980
rect 10647 12940 10692 12968
rect 10686 12928 10692 12940
rect 10744 12968 10750 12980
rect 12161 12971 12219 12977
rect 12161 12968 12173 12971
rect 10744 12940 12173 12968
rect 10744 12928 10750 12940
rect 12161 12937 12173 12940
rect 12207 12968 12219 12971
rect 12250 12968 12256 12980
rect 12207 12940 12256 12968
rect 12207 12937 12219 12940
rect 12161 12931 12219 12937
rect 12250 12928 12256 12940
rect 12308 12928 12314 12980
rect 13906 12968 13912 12980
rect 13867 12940 13912 12968
rect 13906 12928 13912 12940
rect 13964 12928 13970 12980
rect 21269 12971 21327 12977
rect 21269 12937 21281 12971
rect 21315 12968 21327 12971
rect 21450 12968 21456 12980
rect 21315 12940 21456 12968
rect 21315 12937 21327 12940
rect 21269 12931 21327 12937
rect 21450 12928 21456 12940
rect 21508 12928 21514 12980
rect 21634 12968 21640 12980
rect 21595 12940 21640 12968
rect 21634 12928 21640 12940
rect 21692 12928 21698 12980
rect 13538 12900 13544 12912
rect 13499 12872 13544 12900
rect 13538 12860 13544 12872
rect 13596 12860 13602 12912
rect 8573 12835 8631 12841
rect 8573 12801 8585 12835
rect 8619 12832 8631 12835
rect 8938 12832 8944 12844
rect 8619 12804 8944 12832
rect 8619 12801 8631 12804
rect 8573 12795 8631 12801
rect 8938 12792 8944 12804
rect 8996 12792 9002 12844
rect 8662 12764 8668 12776
rect 8623 12736 8668 12764
rect 8662 12724 8668 12736
rect 8720 12724 8726 12776
rect 11054 12724 11060 12776
rect 11112 12764 11118 12776
rect 11149 12767 11207 12773
rect 11149 12764 11161 12767
rect 11112 12736 11161 12764
rect 11112 12724 11118 12736
rect 11149 12733 11161 12736
rect 11195 12764 11207 12767
rect 11609 12767 11667 12773
rect 11609 12764 11621 12767
rect 11195 12736 11621 12764
rect 11195 12733 11207 12736
rect 11149 12727 11207 12733
rect 11609 12733 11621 12736
rect 11655 12733 11667 12767
rect 11609 12727 11667 12733
rect 12437 12767 12495 12773
rect 12437 12733 12449 12767
rect 12483 12764 12495 12767
rect 12897 12767 12955 12773
rect 12897 12764 12909 12767
rect 12483 12736 12909 12764
rect 12483 12733 12495 12736
rect 12437 12727 12495 12733
rect 12897 12733 12909 12736
rect 12943 12733 12955 12767
rect 12897 12727 12955 12733
rect 11330 12628 11336 12640
rect 11243 12600 11336 12628
rect 11330 12588 11336 12600
rect 11388 12628 11394 12640
rect 12452 12628 12480 12727
rect 21266 12724 21272 12776
rect 21324 12764 21330 12776
rect 21726 12764 21732 12776
rect 21324 12736 21732 12764
rect 21324 12724 21330 12736
rect 21726 12724 21732 12736
rect 21784 12724 21790 12776
rect 12618 12628 12624 12640
rect 11388 12600 12480 12628
rect 12579 12600 12624 12628
rect 11388 12588 11394 12600
rect 12618 12588 12624 12600
rect 12676 12588 12682 12640
rect 1104 12538 28888 12560
rect 1104 12486 10982 12538
rect 11034 12486 11046 12538
rect 11098 12486 11110 12538
rect 11162 12486 11174 12538
rect 11226 12486 20982 12538
rect 21034 12486 21046 12538
rect 21098 12486 21110 12538
rect 21162 12486 21174 12538
rect 21226 12486 28888 12538
rect 1104 12464 28888 12486
rect 12529 12427 12587 12433
rect 12529 12393 12541 12427
rect 12575 12424 12587 12427
rect 12618 12424 12624 12436
rect 12575 12396 12624 12424
rect 12575 12393 12587 12396
rect 12529 12387 12587 12393
rect 12618 12384 12624 12396
rect 12676 12424 12682 12436
rect 12805 12427 12863 12433
rect 12805 12424 12817 12427
rect 12676 12396 12817 12424
rect 12676 12384 12682 12396
rect 12805 12393 12817 12396
rect 12851 12424 12863 12427
rect 12851 12396 13768 12424
rect 12851 12393 12863 12396
rect 12805 12387 12863 12393
rect 12342 12356 12348 12368
rect 11624 12328 12348 12356
rect 9769 12291 9827 12297
rect 9769 12257 9781 12291
rect 9815 12288 9827 12291
rect 9858 12288 9864 12300
rect 9815 12260 9864 12288
rect 9815 12257 9827 12260
rect 9769 12251 9827 12257
rect 9858 12248 9864 12260
rect 9916 12248 9922 12300
rect 11624 12297 11652 12328
rect 12342 12316 12348 12328
rect 12400 12316 12406 12368
rect 12986 12316 12992 12368
rect 13044 12356 13050 12368
rect 13044 12328 13676 12356
rect 13044 12316 13050 12328
rect 11609 12291 11667 12297
rect 11609 12257 11621 12291
rect 11655 12257 11667 12291
rect 11609 12251 11667 12257
rect 11698 12248 11704 12300
rect 11756 12288 11762 12300
rect 11793 12291 11851 12297
rect 11793 12288 11805 12291
rect 11756 12260 11805 12288
rect 11756 12248 11762 12260
rect 11793 12257 11805 12260
rect 11839 12257 11851 12291
rect 11974 12288 11980 12300
rect 11935 12260 11980 12288
rect 11793 12251 11851 12257
rect 10318 12180 10324 12232
rect 10376 12220 10382 12232
rect 10594 12220 10600 12232
rect 10376 12192 10600 12220
rect 10376 12180 10382 12192
rect 10594 12180 10600 12192
rect 10652 12180 10658 12232
rect 11808 12220 11836 12251
rect 11974 12248 11980 12260
rect 12032 12248 12038 12300
rect 13173 12291 13231 12297
rect 13173 12257 13185 12291
rect 13219 12257 13231 12291
rect 13173 12251 13231 12257
rect 12526 12220 12532 12232
rect 11808 12192 12532 12220
rect 12526 12180 12532 12192
rect 12584 12220 12590 12232
rect 13188 12220 13216 12251
rect 13262 12248 13268 12300
rect 13320 12288 13326 12300
rect 13648 12297 13676 12328
rect 13740 12297 13768 12396
rect 13633 12291 13691 12297
rect 13320 12260 13365 12288
rect 13320 12248 13326 12260
rect 13633 12257 13645 12291
rect 13679 12257 13691 12291
rect 13633 12251 13691 12257
rect 13725 12291 13783 12297
rect 13725 12257 13737 12291
rect 13771 12257 13783 12291
rect 13725 12251 13783 12257
rect 16209 12291 16267 12297
rect 16209 12257 16221 12291
rect 16255 12288 16267 12291
rect 16942 12288 16948 12300
rect 16255 12260 16948 12288
rect 16255 12257 16267 12260
rect 16209 12251 16267 12257
rect 16942 12248 16948 12260
rect 17000 12248 17006 12300
rect 12584 12192 13216 12220
rect 12584 12180 12590 12192
rect 11422 12152 11428 12164
rect 11383 12124 11428 12152
rect 11422 12112 11428 12124
rect 11480 12112 11486 12164
rect 15286 12112 15292 12164
rect 15344 12152 15350 12164
rect 15746 12152 15752 12164
rect 15344 12124 15752 12152
rect 15344 12112 15350 12124
rect 15746 12112 15752 12124
rect 15804 12152 15810 12164
rect 16025 12155 16083 12161
rect 16025 12152 16037 12155
rect 15804 12124 16037 12152
rect 15804 12112 15810 12124
rect 16025 12121 16037 12124
rect 16071 12121 16083 12155
rect 16025 12115 16083 12121
rect 7926 12044 7932 12096
rect 7984 12084 7990 12096
rect 8662 12084 8668 12096
rect 7984 12056 8668 12084
rect 7984 12044 7990 12056
rect 8662 12044 8668 12056
rect 8720 12044 8726 12096
rect 9950 12084 9956 12096
rect 9911 12056 9956 12084
rect 9950 12044 9956 12056
rect 10008 12044 10014 12096
rect 10410 12084 10416 12096
rect 10371 12056 10416 12084
rect 10410 12044 10416 12056
rect 10468 12044 10474 12096
rect 14182 12084 14188 12096
rect 14143 12056 14188 12084
rect 14182 12044 14188 12056
rect 14240 12044 14246 12096
rect 15562 12084 15568 12096
rect 15523 12056 15568 12084
rect 15562 12044 15568 12056
rect 15620 12044 15626 12096
rect 15838 12084 15844 12096
rect 15799 12056 15844 12084
rect 15838 12044 15844 12056
rect 15896 12044 15902 12096
rect 1104 11994 28888 12016
rect 1104 11942 5982 11994
rect 6034 11942 6046 11994
rect 6098 11942 6110 11994
rect 6162 11942 6174 11994
rect 6226 11942 15982 11994
rect 16034 11942 16046 11994
rect 16098 11942 16110 11994
rect 16162 11942 16174 11994
rect 16226 11942 25982 11994
rect 26034 11942 26046 11994
rect 26098 11942 26110 11994
rect 26162 11942 26174 11994
rect 26226 11942 28888 11994
rect 1104 11920 28888 11942
rect 8938 11840 8944 11892
rect 8996 11880 9002 11892
rect 9125 11883 9183 11889
rect 9125 11880 9137 11883
rect 8996 11852 9137 11880
rect 8996 11840 9002 11852
rect 9125 11849 9137 11852
rect 9171 11849 9183 11883
rect 9490 11880 9496 11892
rect 9451 11852 9496 11880
rect 9125 11843 9183 11849
rect 9140 11676 9168 11843
rect 9490 11840 9496 11852
rect 9548 11840 9554 11892
rect 9858 11880 9864 11892
rect 9819 11852 9864 11880
rect 9858 11840 9864 11852
rect 9916 11840 9922 11892
rect 11701 11883 11759 11889
rect 11701 11849 11713 11883
rect 11747 11880 11759 11883
rect 11974 11880 11980 11892
rect 11747 11852 11980 11880
rect 11747 11849 11759 11852
rect 11701 11843 11759 11849
rect 11974 11840 11980 11852
rect 12032 11840 12038 11892
rect 12986 11840 12992 11892
rect 13044 11880 13050 11892
rect 14093 11883 14151 11889
rect 14093 11880 14105 11883
rect 13044 11852 14105 11880
rect 13044 11840 13050 11852
rect 14093 11849 14105 11852
rect 14139 11849 14151 11883
rect 14918 11880 14924 11892
rect 14879 11852 14924 11880
rect 14093 11843 14151 11849
rect 14918 11840 14924 11852
rect 14976 11840 14982 11892
rect 15378 11880 15384 11892
rect 15339 11852 15384 11880
rect 15378 11840 15384 11852
rect 15436 11840 15442 11892
rect 16942 11880 16948 11892
rect 16903 11852 16948 11880
rect 16942 11840 16948 11852
rect 17000 11840 17006 11892
rect 9508 11812 9536 11840
rect 10137 11815 10195 11821
rect 10137 11812 10149 11815
rect 9508 11784 10149 11812
rect 10137 11781 10149 11784
rect 10183 11812 10195 11815
rect 10183 11784 11192 11812
rect 10183 11781 10195 11784
rect 10137 11775 10195 11781
rect 9309 11679 9367 11685
rect 9309 11676 9321 11679
rect 9140 11648 9321 11676
rect 9309 11645 9321 11648
rect 9355 11645 9367 11679
rect 9309 11639 9367 11645
rect 10410 11636 10416 11688
rect 10468 11676 10474 11688
rect 10781 11679 10839 11685
rect 10781 11676 10793 11679
rect 10468 11648 10793 11676
rect 10468 11636 10474 11648
rect 10781 11645 10793 11648
rect 10827 11645 10839 11679
rect 10781 11639 10839 11645
rect 10318 11608 10324 11620
rect 10279 11580 10324 11608
rect 10318 11568 10324 11580
rect 10376 11568 10382 11620
rect 10796 11608 10824 11639
rect 10870 11636 10876 11688
rect 10928 11676 10934 11688
rect 11164 11685 11192 11784
rect 12526 11772 12532 11824
rect 12584 11812 12590 11824
rect 14461 11815 14519 11821
rect 14461 11812 14473 11815
rect 12584 11784 14473 11812
rect 12584 11772 12590 11784
rect 14461 11781 14473 11784
rect 14507 11781 14519 11815
rect 14936 11812 14964 11840
rect 15746 11812 15752 11824
rect 14936 11784 15752 11812
rect 14461 11775 14519 11781
rect 15746 11772 15752 11784
rect 15804 11812 15810 11824
rect 15804 11784 16068 11812
rect 15804 11772 15810 11784
rect 12158 11744 12164 11756
rect 12119 11716 12164 11744
rect 12158 11704 12164 11716
rect 12216 11744 12222 11756
rect 15562 11744 15568 11756
rect 12216 11716 12848 11744
rect 15523 11716 15568 11744
rect 12216 11704 12222 11716
rect 10965 11679 11023 11685
rect 10965 11676 10977 11679
rect 10928 11648 10977 11676
rect 10928 11636 10934 11648
rect 10965 11645 10977 11648
rect 11011 11645 11023 11679
rect 10965 11639 11023 11645
rect 11149 11679 11207 11685
rect 11149 11645 11161 11679
rect 11195 11645 11207 11679
rect 11149 11639 11207 11645
rect 12434 11636 12440 11688
rect 12492 11676 12498 11688
rect 12618 11676 12624 11688
rect 12492 11648 12537 11676
rect 12579 11648 12624 11676
rect 12492 11636 12498 11648
rect 12618 11636 12624 11648
rect 12676 11636 12682 11688
rect 12820 11676 12848 11716
rect 15562 11704 15568 11716
rect 15620 11704 15626 11756
rect 16040 11753 16068 11784
rect 16025 11747 16083 11753
rect 16025 11713 16037 11747
rect 16071 11713 16083 11747
rect 16025 11707 16083 11713
rect 13081 11679 13139 11685
rect 13081 11676 13093 11679
rect 12820 11648 13093 11676
rect 13081 11645 13093 11648
rect 13127 11645 13139 11679
rect 13081 11639 13139 11645
rect 13173 11679 13231 11685
rect 13173 11645 13185 11679
rect 13219 11645 13231 11679
rect 13173 11639 13231 11645
rect 15749 11679 15807 11685
rect 15749 11645 15761 11679
rect 15795 11676 15807 11679
rect 15930 11676 15936 11688
rect 15795 11648 15936 11676
rect 15795 11645 15807 11648
rect 15749 11639 15807 11645
rect 11330 11608 11336 11620
rect 10796 11580 11336 11608
rect 11330 11568 11336 11580
rect 11388 11568 11394 11620
rect 12636 11608 12664 11636
rect 13188 11608 13216 11639
rect 15930 11636 15936 11648
rect 15988 11636 15994 11688
rect 16117 11679 16175 11685
rect 16117 11645 16129 11679
rect 16163 11645 16175 11679
rect 16117 11639 16175 11645
rect 13722 11608 13728 11620
rect 12636 11580 13216 11608
rect 13683 11580 13728 11608
rect 13722 11568 13728 11580
rect 13780 11568 13786 11620
rect 15654 11568 15660 11620
rect 15712 11608 15718 11620
rect 16132 11608 16160 11639
rect 16577 11611 16635 11617
rect 16577 11608 16589 11611
rect 15712 11580 16589 11608
rect 15712 11568 15718 11580
rect 16577 11577 16589 11580
rect 16623 11577 16635 11611
rect 16577 11571 16635 11577
rect 1104 11450 28888 11472
rect 1104 11398 10982 11450
rect 11034 11398 11046 11450
rect 11098 11398 11110 11450
rect 11162 11398 11174 11450
rect 11226 11398 20982 11450
rect 21034 11398 21046 11450
rect 21098 11398 21110 11450
rect 21162 11398 21174 11450
rect 21226 11398 28888 11450
rect 1104 11376 28888 11398
rect 10413 11339 10471 11345
rect 10413 11305 10425 11339
rect 10459 11336 10471 11339
rect 10870 11336 10876 11348
rect 10459 11308 10876 11336
rect 10459 11305 10471 11308
rect 10413 11299 10471 11305
rect 10870 11296 10876 11308
rect 10928 11336 10934 11348
rect 11609 11339 11667 11345
rect 11609 11336 11621 11339
rect 10928 11308 11621 11336
rect 10928 11296 10934 11308
rect 11609 11305 11621 11308
rect 11655 11336 11667 11339
rect 11698 11336 11704 11348
rect 11655 11308 11704 11336
rect 11655 11305 11667 11308
rect 11609 11299 11667 11305
rect 11698 11296 11704 11308
rect 11756 11296 11762 11348
rect 12069 11339 12127 11345
rect 12069 11305 12081 11339
rect 12115 11336 12127 11339
rect 12342 11336 12348 11348
rect 12115 11308 12348 11336
rect 12115 11305 12127 11308
rect 12069 11299 12127 11305
rect 12342 11296 12348 11308
rect 12400 11296 12406 11348
rect 12434 11296 12440 11348
rect 12492 11336 12498 11348
rect 12492 11308 12537 11336
rect 12492 11296 12498 11308
rect 12618 11296 12624 11348
rect 12676 11336 12682 11348
rect 12805 11339 12863 11345
rect 12805 11336 12817 11339
rect 12676 11308 12817 11336
rect 12676 11296 12682 11308
rect 12805 11305 12817 11308
rect 12851 11336 12863 11339
rect 12851 11308 13216 11336
rect 12851 11305 12863 11308
rect 12805 11299 12863 11305
rect 10778 11228 10784 11280
rect 10836 11268 10842 11280
rect 11330 11268 11336 11280
rect 10836 11240 10916 11268
rect 11291 11240 11336 11268
rect 10836 11228 10842 11240
rect 7006 11160 7012 11212
rect 7064 11200 7070 11212
rect 7834 11200 7840 11212
rect 7064 11172 7840 11200
rect 7064 11160 7070 11172
rect 7834 11160 7840 11172
rect 7892 11200 7898 11212
rect 10888 11209 10916 11240
rect 11330 11228 11336 11240
rect 11388 11228 11394 11280
rect 13188 11268 13216 11308
rect 13262 11296 13268 11348
rect 13320 11336 13326 11348
rect 14645 11339 14703 11345
rect 14645 11336 14657 11339
rect 13320 11308 14657 11336
rect 13320 11296 13326 11308
rect 14645 11305 14657 11308
rect 14691 11305 14703 11339
rect 14645 11299 14703 11305
rect 15930 11296 15936 11348
rect 15988 11336 15994 11348
rect 16669 11339 16727 11345
rect 16669 11336 16681 11339
rect 15988 11308 16681 11336
rect 15988 11296 15994 11308
rect 16669 11305 16681 11308
rect 16715 11305 16727 11339
rect 16669 11299 16727 11305
rect 16942 11296 16948 11348
rect 17000 11336 17006 11348
rect 17773 11339 17831 11345
rect 17773 11336 17785 11339
rect 17000 11308 17785 11336
rect 17000 11296 17006 11308
rect 17773 11305 17785 11308
rect 17819 11336 17831 11339
rect 18046 11336 18052 11348
rect 17819 11308 18052 11336
rect 17819 11305 17831 11308
rect 17773 11299 17831 11305
rect 18046 11296 18052 11308
rect 18104 11296 18110 11348
rect 13354 11268 13360 11280
rect 13188 11240 13360 11268
rect 13188 11209 13216 11240
rect 13354 11228 13360 11240
rect 13412 11268 13418 11280
rect 13412 11240 13768 11268
rect 13412 11228 13418 11240
rect 8021 11203 8079 11209
rect 8021 11200 8033 11203
rect 7892 11172 8033 11200
rect 7892 11160 7898 11172
rect 8021 11169 8033 11172
rect 8067 11169 8079 11203
rect 8021 11163 8079 11169
rect 10873 11203 10931 11209
rect 10873 11169 10885 11203
rect 10919 11169 10931 11203
rect 10873 11163 10931 11169
rect 13173 11203 13231 11209
rect 13173 11169 13185 11203
rect 13219 11169 13231 11203
rect 13630 11200 13636 11212
rect 13591 11172 13636 11200
rect 13173 11163 13231 11169
rect 13630 11160 13636 11172
rect 13688 11160 13694 11212
rect 13740 11209 13768 11240
rect 13725 11203 13783 11209
rect 13725 11169 13737 11203
rect 13771 11169 13783 11203
rect 15565 11203 15623 11209
rect 15565 11200 15577 11203
rect 13725 11163 13783 11169
rect 14292 11172 15577 11200
rect 10781 11135 10839 11141
rect 10781 11101 10793 11135
rect 10827 11132 10839 11135
rect 11514 11132 11520 11144
rect 10827 11104 11520 11132
rect 10827 11101 10839 11104
rect 10781 11095 10839 11101
rect 11514 11092 11520 11104
rect 11572 11092 11578 11144
rect 12802 11092 12808 11144
rect 12860 11132 12866 11144
rect 14292 11141 14320 11172
rect 15565 11169 15577 11172
rect 15611 11200 15623 11203
rect 15654 11200 15660 11212
rect 15611 11172 15660 11200
rect 15611 11169 15623 11172
rect 15565 11163 15623 11169
rect 15654 11160 15660 11172
rect 15712 11160 15718 11212
rect 17954 11200 17960 11212
rect 17915 11172 17960 11200
rect 17954 11160 17960 11172
rect 18012 11160 18018 11212
rect 12989 11135 13047 11141
rect 12989 11132 13001 11135
rect 12860 11104 13001 11132
rect 12860 11092 12866 11104
rect 12989 11101 13001 11104
rect 13035 11101 13047 11135
rect 12989 11095 13047 11101
rect 14277 11135 14335 11141
rect 14277 11101 14289 11135
rect 14323 11101 14335 11135
rect 15286 11132 15292 11144
rect 15247 11104 15292 11132
rect 14277 11095 14335 11101
rect 15286 11092 15292 11104
rect 15344 11092 15350 11144
rect 7837 11067 7895 11073
rect 7837 11033 7849 11067
rect 7883 11064 7895 11067
rect 7926 11064 7932 11076
rect 7883 11036 7932 11064
rect 7883 11033 7895 11036
rect 7837 11027 7895 11033
rect 7926 11024 7932 11036
rect 7984 11024 7990 11076
rect 1104 10906 28888 10928
rect 1104 10854 5982 10906
rect 6034 10854 6046 10906
rect 6098 10854 6110 10906
rect 6162 10854 6174 10906
rect 6226 10854 15982 10906
rect 16034 10854 16046 10906
rect 16098 10854 16110 10906
rect 16162 10854 16174 10906
rect 16226 10854 25982 10906
rect 26034 10854 26046 10906
rect 26098 10854 26110 10906
rect 26162 10854 26174 10906
rect 26226 10854 28888 10906
rect 1104 10832 28888 10854
rect 7834 10792 7840 10804
rect 7795 10764 7840 10792
rect 7834 10752 7840 10764
rect 7892 10752 7898 10804
rect 10778 10792 10784 10804
rect 10739 10764 10784 10792
rect 10778 10752 10784 10764
rect 10836 10752 10842 10804
rect 11241 10795 11299 10801
rect 11241 10761 11253 10795
rect 11287 10792 11299 10795
rect 11330 10792 11336 10804
rect 11287 10764 11336 10792
rect 11287 10761 11299 10764
rect 11241 10755 11299 10761
rect 11330 10752 11336 10764
rect 11388 10792 11394 10804
rect 11514 10792 11520 10804
rect 11388 10764 11520 10792
rect 11388 10752 11394 10764
rect 11514 10752 11520 10764
rect 11572 10752 11578 10804
rect 13081 10795 13139 10801
rect 13081 10761 13093 10795
rect 13127 10792 13139 10795
rect 13446 10792 13452 10804
rect 13127 10764 13452 10792
rect 13127 10761 13139 10764
rect 13081 10755 13139 10761
rect 13446 10752 13452 10764
rect 13504 10792 13510 10804
rect 13630 10792 13636 10804
rect 13504 10764 13636 10792
rect 13504 10752 13510 10764
rect 13630 10752 13636 10764
rect 13688 10752 13694 10804
rect 15381 10795 15439 10801
rect 15381 10761 15393 10795
rect 15427 10792 15439 10795
rect 15654 10792 15660 10804
rect 15427 10764 15660 10792
rect 15427 10761 15439 10764
rect 15381 10755 15439 10761
rect 15654 10752 15660 10764
rect 15712 10752 15718 10804
rect 17862 10792 17868 10804
rect 17823 10764 17868 10792
rect 17862 10752 17868 10764
rect 17920 10752 17926 10804
rect 20809 10795 20867 10801
rect 20809 10761 20821 10795
rect 20855 10792 20867 10795
rect 21358 10792 21364 10804
rect 20855 10764 21364 10792
rect 20855 10761 20867 10764
rect 20809 10755 20867 10761
rect 21358 10752 21364 10764
rect 21416 10752 21422 10804
rect 13354 10724 13360 10736
rect 13315 10696 13360 10724
rect 13354 10684 13360 10696
rect 13412 10724 13418 10736
rect 13725 10727 13783 10733
rect 13725 10724 13737 10727
rect 13412 10696 13737 10724
rect 13412 10684 13418 10696
rect 13725 10693 13737 10696
rect 13771 10693 13783 10727
rect 13725 10687 13783 10693
rect 19242 10656 19248 10668
rect 19155 10628 19248 10656
rect 19242 10616 19248 10628
rect 19300 10656 19306 10668
rect 20530 10656 20536 10668
rect 19300 10628 20536 10656
rect 19300 10616 19306 10628
rect 20530 10616 20536 10628
rect 20588 10616 20594 10668
rect 19521 10591 19579 10597
rect 19521 10588 19533 10591
rect 19352 10560 19533 10588
rect 19058 10520 19064 10532
rect 19019 10492 19064 10520
rect 19058 10480 19064 10492
rect 19116 10520 19122 10532
rect 19352 10520 19380 10560
rect 19521 10557 19533 10560
rect 19567 10557 19579 10591
rect 19521 10551 19579 10557
rect 19116 10492 19380 10520
rect 19116 10480 19122 10492
rect 12713 10455 12771 10461
rect 12713 10421 12725 10455
rect 12759 10452 12771 10455
rect 12802 10452 12808 10464
rect 12759 10424 12808 10452
rect 12759 10421 12771 10424
rect 12713 10415 12771 10421
rect 12802 10412 12808 10424
rect 12860 10412 12866 10464
rect 15286 10412 15292 10464
rect 15344 10452 15350 10464
rect 15657 10455 15715 10461
rect 15657 10452 15669 10455
rect 15344 10424 15669 10452
rect 15344 10412 15350 10424
rect 15657 10421 15669 10424
rect 15703 10421 15715 10455
rect 15657 10415 15715 10421
rect 1104 10362 28888 10384
rect 1104 10310 10982 10362
rect 11034 10310 11046 10362
rect 11098 10310 11110 10362
rect 11162 10310 11174 10362
rect 11226 10310 20982 10362
rect 21034 10310 21046 10362
rect 21098 10310 21110 10362
rect 21162 10310 21174 10362
rect 21226 10310 28888 10362
rect 1104 10288 28888 10310
rect 17954 10208 17960 10260
rect 18012 10248 18018 10260
rect 18785 10251 18843 10257
rect 18785 10248 18797 10251
rect 18012 10220 18797 10248
rect 18012 10208 18018 10220
rect 18785 10217 18797 10220
rect 18831 10248 18843 10251
rect 19242 10248 19248 10260
rect 18831 10220 19248 10248
rect 18831 10217 18843 10220
rect 18785 10211 18843 10217
rect 19242 10208 19248 10220
rect 19300 10208 19306 10260
rect 16390 10112 16396 10124
rect 16351 10084 16396 10112
rect 16390 10072 16396 10084
rect 16448 10072 16454 10124
rect 18046 10072 18052 10124
rect 18104 10112 18110 10124
rect 18782 10112 18788 10124
rect 18104 10084 18788 10112
rect 18104 10072 18110 10084
rect 18782 10072 18788 10084
rect 18840 10112 18846 10124
rect 18969 10115 19027 10121
rect 18969 10112 18981 10115
rect 18840 10084 18981 10112
rect 18840 10072 18846 10084
rect 18969 10081 18981 10084
rect 19015 10081 19027 10115
rect 18969 10075 19027 10081
rect 15746 10004 15752 10056
rect 15804 10044 15810 10056
rect 16301 10047 16359 10053
rect 16301 10044 16313 10047
rect 15804 10016 16313 10044
rect 15804 10004 15810 10016
rect 16301 10013 16313 10016
rect 16347 10044 16359 10047
rect 16482 10044 16488 10056
rect 16347 10016 16488 10044
rect 16347 10013 16359 10016
rect 16301 10007 16359 10013
rect 16482 10004 16488 10016
rect 16540 10004 16546 10056
rect 16574 9908 16580 9920
rect 16535 9880 16580 9908
rect 16574 9868 16580 9880
rect 16632 9868 16638 9920
rect 1104 9818 28888 9840
rect 1104 9766 5982 9818
rect 6034 9766 6046 9818
rect 6098 9766 6110 9818
rect 6162 9766 6174 9818
rect 6226 9766 15982 9818
rect 16034 9766 16046 9818
rect 16098 9766 16110 9818
rect 16162 9766 16174 9818
rect 16226 9766 25982 9818
rect 26034 9766 26046 9818
rect 26098 9766 26110 9818
rect 26162 9766 26174 9818
rect 26226 9766 28888 9818
rect 1104 9744 28888 9766
rect 12618 9664 12624 9716
rect 12676 9704 12682 9716
rect 12805 9707 12863 9713
rect 12805 9704 12817 9707
rect 12676 9676 12817 9704
rect 12676 9664 12682 9676
rect 12805 9673 12817 9676
rect 12851 9673 12863 9707
rect 12805 9667 12863 9673
rect 16390 9664 16396 9716
rect 16448 9704 16454 9716
rect 18782 9704 18788 9716
rect 16448 9676 16620 9704
rect 18743 9676 18788 9704
rect 16448 9664 16454 9676
rect 14918 9528 14924 9580
rect 14976 9568 14982 9580
rect 15013 9571 15071 9577
rect 15013 9568 15025 9571
rect 14976 9540 15025 9568
rect 14976 9528 14982 9540
rect 15013 9537 15025 9540
rect 15059 9568 15071 9571
rect 15470 9568 15476 9580
rect 15059 9540 15476 9568
rect 15059 9537 15071 9540
rect 15013 9531 15071 9537
rect 15470 9528 15476 9540
rect 15528 9528 15534 9580
rect 16592 9568 16620 9676
rect 18782 9664 18788 9676
rect 18840 9664 18846 9716
rect 20530 9596 20536 9648
rect 20588 9636 20594 9648
rect 20714 9636 20720 9648
rect 20588 9608 20720 9636
rect 20588 9596 20594 9608
rect 20714 9596 20720 9608
rect 20772 9596 20778 9648
rect 16853 9571 16911 9577
rect 16853 9568 16865 9571
rect 16592 9540 16865 9568
rect 16853 9537 16865 9540
rect 16899 9568 16911 9571
rect 17497 9571 17555 9577
rect 17497 9568 17509 9571
rect 16899 9540 17509 9568
rect 16899 9537 16911 9540
rect 16853 9531 16911 9537
rect 17497 9537 17509 9540
rect 17543 9537 17555 9571
rect 17497 9531 17555 9537
rect 12253 9503 12311 9509
rect 12253 9469 12265 9503
rect 12299 9500 12311 9503
rect 12434 9500 12440 9512
rect 12299 9472 12440 9500
rect 12299 9469 12311 9472
rect 12253 9463 12311 9469
rect 12434 9460 12440 9472
rect 12492 9500 12498 9512
rect 12529 9503 12587 9509
rect 12529 9500 12541 9503
rect 12492 9472 12541 9500
rect 12492 9460 12498 9472
rect 12529 9469 12541 9472
rect 12575 9469 12587 9503
rect 12529 9463 12587 9469
rect 12621 9503 12679 9509
rect 12621 9469 12633 9503
rect 12667 9500 12679 9503
rect 13449 9503 13507 9509
rect 13449 9500 13461 9503
rect 12667 9472 13461 9500
rect 12667 9469 12679 9472
rect 12621 9463 12679 9469
rect 13449 9469 13461 9472
rect 13495 9500 13507 9503
rect 13909 9503 13967 9509
rect 13909 9500 13921 9503
rect 13495 9472 13921 9500
rect 13495 9469 13507 9472
rect 13449 9463 13507 9469
rect 13909 9469 13921 9472
rect 13955 9500 13967 9503
rect 14458 9500 14464 9512
rect 13955 9472 14464 9500
rect 13955 9469 13967 9472
rect 13909 9463 13967 9469
rect 14458 9460 14464 9472
rect 14516 9460 14522 9512
rect 15197 9503 15255 9509
rect 15197 9469 15209 9503
rect 15243 9500 15255 9503
rect 15286 9500 15292 9512
rect 15243 9472 15292 9500
rect 15243 9469 15255 9472
rect 15197 9463 15255 9469
rect 15286 9460 15292 9472
rect 15344 9460 15350 9512
rect 16482 9460 16488 9512
rect 16540 9500 16546 9512
rect 17129 9503 17187 9509
rect 17129 9500 17141 9503
rect 16540 9472 17141 9500
rect 16540 9460 16546 9472
rect 17129 9469 17141 9472
rect 17175 9469 17187 9503
rect 17129 9463 17187 9469
rect 13262 9324 13268 9376
rect 13320 9364 13326 9376
rect 14093 9367 14151 9373
rect 14093 9364 14105 9367
rect 13320 9336 14105 9364
rect 13320 9324 13326 9336
rect 14093 9333 14105 9336
rect 14139 9333 14151 9367
rect 14093 9327 14151 9333
rect 1104 9274 28888 9296
rect 1104 9222 10982 9274
rect 11034 9222 11046 9274
rect 11098 9222 11110 9274
rect 11162 9222 11174 9274
rect 11226 9222 20982 9274
rect 21034 9222 21046 9274
rect 21098 9222 21110 9274
rect 21162 9222 21174 9274
rect 21226 9222 28888 9274
rect 1104 9200 28888 9222
rect 3050 9092 3056 9104
rect 3011 9064 3056 9092
rect 3050 9052 3056 9064
rect 3108 9052 3114 9104
rect 11606 9052 11612 9104
rect 11664 9092 11670 9104
rect 11664 9064 13124 9092
rect 11664 9052 11670 9064
rect 1397 9027 1455 9033
rect 1397 8993 1409 9027
rect 1443 9024 1455 9027
rect 2038 9024 2044 9036
rect 1443 8996 2044 9024
rect 1443 8993 1455 8996
rect 1397 8987 1455 8993
rect 2038 8984 2044 8996
rect 2096 8984 2102 9036
rect 9674 9024 9680 9036
rect 9635 8996 9680 9024
rect 9674 8984 9680 8996
rect 9732 8984 9738 9036
rect 9953 9027 10011 9033
rect 9953 8993 9965 9027
rect 9999 9024 10011 9027
rect 10318 9024 10324 9036
rect 9999 8996 10324 9024
rect 9999 8993 10011 8996
rect 9953 8987 10011 8993
rect 10318 8984 10324 8996
rect 10376 8984 10382 9036
rect 12618 9024 12624 9036
rect 12579 8996 12624 9024
rect 12618 8984 12624 8996
rect 12676 8984 12682 9036
rect 12986 9024 12992 9036
rect 12947 8996 12992 9024
rect 12986 8984 12992 8996
rect 13044 8984 13050 9036
rect 13096 9033 13124 9064
rect 15470 9052 15476 9104
rect 15528 9092 15534 9104
rect 15528 9064 16896 9092
rect 15528 9052 15534 9064
rect 13081 9027 13139 9033
rect 13081 8993 13093 9027
rect 13127 8993 13139 9027
rect 13081 8987 13139 8993
rect 16574 8984 16580 9036
rect 16632 9024 16638 9036
rect 16868 9033 16896 9064
rect 16669 9027 16727 9033
rect 16669 9024 16681 9027
rect 16632 8996 16681 9024
rect 16632 8984 16638 8996
rect 16669 8993 16681 8996
rect 16715 8993 16727 9027
rect 16669 8987 16727 8993
rect 16853 9027 16911 9033
rect 16853 8993 16865 9027
rect 16899 9024 16911 9027
rect 16942 9024 16948 9036
rect 16899 8996 16948 9024
rect 16899 8993 16911 8996
rect 16853 8987 16911 8993
rect 16942 8984 16948 8996
rect 17000 8984 17006 9036
rect 17034 8984 17040 9036
rect 17092 9024 17098 9036
rect 17586 9024 17592 9036
rect 17092 8996 17592 9024
rect 17092 8984 17098 8996
rect 17586 8984 17592 8996
rect 17644 8984 17650 9036
rect 1578 8916 1584 8968
rect 1636 8956 1642 8968
rect 1673 8959 1731 8965
rect 1673 8956 1685 8959
rect 1636 8928 1685 8956
rect 1636 8916 1642 8928
rect 1673 8925 1685 8928
rect 1719 8925 1731 8959
rect 12158 8956 12164 8968
rect 12119 8928 12164 8956
rect 1673 8919 1731 8925
rect 12158 8916 12164 8928
rect 12216 8916 12222 8968
rect 16482 8888 16488 8900
rect 16443 8860 16488 8888
rect 16482 8848 16488 8860
rect 16540 8848 16546 8900
rect 9125 8823 9183 8829
rect 9125 8789 9137 8823
rect 9171 8820 9183 8823
rect 9674 8820 9680 8832
rect 9171 8792 9680 8820
rect 9171 8789 9183 8792
rect 9125 8783 9183 8789
rect 9674 8780 9680 8792
rect 9732 8820 9738 8832
rect 11057 8823 11115 8829
rect 11057 8820 11069 8823
rect 9732 8792 11069 8820
rect 9732 8780 9738 8792
rect 11057 8789 11069 8792
rect 11103 8789 11115 8823
rect 11057 8783 11115 8789
rect 13541 8823 13599 8829
rect 13541 8789 13553 8823
rect 13587 8820 13599 8823
rect 14090 8820 14096 8832
rect 13587 8792 14096 8820
rect 13587 8789 13599 8792
rect 13541 8783 13599 8789
rect 14090 8780 14096 8792
rect 14148 8780 14154 8832
rect 15470 8820 15476 8832
rect 15431 8792 15476 8820
rect 15470 8780 15476 8792
rect 15528 8780 15534 8832
rect 1104 8730 28888 8752
rect 1104 8678 5982 8730
rect 6034 8678 6046 8730
rect 6098 8678 6110 8730
rect 6162 8678 6174 8730
rect 6226 8678 15982 8730
rect 16034 8678 16046 8730
rect 16098 8678 16110 8730
rect 16162 8678 16174 8730
rect 16226 8678 25982 8730
rect 26034 8678 26046 8730
rect 26098 8678 26110 8730
rect 26162 8678 26174 8730
rect 26226 8678 28888 8730
rect 1104 8656 28888 8678
rect 2038 8616 2044 8628
rect 1999 8588 2044 8616
rect 2038 8576 2044 8588
rect 2096 8576 2102 8628
rect 8846 8616 8852 8628
rect 8807 8588 8852 8616
rect 8846 8576 8852 8588
rect 8904 8616 8910 8628
rect 10226 8616 10232 8628
rect 8904 8588 10232 8616
rect 8904 8576 8910 8588
rect 10226 8576 10232 8588
rect 10284 8576 10290 8628
rect 10318 8576 10324 8628
rect 10376 8616 10382 8628
rect 10505 8619 10563 8625
rect 10505 8616 10517 8619
rect 10376 8588 10517 8616
rect 10376 8576 10382 8588
rect 10505 8585 10517 8588
rect 10551 8585 10563 8619
rect 10505 8579 10563 8585
rect 10594 8576 10600 8628
rect 10652 8616 10658 8628
rect 12161 8619 12219 8625
rect 12161 8616 12173 8619
rect 10652 8588 12173 8616
rect 10652 8576 10658 8588
rect 12161 8585 12173 8588
rect 12207 8585 12219 8619
rect 12618 8616 12624 8628
rect 12579 8588 12624 8616
rect 12161 8579 12219 8585
rect 8573 8551 8631 8557
rect 8573 8517 8585 8551
rect 8619 8548 8631 8551
rect 10336 8548 10364 8576
rect 8619 8520 10364 8548
rect 8619 8517 8631 8520
rect 8573 8511 8631 8517
rect 9493 8415 9551 8421
rect 9493 8381 9505 8415
rect 9539 8381 9551 8415
rect 9674 8412 9680 8424
rect 9635 8384 9680 8412
rect 9493 8375 9551 8381
rect 1578 8344 1584 8356
rect 1539 8316 1584 8344
rect 1578 8304 1584 8316
rect 1636 8304 1642 8356
rect 9030 8344 9036 8356
rect 8991 8316 9036 8344
rect 9030 8304 9036 8316
rect 9088 8304 9094 8356
rect 9508 8344 9536 8375
rect 9674 8372 9680 8384
rect 9732 8372 9738 8424
rect 10060 8421 10088 8520
rect 11606 8508 11612 8560
rect 11664 8548 11670 8560
rect 11793 8551 11851 8557
rect 11793 8548 11805 8551
rect 11664 8520 11805 8548
rect 11664 8508 11670 8520
rect 11793 8517 11805 8520
rect 11839 8517 11851 8551
rect 12176 8548 12204 8579
rect 12618 8576 12624 8588
rect 12676 8576 12682 8628
rect 13998 8576 14004 8628
rect 14056 8616 14062 8628
rect 15562 8616 15568 8628
rect 14056 8588 15568 8616
rect 14056 8576 14062 8588
rect 15562 8576 15568 8588
rect 15620 8576 15626 8628
rect 16574 8616 16580 8628
rect 16535 8588 16580 8616
rect 16574 8576 16580 8588
rect 16632 8576 16638 8628
rect 16942 8616 16948 8628
rect 16903 8588 16948 8616
rect 16942 8576 16948 8588
rect 17000 8576 17006 8628
rect 12986 8548 12992 8560
rect 12176 8520 12992 8548
rect 11793 8511 11851 8517
rect 12986 8508 12992 8520
rect 13044 8508 13050 8560
rect 13262 8508 13268 8560
rect 13320 8548 13326 8560
rect 16301 8551 16359 8557
rect 13320 8520 14412 8548
rect 13320 8508 13326 8520
rect 13722 8480 13728 8492
rect 13683 8452 13728 8480
rect 13722 8440 13728 8452
rect 13780 8440 13786 8492
rect 13998 8480 14004 8492
rect 13959 8452 14004 8480
rect 13998 8440 14004 8452
rect 14056 8440 14062 8492
rect 14384 8489 14412 8520
rect 16301 8517 16313 8551
rect 16347 8548 16359 8551
rect 17034 8548 17040 8560
rect 16347 8520 17040 8548
rect 16347 8517 16359 8520
rect 16301 8511 16359 8517
rect 17034 8508 17040 8520
rect 17092 8508 17098 8560
rect 14369 8483 14427 8489
rect 14369 8449 14381 8483
rect 14415 8449 14427 8483
rect 14369 8443 14427 8449
rect 10016 8415 10088 8421
rect 10016 8381 10028 8415
rect 10062 8384 10088 8415
rect 10226 8412 10232 8424
rect 10187 8384 10232 8412
rect 10062 8381 10074 8384
rect 10016 8375 10074 8381
rect 10226 8372 10232 8384
rect 10284 8412 10290 8424
rect 13262 8412 13268 8424
rect 10284 8384 13268 8412
rect 10284 8372 10290 8384
rect 13262 8372 13268 8384
rect 13320 8372 13326 8424
rect 14090 8412 14096 8424
rect 14051 8384 14096 8412
rect 14090 8372 14096 8384
rect 14148 8372 14154 8424
rect 14461 8415 14519 8421
rect 14461 8381 14473 8415
rect 14507 8381 14519 8415
rect 14461 8375 14519 8381
rect 9858 8344 9864 8356
rect 9508 8316 9864 8344
rect 9122 8236 9128 8288
rect 9180 8276 9186 8288
rect 9508 8276 9536 8316
rect 9858 8304 9864 8316
rect 9916 8304 9922 8356
rect 13814 8304 13820 8356
rect 13872 8344 13878 8356
rect 14476 8344 14504 8375
rect 13872 8316 14504 8344
rect 13872 8304 13878 8316
rect 9180 8248 9536 8276
rect 9180 8236 9186 8248
rect 1104 8186 28888 8208
rect 1104 8134 10982 8186
rect 11034 8134 11046 8186
rect 11098 8134 11110 8186
rect 11162 8134 11174 8186
rect 11226 8134 20982 8186
rect 21034 8134 21046 8186
rect 21098 8134 21110 8186
rect 21162 8134 21174 8186
rect 21226 8134 28888 8186
rect 1104 8112 28888 8134
rect 9122 8072 9128 8084
rect 9083 8044 9128 8072
rect 9122 8032 9128 8044
rect 9180 8032 9186 8084
rect 9766 8032 9772 8084
rect 9824 8072 9830 8084
rect 9861 8075 9919 8081
rect 9861 8072 9873 8075
rect 9824 8044 9873 8072
rect 9824 8032 9830 8044
rect 9861 8041 9873 8044
rect 9907 8041 9919 8075
rect 9861 8035 9919 8041
rect 9876 7936 9904 8035
rect 12434 8032 12440 8084
rect 12492 8072 12498 8084
rect 13814 8072 13820 8084
rect 12492 8044 12537 8072
rect 13775 8044 13820 8072
rect 12492 8032 12498 8044
rect 13814 8032 13820 8044
rect 13872 8032 13878 8084
rect 18138 8072 18144 8084
rect 18099 8044 18144 8072
rect 18138 8032 18144 8044
rect 18196 8032 18202 8084
rect 13446 7964 13452 8016
rect 13504 8004 13510 8016
rect 13541 8007 13599 8013
rect 13541 8004 13553 8007
rect 13504 7976 13553 8004
rect 13504 7964 13510 7976
rect 13541 7973 13553 7976
rect 13587 8004 13599 8007
rect 13998 8004 14004 8016
rect 13587 7976 14004 8004
rect 13587 7973 13599 7976
rect 13541 7967 13599 7973
rect 13998 7964 14004 7976
rect 14056 7964 14062 8016
rect 11054 7936 11060 7948
rect 9876 7908 11060 7936
rect 11054 7896 11060 7908
rect 11112 7896 11118 7948
rect 11333 7939 11391 7945
rect 11333 7905 11345 7939
rect 11379 7936 11391 7939
rect 11606 7936 11612 7948
rect 11379 7908 11612 7936
rect 11379 7905 11391 7908
rect 11333 7899 11391 7905
rect 11606 7896 11612 7908
rect 11664 7896 11670 7948
rect 16850 7936 16856 7948
rect 16811 7908 16856 7936
rect 16850 7896 16856 7908
rect 16908 7896 16914 7948
rect 16577 7871 16635 7877
rect 16577 7837 16589 7871
rect 16623 7868 16635 7871
rect 16942 7868 16948 7880
rect 16623 7840 16948 7868
rect 16623 7837 16635 7840
rect 16577 7831 16635 7837
rect 16942 7828 16948 7840
rect 17000 7828 17006 7880
rect 1104 7642 28888 7664
rect 1104 7590 5982 7642
rect 6034 7590 6046 7642
rect 6098 7590 6110 7642
rect 6162 7590 6174 7642
rect 6226 7590 15982 7642
rect 16034 7590 16046 7642
rect 16098 7590 16110 7642
rect 16162 7590 16174 7642
rect 16226 7590 25982 7642
rect 26034 7590 26046 7642
rect 26098 7590 26110 7642
rect 26162 7590 26174 7642
rect 26226 7590 28888 7642
rect 1104 7568 28888 7590
rect 11149 7531 11207 7537
rect 11149 7497 11161 7531
rect 11195 7528 11207 7531
rect 11606 7528 11612 7540
rect 11195 7500 11612 7528
rect 11195 7497 11207 7500
rect 11149 7491 11207 7497
rect 11606 7488 11612 7500
rect 11664 7488 11670 7540
rect 14090 7488 14096 7540
rect 14148 7528 14154 7540
rect 14461 7531 14519 7537
rect 14461 7528 14473 7531
rect 14148 7500 14473 7528
rect 14148 7488 14154 7500
rect 14461 7497 14473 7500
rect 14507 7497 14519 7531
rect 14461 7491 14519 7497
rect 16669 7531 16727 7537
rect 16669 7497 16681 7531
rect 16715 7528 16727 7531
rect 16850 7528 16856 7540
rect 16715 7500 16856 7528
rect 16715 7497 16727 7500
rect 16669 7491 16727 7497
rect 16850 7488 16856 7500
rect 16908 7488 16914 7540
rect 16942 7488 16948 7540
rect 17000 7528 17006 7540
rect 17037 7531 17095 7537
rect 17037 7528 17049 7531
rect 17000 7500 17049 7528
rect 17000 7488 17006 7500
rect 17037 7497 17049 7500
rect 17083 7528 17095 7531
rect 17862 7528 17868 7540
rect 17083 7500 17868 7528
rect 17083 7497 17095 7500
rect 17037 7491 17095 7497
rect 17862 7488 17868 7500
rect 17920 7488 17926 7540
rect 11054 7420 11060 7472
rect 11112 7460 11118 7472
rect 11425 7463 11483 7469
rect 11425 7460 11437 7463
rect 11112 7432 11437 7460
rect 11112 7420 11118 7432
rect 11425 7429 11437 7432
rect 11471 7429 11483 7463
rect 11425 7423 11483 7429
rect 12989 7395 13047 7401
rect 12989 7361 13001 7395
rect 13035 7392 13047 7395
rect 13357 7395 13415 7401
rect 13357 7392 13369 7395
rect 13035 7364 13369 7392
rect 13035 7361 13047 7364
rect 12989 7355 13047 7361
rect 13357 7361 13369 7364
rect 13403 7392 13415 7395
rect 13814 7392 13820 7404
rect 13403 7364 13820 7392
rect 13403 7361 13415 7364
rect 13357 7355 13415 7361
rect 13814 7352 13820 7364
rect 13872 7352 13878 7404
rect 13078 7324 13084 7336
rect 13039 7296 13084 7324
rect 13078 7284 13084 7296
rect 13136 7284 13142 7336
rect 1104 7098 28888 7120
rect 1104 7046 10982 7098
rect 11034 7046 11046 7098
rect 11098 7046 11110 7098
rect 11162 7046 11174 7098
rect 11226 7046 20982 7098
rect 21034 7046 21046 7098
rect 21098 7046 21110 7098
rect 21162 7046 21174 7098
rect 21226 7046 28888 7098
rect 1104 7024 28888 7046
rect 13078 6644 13084 6656
rect 13039 6616 13084 6644
rect 13078 6604 13084 6616
rect 13136 6644 13142 6656
rect 14550 6644 14556 6656
rect 13136 6616 14556 6644
rect 13136 6604 13142 6616
rect 14550 6604 14556 6616
rect 14608 6604 14614 6656
rect 1104 6554 28888 6576
rect 1104 6502 5982 6554
rect 6034 6502 6046 6554
rect 6098 6502 6110 6554
rect 6162 6502 6174 6554
rect 6226 6502 15982 6554
rect 16034 6502 16046 6554
rect 16098 6502 16110 6554
rect 16162 6502 16174 6554
rect 16226 6502 25982 6554
rect 26034 6502 26046 6554
rect 26098 6502 26110 6554
rect 26162 6502 26174 6554
rect 26226 6502 28888 6554
rect 1104 6480 28888 6502
rect 14182 6400 14188 6452
rect 14240 6440 14246 6452
rect 14369 6443 14427 6449
rect 14369 6440 14381 6443
rect 14240 6412 14381 6440
rect 14240 6400 14246 6412
rect 14369 6409 14381 6412
rect 14415 6409 14427 6443
rect 14369 6403 14427 6409
rect 14384 6304 14412 6403
rect 14829 6307 14887 6313
rect 14829 6304 14841 6307
rect 14384 6276 14841 6304
rect 14829 6273 14841 6276
rect 14875 6304 14887 6307
rect 16298 6304 16304 6316
rect 14875 6276 16304 6304
rect 14875 6273 14887 6276
rect 14829 6267 14887 6273
rect 16298 6264 16304 6276
rect 16356 6264 16362 6316
rect 14550 6236 14556 6248
rect 14511 6208 14556 6236
rect 14550 6196 14556 6208
rect 14608 6196 14614 6248
rect 15930 6100 15936 6112
rect 15891 6072 15936 6100
rect 15930 6060 15936 6072
rect 15988 6060 15994 6112
rect 1104 6010 28888 6032
rect 1104 5958 10982 6010
rect 11034 5958 11046 6010
rect 11098 5958 11110 6010
rect 11162 5958 11174 6010
rect 11226 5958 20982 6010
rect 21034 5958 21046 6010
rect 21098 5958 21110 6010
rect 21162 5958 21174 6010
rect 21226 5958 28888 6010
rect 1104 5936 28888 5958
rect 13354 5788 13360 5840
rect 13412 5828 13418 5840
rect 15286 5828 15292 5840
rect 13412 5800 15292 5828
rect 13412 5788 13418 5800
rect 13814 5760 13820 5772
rect 13775 5732 13820 5760
rect 13814 5720 13820 5732
rect 13872 5720 13878 5772
rect 14182 5760 14188 5772
rect 14143 5732 14188 5760
rect 14182 5720 14188 5732
rect 14240 5720 14246 5772
rect 14384 5769 14412 5800
rect 15286 5788 15292 5800
rect 15344 5828 15350 5840
rect 15746 5828 15752 5840
rect 15344 5800 15752 5828
rect 15344 5788 15350 5800
rect 15746 5788 15752 5800
rect 15804 5828 15810 5840
rect 15804 5800 16436 5828
rect 15804 5788 15810 5800
rect 14369 5763 14427 5769
rect 14369 5729 14381 5763
rect 14415 5729 14427 5763
rect 15930 5760 15936 5772
rect 15891 5732 15936 5760
rect 14369 5723 14427 5729
rect 15930 5720 15936 5732
rect 15988 5720 15994 5772
rect 16298 5760 16304 5772
rect 16259 5732 16304 5760
rect 16298 5720 16304 5732
rect 16356 5720 16362 5772
rect 16408 5769 16436 5800
rect 16393 5763 16451 5769
rect 16393 5729 16405 5763
rect 16439 5729 16451 5763
rect 16393 5723 16451 5729
rect 13722 5652 13728 5704
rect 13780 5692 13786 5704
rect 13909 5695 13967 5701
rect 13909 5692 13921 5695
rect 13780 5664 13921 5692
rect 13780 5652 13786 5664
rect 13909 5661 13921 5664
rect 13955 5692 13967 5695
rect 13998 5692 14004 5704
rect 13955 5664 14004 5692
rect 13955 5661 13967 5664
rect 13909 5655 13967 5661
rect 13998 5652 14004 5664
rect 14056 5652 14062 5704
rect 15749 5695 15807 5701
rect 15749 5661 15761 5695
rect 15795 5661 15807 5695
rect 15749 5655 15807 5661
rect 14016 5624 14044 5652
rect 15654 5624 15660 5636
rect 14016 5596 15660 5624
rect 15654 5584 15660 5596
rect 15712 5624 15718 5636
rect 15764 5624 15792 5655
rect 15712 5596 15792 5624
rect 15712 5584 15718 5596
rect 13078 5556 13084 5568
rect 13039 5528 13084 5556
rect 13078 5516 13084 5528
rect 13136 5516 13142 5568
rect 13446 5556 13452 5568
rect 13407 5528 13452 5556
rect 13446 5516 13452 5528
rect 13504 5516 13510 5568
rect 15562 5556 15568 5568
rect 15523 5528 15568 5556
rect 15562 5516 15568 5528
rect 15620 5516 15626 5568
rect 1104 5466 28888 5488
rect 1104 5414 5982 5466
rect 6034 5414 6046 5466
rect 6098 5414 6110 5466
rect 6162 5414 6174 5466
rect 6226 5414 15982 5466
rect 16034 5414 16046 5466
rect 16098 5414 16110 5466
rect 16162 5414 16174 5466
rect 16226 5414 25982 5466
rect 26034 5414 26046 5466
rect 26098 5414 26110 5466
rect 26162 5414 26174 5466
rect 26226 5414 28888 5466
rect 1104 5392 28888 5414
rect 11422 5312 11428 5364
rect 11480 5352 11486 5364
rect 12161 5355 12219 5361
rect 12161 5352 12173 5355
rect 11480 5324 12173 5352
rect 11480 5312 11486 5324
rect 12161 5321 12173 5324
rect 12207 5321 12219 5355
rect 12161 5315 12219 5321
rect 12989 5355 13047 5361
rect 12989 5321 13001 5355
rect 13035 5352 13047 5355
rect 13354 5352 13360 5364
rect 13035 5324 13360 5352
rect 13035 5321 13047 5324
rect 12989 5315 13047 5321
rect 12176 5216 12204 5315
rect 13354 5312 13360 5324
rect 13412 5312 13418 5364
rect 15286 5352 15292 5364
rect 15247 5324 15292 5352
rect 15286 5312 15292 5324
rect 15344 5312 15350 5364
rect 15654 5352 15660 5364
rect 15615 5324 15660 5352
rect 15654 5312 15660 5324
rect 15712 5312 15718 5364
rect 15838 5312 15844 5364
rect 15896 5352 15902 5364
rect 16025 5355 16083 5361
rect 16025 5352 16037 5355
rect 15896 5324 16037 5352
rect 15896 5312 15902 5324
rect 16025 5321 16037 5324
rect 16071 5321 16083 5355
rect 16025 5315 16083 5321
rect 12176 5188 13400 5216
rect 13078 5148 13084 5160
rect 13039 5120 13084 5148
rect 13078 5108 13084 5120
rect 13136 5108 13142 5160
rect 13372 5157 13400 5188
rect 13357 5151 13415 5157
rect 13357 5117 13369 5151
rect 13403 5148 13415 5151
rect 14182 5148 14188 5160
rect 13403 5120 14188 5148
rect 13403 5117 13415 5120
rect 13357 5111 13415 5117
rect 14182 5108 14188 5120
rect 14240 5108 14246 5160
rect 13630 4972 13636 5024
rect 13688 5012 13694 5024
rect 13814 5012 13820 5024
rect 13688 4984 13820 5012
rect 13688 4972 13694 4984
rect 13814 4972 13820 4984
rect 13872 5012 13878 5024
rect 14461 5015 14519 5021
rect 14461 5012 14473 5015
rect 13872 4984 14473 5012
rect 13872 4972 13878 4984
rect 14461 4981 14473 4984
rect 14507 4981 14519 5015
rect 14461 4975 14519 4981
rect 1104 4922 28888 4944
rect 1104 4870 10982 4922
rect 11034 4870 11046 4922
rect 11098 4870 11110 4922
rect 11162 4870 11174 4922
rect 11226 4870 20982 4922
rect 21034 4870 21046 4922
rect 21098 4870 21110 4922
rect 21162 4870 21174 4922
rect 21226 4870 28888 4922
rect 1104 4848 28888 4870
rect 13630 4808 13636 4820
rect 13591 4780 13636 4808
rect 13630 4768 13636 4780
rect 13688 4768 13694 4820
rect 14001 4811 14059 4817
rect 14001 4777 14013 4811
rect 14047 4808 14059 4811
rect 14182 4808 14188 4820
rect 14047 4780 14188 4808
rect 14047 4777 14059 4780
rect 14001 4771 14059 4777
rect 14182 4768 14188 4780
rect 14240 4768 14246 4820
rect 15565 4811 15623 4817
rect 15565 4777 15577 4811
rect 15611 4808 15623 4811
rect 16298 4808 16304 4820
rect 15611 4780 16304 4808
rect 15611 4777 15623 4780
rect 15565 4771 15623 4777
rect 16298 4768 16304 4780
rect 16356 4768 16362 4820
rect 12621 4743 12679 4749
rect 12621 4709 12633 4743
rect 12667 4740 12679 4743
rect 13538 4740 13544 4752
rect 12667 4712 13544 4740
rect 12667 4709 12679 4712
rect 12621 4703 12679 4709
rect 13538 4700 13544 4712
rect 13596 4700 13602 4752
rect 10870 4632 10876 4684
rect 10928 4672 10934 4684
rect 10965 4675 11023 4681
rect 10965 4672 10977 4675
rect 10928 4644 10977 4672
rect 10928 4632 10934 4644
rect 10965 4641 10977 4644
rect 11011 4641 11023 4675
rect 10965 4635 11023 4641
rect 11241 4675 11299 4681
rect 11241 4641 11253 4675
rect 11287 4672 11299 4675
rect 11514 4672 11520 4684
rect 11287 4644 11520 4672
rect 11287 4641 11299 4644
rect 11241 4635 11299 4641
rect 11514 4632 11520 4644
rect 11572 4632 11578 4684
rect 13265 4675 13323 4681
rect 13265 4641 13277 4675
rect 13311 4672 13323 4675
rect 13722 4672 13728 4684
rect 13311 4644 13728 4672
rect 13311 4641 13323 4644
rect 13265 4635 13323 4641
rect 13722 4632 13728 4644
rect 13780 4632 13786 4684
rect 1104 4378 28888 4400
rect 1104 4326 5982 4378
rect 6034 4326 6046 4378
rect 6098 4326 6110 4378
rect 6162 4326 6174 4378
rect 6226 4326 15982 4378
rect 16034 4326 16046 4378
rect 16098 4326 16110 4378
rect 16162 4326 16174 4378
rect 16226 4326 25982 4378
rect 26034 4326 26046 4378
rect 26098 4326 26110 4378
rect 26162 4326 26174 4378
rect 26226 4326 28888 4378
rect 1104 4304 28888 4326
rect 2774 4088 2780 4140
rect 2832 4128 2838 4140
rect 3694 4128 3700 4140
rect 2832 4100 3700 4128
rect 2832 4088 2838 4100
rect 3694 4088 3700 4100
rect 3752 4088 3758 4140
rect 10870 4088 10876 4140
rect 10928 4128 10934 4140
rect 11333 4131 11391 4137
rect 11333 4128 11345 4131
rect 10928 4100 11345 4128
rect 10928 4088 10934 4100
rect 11333 4097 11345 4100
rect 11379 4097 11391 4131
rect 11333 4091 11391 4097
rect 13814 4088 13820 4140
rect 13872 4128 13878 4140
rect 15102 4128 15108 4140
rect 13872 4100 15108 4128
rect 13872 4088 13878 4100
rect 15102 4088 15108 4100
rect 15160 4088 15166 4140
rect 11057 3995 11115 4001
rect 11057 3961 11069 3995
rect 11103 3992 11115 3995
rect 11514 3992 11520 4004
rect 11103 3964 11520 3992
rect 11103 3961 11115 3964
rect 11057 3955 11115 3961
rect 11514 3952 11520 3964
rect 11572 3952 11578 4004
rect 1104 3834 28888 3856
rect 1104 3782 10982 3834
rect 11034 3782 11046 3834
rect 11098 3782 11110 3834
rect 11162 3782 11174 3834
rect 11226 3782 20982 3834
rect 21034 3782 21046 3834
rect 21098 3782 21110 3834
rect 21162 3782 21174 3834
rect 21226 3782 28888 3834
rect 1104 3760 28888 3782
rect 9858 3680 9864 3732
rect 9916 3720 9922 3732
rect 9953 3723 10011 3729
rect 9953 3720 9965 3723
rect 9916 3692 9965 3720
rect 9916 3680 9922 3692
rect 9953 3689 9965 3692
rect 9999 3720 10011 3723
rect 10778 3720 10784 3732
rect 9999 3692 10784 3720
rect 9999 3689 10011 3692
rect 9953 3683 10011 3689
rect 10428 3593 10456 3692
rect 10778 3680 10784 3692
rect 10836 3680 10842 3732
rect 11790 3720 11796 3732
rect 11751 3692 11796 3720
rect 11790 3680 11796 3692
rect 11848 3680 11854 3732
rect 19426 3720 19432 3732
rect 19387 3692 19432 3720
rect 19426 3680 19432 3692
rect 19484 3680 19490 3732
rect 10413 3587 10471 3593
rect 10413 3553 10425 3587
rect 10459 3553 10471 3587
rect 10413 3547 10471 3553
rect 17865 3587 17923 3593
rect 17865 3553 17877 3587
rect 17911 3584 17923 3587
rect 17954 3584 17960 3596
rect 17911 3556 17960 3584
rect 17911 3553 17923 3556
rect 17865 3547 17923 3553
rect 17954 3544 17960 3556
rect 18012 3544 18018 3596
rect 10594 3476 10600 3528
rect 10652 3516 10658 3528
rect 10689 3519 10747 3525
rect 10689 3516 10701 3519
rect 10652 3488 10701 3516
rect 10652 3476 10658 3488
rect 10689 3485 10701 3488
rect 10735 3485 10747 3519
rect 18138 3516 18144 3528
rect 18099 3488 18144 3516
rect 10689 3479 10747 3485
rect 18138 3476 18144 3488
rect 18196 3476 18202 3528
rect 1104 3290 28888 3312
rect 1104 3238 5982 3290
rect 6034 3238 6046 3290
rect 6098 3238 6110 3290
rect 6162 3238 6174 3290
rect 6226 3238 15982 3290
rect 16034 3238 16046 3290
rect 16098 3238 16110 3290
rect 16162 3238 16174 3290
rect 16226 3238 25982 3290
rect 26034 3238 26046 3290
rect 26098 3238 26110 3290
rect 26162 3238 26174 3290
rect 26226 3238 28888 3290
rect 1104 3216 28888 3238
rect 11330 3136 11336 3188
rect 11388 3176 11394 3188
rect 11425 3179 11483 3185
rect 11425 3176 11437 3179
rect 11388 3148 11437 3176
rect 11388 3136 11394 3148
rect 11425 3145 11437 3148
rect 11471 3145 11483 3179
rect 11425 3139 11483 3145
rect 18138 3136 18144 3188
rect 18196 3176 18202 3188
rect 18233 3179 18291 3185
rect 18233 3176 18245 3179
rect 18196 3148 18245 3176
rect 18196 3136 18202 3148
rect 18233 3145 18245 3148
rect 18279 3176 18291 3179
rect 18414 3176 18420 3188
rect 18279 3148 18420 3176
rect 18279 3145 18291 3148
rect 18233 3139 18291 3145
rect 18414 3136 18420 3148
rect 18472 3136 18478 3188
rect 17954 3068 17960 3120
rect 18012 3108 18018 3120
rect 18601 3111 18659 3117
rect 18601 3108 18613 3111
rect 18012 3080 18613 3108
rect 18012 3068 18018 3080
rect 18601 3077 18613 3080
rect 18647 3077 18659 3111
rect 18601 3071 18659 3077
rect 9769 3043 9827 3049
rect 9769 3009 9781 3043
rect 9815 3040 9827 3043
rect 10134 3040 10140 3052
rect 9815 3012 10140 3040
rect 9815 3009 9827 3012
rect 9769 3003 9827 3009
rect 10134 3000 10140 3012
rect 10192 3000 10198 3052
rect 9858 2972 9864 2984
rect 9819 2944 9864 2972
rect 9858 2932 9864 2944
rect 9916 2932 9922 2984
rect 1104 2746 28888 2768
rect 1104 2694 10982 2746
rect 11034 2694 11046 2746
rect 11098 2694 11110 2746
rect 11162 2694 11174 2746
rect 11226 2694 20982 2746
rect 21034 2694 21046 2746
rect 21098 2694 21110 2746
rect 21162 2694 21174 2746
rect 21226 2694 28888 2746
rect 1104 2672 28888 2694
rect 10778 2632 10784 2644
rect 10739 2604 10784 2632
rect 10778 2592 10784 2604
rect 10836 2592 10842 2644
rect 13998 2632 14004 2644
rect 13959 2604 14004 2632
rect 13998 2592 14004 2604
rect 14056 2592 14062 2644
rect 17773 2635 17831 2641
rect 17773 2601 17785 2635
rect 17819 2632 17831 2635
rect 17954 2632 17960 2644
rect 17819 2604 17960 2632
rect 17819 2601 17831 2604
rect 17773 2595 17831 2601
rect 17954 2592 17960 2604
rect 18012 2632 18018 2644
rect 20533 2635 20591 2641
rect 20533 2632 20545 2635
rect 18012 2604 20545 2632
rect 18012 2592 18018 2604
rect 20533 2601 20545 2604
rect 20579 2632 20591 2635
rect 21450 2632 21456 2644
rect 20579 2604 21456 2632
rect 20579 2601 20591 2604
rect 20533 2595 20591 2601
rect 21450 2592 21456 2604
rect 21508 2592 21514 2644
rect 12434 2456 12440 2508
rect 12492 2496 12498 2508
rect 12897 2499 12955 2505
rect 12897 2496 12909 2499
rect 12492 2468 12909 2496
rect 12492 2456 12498 2468
rect 12897 2465 12909 2468
rect 12943 2465 12955 2499
rect 12897 2459 12955 2465
rect 18141 2499 18199 2505
rect 18141 2465 18153 2499
rect 18187 2496 18199 2499
rect 21729 2499 21787 2505
rect 21729 2496 21741 2499
rect 18187 2468 18644 2496
rect 18187 2465 18199 2468
rect 18141 2459 18199 2465
rect 18616 2440 18644 2468
rect 20916 2468 21741 2496
rect 12069 2431 12127 2437
rect 12069 2397 12081 2431
rect 12115 2428 12127 2431
rect 12621 2431 12679 2437
rect 12621 2428 12633 2431
rect 12115 2400 12633 2428
rect 12115 2397 12127 2400
rect 12069 2391 12127 2397
rect 12621 2397 12633 2400
rect 12667 2428 12679 2431
rect 13078 2428 13084 2440
rect 12667 2400 13084 2428
rect 12667 2397 12679 2400
rect 12621 2391 12679 2397
rect 13078 2388 13084 2400
rect 13136 2388 13142 2440
rect 17954 2388 17960 2440
rect 18012 2428 18018 2440
rect 18325 2431 18383 2437
rect 18325 2428 18337 2431
rect 18012 2400 18337 2428
rect 18012 2388 18018 2400
rect 18325 2397 18337 2400
rect 18371 2397 18383 2431
rect 18598 2428 18604 2440
rect 18559 2400 18604 2428
rect 18325 2391 18383 2397
rect 18598 2388 18604 2400
rect 18656 2388 18662 2440
rect 20916 2372 20944 2468
rect 21729 2465 21741 2468
rect 21775 2465 21787 2499
rect 21729 2459 21787 2465
rect 21450 2428 21456 2440
rect 21411 2400 21456 2428
rect 21450 2388 21456 2400
rect 21508 2388 21514 2440
rect 20254 2320 20260 2372
rect 20312 2360 20318 2372
rect 20622 2360 20628 2372
rect 20312 2332 20628 2360
rect 20312 2320 20318 2332
rect 20622 2320 20628 2332
rect 20680 2320 20686 2372
rect 20898 2360 20904 2372
rect 20859 2332 20904 2360
rect 20898 2320 20904 2332
rect 20956 2320 20962 2372
rect 10505 2295 10563 2301
rect 10505 2261 10517 2295
rect 10551 2292 10563 2295
rect 10594 2292 10600 2304
rect 10551 2264 10600 2292
rect 10551 2261 10563 2264
rect 10505 2255 10563 2261
rect 10594 2252 10600 2264
rect 10652 2252 10658 2304
rect 12434 2292 12440 2304
rect 12395 2264 12440 2292
rect 12434 2252 12440 2264
rect 12492 2252 12498 2304
rect 18138 2252 18144 2304
rect 18196 2292 18202 2304
rect 19705 2295 19763 2301
rect 19705 2292 19717 2295
rect 18196 2264 19717 2292
rect 18196 2252 18202 2264
rect 19705 2261 19717 2264
rect 19751 2261 19763 2295
rect 19705 2255 19763 2261
rect 23017 2295 23075 2301
rect 23017 2261 23029 2295
rect 23063 2292 23075 2295
rect 24854 2292 24860 2304
rect 23063 2264 24860 2292
rect 23063 2261 23075 2264
rect 23017 2255 23075 2261
rect 24854 2252 24860 2264
rect 24912 2252 24918 2304
rect 1104 2202 28888 2224
rect 1104 2150 5982 2202
rect 6034 2150 6046 2202
rect 6098 2150 6110 2202
rect 6162 2150 6174 2202
rect 6226 2150 15982 2202
rect 16034 2150 16046 2202
rect 16098 2150 16110 2202
rect 16162 2150 16174 2202
rect 16226 2150 25982 2202
rect 26034 2150 26046 2202
rect 26098 2150 26110 2202
rect 26162 2150 26174 2202
rect 26226 2150 28888 2202
rect 1104 2128 28888 2150
<< via1 >>
rect 10982 77766 11034 77818
rect 11046 77766 11098 77818
rect 11110 77766 11162 77818
rect 11174 77766 11226 77818
rect 20982 77766 21034 77818
rect 21046 77766 21098 77818
rect 21110 77766 21162 77818
rect 21174 77766 21226 77818
rect 3332 77324 3384 77376
rect 10324 77324 10376 77376
rect 13820 77367 13872 77376
rect 13820 77333 13829 77367
rect 13829 77333 13863 77367
rect 13863 77333 13872 77367
rect 13820 77324 13872 77333
rect 23848 77324 23900 77376
rect 25872 77324 25924 77376
rect 5982 77222 6034 77274
rect 6046 77222 6098 77274
rect 6110 77222 6162 77274
rect 6174 77222 6226 77274
rect 15982 77222 16034 77274
rect 16046 77222 16098 77274
rect 16110 77222 16162 77274
rect 16174 77222 16226 77274
rect 25982 77222 26034 77274
rect 26046 77222 26098 77274
rect 26110 77222 26162 77274
rect 26174 77222 26226 77274
rect 17500 77120 17552 77172
rect 14280 76984 14332 77036
rect 13820 76959 13872 76968
rect 13820 76925 13829 76959
rect 13829 76925 13863 76959
rect 13863 76925 13872 76959
rect 13820 76916 13872 76925
rect 19340 76959 19392 76968
rect 19340 76925 19349 76959
rect 19349 76925 19383 76959
rect 19383 76925 19392 76959
rect 19340 76916 19392 76925
rect 22744 76848 22796 76900
rect 15292 76780 15344 76832
rect 10982 76678 11034 76730
rect 11046 76678 11098 76730
rect 11110 76678 11162 76730
rect 11174 76678 11226 76730
rect 20982 76678 21034 76730
rect 21046 76678 21098 76730
rect 21110 76678 21162 76730
rect 21174 76678 21226 76730
rect 8760 76440 8812 76492
rect 9772 76440 9824 76492
rect 20812 76440 20864 76492
rect 10048 76372 10100 76424
rect 12348 76372 12400 76424
rect 12440 76415 12492 76424
rect 12440 76381 12449 76415
rect 12449 76381 12483 76415
rect 12483 76381 12492 76415
rect 12440 76372 12492 76381
rect 19248 76372 19300 76424
rect 21364 76372 21416 76424
rect 13728 76347 13780 76356
rect 13728 76313 13737 76347
rect 13737 76313 13771 76347
rect 13771 76313 13780 76347
rect 13728 76304 13780 76313
rect 11612 76236 11664 76288
rect 22652 76236 22704 76288
rect 5982 76134 6034 76186
rect 6046 76134 6098 76186
rect 6110 76134 6162 76186
rect 6174 76134 6226 76186
rect 15982 76134 16034 76186
rect 16046 76134 16098 76186
rect 16110 76134 16162 76186
rect 16174 76134 16226 76186
rect 25982 76134 26034 76186
rect 26046 76134 26098 76186
rect 26110 76134 26162 76186
rect 26174 76134 26226 76186
rect 9772 76075 9824 76084
rect 9772 76041 9781 76075
rect 9781 76041 9815 76075
rect 9815 76041 9824 76075
rect 9772 76032 9824 76041
rect 20812 76032 20864 76084
rect 12440 75896 12492 75948
rect 1400 75828 1452 75880
rect 1860 75828 1912 75880
rect 12164 75871 12216 75880
rect 12164 75837 12173 75871
rect 12173 75837 12207 75871
rect 12207 75837 12216 75871
rect 13544 75871 13596 75880
rect 12164 75828 12216 75837
rect 10140 75735 10192 75744
rect 10140 75701 10149 75735
rect 10149 75701 10183 75735
rect 10183 75701 10192 75735
rect 10140 75692 10192 75701
rect 12348 75692 12400 75744
rect 12440 75692 12492 75744
rect 13544 75837 13553 75871
rect 13553 75837 13587 75871
rect 13587 75837 13596 75871
rect 13544 75828 13596 75837
rect 13360 75735 13412 75744
rect 13360 75701 13369 75735
rect 13369 75701 13403 75735
rect 13403 75701 13412 75735
rect 15108 75735 15160 75744
rect 13360 75692 13412 75701
rect 15108 75701 15117 75735
rect 15117 75701 15151 75735
rect 15151 75701 15160 75735
rect 15108 75692 15160 75701
rect 21364 75735 21416 75744
rect 21364 75701 21373 75735
rect 21373 75701 21407 75735
rect 21407 75701 21416 75735
rect 21364 75692 21416 75701
rect 10982 75590 11034 75642
rect 11046 75590 11098 75642
rect 11110 75590 11162 75642
rect 11174 75590 11226 75642
rect 20982 75590 21034 75642
rect 21046 75590 21098 75642
rect 21110 75590 21162 75642
rect 21174 75590 21226 75642
rect 25044 75531 25096 75540
rect 25044 75497 25053 75531
rect 25053 75497 25087 75531
rect 25087 75497 25096 75531
rect 25044 75488 25096 75497
rect 10508 75352 10560 75404
rect 11336 75352 11388 75404
rect 10140 75284 10192 75336
rect 10784 75284 10836 75336
rect 23664 75327 23716 75336
rect 23664 75293 23673 75327
rect 23673 75293 23707 75327
rect 23707 75293 23716 75327
rect 23664 75284 23716 75293
rect 23940 75327 23992 75336
rect 23940 75293 23949 75327
rect 23949 75293 23983 75327
rect 23983 75293 23992 75327
rect 23940 75284 23992 75293
rect 11980 75191 12032 75200
rect 11980 75157 11989 75191
rect 11989 75157 12023 75191
rect 12023 75157 12032 75191
rect 11980 75148 12032 75157
rect 12440 75148 12492 75200
rect 5982 75046 6034 75098
rect 6046 75046 6098 75098
rect 6110 75046 6162 75098
rect 6174 75046 6226 75098
rect 15982 75046 16034 75098
rect 16046 75046 16098 75098
rect 16110 75046 16162 75098
rect 16174 75046 16226 75098
rect 25982 75046 26034 75098
rect 26046 75046 26098 75098
rect 26110 75046 26162 75098
rect 26174 75046 26226 75098
rect 10508 74987 10560 74996
rect 10508 74953 10517 74987
rect 10517 74953 10551 74987
rect 10551 74953 10560 74987
rect 10508 74944 10560 74953
rect 17960 74944 18012 74996
rect 23664 74944 23716 74996
rect 24768 74944 24820 74996
rect 4160 74740 4212 74792
rect 5448 74740 5500 74792
rect 12532 74740 12584 74792
rect 13728 74740 13780 74792
rect 13820 74740 13872 74792
rect 14740 74740 14792 74792
rect 15660 74740 15712 74792
rect 16488 74740 16540 74792
rect 19156 74740 19208 74792
rect 4620 74604 4672 74656
rect 5540 74604 5592 74656
rect 6460 74604 6512 74656
rect 6920 74604 6972 74656
rect 10784 74647 10836 74656
rect 10784 74613 10793 74647
rect 10793 74613 10827 74647
rect 10827 74613 10836 74647
rect 10784 74604 10836 74613
rect 20352 74604 20404 74656
rect 22100 74604 22152 74656
rect 22560 74604 22612 74656
rect 23940 74647 23992 74656
rect 23940 74613 23949 74647
rect 23949 74613 23983 74647
rect 23983 74613 23992 74647
rect 23940 74604 23992 74613
rect 27620 74604 27672 74656
rect 29000 74604 29052 74656
rect 10982 74502 11034 74554
rect 11046 74502 11098 74554
rect 11110 74502 11162 74554
rect 11174 74502 11226 74554
rect 20982 74502 21034 74554
rect 21046 74502 21098 74554
rect 21110 74502 21162 74554
rect 21174 74502 21226 74554
rect 19248 74400 19300 74452
rect 11980 74264 12032 74316
rect 12348 74196 12400 74248
rect 13084 74060 13136 74112
rect 5982 73958 6034 74010
rect 6046 73958 6098 74010
rect 6110 73958 6162 74010
rect 6174 73958 6226 74010
rect 15982 73958 16034 74010
rect 16046 73958 16098 74010
rect 16110 73958 16162 74010
rect 16174 73958 16226 74010
rect 25982 73958 26034 74010
rect 26046 73958 26098 74010
rect 26110 73958 26162 74010
rect 26174 73958 26226 74010
rect 11980 73856 12032 73908
rect 12440 73516 12492 73568
rect 10982 73414 11034 73466
rect 11046 73414 11098 73466
rect 11110 73414 11162 73466
rect 11174 73414 11226 73466
rect 20982 73414 21034 73466
rect 21046 73414 21098 73466
rect 21110 73414 21162 73466
rect 21174 73414 21226 73466
rect 14372 73287 14424 73296
rect 14372 73253 14381 73287
rect 14381 73253 14415 73287
rect 14415 73253 14424 73287
rect 14372 73244 14424 73253
rect 13084 73176 13136 73228
rect 12440 73108 12492 73160
rect 5982 72870 6034 72922
rect 6046 72870 6098 72922
rect 6110 72870 6162 72922
rect 6174 72870 6226 72922
rect 15982 72870 16034 72922
rect 16046 72870 16098 72922
rect 16110 72870 16162 72922
rect 16174 72870 16226 72922
rect 25982 72870 26034 72922
rect 26046 72870 26098 72922
rect 26110 72870 26162 72922
rect 26174 72870 26226 72922
rect 13084 72768 13136 72820
rect 12440 72428 12492 72480
rect 10982 72326 11034 72378
rect 11046 72326 11098 72378
rect 11110 72326 11162 72378
rect 11174 72326 11226 72378
rect 20982 72326 21034 72378
rect 21046 72326 21098 72378
rect 21110 72326 21162 72378
rect 21174 72326 21226 72378
rect 22560 72199 22612 72208
rect 22560 72165 22569 72199
rect 22569 72165 22603 72199
rect 22603 72165 22612 72199
rect 22560 72156 22612 72165
rect 20812 72088 20864 72140
rect 21364 72020 21416 72072
rect 5982 71782 6034 71834
rect 6046 71782 6098 71834
rect 6110 71782 6162 71834
rect 6174 71782 6226 71834
rect 15982 71782 16034 71834
rect 16046 71782 16098 71834
rect 16110 71782 16162 71834
rect 16174 71782 16226 71834
rect 25982 71782 26034 71834
rect 26046 71782 26098 71834
rect 26110 71782 26162 71834
rect 26174 71782 26226 71834
rect 20812 71340 20864 71392
rect 21364 71383 21416 71392
rect 21364 71349 21373 71383
rect 21373 71349 21407 71383
rect 21407 71349 21416 71383
rect 21364 71340 21416 71349
rect 10982 71238 11034 71290
rect 11046 71238 11098 71290
rect 11110 71238 11162 71290
rect 11174 71238 11226 71290
rect 20982 71238 21034 71290
rect 21046 71238 21098 71290
rect 21110 71238 21162 71290
rect 21174 71238 21226 71290
rect 7564 71068 7616 71120
rect 8024 71068 8076 71120
rect 23388 71068 23440 71120
rect 20996 71000 21048 71052
rect 21364 70932 21416 70984
rect 23112 70932 23164 70984
rect 23388 70932 23440 70984
rect 5982 70694 6034 70746
rect 6046 70694 6098 70746
rect 6110 70694 6162 70746
rect 6174 70694 6226 70746
rect 15982 70694 16034 70746
rect 16046 70694 16098 70746
rect 16110 70694 16162 70746
rect 16174 70694 16226 70746
rect 25982 70694 26034 70746
rect 26046 70694 26098 70746
rect 26110 70694 26162 70746
rect 26174 70694 26226 70746
rect 20904 70567 20956 70576
rect 20904 70533 20913 70567
rect 20913 70533 20947 70567
rect 20947 70533 20956 70567
rect 20904 70524 20956 70533
rect 26424 70499 26476 70508
rect 26424 70465 26433 70499
rect 26433 70465 26467 70499
rect 26467 70465 26476 70499
rect 26424 70456 26476 70465
rect 21364 70431 21416 70440
rect 21364 70397 21373 70431
rect 21373 70397 21407 70431
rect 21407 70397 21416 70431
rect 21364 70388 21416 70397
rect 21732 70388 21784 70440
rect 24860 70388 24912 70440
rect 26148 70431 26200 70440
rect 26148 70397 26157 70431
rect 26157 70397 26191 70431
rect 26191 70397 26200 70431
rect 26148 70388 26200 70397
rect 27712 70320 27764 70372
rect 27896 70320 27948 70372
rect 26424 70252 26476 70304
rect 10982 70150 11034 70202
rect 11046 70150 11098 70202
rect 11110 70150 11162 70202
rect 11174 70150 11226 70202
rect 20982 70150 21034 70202
rect 21046 70150 21098 70202
rect 21110 70150 21162 70202
rect 21174 70150 21226 70202
rect 2780 70091 2832 70100
rect 2780 70057 2789 70091
rect 2789 70057 2823 70091
rect 2823 70057 2832 70091
rect 2780 70048 2832 70057
rect 25872 70048 25924 70100
rect 26148 70091 26200 70100
rect 26148 70057 26157 70091
rect 26157 70057 26191 70091
rect 26191 70057 26200 70091
rect 26148 70048 26200 70057
rect 2044 69912 2096 69964
rect 1676 69887 1728 69896
rect 1676 69853 1685 69887
rect 1685 69853 1719 69887
rect 1719 69853 1728 69887
rect 1676 69844 1728 69853
rect 5982 69606 6034 69658
rect 6046 69606 6098 69658
rect 6110 69606 6162 69658
rect 6174 69606 6226 69658
rect 15982 69606 16034 69658
rect 16046 69606 16098 69658
rect 16110 69606 16162 69658
rect 16174 69606 16226 69658
rect 25982 69606 26034 69658
rect 26046 69606 26098 69658
rect 26110 69606 26162 69658
rect 26174 69606 26226 69658
rect 12348 69436 12400 69488
rect 1584 69368 1636 69420
rect 2044 69411 2096 69420
rect 2044 69377 2053 69411
rect 2053 69377 2087 69411
rect 2087 69377 2096 69411
rect 2044 69368 2096 69377
rect 26424 69411 26476 69420
rect 26424 69377 26433 69411
rect 26433 69377 26467 69411
rect 26467 69377 26476 69411
rect 26424 69368 26476 69377
rect 1676 69343 1728 69352
rect 1676 69309 1685 69343
rect 1685 69309 1719 69343
rect 1719 69309 1728 69343
rect 1676 69300 1728 69309
rect 11336 69300 11388 69352
rect 24860 69300 24912 69352
rect 25872 69300 25924 69352
rect 26240 69300 26292 69352
rect 27712 69207 27764 69216
rect 27712 69173 27721 69207
rect 27721 69173 27755 69207
rect 27755 69173 27764 69207
rect 27712 69164 27764 69173
rect 10982 69062 11034 69114
rect 11046 69062 11098 69114
rect 11110 69062 11162 69114
rect 11174 69062 11226 69114
rect 20982 69062 21034 69114
rect 21046 69062 21098 69114
rect 21110 69062 21162 69114
rect 21174 69062 21226 69114
rect 26240 69003 26292 69012
rect 26240 68969 26249 69003
rect 26249 68969 26283 69003
rect 26283 68969 26292 69003
rect 26240 68960 26292 68969
rect 5982 68518 6034 68570
rect 6046 68518 6098 68570
rect 6110 68518 6162 68570
rect 6174 68518 6226 68570
rect 15982 68518 16034 68570
rect 16046 68518 16098 68570
rect 16110 68518 16162 68570
rect 16174 68518 16226 68570
rect 25982 68518 26034 68570
rect 26046 68518 26098 68570
rect 26110 68518 26162 68570
rect 26174 68518 26226 68570
rect 9128 68459 9180 68468
rect 9128 68425 9137 68459
rect 9137 68425 9171 68459
rect 9171 68425 9180 68459
rect 9128 68416 9180 68425
rect 10692 68416 10744 68468
rect 11336 68416 11388 68468
rect 10982 67974 11034 68026
rect 11046 67974 11098 68026
rect 11110 67974 11162 68026
rect 11174 67974 11226 68026
rect 20982 67974 21034 68026
rect 21046 67974 21098 68026
rect 21110 67974 21162 68026
rect 21174 67974 21226 68026
rect 11244 67600 11296 67652
rect 11980 67600 12032 67652
rect 16396 67600 16448 67652
rect 16580 67600 16632 67652
rect 5982 67430 6034 67482
rect 6046 67430 6098 67482
rect 6110 67430 6162 67482
rect 6174 67430 6226 67482
rect 15982 67430 16034 67482
rect 16046 67430 16098 67482
rect 16110 67430 16162 67482
rect 16174 67430 16226 67482
rect 25982 67430 26034 67482
rect 26046 67430 26098 67482
rect 26110 67430 26162 67482
rect 26174 67430 26226 67482
rect 10692 67371 10744 67380
rect 10692 67337 10701 67371
rect 10701 67337 10735 67371
rect 10735 67337 10744 67371
rect 10692 67328 10744 67337
rect 11980 66988 12032 67040
rect 10982 66886 11034 66938
rect 11046 66886 11098 66938
rect 11110 66886 11162 66938
rect 11174 66886 11226 66938
rect 20982 66886 21034 66938
rect 21046 66886 21098 66938
rect 21110 66886 21162 66938
rect 21174 66886 21226 66938
rect 21732 66784 21784 66836
rect 17224 66691 17276 66700
rect 17224 66657 17233 66691
rect 17233 66657 17267 66691
rect 17267 66657 17276 66691
rect 17224 66648 17276 66657
rect 17868 66648 17920 66700
rect 21824 66691 21876 66700
rect 21824 66657 21833 66691
rect 21833 66657 21867 66691
rect 21867 66657 21876 66691
rect 21824 66648 21876 66657
rect 16948 66623 17000 66632
rect 16948 66589 16957 66623
rect 16957 66589 16991 66623
rect 16991 66589 17000 66623
rect 16948 66580 17000 66589
rect 17592 66555 17644 66564
rect 17592 66521 17601 66555
rect 17601 66521 17635 66555
rect 17635 66521 17644 66555
rect 17592 66512 17644 66521
rect 18052 66444 18104 66496
rect 18880 66444 18932 66496
rect 5982 66342 6034 66394
rect 6046 66342 6098 66394
rect 6110 66342 6162 66394
rect 6174 66342 6226 66394
rect 15982 66342 16034 66394
rect 16046 66342 16098 66394
rect 16110 66342 16162 66394
rect 16174 66342 16226 66394
rect 25982 66342 26034 66394
rect 26046 66342 26098 66394
rect 26110 66342 26162 66394
rect 26174 66342 26226 66394
rect 21824 66240 21876 66292
rect 27712 66240 27764 66292
rect 27988 66240 28040 66292
rect 18052 66147 18104 66156
rect 18052 66113 18061 66147
rect 18061 66113 18095 66147
rect 18095 66113 18104 66147
rect 18052 66104 18104 66113
rect 16948 65968 17000 66020
rect 17592 65968 17644 66020
rect 17776 66011 17828 66020
rect 17776 65977 17785 66011
rect 17785 65977 17819 66011
rect 17819 65977 17828 66011
rect 17776 65968 17828 65977
rect 20536 65968 20588 66020
rect 15476 65900 15528 65952
rect 17224 65943 17276 65952
rect 17224 65909 17233 65943
rect 17233 65909 17267 65943
rect 17267 65909 17276 65943
rect 17224 65900 17276 65909
rect 10982 65798 11034 65850
rect 11046 65798 11098 65850
rect 11110 65798 11162 65850
rect 11174 65798 11226 65850
rect 20982 65798 21034 65850
rect 21046 65798 21098 65850
rect 21110 65798 21162 65850
rect 21174 65798 21226 65850
rect 18604 65671 18656 65680
rect 18604 65637 18613 65671
rect 18613 65637 18647 65671
rect 18647 65637 18656 65671
rect 18604 65628 18656 65637
rect 14372 65560 14424 65612
rect 15660 65603 15712 65612
rect 15660 65569 15669 65603
rect 15669 65569 15703 65603
rect 15703 65569 15712 65603
rect 15660 65560 15712 65569
rect 15844 65560 15896 65612
rect 17868 65603 17920 65612
rect 17868 65569 17877 65603
rect 17877 65569 17911 65603
rect 17911 65569 17920 65603
rect 17868 65560 17920 65569
rect 17960 65560 18012 65612
rect 18236 65560 18288 65612
rect 17592 65535 17644 65544
rect 17592 65501 17601 65535
rect 17601 65501 17635 65535
rect 17635 65501 17644 65535
rect 17592 65492 17644 65501
rect 24952 65492 25004 65544
rect 25780 65492 25832 65544
rect 15200 65424 15252 65476
rect 5982 65254 6034 65306
rect 6046 65254 6098 65306
rect 6110 65254 6162 65306
rect 6174 65254 6226 65306
rect 15982 65254 16034 65306
rect 16046 65254 16098 65306
rect 16110 65254 16162 65306
rect 16174 65254 16226 65306
rect 25982 65254 26034 65306
rect 26046 65254 26098 65306
rect 26110 65254 26162 65306
rect 26174 65254 26226 65306
rect 14372 65016 14424 65068
rect 17868 65152 17920 65204
rect 21824 65152 21876 65204
rect 24768 65152 24820 65204
rect 15384 65084 15436 65136
rect 17224 65016 17276 65068
rect 15844 64948 15896 65000
rect 15660 64880 15712 64932
rect 17592 64923 17644 64932
rect 17592 64889 17601 64923
rect 17601 64889 17635 64923
rect 17635 64889 17644 64923
rect 17592 64880 17644 64889
rect 18236 64923 18288 64932
rect 18236 64889 18245 64923
rect 18245 64889 18279 64923
rect 18279 64889 18288 64923
rect 18236 64880 18288 64889
rect 22468 64880 22520 64932
rect 10982 64710 11034 64762
rect 11046 64710 11098 64762
rect 11110 64710 11162 64762
rect 11174 64710 11226 64762
rect 20982 64710 21034 64762
rect 21046 64710 21098 64762
rect 21110 64710 21162 64762
rect 21174 64710 21226 64762
rect 20720 64472 20772 64524
rect 21548 64472 21600 64524
rect 21640 64404 21692 64456
rect 15844 64336 15896 64388
rect 15660 64268 15712 64320
rect 23480 64268 23532 64320
rect 5982 64166 6034 64218
rect 6046 64166 6098 64218
rect 6110 64166 6162 64218
rect 6174 64166 6226 64218
rect 15982 64166 16034 64218
rect 16046 64166 16098 64218
rect 16110 64166 16162 64218
rect 16174 64166 16226 64218
rect 25982 64166 26034 64218
rect 26046 64166 26098 64218
rect 26110 64166 26162 64218
rect 26174 64166 26226 64218
rect 21548 64107 21600 64116
rect 21548 64073 21557 64107
rect 21557 64073 21591 64107
rect 21591 64073 21600 64107
rect 21548 64064 21600 64073
rect 21640 64064 21692 64116
rect 15660 63928 15712 63980
rect 17040 63971 17092 63980
rect 16212 63860 16264 63912
rect 17040 63937 17049 63971
rect 17049 63937 17083 63971
rect 17083 63937 17092 63971
rect 17040 63928 17092 63937
rect 18604 63971 18656 63980
rect 18604 63937 18613 63971
rect 18613 63937 18647 63971
rect 18647 63937 18656 63971
rect 18604 63928 18656 63937
rect 18880 63860 18932 63912
rect 20444 63835 20496 63844
rect 20444 63801 20453 63835
rect 20453 63801 20487 63835
rect 20487 63801 20496 63835
rect 20444 63792 20496 63801
rect 15752 63724 15804 63776
rect 10982 63622 11034 63674
rect 11046 63622 11098 63674
rect 11110 63622 11162 63674
rect 11174 63622 11226 63674
rect 20982 63622 21034 63674
rect 21046 63622 21098 63674
rect 21110 63622 21162 63674
rect 21174 63622 21226 63674
rect 18880 63563 18932 63572
rect 18880 63529 18889 63563
rect 18889 63529 18923 63563
rect 18923 63529 18932 63563
rect 18880 63520 18932 63529
rect 23664 63495 23716 63504
rect 23664 63461 23673 63495
rect 23673 63461 23707 63495
rect 23707 63461 23716 63495
rect 23664 63452 23716 63461
rect 15660 63427 15712 63436
rect 15660 63393 15669 63427
rect 15669 63393 15703 63427
rect 15703 63393 15712 63427
rect 15660 63384 15712 63393
rect 15752 63384 15804 63436
rect 24216 63384 24268 63436
rect 24400 63427 24452 63436
rect 24400 63393 24409 63427
rect 24409 63393 24443 63427
rect 24443 63393 24452 63427
rect 24400 63384 24452 63393
rect 15568 63316 15620 63368
rect 24032 63316 24084 63368
rect 15108 63248 15160 63300
rect 5982 63078 6034 63130
rect 6046 63078 6098 63130
rect 6110 63078 6162 63130
rect 6174 63078 6226 63130
rect 15982 63078 16034 63130
rect 16046 63078 16098 63130
rect 16110 63078 16162 63130
rect 16174 63078 16226 63130
rect 25982 63078 26034 63130
rect 26046 63078 26098 63130
rect 26110 63078 26162 63130
rect 26174 63078 26226 63130
rect 23480 63019 23532 63028
rect 23480 62985 23489 63019
rect 23489 62985 23523 63019
rect 23523 62985 23532 63019
rect 23480 62976 23532 62985
rect 24400 62976 24452 63028
rect 25872 62840 25924 62892
rect 27620 62840 27672 62892
rect 27804 62840 27856 62892
rect 14096 62772 14148 62824
rect 15660 62815 15712 62824
rect 15660 62781 15669 62815
rect 15669 62781 15703 62815
rect 15703 62781 15712 62815
rect 15660 62772 15712 62781
rect 24216 62772 24268 62824
rect 24860 62772 24912 62824
rect 26148 62815 26200 62824
rect 26148 62781 26157 62815
rect 26157 62781 26191 62815
rect 26191 62781 26200 62815
rect 26148 62772 26200 62781
rect 13360 62704 13412 62756
rect 15752 62704 15804 62756
rect 27804 62747 27856 62756
rect 27804 62713 27813 62747
rect 27813 62713 27847 62747
rect 27847 62713 27856 62747
rect 27804 62704 27856 62713
rect 15568 62636 15620 62688
rect 24032 62636 24084 62688
rect 10982 62534 11034 62586
rect 11046 62534 11098 62586
rect 11110 62534 11162 62586
rect 11174 62534 11226 62586
rect 20982 62534 21034 62586
rect 21046 62534 21098 62586
rect 21110 62534 21162 62586
rect 21174 62534 21226 62586
rect 15476 62432 15528 62484
rect 15660 62432 15712 62484
rect 25872 62432 25924 62484
rect 26148 62475 26200 62484
rect 26148 62441 26157 62475
rect 26157 62441 26191 62475
rect 26191 62441 26200 62475
rect 26148 62432 26200 62441
rect 15844 62364 15896 62416
rect 13728 62296 13780 62348
rect 15476 62296 15528 62348
rect 16304 62296 16356 62348
rect 16672 62228 16724 62280
rect 16580 62160 16632 62212
rect 17868 62160 17920 62212
rect 19248 62092 19300 62144
rect 5982 61990 6034 62042
rect 6046 61990 6098 62042
rect 6110 61990 6162 62042
rect 6174 61990 6226 62042
rect 15982 61990 16034 62042
rect 16046 61990 16098 62042
rect 16110 61990 16162 62042
rect 16174 61990 16226 62042
rect 25982 61990 26034 62042
rect 26046 61990 26098 62042
rect 26110 61990 26162 62042
rect 26174 61990 26226 62042
rect 13820 61931 13872 61940
rect 13820 61897 13829 61931
rect 13829 61897 13863 61931
rect 13863 61897 13872 61931
rect 13820 61888 13872 61897
rect 12440 61795 12492 61804
rect 12440 61761 12449 61795
rect 12449 61761 12483 61795
rect 12483 61761 12492 61795
rect 20076 61795 20128 61804
rect 12440 61752 12492 61761
rect 20076 61761 20085 61795
rect 20085 61761 20119 61795
rect 20119 61761 20128 61795
rect 20076 61752 20128 61761
rect 25780 61752 25832 61804
rect 12164 61727 12216 61736
rect 12164 61693 12173 61727
rect 12173 61693 12207 61727
rect 12207 61693 12216 61727
rect 12164 61684 12216 61693
rect 15844 61548 15896 61600
rect 16580 61616 16632 61668
rect 19248 61684 19300 61736
rect 19432 61684 19484 61736
rect 19800 61727 19852 61736
rect 19800 61693 19809 61727
rect 19809 61693 19843 61727
rect 19843 61693 19852 61727
rect 19800 61684 19852 61693
rect 25872 61684 25924 61736
rect 28080 61616 28132 61668
rect 16304 61591 16356 61600
rect 16304 61557 16313 61591
rect 16313 61557 16347 61591
rect 16347 61557 16356 61591
rect 16304 61548 16356 61557
rect 16672 61591 16724 61600
rect 16672 61557 16681 61591
rect 16681 61557 16715 61591
rect 16715 61557 16724 61591
rect 16672 61548 16724 61557
rect 17684 61548 17736 61600
rect 18052 61548 18104 61600
rect 18788 61591 18840 61600
rect 18788 61557 18797 61591
rect 18797 61557 18831 61591
rect 18831 61557 18840 61591
rect 18788 61548 18840 61557
rect 10982 61446 11034 61498
rect 11046 61446 11098 61498
rect 11110 61446 11162 61498
rect 11174 61446 11226 61498
rect 20982 61446 21034 61498
rect 21046 61446 21098 61498
rect 21110 61446 21162 61498
rect 21174 61446 21226 61498
rect 1584 61387 1636 61396
rect 1584 61353 1593 61387
rect 1593 61353 1627 61387
rect 1627 61353 1636 61387
rect 1584 61344 1636 61353
rect 12440 61387 12492 61396
rect 12440 61353 12449 61387
rect 12449 61353 12483 61387
rect 12483 61353 12492 61387
rect 20720 61387 20772 61396
rect 12440 61344 12492 61353
rect 20720 61353 20729 61387
rect 20729 61353 20763 61387
rect 20763 61353 20772 61387
rect 20720 61344 20772 61353
rect 25872 61344 25924 61396
rect 17868 61276 17920 61328
rect 21456 61319 21508 61328
rect 21456 61285 21465 61319
rect 21465 61285 21499 61319
rect 21499 61285 21508 61319
rect 21456 61276 21508 61285
rect 26700 61319 26752 61328
rect 26700 61285 26709 61319
rect 26709 61285 26743 61319
rect 26743 61285 26752 61319
rect 26700 61276 26752 61285
rect 18052 61251 18104 61260
rect 17500 61140 17552 61192
rect 18052 61217 18061 61251
rect 18061 61217 18095 61251
rect 18095 61217 18104 61251
rect 18052 61208 18104 61217
rect 19156 61251 19208 61260
rect 19156 61217 19165 61251
rect 19165 61217 19199 61251
rect 19199 61217 19208 61251
rect 19156 61208 19208 61217
rect 22008 61208 22060 61260
rect 27344 61208 27396 61260
rect 27804 61208 27856 61260
rect 21364 61183 21416 61192
rect 17960 61072 18012 61124
rect 21364 61149 21373 61183
rect 21373 61149 21407 61183
rect 21407 61149 21416 61183
rect 21364 61140 21416 61149
rect 22836 61140 22888 61192
rect 26516 61140 26568 61192
rect 26884 61140 26936 61192
rect 19248 61072 19300 61124
rect 21272 61072 21324 61124
rect 16580 61004 16632 61056
rect 18604 61047 18656 61056
rect 18604 61013 18613 61047
rect 18613 61013 18647 61047
rect 18647 61013 18656 61047
rect 18604 61004 18656 61013
rect 19616 61004 19668 61056
rect 20812 61004 20864 61056
rect 21456 61004 21508 61056
rect 5982 60902 6034 60954
rect 6046 60902 6098 60954
rect 6110 60902 6162 60954
rect 6174 60902 6226 60954
rect 15982 60902 16034 60954
rect 16046 60902 16098 60954
rect 16110 60902 16162 60954
rect 16174 60902 16226 60954
rect 25982 60902 26034 60954
rect 26046 60902 26098 60954
rect 26110 60902 26162 60954
rect 26174 60902 26226 60954
rect 2780 60843 2832 60852
rect 2780 60809 2789 60843
rect 2789 60809 2823 60843
rect 2823 60809 2832 60843
rect 2780 60800 2832 60809
rect 19064 60800 19116 60852
rect 19248 60800 19300 60852
rect 22008 60843 22060 60852
rect 22008 60809 22017 60843
rect 22017 60809 22051 60843
rect 22051 60809 22060 60843
rect 22008 60800 22060 60809
rect 22836 60800 22888 60852
rect 25504 60800 25556 60852
rect 26884 60843 26936 60852
rect 26884 60809 26893 60843
rect 26893 60809 26927 60843
rect 26927 60809 26936 60843
rect 26884 60800 26936 60809
rect 27344 60843 27396 60852
rect 27344 60809 27353 60843
rect 27353 60809 27387 60843
rect 27387 60809 27396 60843
rect 27344 60800 27396 60809
rect 18880 60775 18932 60784
rect 18880 60741 18889 60775
rect 18889 60741 18923 60775
rect 18923 60741 18932 60775
rect 18880 60732 18932 60741
rect 19156 60732 19208 60784
rect 1584 60664 1636 60716
rect 15660 60664 15712 60716
rect 1676 60639 1728 60648
rect 1676 60605 1685 60639
rect 1685 60605 1719 60639
rect 1719 60605 1728 60639
rect 1676 60596 1728 60605
rect 17040 60664 17092 60716
rect 17500 60707 17552 60716
rect 17500 60673 17509 60707
rect 17509 60673 17543 60707
rect 17543 60673 17552 60707
rect 17500 60664 17552 60673
rect 20628 60707 20680 60716
rect 20628 60673 20637 60707
rect 20637 60673 20671 60707
rect 20671 60673 20680 60707
rect 20628 60664 20680 60673
rect 21272 60664 21324 60716
rect 21364 60664 21416 60716
rect 26516 60707 26568 60716
rect 26516 60673 26525 60707
rect 26525 60673 26559 60707
rect 26559 60673 26568 60707
rect 26516 60664 26568 60673
rect 16580 60596 16632 60648
rect 18236 60639 18288 60648
rect 16212 60528 16264 60580
rect 18236 60605 18245 60639
rect 18245 60605 18279 60639
rect 18279 60605 18288 60639
rect 18236 60596 18288 60605
rect 18604 60639 18656 60648
rect 18604 60605 18613 60639
rect 18613 60605 18647 60639
rect 18647 60605 18656 60639
rect 18604 60596 18656 60605
rect 18880 60639 18932 60648
rect 18880 60605 18889 60639
rect 18889 60605 18923 60639
rect 18923 60605 18932 60639
rect 18880 60596 18932 60605
rect 20720 60596 20772 60648
rect 21548 60596 21600 60648
rect 19340 60528 19392 60580
rect 10982 60358 11034 60410
rect 11046 60358 11098 60410
rect 11110 60358 11162 60410
rect 11174 60358 11226 60410
rect 20982 60358 21034 60410
rect 21046 60358 21098 60410
rect 21110 60358 21162 60410
rect 21174 60358 21226 60410
rect 15660 60256 15712 60308
rect 16212 60299 16264 60308
rect 16212 60265 16221 60299
rect 16221 60265 16255 60299
rect 16255 60265 16264 60299
rect 16212 60256 16264 60265
rect 17684 60256 17736 60308
rect 18880 60256 18932 60308
rect 19432 60256 19484 60308
rect 16856 60231 16908 60240
rect 16856 60197 16865 60231
rect 16865 60197 16899 60231
rect 16899 60197 16908 60231
rect 16856 60188 16908 60197
rect 17040 60120 17092 60172
rect 17224 60120 17276 60172
rect 19524 60120 19576 60172
rect 19800 60120 19852 60172
rect 20628 60163 20680 60172
rect 20628 60129 20637 60163
rect 20637 60129 20671 60163
rect 20671 60129 20680 60163
rect 20628 60120 20680 60129
rect 21548 60120 21600 60172
rect 22744 60120 22796 60172
rect 22928 60163 22980 60172
rect 22928 60129 22937 60163
rect 22937 60129 22971 60163
rect 22971 60129 22980 60163
rect 22928 60120 22980 60129
rect 17684 59984 17736 60036
rect 1676 59959 1728 59968
rect 1676 59925 1685 59959
rect 1685 59925 1719 59959
rect 1719 59925 1728 59959
rect 1676 59916 1728 59925
rect 2044 59916 2096 59968
rect 17316 59916 17368 59968
rect 18236 60052 18288 60104
rect 18788 60052 18840 60104
rect 21824 60095 21876 60104
rect 19708 60027 19760 60036
rect 19708 59993 19717 60027
rect 19717 59993 19751 60027
rect 19751 59993 19760 60027
rect 19708 59984 19760 59993
rect 21824 60061 21833 60095
rect 21833 60061 21867 60095
rect 21867 60061 21876 60095
rect 21824 60052 21876 60061
rect 22836 60095 22888 60104
rect 22836 60061 22845 60095
rect 22845 60061 22879 60095
rect 22879 60061 22888 60095
rect 22836 60052 22888 60061
rect 22192 59984 22244 60036
rect 5982 59814 6034 59866
rect 6046 59814 6098 59866
rect 6110 59814 6162 59866
rect 6174 59814 6226 59866
rect 15982 59814 16034 59866
rect 16046 59814 16098 59866
rect 16110 59814 16162 59866
rect 16174 59814 16226 59866
rect 25982 59814 26034 59866
rect 26046 59814 26098 59866
rect 26110 59814 26162 59866
rect 26174 59814 26226 59866
rect 17500 59712 17552 59764
rect 19064 59712 19116 59764
rect 17684 59644 17736 59696
rect 18880 59576 18932 59628
rect 22836 59644 22888 59696
rect 16212 59508 16264 59560
rect 15752 59483 15804 59492
rect 15752 59449 15761 59483
rect 15761 59449 15795 59483
rect 15795 59449 15804 59483
rect 15752 59440 15804 59449
rect 14556 59372 14608 59424
rect 15568 59415 15620 59424
rect 15568 59381 15577 59415
rect 15577 59381 15611 59415
rect 15611 59381 15620 59415
rect 17316 59508 17368 59560
rect 18788 59551 18840 59560
rect 18788 59517 18797 59551
rect 18797 59517 18831 59551
rect 18831 59517 18840 59551
rect 18788 59508 18840 59517
rect 19064 59551 19116 59560
rect 19064 59517 19073 59551
rect 19073 59517 19107 59551
rect 19107 59517 19116 59551
rect 19064 59508 19116 59517
rect 21916 59576 21968 59628
rect 21272 59551 21324 59560
rect 21272 59517 21281 59551
rect 21281 59517 21315 59551
rect 21315 59517 21324 59551
rect 21272 59508 21324 59517
rect 21364 59508 21416 59560
rect 21640 59508 21692 59560
rect 19800 59483 19852 59492
rect 19800 59449 19809 59483
rect 19809 59449 19843 59483
rect 19843 59449 19852 59483
rect 19800 59440 19852 59449
rect 17040 59415 17092 59424
rect 15568 59372 15620 59381
rect 17040 59381 17049 59415
rect 17049 59381 17083 59415
rect 17083 59381 17092 59415
rect 17040 59372 17092 59381
rect 22192 59415 22244 59424
rect 22192 59381 22201 59415
rect 22201 59381 22235 59415
rect 22235 59381 22244 59415
rect 22192 59372 22244 59381
rect 22744 59372 22796 59424
rect 10982 59270 11034 59322
rect 11046 59270 11098 59322
rect 11110 59270 11162 59322
rect 11174 59270 11226 59322
rect 20982 59270 21034 59322
rect 21046 59270 21098 59322
rect 21110 59270 21162 59322
rect 21174 59270 21226 59322
rect 19340 59168 19392 59220
rect 17592 59143 17644 59152
rect 14740 59032 14792 59084
rect 15660 59032 15712 59084
rect 17592 59109 17601 59143
rect 17601 59109 17635 59143
rect 17635 59109 17644 59143
rect 17592 59100 17644 59109
rect 16856 59032 16908 59084
rect 17684 59032 17736 59084
rect 21364 59100 21416 59152
rect 19616 59075 19668 59084
rect 19616 59041 19625 59075
rect 19625 59041 19659 59075
rect 19659 59041 19668 59075
rect 19616 59032 19668 59041
rect 21824 59032 21876 59084
rect 22836 59032 22888 59084
rect 23480 59075 23532 59084
rect 23480 59041 23489 59075
rect 23489 59041 23523 59075
rect 23523 59041 23532 59075
rect 23480 59032 23532 59041
rect 15568 58964 15620 59016
rect 17960 58964 18012 59016
rect 18144 58964 18196 59016
rect 16672 58939 16724 58948
rect 16672 58905 16681 58939
rect 16681 58905 16715 58939
rect 16715 58905 16724 58939
rect 16672 58896 16724 58905
rect 17316 58939 17368 58948
rect 17316 58905 17325 58939
rect 17325 58905 17359 58939
rect 17359 58905 17368 58939
rect 18972 58964 19024 59016
rect 22100 58964 22152 59016
rect 23296 59007 23348 59016
rect 23296 58973 23305 59007
rect 23305 58973 23339 59007
rect 23339 58973 23348 59007
rect 23296 58964 23348 58973
rect 17316 58896 17368 58905
rect 19156 58896 19208 58948
rect 20996 58896 21048 58948
rect 14648 58871 14700 58880
rect 14648 58837 14657 58871
rect 14657 58837 14691 58871
rect 14691 58837 14700 58871
rect 14648 58828 14700 58837
rect 18788 58828 18840 58880
rect 19524 58871 19576 58880
rect 19524 58837 19533 58871
rect 19533 58837 19567 58871
rect 19567 58837 19576 58871
rect 19524 58828 19576 58837
rect 24308 58871 24360 58880
rect 24308 58837 24317 58871
rect 24317 58837 24351 58871
rect 24351 58837 24360 58871
rect 24308 58828 24360 58837
rect 5982 58726 6034 58778
rect 6046 58726 6098 58778
rect 6110 58726 6162 58778
rect 6174 58726 6226 58778
rect 15982 58726 16034 58778
rect 16046 58726 16098 58778
rect 16110 58726 16162 58778
rect 16174 58726 16226 58778
rect 25982 58726 26034 58778
rect 26046 58726 26098 58778
rect 26110 58726 26162 58778
rect 26174 58726 26226 58778
rect 2872 58624 2924 58676
rect 14464 58667 14516 58676
rect 14464 58633 14473 58667
rect 14473 58633 14507 58667
rect 14507 58633 14516 58667
rect 14464 58624 14516 58633
rect 15568 58624 15620 58676
rect 19064 58624 19116 58676
rect 21824 58667 21876 58676
rect 16488 58488 16540 58540
rect 18880 58488 18932 58540
rect 18972 58488 19024 58540
rect 21824 58633 21833 58667
rect 21833 58633 21867 58667
rect 21867 58633 21876 58667
rect 21824 58624 21876 58633
rect 22836 58624 22888 58676
rect 23296 58624 23348 58676
rect 23756 58624 23808 58676
rect 23664 58531 23716 58540
rect 3148 58463 3200 58472
rect 3148 58429 3157 58463
rect 3157 58429 3191 58463
rect 3191 58429 3200 58463
rect 3148 58420 3200 58429
rect 5448 58352 5500 58404
rect 14740 58352 14792 58404
rect 15660 58463 15712 58472
rect 14832 58327 14884 58336
rect 14832 58293 14841 58327
rect 14841 58293 14875 58327
rect 14875 58293 14884 58327
rect 14832 58284 14884 58293
rect 15660 58429 15669 58463
rect 15669 58429 15703 58463
rect 15703 58429 15712 58463
rect 15660 58420 15712 58429
rect 16212 58463 16264 58472
rect 16212 58429 16221 58463
rect 16221 58429 16255 58463
rect 16255 58429 16264 58463
rect 16212 58420 16264 58429
rect 19616 58463 19668 58472
rect 16488 58352 16540 58404
rect 17132 58352 17184 58404
rect 15568 58284 15620 58336
rect 17224 58327 17276 58336
rect 17224 58293 17233 58327
rect 17233 58293 17267 58327
rect 17267 58293 17276 58327
rect 17224 58284 17276 58293
rect 17684 58352 17736 58404
rect 19616 58429 19625 58463
rect 19625 58429 19659 58463
rect 19659 58429 19668 58463
rect 19616 58420 19668 58429
rect 20076 58420 20128 58472
rect 20996 58463 21048 58472
rect 19524 58352 19576 58404
rect 19708 58352 19760 58404
rect 20996 58429 21005 58463
rect 21005 58429 21039 58463
rect 21039 58429 21048 58463
rect 20996 58420 21048 58429
rect 23664 58497 23673 58531
rect 23673 58497 23707 58531
rect 23707 58497 23716 58531
rect 23664 58488 23716 58497
rect 24584 58488 24636 58540
rect 22560 58420 22612 58472
rect 23296 58420 23348 58472
rect 24308 58420 24360 58472
rect 21824 58284 21876 58336
rect 23572 58284 23624 58336
rect 10982 58182 11034 58234
rect 11046 58182 11098 58234
rect 11110 58182 11162 58234
rect 11174 58182 11226 58234
rect 20982 58182 21034 58234
rect 21046 58182 21098 58234
rect 21110 58182 21162 58234
rect 21174 58182 21226 58234
rect 11704 58080 11756 58132
rect 11980 58123 12032 58132
rect 11980 58089 11989 58123
rect 11989 58089 12023 58123
rect 12023 58089 12032 58123
rect 11980 58080 12032 58089
rect 14372 58123 14424 58132
rect 14372 58089 14381 58123
rect 14381 58089 14415 58123
rect 14415 58089 14424 58123
rect 14372 58080 14424 58089
rect 15752 58080 15804 58132
rect 15660 58012 15712 58064
rect 12072 57944 12124 57996
rect 3148 57876 3200 57928
rect 3332 57876 3384 57928
rect 13452 57876 13504 57928
rect 15108 57944 15160 57996
rect 20720 58080 20772 58132
rect 23112 58080 23164 58132
rect 23480 58080 23532 58132
rect 17040 58012 17092 58064
rect 17592 58012 17644 58064
rect 20628 58012 20680 58064
rect 20996 58012 21048 58064
rect 16856 57944 16908 57996
rect 14372 57876 14424 57928
rect 15384 57919 15436 57928
rect 15384 57885 15393 57919
rect 15393 57885 15427 57919
rect 15427 57885 15436 57919
rect 15384 57876 15436 57885
rect 18144 57944 18196 57996
rect 19340 57987 19392 57996
rect 19340 57953 19349 57987
rect 19349 57953 19383 57987
rect 19383 57953 19392 57987
rect 19708 57987 19760 57996
rect 19340 57944 19392 57953
rect 19708 57953 19717 57987
rect 19717 57953 19751 57987
rect 19751 57953 19760 57987
rect 19708 57944 19760 57953
rect 23756 57987 23808 57996
rect 23756 57953 23765 57987
rect 23765 57953 23799 57987
rect 23799 57953 23808 57987
rect 23756 57944 23808 57953
rect 23940 57987 23992 57996
rect 23940 57953 23949 57987
rect 23949 57953 23983 57987
rect 23983 57953 23992 57987
rect 23940 57944 23992 57953
rect 24584 57944 24636 57996
rect 17592 57919 17644 57928
rect 17592 57885 17601 57919
rect 17601 57885 17635 57919
rect 17635 57885 17644 57919
rect 17776 57919 17828 57928
rect 17592 57876 17644 57885
rect 17776 57885 17785 57919
rect 17785 57885 17819 57919
rect 17819 57885 17828 57919
rect 17776 57876 17828 57885
rect 18512 57876 18564 57928
rect 20720 57876 20772 57928
rect 21364 57876 21416 57928
rect 3608 57808 3660 57860
rect 13728 57808 13780 57860
rect 15752 57808 15804 57860
rect 13544 57783 13596 57792
rect 13544 57749 13553 57783
rect 13553 57749 13587 57783
rect 13587 57749 13596 57783
rect 13544 57740 13596 57749
rect 14740 57783 14792 57792
rect 14740 57749 14749 57783
rect 14749 57749 14783 57783
rect 14783 57749 14792 57783
rect 14740 57740 14792 57749
rect 15384 57740 15436 57792
rect 19616 57808 19668 57860
rect 20260 57808 20312 57860
rect 22100 57876 22152 57928
rect 22376 57808 22428 57860
rect 24400 57851 24452 57860
rect 24400 57817 24409 57851
rect 24409 57817 24443 57851
rect 24443 57817 24452 57851
rect 24400 57808 24452 57817
rect 17040 57783 17092 57792
rect 17040 57749 17049 57783
rect 17049 57749 17083 57783
rect 17083 57749 17092 57783
rect 17040 57740 17092 57749
rect 17132 57740 17184 57792
rect 17592 57740 17644 57792
rect 18328 57783 18380 57792
rect 18328 57749 18337 57783
rect 18337 57749 18371 57783
rect 18371 57749 18380 57783
rect 18328 57740 18380 57749
rect 18604 57783 18656 57792
rect 18604 57749 18613 57783
rect 18613 57749 18647 57783
rect 18647 57749 18656 57783
rect 18604 57740 18656 57749
rect 20076 57740 20128 57792
rect 22560 57783 22612 57792
rect 22560 57749 22569 57783
rect 22569 57749 22603 57783
rect 22603 57749 22612 57783
rect 22560 57740 22612 57749
rect 23020 57783 23072 57792
rect 23020 57749 23029 57783
rect 23029 57749 23063 57783
rect 23063 57749 23072 57783
rect 23020 57740 23072 57749
rect 5982 57638 6034 57690
rect 6046 57638 6098 57690
rect 6110 57638 6162 57690
rect 6174 57638 6226 57690
rect 15982 57638 16034 57690
rect 16046 57638 16098 57690
rect 16110 57638 16162 57690
rect 16174 57638 16226 57690
rect 25982 57638 26034 57690
rect 26046 57638 26098 57690
rect 26110 57638 26162 57690
rect 26174 57638 26226 57690
rect 5540 57536 5592 57588
rect 13452 57579 13504 57588
rect 2688 57443 2740 57452
rect 2688 57409 2697 57443
rect 2697 57409 2731 57443
rect 2731 57409 2740 57443
rect 2688 57400 2740 57409
rect 2964 57400 3016 57452
rect 13452 57545 13461 57579
rect 13461 57545 13495 57579
rect 13495 57545 13504 57579
rect 13452 57536 13504 57545
rect 17684 57536 17736 57588
rect 18696 57579 18748 57588
rect 18696 57545 18705 57579
rect 18705 57545 18739 57579
rect 18739 57545 18748 57579
rect 18696 57536 18748 57545
rect 19524 57579 19576 57588
rect 19524 57545 19533 57579
rect 19533 57545 19567 57579
rect 19567 57545 19576 57579
rect 19524 57536 19576 57545
rect 20444 57536 20496 57588
rect 20812 57536 20864 57588
rect 22100 57536 22152 57588
rect 22376 57536 22428 57588
rect 23664 57536 23716 57588
rect 23756 57536 23808 57588
rect 18328 57511 18380 57520
rect 18328 57477 18337 57511
rect 18337 57477 18371 57511
rect 18371 57477 18380 57511
rect 18328 57468 18380 57477
rect 13452 57400 13504 57452
rect 14648 57443 14700 57452
rect 14648 57409 14657 57443
rect 14657 57409 14691 57443
rect 14691 57409 14700 57443
rect 14648 57400 14700 57409
rect 17040 57400 17092 57452
rect 18604 57400 18656 57452
rect 3608 57375 3660 57384
rect 3608 57341 3617 57375
rect 3617 57341 3651 57375
rect 3651 57341 3660 57375
rect 7012 57375 7064 57384
rect 3608 57332 3660 57341
rect 7012 57341 7021 57375
rect 7021 57341 7055 57375
rect 7055 57341 7064 57375
rect 7012 57332 7064 57341
rect 13544 57375 13596 57384
rect 13544 57341 13553 57375
rect 13553 57341 13587 57375
rect 13587 57341 13596 57375
rect 13544 57332 13596 57341
rect 9680 57264 9732 57316
rect 14740 57332 14792 57384
rect 15752 57332 15804 57384
rect 16948 57375 17000 57384
rect 16948 57341 16957 57375
rect 16957 57341 16991 57375
rect 16991 57341 17000 57375
rect 16948 57332 17000 57341
rect 15660 57307 15712 57316
rect 15660 57273 15669 57307
rect 15669 57273 15703 57307
rect 15703 57273 15712 57307
rect 15660 57264 15712 57273
rect 17040 57264 17092 57316
rect 2136 57239 2188 57248
rect 2136 57205 2145 57239
rect 2145 57205 2179 57239
rect 2179 57205 2188 57239
rect 2136 57196 2188 57205
rect 12072 57239 12124 57248
rect 12072 57205 12081 57239
rect 12081 57205 12115 57239
rect 12115 57205 12124 57239
rect 12072 57196 12124 57205
rect 14004 57196 14056 57248
rect 14372 57239 14424 57248
rect 14372 57205 14381 57239
rect 14381 57205 14415 57239
rect 14415 57205 14424 57239
rect 14372 57196 14424 57205
rect 16212 57239 16264 57248
rect 16212 57205 16221 57239
rect 16221 57205 16255 57239
rect 16255 57205 16264 57239
rect 16212 57196 16264 57205
rect 16856 57239 16908 57248
rect 16856 57205 16865 57239
rect 16865 57205 16899 57239
rect 16899 57205 16908 57239
rect 16856 57196 16908 57205
rect 17132 57196 17184 57248
rect 17592 57196 17644 57248
rect 19524 57332 19576 57384
rect 20076 57332 20128 57384
rect 20352 57332 20404 57384
rect 21640 57468 21692 57520
rect 23940 57511 23992 57520
rect 23940 57477 23949 57511
rect 23949 57477 23983 57511
rect 23983 57477 23992 57511
rect 23940 57468 23992 57477
rect 18052 57307 18104 57316
rect 18052 57273 18061 57307
rect 18061 57273 18095 57307
rect 18095 57273 18104 57307
rect 18052 57264 18104 57273
rect 20720 57332 20772 57384
rect 22376 57375 22428 57384
rect 22376 57341 22385 57375
rect 22385 57341 22419 57375
rect 22419 57341 22428 57375
rect 22376 57332 22428 57341
rect 21824 57264 21876 57316
rect 19064 57239 19116 57248
rect 19064 57205 19073 57239
rect 19073 57205 19107 57239
rect 19107 57205 19116 57239
rect 19064 57196 19116 57205
rect 20628 57196 20680 57248
rect 10982 57094 11034 57146
rect 11046 57094 11098 57146
rect 11110 57094 11162 57146
rect 11174 57094 11226 57146
rect 20982 57094 21034 57146
rect 21046 57094 21098 57146
rect 21110 57094 21162 57146
rect 21174 57094 21226 57146
rect 2136 56992 2188 57044
rect 7012 57035 7064 57044
rect 7012 57001 7021 57035
rect 7021 57001 7055 57035
rect 7055 57001 7064 57035
rect 7012 56992 7064 57001
rect 13452 56992 13504 57044
rect 13728 57035 13780 57044
rect 13728 57001 13737 57035
rect 13737 57001 13771 57035
rect 13771 57001 13780 57035
rect 13728 56992 13780 57001
rect 14372 57035 14424 57044
rect 14372 57001 14381 57035
rect 14381 57001 14415 57035
rect 14415 57001 14424 57035
rect 14372 56992 14424 57001
rect 16580 56992 16632 57044
rect 20720 57035 20772 57044
rect 20720 57001 20729 57035
rect 20729 57001 20763 57035
rect 20763 57001 20772 57035
rect 20720 56992 20772 57001
rect 21640 56992 21692 57044
rect 23296 56992 23348 57044
rect 17224 56967 17276 56976
rect 1676 56899 1728 56908
rect 1676 56865 1685 56899
rect 1685 56865 1719 56899
rect 1719 56865 1728 56899
rect 1676 56856 1728 56865
rect 13268 56856 13320 56908
rect 14188 56899 14240 56908
rect 14188 56865 14197 56899
rect 14197 56865 14231 56899
rect 14231 56865 14240 56899
rect 14188 56856 14240 56865
rect 14740 56856 14792 56908
rect 17224 56933 17233 56967
rect 17233 56933 17267 56967
rect 17267 56933 17276 56967
rect 17224 56924 17276 56933
rect 16488 56856 16540 56908
rect 16580 56856 16632 56908
rect 18512 56856 18564 56908
rect 19984 56924 20036 56976
rect 19340 56899 19392 56908
rect 19340 56865 19349 56899
rect 19349 56865 19383 56899
rect 19383 56865 19392 56899
rect 19340 56856 19392 56865
rect 19708 56856 19760 56908
rect 20444 56856 20496 56908
rect 20996 56856 21048 56908
rect 22744 56856 22796 56908
rect 1584 56788 1636 56840
rect 2136 56788 2188 56840
rect 14924 56788 14976 56840
rect 17776 56788 17828 56840
rect 20076 56788 20128 56840
rect 21364 56788 21416 56840
rect 21824 56788 21876 56840
rect 15752 56720 15804 56772
rect 16212 56720 16264 56772
rect 16672 56720 16724 56772
rect 16948 56720 17000 56772
rect 17960 56720 18012 56772
rect 18052 56720 18104 56772
rect 19064 56720 19116 56772
rect 19524 56720 19576 56772
rect 19708 56720 19760 56772
rect 15108 56695 15160 56704
rect 15108 56661 15117 56695
rect 15117 56661 15151 56695
rect 15151 56661 15160 56695
rect 15108 56652 15160 56661
rect 17224 56652 17276 56704
rect 17500 56695 17552 56704
rect 17500 56661 17509 56695
rect 17509 56661 17543 56695
rect 17543 56661 17552 56695
rect 17500 56652 17552 56661
rect 17592 56652 17644 56704
rect 23296 56652 23348 56704
rect 23940 56652 23992 56704
rect 5982 56550 6034 56602
rect 6046 56550 6098 56602
rect 6110 56550 6162 56602
rect 6174 56550 6226 56602
rect 15982 56550 16034 56602
rect 16046 56550 16098 56602
rect 16110 56550 16162 56602
rect 16174 56550 16226 56602
rect 25982 56550 26034 56602
rect 26046 56550 26098 56602
rect 26110 56550 26162 56602
rect 26174 56550 26226 56602
rect 1676 56491 1728 56500
rect 1676 56457 1685 56491
rect 1685 56457 1719 56491
rect 1719 56457 1728 56491
rect 1676 56448 1728 56457
rect 2228 56448 2280 56500
rect 15200 56491 15252 56500
rect 15200 56457 15209 56491
rect 15209 56457 15243 56491
rect 15243 56457 15252 56491
rect 15200 56448 15252 56457
rect 17960 56448 18012 56500
rect 20720 56448 20772 56500
rect 20996 56448 21048 56500
rect 23020 56448 23072 56500
rect 25780 56448 25832 56500
rect 13728 56423 13780 56432
rect 13728 56389 13737 56423
rect 13737 56389 13771 56423
rect 13771 56389 13780 56423
rect 13728 56380 13780 56389
rect 15016 56380 15068 56432
rect 15108 56380 15160 56432
rect 16580 56423 16632 56432
rect 14280 56312 14332 56364
rect 15200 56312 15252 56364
rect 16120 56312 16172 56364
rect 16580 56389 16589 56423
rect 16589 56389 16623 56423
rect 16623 56389 16632 56423
rect 16580 56380 16632 56389
rect 17500 56380 17552 56432
rect 18328 56423 18380 56432
rect 18328 56389 18337 56423
rect 18337 56389 18371 56423
rect 18371 56389 18380 56423
rect 18328 56380 18380 56389
rect 19064 56380 19116 56432
rect 19340 56380 19392 56432
rect 15108 56176 15160 56228
rect 16488 56176 16540 56228
rect 13268 56151 13320 56160
rect 13268 56117 13277 56151
rect 13277 56117 13311 56151
rect 13311 56117 13320 56151
rect 13268 56108 13320 56117
rect 14280 56108 14332 56160
rect 15016 56108 15068 56160
rect 15568 56151 15620 56160
rect 15568 56117 15577 56151
rect 15577 56117 15611 56151
rect 15611 56117 15620 56151
rect 15568 56108 15620 56117
rect 16212 56108 16264 56160
rect 16672 56312 16724 56364
rect 17776 56312 17828 56364
rect 19616 56355 19668 56364
rect 16948 56108 17000 56160
rect 19616 56321 19625 56355
rect 19625 56321 19659 56355
rect 19659 56321 19668 56355
rect 19616 56312 19668 56321
rect 20352 56287 20404 56296
rect 18052 56219 18104 56228
rect 18052 56185 18061 56219
rect 18061 56185 18095 56219
rect 18095 56185 18104 56219
rect 18052 56176 18104 56185
rect 18420 56176 18472 56228
rect 20352 56253 20361 56287
rect 20361 56253 20395 56287
rect 20395 56253 20404 56287
rect 20352 56244 20404 56253
rect 20720 56244 20772 56296
rect 25872 56312 25924 56364
rect 21364 56244 21416 56296
rect 25780 56244 25832 56296
rect 21272 56176 21324 56228
rect 22468 56176 22520 56228
rect 22836 56176 22888 56228
rect 21640 56108 21692 56160
rect 22100 56151 22152 56160
rect 22100 56117 22109 56151
rect 22109 56117 22143 56151
rect 22143 56117 22152 56151
rect 22744 56151 22796 56160
rect 22100 56108 22152 56117
rect 22744 56117 22753 56151
rect 22753 56117 22787 56151
rect 22787 56117 22796 56151
rect 22744 56108 22796 56117
rect 24308 56108 24360 56160
rect 24676 56108 24728 56160
rect 27712 56151 27764 56160
rect 27712 56117 27721 56151
rect 27721 56117 27755 56151
rect 27755 56117 27764 56151
rect 27712 56108 27764 56117
rect 10982 56006 11034 56058
rect 11046 56006 11098 56058
rect 11110 56006 11162 56058
rect 11174 56006 11226 56058
rect 20982 56006 21034 56058
rect 21046 56006 21098 56058
rect 21110 56006 21162 56058
rect 21174 56006 21226 56058
rect 14004 55947 14056 55956
rect 14004 55913 14013 55947
rect 14013 55913 14047 55947
rect 14047 55913 14056 55947
rect 14004 55904 14056 55913
rect 14280 55904 14332 55956
rect 16120 55904 16172 55956
rect 17500 55904 17552 55956
rect 19984 55904 20036 55956
rect 20260 55904 20312 55956
rect 20444 55947 20496 55956
rect 20444 55913 20453 55947
rect 20453 55913 20487 55947
rect 20487 55913 20496 55947
rect 20444 55904 20496 55913
rect 21640 55904 21692 55956
rect 25872 55904 25924 55956
rect 14832 55836 14884 55888
rect 16212 55836 16264 55888
rect 17776 55836 17828 55888
rect 18788 55879 18840 55888
rect 18788 55845 18797 55879
rect 18797 55845 18831 55879
rect 18831 55845 18840 55879
rect 18788 55836 18840 55845
rect 19340 55836 19392 55888
rect 9680 55768 9732 55820
rect 10600 55768 10652 55820
rect 13176 55811 13228 55820
rect 13176 55777 13185 55811
rect 13185 55777 13219 55811
rect 13219 55777 13228 55811
rect 13176 55768 13228 55777
rect 14004 55768 14056 55820
rect 10876 55700 10928 55752
rect 14372 55632 14424 55684
rect 12072 55607 12124 55616
rect 12072 55573 12081 55607
rect 12081 55573 12115 55607
rect 12115 55573 12124 55607
rect 12072 55564 12124 55573
rect 13084 55564 13136 55616
rect 16856 55768 16908 55820
rect 16948 55743 17000 55752
rect 16948 55709 16957 55743
rect 16957 55709 16991 55743
rect 16991 55709 17000 55743
rect 16948 55700 17000 55709
rect 19064 55700 19116 55752
rect 20904 55811 20956 55820
rect 20904 55777 20913 55811
rect 20913 55777 20947 55811
rect 20947 55777 20956 55811
rect 20904 55768 20956 55777
rect 21640 55768 21692 55820
rect 22744 55836 22796 55888
rect 22376 55811 22428 55820
rect 22376 55777 22385 55811
rect 22385 55777 22419 55811
rect 22419 55777 22428 55811
rect 22376 55768 22428 55777
rect 23848 55768 23900 55820
rect 17040 55632 17092 55684
rect 20352 55700 20404 55752
rect 22744 55700 22796 55752
rect 26332 55700 26384 55752
rect 20168 55632 20220 55684
rect 14924 55564 14976 55616
rect 15108 55607 15160 55616
rect 15108 55573 15117 55607
rect 15117 55573 15151 55607
rect 15151 55573 15160 55607
rect 15108 55564 15160 55573
rect 15568 55564 15620 55616
rect 16488 55607 16540 55616
rect 16488 55573 16497 55607
rect 16497 55573 16531 55607
rect 16531 55573 16540 55607
rect 16488 55564 16540 55573
rect 17132 55564 17184 55616
rect 21088 55607 21140 55616
rect 21088 55573 21097 55607
rect 21097 55573 21131 55607
rect 21131 55573 21140 55607
rect 21088 55564 21140 55573
rect 22652 55564 22704 55616
rect 24860 55607 24912 55616
rect 24860 55573 24869 55607
rect 24869 55573 24903 55607
rect 24903 55573 24912 55607
rect 24860 55564 24912 55573
rect 5982 55462 6034 55514
rect 6046 55462 6098 55514
rect 6110 55462 6162 55514
rect 6174 55462 6226 55514
rect 15982 55462 16034 55514
rect 16046 55462 16098 55514
rect 16110 55462 16162 55514
rect 16174 55462 16226 55514
rect 25982 55462 26034 55514
rect 26046 55462 26098 55514
rect 26110 55462 26162 55514
rect 26174 55462 26226 55514
rect 10600 55403 10652 55412
rect 10600 55369 10609 55403
rect 10609 55369 10643 55403
rect 10643 55369 10652 55403
rect 10600 55360 10652 55369
rect 10876 55403 10928 55412
rect 10876 55369 10885 55403
rect 10885 55369 10919 55403
rect 10919 55369 10928 55403
rect 10876 55360 10928 55369
rect 13176 55360 13228 55412
rect 15016 55360 15068 55412
rect 16488 55360 16540 55412
rect 16672 55403 16724 55412
rect 16672 55369 16681 55403
rect 16681 55369 16715 55403
rect 16715 55369 16724 55403
rect 16672 55360 16724 55369
rect 16948 55360 17000 55412
rect 14740 55335 14792 55344
rect 14740 55301 14749 55335
rect 14749 55301 14783 55335
rect 14783 55301 14792 55335
rect 14740 55292 14792 55301
rect 15200 55292 15252 55344
rect 15936 55292 15988 55344
rect 17040 55335 17092 55344
rect 17040 55301 17049 55335
rect 17049 55301 17083 55335
rect 17083 55301 17092 55335
rect 17040 55292 17092 55301
rect 14648 55267 14700 55276
rect 14648 55233 14654 55267
rect 14654 55233 14700 55267
rect 14648 55224 14700 55233
rect 14832 55267 14884 55276
rect 14832 55233 14841 55267
rect 14841 55233 14875 55267
rect 14875 55233 14884 55267
rect 14832 55224 14884 55233
rect 17960 55360 18012 55412
rect 23112 55403 23164 55412
rect 23112 55369 23121 55403
rect 23121 55369 23155 55403
rect 23155 55369 23164 55403
rect 23112 55360 23164 55369
rect 23848 55403 23900 55412
rect 23848 55369 23857 55403
rect 23857 55369 23891 55403
rect 23891 55369 23900 55403
rect 23848 55360 23900 55369
rect 22376 55292 22428 55344
rect 22652 55267 22704 55276
rect 22652 55233 22661 55267
rect 22661 55233 22695 55267
rect 22695 55233 22704 55267
rect 22652 55224 22704 55233
rect 24032 55224 24084 55276
rect 27528 55224 27580 55276
rect 14464 55199 14516 55208
rect 14464 55165 14473 55199
rect 14473 55165 14507 55199
rect 14507 55165 14516 55199
rect 14464 55156 14516 55165
rect 16580 55156 16632 55208
rect 16856 55156 16908 55208
rect 18052 55199 18104 55208
rect 18052 55165 18061 55199
rect 18061 55165 18095 55199
rect 18095 55165 18104 55199
rect 18052 55156 18104 55165
rect 20628 55199 20680 55208
rect 20628 55165 20637 55199
rect 20637 55165 20671 55199
rect 20671 55165 20680 55199
rect 20628 55156 20680 55165
rect 22008 55156 22060 55208
rect 13268 55063 13320 55072
rect 13268 55029 13277 55063
rect 13277 55029 13311 55063
rect 13311 55029 13320 55063
rect 13268 55020 13320 55029
rect 17040 55088 17092 55140
rect 17500 55088 17552 55140
rect 18788 55131 18840 55140
rect 18788 55097 18797 55131
rect 18797 55097 18831 55131
rect 18831 55097 18840 55131
rect 18788 55088 18840 55097
rect 23112 55156 23164 55208
rect 24124 55156 24176 55208
rect 24492 55156 24544 55208
rect 14004 55020 14056 55072
rect 15108 55020 15160 55072
rect 15936 55063 15988 55072
rect 15936 55029 15945 55063
rect 15945 55029 15979 55063
rect 15979 55029 15988 55063
rect 15936 55020 15988 55029
rect 18052 55020 18104 55072
rect 19156 55020 19208 55072
rect 19984 55020 20036 55072
rect 24676 55088 24728 55140
rect 26240 55156 26292 55208
rect 21640 55063 21692 55072
rect 21640 55029 21649 55063
rect 21649 55029 21683 55063
rect 21683 55029 21692 55063
rect 21640 55020 21692 55029
rect 21916 55020 21968 55072
rect 24032 55020 24084 55072
rect 10982 54918 11034 54970
rect 11046 54918 11098 54970
rect 11110 54918 11162 54970
rect 11174 54918 11226 54970
rect 20982 54918 21034 54970
rect 21046 54918 21098 54970
rect 21110 54918 21162 54970
rect 21174 54918 21226 54970
rect 14464 54816 14516 54868
rect 15292 54816 15344 54868
rect 15568 54816 15620 54868
rect 17132 54859 17184 54868
rect 12072 54791 12124 54800
rect 12072 54757 12081 54791
rect 12081 54757 12115 54791
rect 12115 54757 12124 54791
rect 12072 54748 12124 54757
rect 12256 54680 12308 54732
rect 13820 54680 13872 54732
rect 14648 54748 14700 54800
rect 15016 54748 15068 54800
rect 17132 54825 17141 54859
rect 17141 54825 17175 54859
rect 17175 54825 17184 54859
rect 17132 54816 17184 54825
rect 17592 54816 17644 54868
rect 19340 54859 19392 54868
rect 19340 54825 19349 54859
rect 19349 54825 19383 54859
rect 19383 54825 19392 54859
rect 19340 54816 19392 54825
rect 19616 54859 19668 54868
rect 19616 54825 19625 54859
rect 19625 54825 19659 54859
rect 19659 54825 19668 54859
rect 19616 54816 19668 54825
rect 20168 54816 20220 54868
rect 21824 54816 21876 54868
rect 22376 54859 22428 54868
rect 22376 54825 22385 54859
rect 22385 54825 22419 54859
rect 22419 54825 22428 54859
rect 22376 54816 22428 54825
rect 24124 54816 24176 54868
rect 24676 54859 24728 54868
rect 24676 54825 24685 54859
rect 24685 54825 24719 54859
rect 24719 54825 24728 54859
rect 24676 54816 24728 54825
rect 16672 54791 16724 54800
rect 16672 54757 16681 54791
rect 16681 54757 16715 54791
rect 16715 54757 16724 54791
rect 16672 54748 16724 54757
rect 16856 54748 16908 54800
rect 17684 54748 17736 54800
rect 23204 54748 23256 54800
rect 14832 54680 14884 54732
rect 15292 54680 15344 54732
rect 11980 54544 12032 54596
rect 13084 54544 13136 54596
rect 14740 54612 14792 54664
rect 15200 54612 15252 54664
rect 16304 54612 16356 54664
rect 16488 54612 16540 54664
rect 17500 54612 17552 54664
rect 17960 54612 18012 54664
rect 18788 54680 18840 54732
rect 21088 54723 21140 54732
rect 21088 54689 21097 54723
rect 21097 54689 21131 54723
rect 21131 54689 21140 54723
rect 21088 54680 21140 54689
rect 21824 54723 21876 54732
rect 21824 54689 21833 54723
rect 21833 54689 21867 54723
rect 21867 54689 21876 54723
rect 21824 54680 21876 54689
rect 21916 54723 21968 54732
rect 21916 54689 21925 54723
rect 21925 54689 21959 54723
rect 21959 54689 21968 54723
rect 24768 54748 24820 54800
rect 21916 54680 21968 54689
rect 24216 54680 24268 54732
rect 24676 54680 24728 54732
rect 27712 54680 27764 54732
rect 18236 54612 18288 54664
rect 19156 54612 19208 54664
rect 20720 54612 20772 54664
rect 21364 54612 21416 54664
rect 23112 54612 23164 54664
rect 23572 54612 23624 54664
rect 26608 54655 26660 54664
rect 26608 54621 26617 54655
rect 26617 54621 26651 54655
rect 26651 54621 26660 54655
rect 26608 54612 26660 54621
rect 26976 54612 27028 54664
rect 27528 54655 27580 54664
rect 27528 54621 27537 54655
rect 27537 54621 27571 54655
rect 27571 54621 27580 54655
rect 27528 54612 27580 54621
rect 14924 54544 14976 54596
rect 15936 54587 15988 54596
rect 12348 54519 12400 54528
rect 12348 54485 12357 54519
rect 12357 54485 12391 54519
rect 12391 54485 12400 54519
rect 12348 54476 12400 54485
rect 13912 54476 13964 54528
rect 15108 54476 15160 54528
rect 15936 54553 15945 54587
rect 15945 54553 15979 54587
rect 15979 54553 15988 54587
rect 15936 54544 15988 54553
rect 16672 54544 16724 54596
rect 16304 54519 16356 54528
rect 16304 54485 16313 54519
rect 16313 54485 16347 54519
rect 16347 54485 16356 54519
rect 16304 54476 16356 54485
rect 20352 54519 20404 54528
rect 20352 54485 20361 54519
rect 20361 54485 20395 54519
rect 20395 54485 20404 54519
rect 20352 54476 20404 54485
rect 26332 54476 26384 54528
rect 5982 54374 6034 54426
rect 6046 54374 6098 54426
rect 6110 54374 6162 54426
rect 6174 54374 6226 54426
rect 15982 54374 16034 54426
rect 16046 54374 16098 54426
rect 16110 54374 16162 54426
rect 16174 54374 16226 54426
rect 25982 54374 26034 54426
rect 26046 54374 26098 54426
rect 26110 54374 26162 54426
rect 26174 54374 26226 54426
rect 12256 54315 12308 54324
rect 12256 54281 12265 54315
rect 12265 54281 12299 54315
rect 12299 54281 12308 54315
rect 12256 54272 12308 54281
rect 13820 54272 13872 54324
rect 16580 54315 16632 54324
rect 16580 54281 16589 54315
rect 16589 54281 16623 54315
rect 16623 54281 16632 54315
rect 16580 54272 16632 54281
rect 18512 54315 18564 54324
rect 18512 54281 18521 54315
rect 18521 54281 18555 54315
rect 18555 54281 18564 54315
rect 18512 54272 18564 54281
rect 19340 54272 19392 54324
rect 11888 54179 11940 54188
rect 11888 54145 11897 54179
rect 11897 54145 11931 54179
rect 11931 54145 11940 54179
rect 11888 54136 11940 54145
rect 15108 54204 15160 54256
rect 16028 54247 16080 54256
rect 16028 54213 16037 54247
rect 16037 54213 16071 54247
rect 16071 54213 16080 54247
rect 16028 54204 16080 54213
rect 12348 54068 12400 54120
rect 13452 54111 13504 54120
rect 13452 54077 13461 54111
rect 13461 54077 13495 54111
rect 13495 54077 13504 54111
rect 13452 54068 13504 54077
rect 13912 54068 13964 54120
rect 17960 54136 18012 54188
rect 18788 54136 18840 54188
rect 14832 54068 14884 54120
rect 14004 54043 14056 54052
rect 14004 54009 14013 54043
rect 14013 54009 14047 54043
rect 14047 54009 14056 54043
rect 14004 54000 14056 54009
rect 15016 54043 15068 54052
rect 15016 54009 15025 54043
rect 15025 54009 15059 54043
rect 15059 54009 15068 54043
rect 15016 54000 15068 54009
rect 15200 54000 15252 54052
rect 16120 54068 16172 54120
rect 16212 54000 16264 54052
rect 11520 53975 11572 53984
rect 11520 53941 11529 53975
rect 11529 53941 11563 53975
rect 11563 53941 11572 53975
rect 11520 53932 11572 53941
rect 13820 53975 13872 53984
rect 13820 53941 13829 53975
rect 13829 53941 13863 53975
rect 13863 53941 13872 53975
rect 13820 53932 13872 53941
rect 16856 53932 16908 53984
rect 21916 54272 21968 54324
rect 27712 54272 27764 54324
rect 25872 54179 25924 54188
rect 22192 54111 22244 54120
rect 22192 54077 22201 54111
rect 22201 54077 22235 54111
rect 22235 54077 22244 54111
rect 22192 54068 22244 54077
rect 22376 54068 22428 54120
rect 22652 54111 22704 54120
rect 22652 54077 22661 54111
rect 22661 54077 22695 54111
rect 22695 54077 22704 54111
rect 22652 54068 22704 54077
rect 23572 54068 23624 54120
rect 23664 54111 23716 54120
rect 23664 54077 23673 54111
rect 23673 54077 23707 54111
rect 23707 54077 23716 54111
rect 25872 54145 25881 54179
rect 25881 54145 25915 54179
rect 25915 54145 25924 54179
rect 25872 54136 25924 54145
rect 23664 54068 23716 54077
rect 25964 54111 26016 54120
rect 25964 54077 25973 54111
rect 25973 54077 26007 54111
rect 26007 54077 26016 54111
rect 25964 54068 26016 54077
rect 26332 54068 26384 54120
rect 18236 54043 18288 54052
rect 18236 54009 18245 54043
rect 18245 54009 18279 54043
rect 18279 54009 18288 54043
rect 18236 54000 18288 54009
rect 19340 54000 19392 54052
rect 19708 54000 19760 54052
rect 20628 54000 20680 54052
rect 23112 54000 23164 54052
rect 17684 53932 17736 53984
rect 18788 53932 18840 53984
rect 22468 53932 22520 53984
rect 23020 53932 23072 53984
rect 23664 53932 23716 53984
rect 27344 53975 27396 53984
rect 27344 53941 27353 53975
rect 27353 53941 27387 53975
rect 27387 53941 27396 53975
rect 27344 53932 27396 53941
rect 10982 53830 11034 53882
rect 11046 53830 11098 53882
rect 11110 53830 11162 53882
rect 11174 53830 11226 53882
rect 20982 53830 21034 53882
rect 21046 53830 21098 53882
rect 21110 53830 21162 53882
rect 21174 53830 21226 53882
rect 12072 53728 12124 53780
rect 18144 53728 18196 53780
rect 13912 53703 13964 53712
rect 13912 53669 13921 53703
rect 13921 53669 13955 53703
rect 13955 53669 13964 53703
rect 13912 53660 13964 53669
rect 17776 53660 17828 53712
rect 11244 53635 11296 53644
rect 11244 53601 11253 53635
rect 11253 53601 11287 53635
rect 11287 53601 11296 53635
rect 11244 53592 11296 53601
rect 12072 53592 12124 53644
rect 16212 53635 16264 53644
rect 16212 53601 16221 53635
rect 16221 53601 16255 53635
rect 16255 53601 16264 53635
rect 18052 53635 18104 53644
rect 16212 53592 16264 53601
rect 18052 53601 18061 53635
rect 18061 53601 18095 53635
rect 18095 53601 18104 53635
rect 18052 53592 18104 53601
rect 18236 53635 18288 53644
rect 18236 53601 18245 53635
rect 18245 53601 18279 53635
rect 18279 53601 18288 53635
rect 18236 53592 18288 53601
rect 12440 53524 12492 53576
rect 15200 53524 15252 53576
rect 16948 53524 17000 53576
rect 17316 53524 17368 53576
rect 17592 53567 17644 53576
rect 17592 53533 17601 53567
rect 17601 53533 17635 53567
rect 17635 53533 17644 53567
rect 17592 53524 17644 53533
rect 18144 53524 18196 53576
rect 18696 53728 18748 53780
rect 19156 53728 19208 53780
rect 20720 53771 20772 53780
rect 19616 53660 19668 53712
rect 20720 53737 20729 53771
rect 20729 53737 20763 53771
rect 20763 53737 20772 53771
rect 20720 53728 20772 53737
rect 21824 53728 21876 53780
rect 22376 53771 22428 53780
rect 22376 53737 22385 53771
rect 22385 53737 22419 53771
rect 22419 53737 22428 53771
rect 22376 53728 22428 53737
rect 23940 53728 23992 53780
rect 26608 53728 26660 53780
rect 18696 53592 18748 53644
rect 19432 53592 19484 53644
rect 19708 53635 19760 53644
rect 19708 53601 19717 53635
rect 19717 53601 19751 53635
rect 19751 53601 19760 53635
rect 19708 53592 19760 53601
rect 20168 53592 20220 53644
rect 21088 53592 21140 53644
rect 23112 53635 23164 53644
rect 23112 53601 23121 53635
rect 23121 53601 23155 53635
rect 23155 53601 23164 53635
rect 23112 53592 23164 53601
rect 23940 53635 23992 53644
rect 23940 53601 23949 53635
rect 23949 53601 23983 53635
rect 23983 53601 23992 53635
rect 23940 53592 23992 53601
rect 27528 53660 27580 53712
rect 21364 53567 21416 53576
rect 21364 53533 21373 53567
rect 21373 53533 21407 53567
rect 21407 53533 21416 53567
rect 21364 53524 21416 53533
rect 22376 53524 22428 53576
rect 25964 53567 26016 53576
rect 15292 53456 15344 53508
rect 16120 53456 16172 53508
rect 16672 53456 16724 53508
rect 20352 53456 20404 53508
rect 25964 53533 25973 53567
rect 25973 53533 26007 53567
rect 26007 53533 26016 53567
rect 25964 53524 26016 53533
rect 11428 53431 11480 53440
rect 11428 53397 11437 53431
rect 11437 53397 11471 53431
rect 11471 53397 11480 53431
rect 11428 53388 11480 53397
rect 11980 53388 12032 53440
rect 14004 53388 14056 53440
rect 14740 53388 14792 53440
rect 15108 53388 15160 53440
rect 16580 53388 16632 53440
rect 17040 53388 17092 53440
rect 17776 53388 17828 53440
rect 21824 53388 21876 53440
rect 22100 53388 22152 53440
rect 24768 53388 24820 53440
rect 5982 53286 6034 53338
rect 6046 53286 6098 53338
rect 6110 53286 6162 53338
rect 6174 53286 6226 53338
rect 15982 53286 16034 53338
rect 16046 53286 16098 53338
rect 16110 53286 16162 53338
rect 16174 53286 16226 53338
rect 25982 53286 26034 53338
rect 26046 53286 26098 53338
rect 26110 53286 26162 53338
rect 26174 53286 26226 53338
rect 10416 53184 10468 53236
rect 10876 53227 10928 53236
rect 10876 53193 10885 53227
rect 10885 53193 10919 53227
rect 10919 53193 10928 53227
rect 10876 53184 10928 53193
rect 11888 53227 11940 53236
rect 11888 53193 11897 53227
rect 11897 53193 11931 53227
rect 11931 53193 11940 53227
rect 11888 53184 11940 53193
rect 14464 53227 14516 53236
rect 14464 53193 14473 53227
rect 14473 53193 14507 53227
rect 14507 53193 14516 53227
rect 14464 53184 14516 53193
rect 15200 53184 15252 53236
rect 16488 53184 16540 53236
rect 17040 53227 17092 53236
rect 17040 53193 17049 53227
rect 17049 53193 17083 53227
rect 17083 53193 17092 53227
rect 17040 53184 17092 53193
rect 17776 53184 17828 53236
rect 16948 53116 17000 53168
rect 12440 53091 12492 53100
rect 12440 53057 12449 53091
rect 12449 53057 12483 53091
rect 12483 53057 12492 53091
rect 12440 53048 12492 53057
rect 12808 53048 12860 53100
rect 18788 53116 18840 53168
rect 11888 52980 11940 53032
rect 12164 52980 12216 53032
rect 12532 52980 12584 53032
rect 14004 52980 14056 53032
rect 16304 52980 16356 53032
rect 18420 53048 18472 53100
rect 20720 53184 20772 53236
rect 23112 53227 23164 53236
rect 19064 53048 19116 53100
rect 19616 53048 19668 53100
rect 20628 53091 20680 53100
rect 20628 53057 20637 53091
rect 20637 53057 20671 53091
rect 20671 53057 20680 53091
rect 20628 53048 20680 53057
rect 23112 53193 23121 53227
rect 23121 53193 23155 53227
rect 23155 53193 23164 53227
rect 23112 53184 23164 53193
rect 22744 53116 22796 53168
rect 23848 53184 23900 53236
rect 24492 53091 24544 53100
rect 24492 53057 24501 53091
rect 24501 53057 24535 53091
rect 24535 53057 24544 53091
rect 24492 53048 24544 53057
rect 11244 52955 11296 52964
rect 11244 52921 11253 52955
rect 11253 52921 11287 52955
rect 11287 52921 11296 52955
rect 11244 52912 11296 52921
rect 11428 52912 11480 52964
rect 11520 52887 11572 52896
rect 11520 52853 11529 52887
rect 11529 52853 11563 52887
rect 11563 52853 11572 52887
rect 11520 52844 11572 52853
rect 11888 52844 11940 52896
rect 12072 52844 12124 52896
rect 14004 52887 14056 52896
rect 14004 52853 14013 52887
rect 14013 52853 14047 52887
rect 14047 52853 14056 52887
rect 14004 52844 14056 52853
rect 15016 52844 15068 52896
rect 15200 52887 15252 52896
rect 15200 52853 15209 52887
rect 15209 52853 15243 52887
rect 15243 52853 15252 52887
rect 15200 52844 15252 52853
rect 17224 52844 17276 52896
rect 17592 52912 17644 52964
rect 18236 52887 18288 52896
rect 18236 52853 18245 52887
rect 18245 52853 18279 52887
rect 18279 52853 18288 52887
rect 18236 52844 18288 52853
rect 18880 52844 18932 52896
rect 19432 52912 19484 52964
rect 20720 52912 20772 52964
rect 21088 52955 21140 52964
rect 21088 52921 21097 52955
rect 21097 52921 21131 52955
rect 21131 52921 21140 52955
rect 21088 52912 21140 52921
rect 19708 52844 19760 52896
rect 20076 52844 20128 52896
rect 21916 52980 21968 53032
rect 24768 52980 24820 53032
rect 22192 52955 22244 52964
rect 22192 52921 22201 52955
rect 22201 52921 22235 52955
rect 22235 52921 22244 52955
rect 22192 52912 22244 52921
rect 22560 52844 22612 52896
rect 23940 52844 23992 52896
rect 10982 52742 11034 52794
rect 11046 52742 11098 52794
rect 11110 52742 11162 52794
rect 11174 52742 11226 52794
rect 20982 52742 21034 52794
rect 21046 52742 21098 52794
rect 21110 52742 21162 52794
rect 21174 52742 21226 52794
rect 10876 52640 10928 52692
rect 11796 52683 11848 52692
rect 11796 52649 11805 52683
rect 11805 52649 11839 52683
rect 11839 52649 11848 52683
rect 11796 52640 11848 52649
rect 13820 52683 13872 52692
rect 13820 52649 13829 52683
rect 13829 52649 13863 52683
rect 13863 52649 13872 52683
rect 13820 52640 13872 52649
rect 15108 52640 15160 52692
rect 16304 52640 16356 52692
rect 18420 52640 18472 52692
rect 19156 52683 19208 52692
rect 19156 52649 19165 52683
rect 19165 52649 19199 52683
rect 19199 52649 19208 52683
rect 19156 52640 19208 52649
rect 19984 52640 20036 52692
rect 20168 52640 20220 52692
rect 20720 52640 20772 52692
rect 23940 52640 23992 52692
rect 11888 52572 11940 52624
rect 14280 52572 14332 52624
rect 14464 52572 14516 52624
rect 14740 52615 14792 52624
rect 14740 52581 14749 52615
rect 14749 52581 14783 52615
rect 14783 52581 14792 52615
rect 14740 52572 14792 52581
rect 15016 52615 15068 52624
rect 15016 52581 15025 52615
rect 15025 52581 15059 52615
rect 15059 52581 15068 52615
rect 15016 52572 15068 52581
rect 18052 52572 18104 52624
rect 1676 52547 1728 52556
rect 1676 52513 1685 52547
rect 1685 52513 1719 52547
rect 1719 52513 1728 52547
rect 1676 52504 1728 52513
rect 4068 52504 4120 52556
rect 1584 52436 1636 52488
rect 11428 52504 11480 52556
rect 12256 52504 12308 52556
rect 12624 52547 12676 52556
rect 12624 52513 12633 52547
rect 12633 52513 12667 52547
rect 12667 52513 12676 52547
rect 12624 52504 12676 52513
rect 13912 52547 13964 52556
rect 13912 52513 13921 52547
rect 13921 52513 13955 52547
rect 13955 52513 13964 52547
rect 13912 52504 13964 52513
rect 12440 52479 12492 52488
rect 12440 52445 12449 52479
rect 12449 52445 12483 52479
rect 12483 52445 12492 52479
rect 12440 52436 12492 52445
rect 11336 52368 11388 52420
rect 11980 52300 12032 52352
rect 12992 52300 13044 52352
rect 14372 52436 14424 52488
rect 14740 52436 14792 52488
rect 15200 52436 15252 52488
rect 16304 52504 16356 52556
rect 17040 52547 17092 52556
rect 17040 52513 17049 52547
rect 17049 52513 17083 52547
rect 17083 52513 17092 52547
rect 17040 52504 17092 52513
rect 17776 52504 17828 52556
rect 21732 52572 21784 52624
rect 18788 52504 18840 52556
rect 21364 52504 21416 52556
rect 16488 52436 16540 52488
rect 17224 52436 17276 52488
rect 19340 52436 19392 52488
rect 20168 52436 20220 52488
rect 20720 52436 20772 52488
rect 22560 52504 22612 52556
rect 23296 52547 23348 52556
rect 23296 52513 23305 52547
rect 23305 52513 23339 52547
rect 23339 52513 23348 52547
rect 23296 52504 23348 52513
rect 21732 52479 21784 52488
rect 21732 52445 21741 52479
rect 21741 52445 21775 52479
rect 21775 52445 21784 52479
rect 21732 52436 21784 52445
rect 23112 52479 23164 52488
rect 23112 52445 23121 52479
rect 23121 52445 23155 52479
rect 23155 52445 23164 52479
rect 23112 52436 23164 52445
rect 24124 52504 24176 52556
rect 13728 52368 13780 52420
rect 15568 52368 15620 52420
rect 19432 52368 19484 52420
rect 19984 52368 20036 52420
rect 23204 52368 23256 52420
rect 23756 52411 23808 52420
rect 23756 52377 23765 52411
rect 23765 52377 23799 52411
rect 23799 52377 23808 52411
rect 23756 52368 23808 52377
rect 14832 52300 14884 52352
rect 16580 52300 16632 52352
rect 18236 52300 18288 52352
rect 20352 52343 20404 52352
rect 20352 52309 20361 52343
rect 20361 52309 20395 52343
rect 20395 52309 20404 52343
rect 20352 52300 20404 52309
rect 22192 52300 22244 52352
rect 23848 52300 23900 52352
rect 5982 52198 6034 52250
rect 6046 52198 6098 52250
rect 6110 52198 6162 52250
rect 6174 52198 6226 52250
rect 15982 52198 16034 52250
rect 16046 52198 16098 52250
rect 16110 52198 16162 52250
rect 16174 52198 16226 52250
rect 25982 52198 26034 52250
rect 26046 52198 26098 52250
rect 26110 52198 26162 52250
rect 26174 52198 26226 52250
rect 1676 52139 1728 52148
rect 1676 52105 1685 52139
rect 1685 52105 1719 52139
rect 1719 52105 1728 52139
rect 1676 52096 1728 52105
rect 8392 52139 8444 52148
rect 8392 52105 8401 52139
rect 8401 52105 8435 52139
rect 8435 52105 8444 52139
rect 8392 52096 8444 52105
rect 8392 51892 8444 51944
rect 10968 52096 11020 52148
rect 11336 52096 11388 52148
rect 12256 52139 12308 52148
rect 12256 52105 12265 52139
rect 12265 52105 12299 52139
rect 12299 52105 12308 52139
rect 12256 52096 12308 52105
rect 14832 52139 14884 52148
rect 14832 52105 14841 52139
rect 14841 52105 14875 52139
rect 14875 52105 14884 52139
rect 14832 52096 14884 52105
rect 15108 52096 15160 52148
rect 15568 52096 15620 52148
rect 18512 52096 18564 52148
rect 18604 52096 18656 52148
rect 18788 52096 18840 52148
rect 20720 52096 20772 52148
rect 21364 52096 21416 52148
rect 21548 52096 21600 52148
rect 22468 52096 22520 52148
rect 23112 52096 23164 52148
rect 13912 52028 13964 52080
rect 18420 52028 18472 52080
rect 18972 52028 19024 52080
rect 11980 51960 12032 52012
rect 15292 52003 15344 52012
rect 12808 51935 12860 51944
rect 12808 51901 12817 51935
rect 12817 51901 12851 51935
rect 12851 51901 12860 51935
rect 12808 51892 12860 51901
rect 1584 51756 1636 51808
rect 7840 51799 7892 51808
rect 7840 51765 7849 51799
rect 7849 51765 7883 51799
rect 7883 51765 7892 51799
rect 7840 51756 7892 51765
rect 10508 51799 10560 51808
rect 10508 51765 10517 51799
rect 10517 51765 10551 51799
rect 10551 51765 10560 51799
rect 10508 51756 10560 51765
rect 12348 51756 12400 51808
rect 12624 51799 12676 51808
rect 12624 51765 12633 51799
rect 12633 51765 12667 51799
rect 12667 51765 12676 51799
rect 15292 51969 15301 52003
rect 15301 51969 15335 52003
rect 15335 51969 15344 52003
rect 15292 51960 15344 51969
rect 16120 51960 16172 52012
rect 19156 52003 19208 52012
rect 19156 51969 19165 52003
rect 19165 51969 19199 52003
rect 19199 51969 19208 52003
rect 19156 51960 19208 51969
rect 24860 52096 24912 52148
rect 23756 52028 23808 52080
rect 23940 52028 23992 52080
rect 24124 52028 24176 52080
rect 16672 51892 16724 51944
rect 17040 51892 17092 51944
rect 18512 51935 18564 51944
rect 16028 51824 16080 51876
rect 16488 51824 16540 51876
rect 18052 51824 18104 51876
rect 18512 51901 18521 51935
rect 18521 51901 18555 51935
rect 18555 51901 18564 51935
rect 18512 51892 18564 51901
rect 18604 51892 18656 51944
rect 19340 51892 19392 51944
rect 20168 51892 20220 51944
rect 23296 51960 23348 52012
rect 23480 51960 23532 52012
rect 21364 51935 21416 51944
rect 12624 51756 12676 51765
rect 15292 51756 15344 51808
rect 16304 51799 16356 51808
rect 16304 51765 16313 51799
rect 16313 51765 16347 51799
rect 16347 51765 16356 51799
rect 16304 51756 16356 51765
rect 18512 51756 18564 51808
rect 18972 51756 19024 51808
rect 20352 51756 20404 51808
rect 21364 51901 21373 51935
rect 21373 51901 21407 51935
rect 21407 51901 21416 51935
rect 21364 51892 21416 51901
rect 21732 51892 21784 51944
rect 21732 51756 21784 51808
rect 23664 51867 23716 51876
rect 23664 51833 23673 51867
rect 23673 51833 23707 51867
rect 23707 51833 23716 51867
rect 23664 51824 23716 51833
rect 23848 51867 23900 51876
rect 23848 51833 23857 51867
rect 23857 51833 23891 51867
rect 23891 51833 23900 51867
rect 23848 51824 23900 51833
rect 24860 51824 24912 51876
rect 23940 51799 23992 51808
rect 23940 51765 23949 51799
rect 23949 51765 23983 51799
rect 23983 51765 23992 51799
rect 23940 51756 23992 51765
rect 10982 51654 11034 51706
rect 11046 51654 11098 51706
rect 11110 51654 11162 51706
rect 11174 51654 11226 51706
rect 20982 51654 21034 51706
rect 21046 51654 21098 51706
rect 21110 51654 21162 51706
rect 21174 51654 21226 51706
rect 10416 51595 10468 51604
rect 10416 51561 10425 51595
rect 10425 51561 10459 51595
rect 10459 51561 10468 51595
rect 10416 51552 10468 51561
rect 10784 51552 10836 51604
rect 11980 51552 12032 51604
rect 12716 51552 12768 51604
rect 13544 51552 13596 51604
rect 14832 51595 14884 51604
rect 14832 51561 14841 51595
rect 14841 51561 14875 51595
rect 14875 51561 14884 51595
rect 14832 51552 14884 51561
rect 16672 51595 16724 51604
rect 16672 51561 16681 51595
rect 16681 51561 16715 51595
rect 16715 51561 16724 51595
rect 16672 51552 16724 51561
rect 17960 51552 18012 51604
rect 19064 51595 19116 51604
rect 19064 51561 19073 51595
rect 19073 51561 19107 51595
rect 19107 51561 19116 51595
rect 19064 51552 19116 51561
rect 19524 51552 19576 51604
rect 21364 51552 21416 51604
rect 13268 51484 13320 51536
rect 13912 51484 13964 51536
rect 6276 51416 6328 51468
rect 10416 51416 10468 51468
rect 12256 51416 12308 51468
rect 12716 51416 12768 51468
rect 12992 51416 13044 51468
rect 14924 51484 14976 51536
rect 17040 51484 17092 51536
rect 19432 51484 19484 51536
rect 21732 51484 21784 51536
rect 16028 51459 16080 51468
rect 16028 51425 16037 51459
rect 16037 51425 16071 51459
rect 16071 51425 16080 51459
rect 16028 51416 16080 51425
rect 16120 51416 16172 51468
rect 14004 51391 14056 51400
rect 11520 51280 11572 51332
rect 14004 51357 14013 51391
rect 14013 51357 14047 51391
rect 14047 51357 14056 51391
rect 14004 51348 14056 51357
rect 14188 51348 14240 51400
rect 15476 51348 15528 51400
rect 16304 51348 16356 51400
rect 17776 51459 17828 51468
rect 17776 51425 17785 51459
rect 17785 51425 17819 51459
rect 17819 51425 17828 51459
rect 17776 51416 17828 51425
rect 18052 51459 18104 51468
rect 18052 51425 18061 51459
rect 18061 51425 18095 51459
rect 18095 51425 18104 51459
rect 18052 51416 18104 51425
rect 18604 51416 18656 51468
rect 19340 51416 19392 51468
rect 21548 51459 21600 51468
rect 21548 51425 21557 51459
rect 21557 51425 21591 51459
rect 21591 51425 21600 51459
rect 21548 51416 21600 51425
rect 21916 51459 21968 51468
rect 21916 51425 21925 51459
rect 21925 51425 21959 51459
rect 21959 51425 21968 51459
rect 21916 51416 21968 51425
rect 22100 51484 22152 51536
rect 16672 51348 16724 51400
rect 18144 51348 18196 51400
rect 18972 51348 19024 51400
rect 20352 51348 20404 51400
rect 22100 51348 22152 51400
rect 13452 51280 13504 51332
rect 5816 51212 5868 51264
rect 11980 51212 12032 51264
rect 13084 51212 13136 51264
rect 14280 51255 14332 51264
rect 14280 51221 14289 51255
rect 14289 51221 14323 51255
rect 14323 51221 14332 51255
rect 14280 51212 14332 51221
rect 14832 51212 14884 51264
rect 15200 51212 15252 51264
rect 16580 51280 16632 51332
rect 17040 51280 17092 51332
rect 17592 51280 17644 51332
rect 16488 51212 16540 51264
rect 19156 51212 19208 51264
rect 21548 51280 21600 51332
rect 23204 51459 23256 51468
rect 23204 51425 23213 51459
rect 23213 51425 23247 51459
rect 23247 51425 23256 51459
rect 23204 51416 23256 51425
rect 23848 51552 23900 51604
rect 23940 51552 23992 51604
rect 25504 51552 25556 51604
rect 25688 51552 25740 51604
rect 23756 51484 23808 51536
rect 23112 51348 23164 51400
rect 23296 51348 23348 51400
rect 19984 51212 20036 51264
rect 21732 51212 21784 51264
rect 23296 51212 23348 51264
rect 24124 51416 24176 51468
rect 23480 51348 23532 51400
rect 23848 51280 23900 51332
rect 24032 51280 24084 51332
rect 24768 51212 24820 51264
rect 25780 51212 25832 51264
rect 5982 51110 6034 51162
rect 6046 51110 6098 51162
rect 6110 51110 6162 51162
rect 6174 51110 6226 51162
rect 15982 51110 16034 51162
rect 16046 51110 16098 51162
rect 16110 51110 16162 51162
rect 16174 51110 16226 51162
rect 25982 51110 26034 51162
rect 26046 51110 26098 51162
rect 26110 51110 26162 51162
rect 26174 51110 26226 51162
rect 6276 51008 6328 51060
rect 10416 51051 10468 51060
rect 10416 51017 10425 51051
rect 10425 51017 10459 51051
rect 10459 51017 10468 51051
rect 10416 51008 10468 51017
rect 11888 51008 11940 51060
rect 12256 51051 12308 51060
rect 12256 51017 12265 51051
rect 12265 51017 12299 51051
rect 12299 51017 12308 51051
rect 12256 51008 12308 51017
rect 12992 51008 13044 51060
rect 11520 50983 11572 50992
rect 11520 50949 11529 50983
rect 11529 50949 11563 50983
rect 11563 50949 11572 50983
rect 11520 50940 11572 50949
rect 14004 51008 14056 51060
rect 11060 50804 11112 50856
rect 13452 50872 13504 50924
rect 14924 51008 14976 51060
rect 17592 51008 17644 51060
rect 18604 51008 18656 51060
rect 19524 51008 19576 51060
rect 14648 50940 14700 50992
rect 16304 50940 16356 50992
rect 19432 50940 19484 50992
rect 17132 50915 17184 50924
rect 13544 50847 13596 50856
rect 13544 50813 13553 50847
rect 13553 50813 13587 50847
rect 13587 50813 13596 50847
rect 13544 50804 13596 50813
rect 13912 50804 13964 50856
rect 15108 50804 15160 50856
rect 16580 50847 16632 50856
rect 16580 50813 16589 50847
rect 16589 50813 16623 50847
rect 16623 50813 16632 50847
rect 16580 50804 16632 50813
rect 17132 50881 17141 50915
rect 17141 50881 17175 50915
rect 17175 50881 17184 50915
rect 17132 50872 17184 50881
rect 19064 50872 19116 50924
rect 19340 50872 19392 50924
rect 16948 50804 17000 50856
rect 18512 50804 18564 50856
rect 22100 51008 22152 51060
rect 23480 51008 23532 51060
rect 24308 51051 24360 51060
rect 24308 51017 24317 51051
rect 24317 51017 24351 51051
rect 24351 51017 24360 51051
rect 24308 51008 24360 51017
rect 20812 50940 20864 50992
rect 21456 50940 21508 50992
rect 24124 50940 24176 50992
rect 22008 50872 22060 50924
rect 22560 50872 22612 50924
rect 15292 50736 15344 50788
rect 19340 50736 19392 50788
rect 14464 50668 14516 50720
rect 15476 50711 15528 50720
rect 15476 50677 15485 50711
rect 15485 50677 15519 50711
rect 15519 50677 15528 50711
rect 15476 50668 15528 50677
rect 19064 50668 19116 50720
rect 19432 50668 19484 50720
rect 19984 50804 20036 50856
rect 20444 50668 20496 50720
rect 23020 50804 23072 50856
rect 20812 50736 20864 50788
rect 21180 50779 21232 50788
rect 21180 50745 21189 50779
rect 21189 50745 21223 50779
rect 21223 50745 21232 50779
rect 21180 50736 21232 50745
rect 21548 50779 21600 50788
rect 21548 50745 21557 50779
rect 21557 50745 21591 50779
rect 21591 50745 21600 50779
rect 21548 50736 21600 50745
rect 22008 50736 22060 50788
rect 24768 50872 24820 50924
rect 23756 50847 23808 50856
rect 23756 50813 23765 50847
rect 23765 50813 23799 50847
rect 23799 50813 23808 50847
rect 23756 50804 23808 50813
rect 24308 50804 24360 50856
rect 24492 50736 24544 50788
rect 20720 50668 20772 50720
rect 22744 50668 22796 50720
rect 23020 50668 23072 50720
rect 23296 50668 23348 50720
rect 24308 50668 24360 50720
rect 25136 50668 25188 50720
rect 10982 50566 11034 50618
rect 11046 50566 11098 50618
rect 11110 50566 11162 50618
rect 11174 50566 11226 50618
rect 20982 50566 21034 50618
rect 21046 50566 21098 50618
rect 21110 50566 21162 50618
rect 21174 50566 21226 50618
rect 12716 50464 12768 50516
rect 12992 50507 13044 50516
rect 12992 50473 13001 50507
rect 13001 50473 13035 50507
rect 13035 50473 13044 50507
rect 12992 50464 13044 50473
rect 13544 50464 13596 50516
rect 14648 50464 14700 50516
rect 15292 50464 15344 50516
rect 15752 50464 15804 50516
rect 16304 50464 16356 50516
rect 16672 50464 16724 50516
rect 18512 50507 18564 50516
rect 18512 50473 18521 50507
rect 18521 50473 18555 50507
rect 18555 50473 18564 50507
rect 18512 50464 18564 50473
rect 20352 50507 20404 50516
rect 20352 50473 20361 50507
rect 20361 50473 20395 50507
rect 20395 50473 20404 50507
rect 20352 50464 20404 50473
rect 21272 50464 21324 50516
rect 21456 50464 21508 50516
rect 24308 50507 24360 50516
rect 24308 50473 24317 50507
rect 24317 50473 24351 50507
rect 24351 50473 24360 50507
rect 24308 50464 24360 50473
rect 12348 50396 12400 50448
rect 14924 50396 14976 50448
rect 10784 50328 10836 50380
rect 11428 50328 11480 50380
rect 14004 50328 14056 50380
rect 14188 50371 14240 50380
rect 14188 50337 14197 50371
rect 14197 50337 14231 50371
rect 14231 50337 14240 50371
rect 14188 50328 14240 50337
rect 15200 50396 15252 50448
rect 17500 50396 17552 50448
rect 17776 50439 17828 50448
rect 17776 50405 17785 50439
rect 17785 50405 17819 50439
rect 17819 50405 17828 50439
rect 17776 50396 17828 50405
rect 22008 50396 22060 50448
rect 22468 50439 22520 50448
rect 10876 50260 10928 50312
rect 15108 50260 15160 50312
rect 15752 50371 15804 50380
rect 15752 50337 15761 50371
rect 15761 50337 15795 50371
rect 15795 50337 15804 50371
rect 15752 50328 15804 50337
rect 16488 50260 16540 50312
rect 16672 50260 16724 50312
rect 17316 50371 17368 50380
rect 17316 50337 17325 50371
rect 17325 50337 17359 50371
rect 17359 50337 17368 50371
rect 17316 50328 17368 50337
rect 17960 50328 18012 50380
rect 19340 50328 19392 50380
rect 11796 50167 11848 50176
rect 11796 50133 11805 50167
rect 11805 50133 11839 50167
rect 11839 50133 11848 50167
rect 11796 50124 11848 50133
rect 15752 50124 15804 50176
rect 18420 50260 18472 50312
rect 19156 50260 19208 50312
rect 19708 50303 19760 50312
rect 19708 50269 19717 50303
rect 19717 50269 19751 50303
rect 19751 50269 19760 50303
rect 19708 50260 19760 50269
rect 20352 50260 20404 50312
rect 22008 50260 22060 50312
rect 22468 50405 22477 50439
rect 22477 50405 22511 50439
rect 22511 50405 22520 50439
rect 22468 50396 22520 50405
rect 22836 50439 22888 50448
rect 22836 50405 22845 50439
rect 22845 50405 22879 50439
rect 22879 50405 22888 50439
rect 22836 50396 22888 50405
rect 23204 50439 23256 50448
rect 23204 50405 23213 50439
rect 23213 50405 23247 50439
rect 23247 50405 23256 50439
rect 23204 50396 23256 50405
rect 22192 50328 22244 50380
rect 22744 50371 22796 50380
rect 22744 50337 22753 50371
rect 22753 50337 22787 50371
rect 22787 50337 22796 50371
rect 24308 50371 24360 50380
rect 22744 50328 22796 50337
rect 24308 50337 24317 50371
rect 24317 50337 24351 50371
rect 24351 50337 24360 50371
rect 24308 50328 24360 50337
rect 18144 50167 18196 50176
rect 18144 50133 18153 50167
rect 18153 50133 18187 50167
rect 18187 50133 18196 50167
rect 18144 50124 18196 50133
rect 21548 50124 21600 50176
rect 22284 50167 22336 50176
rect 22284 50133 22293 50167
rect 22293 50133 22327 50167
rect 22327 50133 22336 50167
rect 22284 50124 22336 50133
rect 5982 50022 6034 50074
rect 6046 50022 6098 50074
rect 6110 50022 6162 50074
rect 6174 50022 6226 50074
rect 15982 50022 16034 50074
rect 16046 50022 16098 50074
rect 16110 50022 16162 50074
rect 16174 50022 16226 50074
rect 25982 50022 26034 50074
rect 26046 50022 26098 50074
rect 26110 50022 26162 50074
rect 26174 50022 26226 50074
rect 8944 49963 8996 49972
rect 8944 49929 8953 49963
rect 8953 49929 8987 49963
rect 8987 49929 8996 49963
rect 8944 49920 8996 49929
rect 10876 49920 10928 49972
rect 12256 49963 12308 49972
rect 7380 49827 7432 49836
rect 7380 49793 7389 49827
rect 7389 49793 7423 49827
rect 7423 49793 7432 49827
rect 7380 49784 7432 49793
rect 10324 49827 10376 49836
rect 10324 49793 10333 49827
rect 10333 49793 10367 49827
rect 10367 49793 10376 49827
rect 10324 49784 10376 49793
rect 10784 49759 10836 49768
rect 10784 49725 10793 49759
rect 10793 49725 10827 49759
rect 10827 49725 10836 49759
rect 10784 49716 10836 49725
rect 12256 49929 12265 49963
rect 12265 49929 12299 49963
rect 12299 49929 12308 49963
rect 12256 49920 12308 49929
rect 13452 49920 13504 49972
rect 14004 49920 14056 49972
rect 15292 49920 15344 49972
rect 17500 49963 17552 49972
rect 15568 49852 15620 49904
rect 12164 49784 12216 49836
rect 12808 49784 12860 49836
rect 13268 49827 13320 49836
rect 13268 49793 13277 49827
rect 13277 49793 13311 49827
rect 13311 49793 13320 49827
rect 13268 49784 13320 49793
rect 13728 49784 13780 49836
rect 13912 49784 13964 49836
rect 17500 49929 17509 49963
rect 17509 49929 17543 49963
rect 17543 49929 17552 49963
rect 17500 49920 17552 49929
rect 17960 49920 18012 49972
rect 18420 49963 18472 49972
rect 18420 49929 18429 49963
rect 18429 49929 18463 49963
rect 18463 49929 18472 49963
rect 18420 49920 18472 49929
rect 20352 49920 20404 49972
rect 22192 49963 22244 49972
rect 22192 49929 22201 49963
rect 22201 49929 22235 49963
rect 22235 49929 22244 49963
rect 22192 49920 22244 49929
rect 22468 49963 22520 49972
rect 22468 49929 22477 49963
rect 22477 49929 22511 49963
rect 22511 49929 22520 49963
rect 22468 49920 22520 49929
rect 22744 49920 22796 49972
rect 23572 49920 23624 49972
rect 16856 49852 16908 49904
rect 17316 49852 17368 49904
rect 18880 49852 18932 49904
rect 20904 49852 20956 49904
rect 22008 49852 22060 49904
rect 11704 49716 11756 49768
rect 14648 49716 14700 49768
rect 15292 49716 15344 49768
rect 16028 49759 16080 49768
rect 16028 49725 16037 49759
rect 16037 49725 16071 49759
rect 16071 49725 16080 49759
rect 16028 49716 16080 49725
rect 16488 49716 16540 49768
rect 15016 49648 15068 49700
rect 18144 49784 18196 49836
rect 19340 49784 19392 49836
rect 17776 49716 17828 49768
rect 18696 49759 18748 49768
rect 18696 49725 18705 49759
rect 18705 49725 18739 49759
rect 18739 49725 18748 49759
rect 18696 49716 18748 49725
rect 18972 49759 19024 49768
rect 18972 49725 18981 49759
rect 18981 49725 19015 49759
rect 19015 49725 19024 49759
rect 18972 49716 19024 49725
rect 22560 49784 22612 49836
rect 22744 49784 22796 49836
rect 23204 49784 23256 49836
rect 24492 49784 24544 49836
rect 20444 49716 20496 49768
rect 23572 49716 23624 49768
rect 24308 49716 24360 49768
rect 17316 49648 17368 49700
rect 19524 49648 19576 49700
rect 20812 49648 20864 49700
rect 21456 49691 21508 49700
rect 21456 49657 21465 49691
rect 21465 49657 21499 49691
rect 21499 49657 21508 49691
rect 21456 49648 21508 49657
rect 7196 49623 7248 49632
rect 7196 49589 7205 49623
rect 7205 49589 7239 49623
rect 7239 49589 7248 49623
rect 7196 49580 7248 49589
rect 11428 49580 11480 49632
rect 20720 49580 20772 49632
rect 21272 49580 21324 49632
rect 22376 49580 22428 49632
rect 25228 49580 25280 49632
rect 10982 49478 11034 49530
rect 11046 49478 11098 49530
rect 11110 49478 11162 49530
rect 11174 49478 11226 49530
rect 20982 49478 21034 49530
rect 21046 49478 21098 49530
rect 21110 49478 21162 49530
rect 21174 49478 21226 49530
rect 7380 49419 7432 49428
rect 7380 49385 7389 49419
rect 7389 49385 7423 49419
rect 7423 49385 7432 49419
rect 7380 49376 7432 49385
rect 10876 49376 10928 49428
rect 13268 49376 13320 49428
rect 16488 49419 16540 49428
rect 16488 49385 16497 49419
rect 16497 49385 16531 49419
rect 16531 49385 16540 49419
rect 16488 49376 16540 49385
rect 17776 49419 17828 49428
rect 17776 49385 17785 49419
rect 17785 49385 17819 49419
rect 17819 49385 17828 49419
rect 17776 49376 17828 49385
rect 18144 49419 18196 49428
rect 18144 49385 18153 49419
rect 18153 49385 18187 49419
rect 18187 49385 18196 49419
rect 18144 49376 18196 49385
rect 18512 49376 18564 49428
rect 19800 49376 19852 49428
rect 14924 49308 14976 49360
rect 15752 49308 15804 49360
rect 16304 49308 16356 49360
rect 11796 49240 11848 49292
rect 12256 49240 12308 49292
rect 13728 49240 13780 49292
rect 15292 49240 15344 49292
rect 16580 49240 16632 49292
rect 17592 49308 17644 49360
rect 16856 49283 16908 49292
rect 16856 49249 16865 49283
rect 16865 49249 16899 49283
rect 16899 49249 16908 49283
rect 16856 49240 16908 49249
rect 17224 49283 17276 49292
rect 17224 49249 17233 49283
rect 17233 49249 17267 49283
rect 17267 49249 17276 49283
rect 17224 49240 17276 49249
rect 17960 49240 18012 49292
rect 18972 49240 19024 49292
rect 19432 49240 19484 49292
rect 20352 49240 20404 49292
rect 21272 49376 21324 49428
rect 21916 49308 21968 49360
rect 23940 49308 23992 49360
rect 22376 49283 22428 49292
rect 22376 49249 22385 49283
rect 22385 49249 22419 49283
rect 22419 49249 22428 49283
rect 22376 49240 22428 49249
rect 22560 49283 22612 49292
rect 22560 49249 22569 49283
rect 22569 49249 22603 49283
rect 22603 49249 22612 49283
rect 22560 49240 22612 49249
rect 24768 49283 24820 49292
rect 24768 49249 24777 49283
rect 24777 49249 24811 49283
rect 24811 49249 24820 49283
rect 24768 49240 24820 49249
rect 25136 49240 25188 49292
rect 11336 49215 11388 49224
rect 11336 49181 11345 49215
rect 11345 49181 11379 49215
rect 11379 49181 11388 49215
rect 11336 49172 11388 49181
rect 11520 49172 11572 49224
rect 12716 49215 12768 49224
rect 12716 49181 12725 49215
rect 12725 49181 12759 49215
rect 12759 49181 12768 49215
rect 12716 49172 12768 49181
rect 18144 49172 18196 49224
rect 18420 49172 18472 49224
rect 19340 49215 19392 49224
rect 19340 49181 19349 49215
rect 19349 49181 19383 49215
rect 19383 49181 19392 49215
rect 19340 49172 19392 49181
rect 23940 49172 23992 49224
rect 24400 49172 24452 49224
rect 10784 49104 10836 49156
rect 11428 49036 11480 49088
rect 21640 49104 21692 49156
rect 13912 49036 13964 49088
rect 14832 49036 14884 49088
rect 15292 49036 15344 49088
rect 15660 49036 15712 49088
rect 19064 49036 19116 49088
rect 19340 49036 19392 49088
rect 19984 49036 20036 49088
rect 22100 49104 22152 49156
rect 22836 49036 22888 49088
rect 23480 49036 23532 49088
rect 24400 49079 24452 49088
rect 24400 49045 24409 49079
rect 24409 49045 24443 49079
rect 24443 49045 24452 49079
rect 24400 49036 24452 49045
rect 5982 48934 6034 48986
rect 6046 48934 6098 48986
rect 6110 48934 6162 48986
rect 6174 48934 6226 48986
rect 15982 48934 16034 48986
rect 16046 48934 16098 48986
rect 16110 48934 16162 48986
rect 16174 48934 16226 48986
rect 25982 48934 26034 48986
rect 26046 48934 26098 48986
rect 26110 48934 26162 48986
rect 26174 48934 26226 48986
rect 11796 48875 11848 48884
rect 11796 48841 11805 48875
rect 11805 48841 11839 48875
rect 11839 48841 11848 48875
rect 11796 48832 11848 48841
rect 12256 48875 12308 48884
rect 12256 48841 12265 48875
rect 12265 48841 12299 48875
rect 12299 48841 12308 48875
rect 12256 48832 12308 48841
rect 12900 48832 12952 48884
rect 13544 48875 13596 48884
rect 13544 48841 13553 48875
rect 13553 48841 13587 48875
rect 13587 48841 13596 48875
rect 13544 48832 13596 48841
rect 15200 48832 15252 48884
rect 16856 48832 16908 48884
rect 18420 48832 18472 48884
rect 19432 48875 19484 48884
rect 19432 48841 19441 48875
rect 19441 48841 19475 48875
rect 19475 48841 19484 48875
rect 19432 48832 19484 48841
rect 15476 48807 15528 48816
rect 15476 48773 15485 48807
rect 15485 48773 15519 48807
rect 15519 48773 15528 48807
rect 15476 48764 15528 48773
rect 16580 48764 16632 48816
rect 12900 48628 12952 48680
rect 13636 48671 13688 48680
rect 13636 48637 13645 48671
rect 13645 48637 13679 48671
rect 13679 48637 13688 48671
rect 13636 48628 13688 48637
rect 14648 48671 14700 48680
rect 14648 48637 14657 48671
rect 14657 48637 14691 48671
rect 14691 48637 14700 48671
rect 14648 48628 14700 48637
rect 14740 48628 14792 48680
rect 16304 48696 16356 48748
rect 17132 48696 17184 48748
rect 21272 48832 21324 48884
rect 22376 48832 22428 48884
rect 24768 48875 24820 48884
rect 24768 48841 24777 48875
rect 24777 48841 24811 48875
rect 24811 48841 24820 48875
rect 24768 48832 24820 48841
rect 25412 48875 25464 48884
rect 25412 48841 25421 48875
rect 25421 48841 25455 48875
rect 25455 48841 25464 48875
rect 25412 48832 25464 48841
rect 19984 48739 20036 48748
rect 19984 48705 19993 48739
rect 19993 48705 20027 48739
rect 20027 48705 20036 48739
rect 19984 48696 20036 48705
rect 22928 48696 22980 48748
rect 23664 48739 23716 48748
rect 23664 48705 23673 48739
rect 23673 48705 23707 48739
rect 23707 48705 23716 48739
rect 23664 48696 23716 48705
rect 16488 48628 16540 48680
rect 16948 48671 17000 48680
rect 16948 48637 16957 48671
rect 16957 48637 16991 48671
rect 16991 48637 17000 48671
rect 18052 48671 18104 48680
rect 16948 48628 17000 48637
rect 15108 48560 15160 48612
rect 11336 48492 11388 48544
rect 12808 48535 12860 48544
rect 12808 48501 12817 48535
rect 12817 48501 12851 48535
rect 12851 48501 12860 48535
rect 12808 48492 12860 48501
rect 13820 48535 13872 48544
rect 13820 48501 13829 48535
rect 13829 48501 13863 48535
rect 13863 48501 13872 48535
rect 13820 48492 13872 48501
rect 17316 48492 17368 48544
rect 18052 48637 18061 48671
rect 18061 48637 18095 48671
rect 18095 48637 18104 48671
rect 18052 48628 18104 48637
rect 18236 48628 18288 48680
rect 18604 48628 18656 48680
rect 19064 48671 19116 48680
rect 19064 48637 19073 48671
rect 19073 48637 19107 48671
rect 19107 48637 19116 48671
rect 19064 48628 19116 48637
rect 19800 48628 19852 48680
rect 21456 48628 21508 48680
rect 22008 48628 22060 48680
rect 17684 48560 17736 48612
rect 17776 48492 17828 48544
rect 18328 48535 18380 48544
rect 18328 48501 18337 48535
rect 18337 48501 18371 48535
rect 18371 48501 18380 48535
rect 18328 48492 18380 48501
rect 19156 48560 19208 48612
rect 22468 48671 22520 48680
rect 22468 48637 22477 48671
rect 22477 48637 22511 48671
rect 22511 48637 22520 48671
rect 22468 48628 22520 48637
rect 25228 48671 25280 48680
rect 25228 48637 25237 48671
rect 25237 48637 25271 48671
rect 25271 48637 25280 48671
rect 25228 48628 25280 48637
rect 21456 48492 21508 48544
rect 10982 48390 11034 48442
rect 11046 48390 11098 48442
rect 11110 48390 11162 48442
rect 11174 48390 11226 48442
rect 20982 48390 21034 48442
rect 21046 48390 21098 48442
rect 21110 48390 21162 48442
rect 21174 48390 21226 48442
rect 11428 48288 11480 48340
rect 13636 48288 13688 48340
rect 14740 48331 14792 48340
rect 14740 48297 14749 48331
rect 14749 48297 14783 48331
rect 14783 48297 14792 48331
rect 14740 48288 14792 48297
rect 13176 48220 13228 48272
rect 13360 48263 13412 48272
rect 13360 48229 13369 48263
rect 13369 48229 13403 48263
rect 13403 48229 13412 48263
rect 13360 48220 13412 48229
rect 15660 48288 15712 48340
rect 14188 48195 14240 48204
rect 14188 48161 14197 48195
rect 14197 48161 14231 48195
rect 14231 48161 14240 48195
rect 14188 48152 14240 48161
rect 13728 48084 13780 48136
rect 14832 48152 14884 48204
rect 15752 48220 15804 48272
rect 17224 48220 17276 48272
rect 17684 48195 17736 48204
rect 13452 48016 13504 48068
rect 15752 48084 15804 48136
rect 14648 48016 14700 48068
rect 15016 48059 15068 48068
rect 15016 48025 15025 48059
rect 15025 48025 15059 48059
rect 15059 48025 15068 48059
rect 15016 48016 15068 48025
rect 15108 48016 15160 48068
rect 15292 48016 15344 48068
rect 15476 48016 15528 48068
rect 17684 48161 17693 48195
rect 17693 48161 17727 48195
rect 17727 48161 17736 48195
rect 19064 48288 19116 48340
rect 19800 48288 19852 48340
rect 18880 48263 18932 48272
rect 18880 48229 18889 48263
rect 18889 48229 18923 48263
rect 18923 48229 18932 48263
rect 18880 48220 18932 48229
rect 18972 48220 19024 48272
rect 18052 48195 18104 48204
rect 17684 48152 17736 48161
rect 18052 48161 18061 48195
rect 18061 48161 18095 48195
rect 18095 48161 18104 48195
rect 18052 48152 18104 48161
rect 18236 48195 18288 48204
rect 18236 48161 18245 48195
rect 18245 48161 18279 48195
rect 18279 48161 18288 48195
rect 18236 48152 18288 48161
rect 19892 48152 19944 48204
rect 20076 48152 20128 48204
rect 16672 48084 16724 48136
rect 19156 48084 19208 48136
rect 19800 48084 19852 48136
rect 19984 48127 20036 48136
rect 19984 48093 19993 48127
rect 19993 48093 20027 48127
rect 20027 48093 20036 48127
rect 19984 48084 20036 48093
rect 18880 48016 18932 48068
rect 16856 47948 16908 48000
rect 19156 47991 19208 48000
rect 19156 47957 19165 47991
rect 19165 47957 19199 47991
rect 19199 47957 19208 47991
rect 19156 47948 19208 47957
rect 21548 48220 21600 48272
rect 22560 48288 22612 48340
rect 22652 48195 22704 48204
rect 21548 48084 21600 48136
rect 21548 47948 21600 48000
rect 22652 48161 22661 48195
rect 22661 48161 22695 48195
rect 22695 48161 22704 48195
rect 22652 48152 22704 48161
rect 22928 48220 22980 48272
rect 25136 48263 25188 48272
rect 25136 48229 25145 48263
rect 25145 48229 25179 48263
rect 25179 48229 25188 48263
rect 25136 48220 25188 48229
rect 23572 48152 23624 48204
rect 24676 48195 24728 48204
rect 24676 48161 24685 48195
rect 24685 48161 24719 48195
rect 24719 48161 24728 48195
rect 24676 48152 24728 48161
rect 23756 48127 23808 48136
rect 22836 48016 22888 48068
rect 23756 48093 23765 48127
rect 23765 48093 23799 48127
rect 23799 48093 23808 48127
rect 23756 48084 23808 48093
rect 23480 47948 23532 48000
rect 24860 47991 24912 48000
rect 24860 47957 24869 47991
rect 24869 47957 24903 47991
rect 24903 47957 24912 47991
rect 24860 47948 24912 47957
rect 26332 47948 26384 48000
rect 5982 47846 6034 47898
rect 6046 47846 6098 47898
rect 6110 47846 6162 47898
rect 6174 47846 6226 47898
rect 15982 47846 16034 47898
rect 16046 47846 16098 47898
rect 16110 47846 16162 47898
rect 16174 47846 16226 47898
rect 25982 47846 26034 47898
rect 26046 47846 26098 47898
rect 26110 47846 26162 47898
rect 26174 47846 26226 47898
rect 7840 47744 7892 47796
rect 13084 47787 13136 47796
rect 13084 47753 13093 47787
rect 13093 47753 13127 47787
rect 13127 47753 13136 47787
rect 13084 47744 13136 47753
rect 13452 47787 13504 47796
rect 13452 47753 13461 47787
rect 13461 47753 13495 47787
rect 13495 47753 13504 47787
rect 13452 47744 13504 47753
rect 13820 47744 13872 47796
rect 14464 47744 14516 47796
rect 14648 47787 14700 47796
rect 14648 47753 14657 47787
rect 14657 47753 14691 47787
rect 14691 47753 14700 47787
rect 14648 47744 14700 47753
rect 15200 47744 15252 47796
rect 16856 47787 16908 47796
rect 13728 47676 13780 47728
rect 14188 47608 14240 47660
rect 16856 47753 16865 47787
rect 16865 47753 16899 47787
rect 16899 47753 16908 47787
rect 16856 47744 16908 47753
rect 17040 47744 17092 47796
rect 19800 47787 19852 47796
rect 19800 47753 19809 47787
rect 19809 47753 19843 47787
rect 19843 47753 19852 47787
rect 19800 47744 19852 47753
rect 19892 47744 19944 47796
rect 23112 47787 23164 47796
rect 23112 47753 23121 47787
rect 23121 47753 23155 47787
rect 23155 47753 23164 47787
rect 23112 47744 23164 47753
rect 24492 47744 24544 47796
rect 24676 47744 24728 47796
rect 27712 47787 27764 47796
rect 27712 47753 27721 47787
rect 27721 47753 27755 47787
rect 27755 47753 27764 47787
rect 27712 47744 27764 47753
rect 17316 47676 17368 47728
rect 17592 47676 17644 47728
rect 16488 47651 16540 47660
rect 16488 47617 16497 47651
rect 16497 47617 16531 47651
rect 16531 47617 16540 47651
rect 16488 47608 16540 47617
rect 18052 47608 18104 47660
rect 19984 47676 20036 47728
rect 20352 47676 20404 47728
rect 22652 47676 22704 47728
rect 23572 47676 23624 47728
rect 23756 47676 23808 47728
rect 8208 47583 8260 47592
rect 8208 47549 8217 47583
rect 8217 47549 8251 47583
rect 8251 47549 8260 47583
rect 8208 47540 8260 47549
rect 15660 47540 15712 47592
rect 16304 47583 16356 47592
rect 16304 47549 16313 47583
rect 16313 47549 16347 47583
rect 16347 47549 16356 47583
rect 16304 47540 16356 47549
rect 17592 47583 17644 47592
rect 17592 47549 17601 47583
rect 17601 47549 17635 47583
rect 17635 47549 17644 47583
rect 17592 47540 17644 47549
rect 18788 47540 18840 47592
rect 18972 47583 19024 47592
rect 18972 47549 18981 47583
rect 18981 47549 19015 47583
rect 19015 47549 19024 47583
rect 19616 47608 19668 47660
rect 24400 47608 24452 47660
rect 18972 47540 19024 47549
rect 19156 47540 19208 47592
rect 20720 47540 20772 47592
rect 21272 47540 21324 47592
rect 21456 47583 21508 47592
rect 21456 47549 21465 47583
rect 21465 47549 21499 47583
rect 21499 47549 21508 47583
rect 21456 47540 21508 47549
rect 21640 47540 21692 47592
rect 23480 47583 23532 47592
rect 23480 47549 23489 47583
rect 23489 47549 23523 47583
rect 23523 47549 23532 47583
rect 23480 47540 23532 47549
rect 23756 47540 23808 47592
rect 24492 47583 24544 47592
rect 24492 47549 24501 47583
rect 24501 47549 24535 47583
rect 24535 47549 24544 47583
rect 24492 47540 24544 47549
rect 16212 47472 16264 47524
rect 22560 47472 22612 47524
rect 23204 47472 23256 47524
rect 24124 47472 24176 47524
rect 9772 47447 9824 47456
rect 9772 47413 9781 47447
rect 9781 47413 9815 47447
rect 9815 47413 9824 47447
rect 9772 47404 9824 47413
rect 11980 47404 12032 47456
rect 15016 47447 15068 47456
rect 15016 47413 15025 47447
rect 15025 47413 15059 47447
rect 15059 47413 15068 47447
rect 15016 47404 15068 47413
rect 20444 47404 20496 47456
rect 21548 47447 21600 47456
rect 21548 47413 21557 47447
rect 21557 47413 21591 47447
rect 21591 47413 21600 47447
rect 21548 47404 21600 47413
rect 25780 47608 25832 47660
rect 26332 47608 26384 47660
rect 26884 47608 26936 47660
rect 25872 47540 25924 47592
rect 25412 47404 25464 47456
rect 10982 47302 11034 47354
rect 11046 47302 11098 47354
rect 11110 47302 11162 47354
rect 11174 47302 11226 47354
rect 20982 47302 21034 47354
rect 21046 47302 21098 47354
rect 21110 47302 21162 47354
rect 21174 47302 21226 47354
rect 8208 47243 8260 47252
rect 8208 47209 8217 47243
rect 8217 47209 8251 47243
rect 8251 47209 8260 47243
rect 8208 47200 8260 47209
rect 13728 47243 13780 47252
rect 13728 47209 13737 47243
rect 13737 47209 13771 47243
rect 13771 47209 13780 47243
rect 13728 47200 13780 47209
rect 14004 47243 14056 47252
rect 14004 47209 14013 47243
rect 14013 47209 14047 47243
rect 14047 47209 14056 47243
rect 14004 47200 14056 47209
rect 14096 47200 14148 47252
rect 14740 47243 14792 47252
rect 14740 47209 14749 47243
rect 14749 47209 14783 47243
rect 14783 47209 14792 47243
rect 14740 47200 14792 47209
rect 17500 47200 17552 47252
rect 17960 47200 18012 47252
rect 21640 47200 21692 47252
rect 22652 47200 22704 47252
rect 22744 47200 22796 47252
rect 23664 47200 23716 47252
rect 24124 47243 24176 47252
rect 24124 47209 24133 47243
rect 24133 47209 24167 47243
rect 24167 47209 24176 47243
rect 26700 47243 26752 47252
rect 24124 47200 24176 47209
rect 14924 47132 14976 47184
rect 12532 47107 12584 47116
rect 12532 47073 12541 47107
rect 12541 47073 12575 47107
rect 12575 47073 12584 47107
rect 12532 47064 12584 47073
rect 13728 47064 13780 47116
rect 14188 47107 14240 47116
rect 14188 47073 14197 47107
rect 14197 47073 14231 47107
rect 14231 47073 14240 47107
rect 14188 47064 14240 47073
rect 14464 47064 14516 47116
rect 15476 47064 15528 47116
rect 17132 47132 17184 47184
rect 16304 47064 16356 47116
rect 17316 47064 17368 47116
rect 17776 47132 17828 47184
rect 18328 47132 18380 47184
rect 22468 47175 22520 47184
rect 22468 47141 22477 47175
rect 22477 47141 22511 47175
rect 22511 47141 22520 47175
rect 22468 47132 22520 47141
rect 17960 47064 18012 47116
rect 18972 47107 19024 47116
rect 18972 47073 18981 47107
rect 18981 47073 19015 47107
rect 19015 47073 19024 47107
rect 18972 47064 19024 47073
rect 19156 47064 19208 47116
rect 19708 47064 19760 47116
rect 20996 47107 21048 47116
rect 20996 47073 21005 47107
rect 21005 47073 21039 47107
rect 21039 47073 21048 47107
rect 20996 47064 21048 47073
rect 21640 47064 21692 47116
rect 22008 47064 22060 47116
rect 22744 47064 22796 47116
rect 23204 47132 23256 47184
rect 23296 47107 23348 47116
rect 23296 47073 23305 47107
rect 23305 47073 23339 47107
rect 23339 47073 23348 47107
rect 23296 47064 23348 47073
rect 26700 47209 26709 47243
rect 26709 47209 26743 47243
rect 26743 47209 26752 47243
rect 26700 47200 26752 47209
rect 24768 47064 24820 47116
rect 25320 47107 25372 47116
rect 25320 47073 25329 47107
rect 25329 47073 25363 47107
rect 25363 47073 25372 47107
rect 25320 47064 25372 47073
rect 25688 47064 25740 47116
rect 26516 47107 26568 47116
rect 26516 47073 26525 47107
rect 26525 47073 26559 47107
rect 26559 47073 26568 47107
rect 26516 47064 26568 47073
rect 12624 47039 12676 47048
rect 12624 47005 12633 47039
rect 12633 47005 12667 47039
rect 12667 47005 12676 47039
rect 12624 46996 12676 47005
rect 15200 46996 15252 47048
rect 16672 46996 16724 47048
rect 24308 46996 24360 47048
rect 16120 46971 16172 46980
rect 16120 46937 16129 46971
rect 16129 46937 16163 46971
rect 16163 46937 16172 46971
rect 16120 46928 16172 46937
rect 17592 46971 17644 46980
rect 17592 46937 17601 46971
rect 17601 46937 17635 46971
rect 17635 46937 17644 46971
rect 17592 46928 17644 46937
rect 18236 46928 18288 46980
rect 24492 46928 24544 46980
rect 19892 46903 19944 46912
rect 19892 46869 19901 46903
rect 19901 46869 19935 46903
rect 19935 46869 19944 46903
rect 19892 46860 19944 46869
rect 21456 46860 21508 46912
rect 21732 46860 21784 46912
rect 22008 46903 22060 46912
rect 22008 46869 22017 46903
rect 22017 46869 22051 46903
rect 22051 46869 22060 46903
rect 22008 46860 22060 46869
rect 25872 46860 25924 46912
rect 5982 46758 6034 46810
rect 6046 46758 6098 46810
rect 6110 46758 6162 46810
rect 6174 46758 6226 46810
rect 15982 46758 16034 46810
rect 16046 46758 16098 46810
rect 16110 46758 16162 46810
rect 16174 46758 16226 46810
rect 25982 46758 26034 46810
rect 26046 46758 26098 46810
rect 26110 46758 26162 46810
rect 26174 46758 26226 46810
rect 13728 46656 13780 46708
rect 14464 46699 14516 46708
rect 14464 46665 14473 46699
rect 14473 46665 14507 46699
rect 14507 46665 14516 46699
rect 14464 46656 14516 46665
rect 14924 46699 14976 46708
rect 14924 46665 14933 46699
rect 14933 46665 14967 46699
rect 14967 46665 14976 46699
rect 14924 46656 14976 46665
rect 15016 46656 15068 46708
rect 17316 46656 17368 46708
rect 17684 46656 17736 46708
rect 18052 46656 18104 46708
rect 12532 46631 12584 46640
rect 12532 46597 12541 46631
rect 12541 46597 12575 46631
rect 12575 46597 12584 46631
rect 12532 46588 12584 46597
rect 15200 46520 15252 46572
rect 16120 46520 16172 46572
rect 12440 46495 12492 46504
rect 12440 46461 12449 46495
rect 12449 46461 12483 46495
rect 12483 46461 12492 46495
rect 12716 46495 12768 46504
rect 12440 46452 12492 46461
rect 12716 46461 12725 46495
rect 12725 46461 12759 46495
rect 12759 46461 12768 46495
rect 12716 46452 12768 46461
rect 16212 46495 16264 46504
rect 16212 46461 16221 46495
rect 16221 46461 16255 46495
rect 16255 46461 16264 46495
rect 16212 46452 16264 46461
rect 17960 46520 18012 46572
rect 19064 46520 19116 46572
rect 19708 46563 19760 46572
rect 19708 46529 19717 46563
rect 19717 46529 19751 46563
rect 19751 46529 19760 46563
rect 19708 46520 19760 46529
rect 23572 46656 23624 46708
rect 20720 46563 20772 46572
rect 20720 46529 20729 46563
rect 20729 46529 20763 46563
rect 20763 46529 20772 46563
rect 20720 46520 20772 46529
rect 21732 46588 21784 46640
rect 22100 46588 22152 46640
rect 22468 46588 22520 46640
rect 23204 46588 23256 46640
rect 23480 46588 23532 46640
rect 22376 46520 22428 46572
rect 24400 46588 24452 46640
rect 26516 46656 26568 46708
rect 18328 46495 18380 46504
rect 15752 46384 15804 46436
rect 18328 46461 18337 46495
rect 18337 46461 18371 46495
rect 18371 46461 18380 46495
rect 18328 46452 18380 46461
rect 19892 46452 19944 46504
rect 17132 46427 17184 46436
rect 17132 46393 17141 46427
rect 17141 46393 17175 46427
rect 17175 46393 17184 46427
rect 17132 46384 17184 46393
rect 18788 46384 18840 46436
rect 19340 46384 19392 46436
rect 19708 46384 19760 46436
rect 19800 46384 19852 46436
rect 20996 46427 21048 46436
rect 20996 46393 21005 46427
rect 21005 46393 21039 46427
rect 21039 46393 21048 46427
rect 20996 46384 21048 46393
rect 23480 46452 23532 46504
rect 24860 46495 24912 46504
rect 24860 46461 24869 46495
rect 24869 46461 24903 46495
rect 24903 46461 24912 46495
rect 24860 46452 24912 46461
rect 25964 46495 26016 46504
rect 25964 46461 25973 46495
rect 25973 46461 26007 46495
rect 26007 46461 26016 46495
rect 25964 46452 26016 46461
rect 11888 46359 11940 46368
rect 11888 46325 11897 46359
rect 11897 46325 11931 46359
rect 11931 46325 11940 46359
rect 11888 46316 11940 46325
rect 12348 46316 12400 46368
rect 14188 46359 14240 46368
rect 14188 46325 14197 46359
rect 14197 46325 14231 46359
rect 14231 46325 14240 46359
rect 14188 46316 14240 46325
rect 15568 46359 15620 46368
rect 15568 46325 15577 46359
rect 15577 46325 15611 46359
rect 15611 46325 15620 46359
rect 15568 46316 15620 46325
rect 19156 46359 19208 46368
rect 19156 46325 19165 46359
rect 19165 46325 19199 46359
rect 19199 46325 19208 46359
rect 19156 46316 19208 46325
rect 20352 46316 20404 46368
rect 22744 46427 22796 46436
rect 22744 46393 22753 46427
rect 22753 46393 22787 46427
rect 22787 46393 22796 46427
rect 22744 46384 22796 46393
rect 25136 46427 25188 46436
rect 22100 46316 22152 46368
rect 22192 46316 22244 46368
rect 22468 46316 22520 46368
rect 23572 46316 23624 46368
rect 23940 46316 23992 46368
rect 24768 46316 24820 46368
rect 25136 46393 25145 46427
rect 25145 46393 25179 46427
rect 25179 46393 25188 46427
rect 25136 46384 25188 46393
rect 25044 46316 25096 46368
rect 26516 46427 26568 46436
rect 26516 46393 26525 46427
rect 26525 46393 26559 46427
rect 26559 46393 26568 46427
rect 26516 46384 26568 46393
rect 26332 46316 26384 46368
rect 10982 46214 11034 46266
rect 11046 46214 11098 46266
rect 11110 46214 11162 46266
rect 11174 46214 11226 46266
rect 20982 46214 21034 46266
rect 21046 46214 21098 46266
rect 21110 46214 21162 46266
rect 21174 46214 21226 46266
rect 11888 46155 11940 46164
rect 11888 46121 11897 46155
rect 11897 46121 11931 46155
rect 11931 46121 11940 46155
rect 11888 46112 11940 46121
rect 14096 46112 14148 46164
rect 16120 46112 16172 46164
rect 16212 46112 16264 46164
rect 17224 46112 17276 46164
rect 17500 46155 17552 46164
rect 17500 46121 17509 46155
rect 17509 46121 17543 46155
rect 17543 46121 17552 46155
rect 17500 46112 17552 46121
rect 18788 46112 18840 46164
rect 19800 46112 19852 46164
rect 23204 46112 23256 46164
rect 13268 46044 13320 46096
rect 15568 46044 15620 46096
rect 12440 46019 12492 46028
rect 12440 45985 12449 46019
rect 12449 45985 12483 46019
rect 12483 45985 12492 46019
rect 12440 45976 12492 45985
rect 12716 46019 12768 46028
rect 12716 45985 12725 46019
rect 12725 45985 12759 46019
rect 12759 45985 12768 46019
rect 12716 45976 12768 45985
rect 13452 45976 13504 46028
rect 15476 46019 15528 46028
rect 15476 45985 15485 46019
rect 15485 45985 15519 46019
rect 15519 45985 15528 46019
rect 15476 45976 15528 45985
rect 13820 45908 13872 45960
rect 14188 45908 14240 45960
rect 15752 45976 15804 46028
rect 16580 45976 16632 46028
rect 17040 45976 17092 46028
rect 22744 46044 22796 46096
rect 19064 45976 19116 46028
rect 19432 45976 19484 46028
rect 20720 45976 20772 46028
rect 21088 46019 21140 46028
rect 21088 45985 21097 46019
rect 21097 45985 21131 46019
rect 21131 45985 21140 46019
rect 21088 45976 21140 45985
rect 23204 45976 23256 46028
rect 23480 46112 23532 46164
rect 24400 46112 24452 46164
rect 24676 46112 24728 46164
rect 25320 46112 25372 46164
rect 25780 46044 25832 46096
rect 16488 45908 16540 45960
rect 19156 45951 19208 45960
rect 19156 45917 19165 45951
rect 19165 45917 19199 45951
rect 19199 45917 19208 45951
rect 19156 45908 19208 45917
rect 22560 45908 22612 45960
rect 23480 45976 23532 46028
rect 24124 45976 24176 46028
rect 24492 45908 24544 45960
rect 12624 45840 12676 45892
rect 16120 45883 16172 45892
rect 16120 45849 16129 45883
rect 16129 45849 16163 45883
rect 16163 45849 16172 45883
rect 16120 45840 16172 45849
rect 16672 45840 16724 45892
rect 24860 45840 24912 45892
rect 25964 45976 26016 46028
rect 1584 45815 1636 45824
rect 1584 45781 1593 45815
rect 1593 45781 1627 45815
rect 1627 45781 1636 45815
rect 1584 45772 1636 45781
rect 14464 45815 14516 45824
rect 14464 45781 14473 45815
rect 14473 45781 14507 45815
rect 14507 45781 14516 45815
rect 14464 45772 14516 45781
rect 18328 45815 18380 45824
rect 18328 45781 18337 45815
rect 18337 45781 18371 45815
rect 18371 45781 18380 45815
rect 18328 45772 18380 45781
rect 20076 45772 20128 45824
rect 20904 45772 20956 45824
rect 22100 45772 22152 45824
rect 23296 45772 23348 45824
rect 23940 45772 23992 45824
rect 24400 45772 24452 45824
rect 25872 45772 25924 45824
rect 5982 45670 6034 45722
rect 6046 45670 6098 45722
rect 6110 45670 6162 45722
rect 6174 45670 6226 45722
rect 15982 45670 16034 45722
rect 16046 45670 16098 45722
rect 16110 45670 16162 45722
rect 16174 45670 16226 45722
rect 25982 45670 26034 45722
rect 26046 45670 26098 45722
rect 26110 45670 26162 45722
rect 26174 45670 26226 45722
rect 12256 45568 12308 45620
rect 15476 45611 15528 45620
rect 1584 45432 1636 45484
rect 1768 45432 1820 45484
rect 12348 45500 12400 45552
rect 13912 45500 13964 45552
rect 15476 45577 15485 45611
rect 15485 45577 15519 45611
rect 15519 45577 15528 45611
rect 15476 45568 15528 45577
rect 17224 45568 17276 45620
rect 17684 45568 17736 45620
rect 18696 45568 18748 45620
rect 18880 45568 18932 45620
rect 20720 45568 20772 45620
rect 21088 45568 21140 45620
rect 22744 45568 22796 45620
rect 23480 45568 23532 45620
rect 23664 45568 23716 45620
rect 24492 45568 24544 45620
rect 17776 45500 17828 45552
rect 12440 45364 12492 45416
rect 13636 45432 13688 45484
rect 12624 45364 12676 45416
rect 13452 45407 13504 45416
rect 13452 45373 13461 45407
rect 13461 45373 13495 45407
rect 13495 45373 13504 45407
rect 13452 45364 13504 45373
rect 14096 45364 14148 45416
rect 14464 45407 14516 45416
rect 14464 45373 14473 45407
rect 14473 45373 14507 45407
rect 14507 45373 14516 45407
rect 14464 45364 14516 45373
rect 17408 45432 17460 45484
rect 19800 45500 19852 45552
rect 18972 45432 19024 45484
rect 16488 45364 16540 45416
rect 17224 45364 17276 45416
rect 18328 45407 18380 45416
rect 4068 45296 4120 45348
rect 14004 45296 14056 45348
rect 14556 45296 14608 45348
rect 17592 45296 17644 45348
rect 18328 45373 18337 45407
rect 18337 45373 18371 45407
rect 18371 45373 18380 45407
rect 18328 45364 18380 45373
rect 19432 45364 19484 45416
rect 19984 45407 20036 45416
rect 19984 45373 19993 45407
rect 19993 45373 20027 45407
rect 20027 45373 20036 45407
rect 19984 45364 20036 45373
rect 20352 45407 20404 45416
rect 20352 45373 20361 45407
rect 20361 45373 20395 45407
rect 20395 45373 20404 45407
rect 20352 45364 20404 45373
rect 20904 45407 20956 45416
rect 20904 45373 20913 45407
rect 20913 45373 20947 45407
rect 20947 45373 20956 45407
rect 20904 45364 20956 45373
rect 19064 45296 19116 45348
rect 22008 45364 22060 45416
rect 22376 45407 22428 45416
rect 22376 45373 22385 45407
rect 22385 45373 22419 45407
rect 22419 45373 22428 45407
rect 22376 45364 22428 45373
rect 22652 45339 22704 45348
rect 22652 45305 22661 45339
rect 22661 45305 22695 45339
rect 22695 45305 22704 45339
rect 22652 45296 22704 45305
rect 11520 45271 11572 45280
rect 11520 45237 11529 45271
rect 11529 45237 11563 45271
rect 11563 45237 11572 45271
rect 11520 45228 11572 45237
rect 19340 45271 19392 45280
rect 19340 45237 19349 45271
rect 19349 45237 19383 45271
rect 19383 45237 19392 45271
rect 19340 45228 19392 45237
rect 21732 45271 21784 45280
rect 21732 45237 21741 45271
rect 21741 45237 21775 45271
rect 21775 45237 21784 45271
rect 21732 45228 21784 45237
rect 23664 45432 23716 45484
rect 24676 45500 24728 45552
rect 24492 45364 24544 45416
rect 23848 45339 23900 45348
rect 23848 45305 23857 45339
rect 23857 45305 23891 45339
rect 23891 45305 23900 45339
rect 23848 45296 23900 45305
rect 25044 45364 25096 45416
rect 25136 45296 25188 45348
rect 24676 45228 24728 45280
rect 25044 45228 25096 45280
rect 25228 45228 25280 45280
rect 25780 45271 25832 45280
rect 25780 45237 25789 45271
rect 25789 45237 25823 45271
rect 25823 45237 25832 45271
rect 25780 45228 25832 45237
rect 26332 45339 26384 45348
rect 26332 45305 26341 45339
rect 26341 45305 26375 45339
rect 26375 45305 26384 45339
rect 26332 45296 26384 45305
rect 26056 45228 26108 45280
rect 26608 45271 26660 45280
rect 26608 45237 26617 45271
rect 26617 45237 26651 45271
rect 26651 45237 26660 45271
rect 26608 45228 26660 45237
rect 10982 45126 11034 45178
rect 11046 45126 11098 45178
rect 11110 45126 11162 45178
rect 11174 45126 11226 45178
rect 20982 45126 21034 45178
rect 21046 45126 21098 45178
rect 21110 45126 21162 45178
rect 21174 45126 21226 45178
rect 1768 45024 1820 45076
rect 1952 45067 2004 45076
rect 1952 45033 1961 45067
rect 1961 45033 1995 45067
rect 1995 45033 2004 45067
rect 1952 45024 2004 45033
rect 12624 45024 12676 45076
rect 14556 45067 14608 45076
rect 14556 45033 14565 45067
rect 14565 45033 14599 45067
rect 14599 45033 14608 45067
rect 14556 45024 14608 45033
rect 15752 45024 15804 45076
rect 16856 45067 16908 45076
rect 16856 45033 16865 45067
rect 16865 45033 16899 45067
rect 16899 45033 16908 45067
rect 16856 45024 16908 45033
rect 17040 45024 17092 45076
rect 18144 45067 18196 45076
rect 18144 45033 18153 45067
rect 18153 45033 18187 45067
rect 18187 45033 18196 45067
rect 18144 45024 18196 45033
rect 20352 45024 20404 45076
rect 21548 45024 21600 45076
rect 22008 45024 22060 45076
rect 23296 45067 23348 45076
rect 23296 45033 23305 45067
rect 23305 45033 23339 45067
rect 23339 45033 23348 45067
rect 23296 45024 23348 45033
rect 23664 45067 23716 45076
rect 23664 45033 23673 45067
rect 23673 45033 23707 45067
rect 23707 45033 23716 45067
rect 23664 45024 23716 45033
rect 24860 45067 24912 45076
rect 24860 45033 24869 45067
rect 24869 45033 24903 45067
rect 24903 45033 24912 45067
rect 24860 45024 24912 45033
rect 25780 45024 25832 45076
rect 26700 45067 26752 45076
rect 26700 45033 26709 45067
rect 26709 45033 26743 45067
rect 26743 45033 26752 45067
rect 26700 45024 26752 45033
rect 13636 44999 13688 45008
rect 13636 44965 13645 44999
rect 13645 44965 13679 44999
rect 13679 44965 13688 44999
rect 13636 44956 13688 44965
rect 19064 44956 19116 45008
rect 19984 44956 20036 45008
rect 21272 44956 21324 45008
rect 11796 44931 11848 44940
rect 11796 44897 11805 44931
rect 11805 44897 11839 44931
rect 11839 44897 11848 44931
rect 11796 44888 11848 44897
rect 13452 44931 13504 44940
rect 13452 44897 13461 44931
rect 13461 44897 13495 44931
rect 13495 44897 13504 44931
rect 13452 44888 13504 44897
rect 16672 44931 16724 44940
rect 16672 44897 16681 44931
rect 16681 44897 16715 44931
rect 16715 44897 16724 44931
rect 16672 44888 16724 44897
rect 17684 44931 17736 44940
rect 17684 44897 17693 44931
rect 17693 44897 17727 44931
rect 17727 44897 17736 44931
rect 17684 44888 17736 44897
rect 18052 44888 18104 44940
rect 18604 44888 18656 44940
rect 19432 44888 19484 44940
rect 21548 44888 21600 44940
rect 22192 44888 22244 44940
rect 23112 44956 23164 45008
rect 22560 44888 22612 44940
rect 26608 44956 26660 45008
rect 23572 44888 23624 44940
rect 25412 44931 25464 44940
rect 25412 44897 25421 44931
rect 25421 44897 25455 44931
rect 25455 44897 25464 44931
rect 25412 44888 25464 44897
rect 26056 44888 26108 44940
rect 26792 44931 26844 44940
rect 26792 44897 26801 44931
rect 26801 44897 26835 44931
rect 26835 44897 26844 44931
rect 26792 44888 26844 44897
rect 11980 44820 12032 44872
rect 18328 44820 18380 44872
rect 19708 44863 19760 44872
rect 19708 44829 19717 44863
rect 19717 44829 19751 44863
rect 19751 44829 19760 44863
rect 19708 44820 19760 44829
rect 20352 44820 20404 44872
rect 20904 44820 20956 44872
rect 21180 44863 21232 44872
rect 21180 44829 21189 44863
rect 21189 44829 21223 44863
rect 21223 44829 21232 44863
rect 21180 44820 21232 44829
rect 22100 44820 22152 44872
rect 17776 44795 17828 44804
rect 17776 44761 17785 44795
rect 17785 44761 17819 44795
rect 17819 44761 17828 44795
rect 17776 44752 17828 44761
rect 19800 44752 19852 44804
rect 20720 44752 20772 44804
rect 22468 44752 22520 44804
rect 23664 44820 23716 44872
rect 25136 44820 25188 44872
rect 26516 44863 26568 44872
rect 26516 44829 26525 44863
rect 26525 44829 26559 44863
rect 26559 44829 26568 44863
rect 26516 44820 26568 44829
rect 27068 44820 27120 44872
rect 1584 44684 1636 44736
rect 19156 44684 19208 44736
rect 19984 44684 20036 44736
rect 22284 44684 22336 44736
rect 26884 44684 26936 44736
rect 5982 44582 6034 44634
rect 6046 44582 6098 44634
rect 6110 44582 6162 44634
rect 6174 44582 6226 44634
rect 15982 44582 16034 44634
rect 16046 44582 16098 44634
rect 16110 44582 16162 44634
rect 16174 44582 16226 44634
rect 25982 44582 26034 44634
rect 26046 44582 26098 44634
rect 26110 44582 26162 44634
rect 26174 44582 26226 44634
rect 2964 44523 3016 44532
rect 2964 44489 2973 44523
rect 2973 44489 3007 44523
rect 3007 44489 3016 44523
rect 2964 44480 3016 44489
rect 11796 44480 11848 44532
rect 15568 44480 15620 44532
rect 12624 44412 12676 44464
rect 1584 44344 1636 44396
rect 1952 44276 2004 44328
rect 11520 44276 11572 44328
rect 12624 44319 12676 44328
rect 12624 44285 12630 44319
rect 12630 44285 12676 44319
rect 12624 44276 12676 44285
rect 10784 44183 10836 44192
rect 10784 44149 10793 44183
rect 10793 44149 10827 44183
rect 10827 44149 10836 44183
rect 10784 44140 10836 44149
rect 11796 44140 11848 44192
rect 13084 44183 13136 44192
rect 13084 44149 13093 44183
rect 13093 44149 13127 44183
rect 13127 44149 13136 44183
rect 13084 44140 13136 44149
rect 13452 44183 13504 44192
rect 13452 44149 13461 44183
rect 13461 44149 13495 44183
rect 13495 44149 13504 44183
rect 13452 44140 13504 44149
rect 13820 44276 13872 44328
rect 19800 44480 19852 44532
rect 17960 44412 18012 44464
rect 16672 44344 16724 44396
rect 17500 44344 17552 44396
rect 18328 44344 18380 44396
rect 20904 44480 20956 44532
rect 22468 44480 22520 44532
rect 23112 44523 23164 44532
rect 23112 44489 23121 44523
rect 23121 44489 23155 44523
rect 23155 44489 23164 44523
rect 23112 44480 23164 44489
rect 25136 44480 25188 44532
rect 16488 44276 16540 44328
rect 16580 44276 16632 44328
rect 18512 44319 18564 44328
rect 14004 44140 14056 44192
rect 16120 44183 16172 44192
rect 16120 44149 16129 44183
rect 16129 44149 16163 44183
rect 16163 44149 16172 44183
rect 16120 44140 16172 44149
rect 16672 44140 16724 44192
rect 16948 44140 17000 44192
rect 18512 44285 18521 44319
rect 18521 44285 18555 44319
rect 18555 44285 18564 44319
rect 18512 44276 18564 44285
rect 19340 44276 19392 44328
rect 20352 44412 20404 44464
rect 20444 44412 20496 44464
rect 24676 44412 24728 44464
rect 24768 44412 24820 44464
rect 25044 44412 25096 44464
rect 21180 44344 21232 44396
rect 24032 44344 24084 44396
rect 24216 44344 24268 44396
rect 24860 44387 24912 44396
rect 24860 44353 24869 44387
rect 24869 44353 24903 44387
rect 24903 44353 24912 44387
rect 24860 44344 24912 44353
rect 26424 44387 26476 44396
rect 26424 44353 26433 44387
rect 26433 44353 26467 44387
rect 26467 44353 26476 44387
rect 26424 44344 26476 44353
rect 20444 44276 20496 44328
rect 22100 44276 22152 44328
rect 22284 44276 22336 44328
rect 22560 44319 22612 44328
rect 22560 44285 22569 44319
rect 22569 44285 22603 44319
rect 22603 44285 22612 44319
rect 22560 44276 22612 44285
rect 22652 44276 22704 44328
rect 23848 44276 23900 44328
rect 24676 44276 24728 44328
rect 26608 44344 26660 44396
rect 26884 44344 26936 44396
rect 26700 44276 26752 44328
rect 21824 44208 21876 44260
rect 25136 44208 25188 44260
rect 17684 44140 17736 44192
rect 20076 44140 20128 44192
rect 22468 44140 22520 44192
rect 22652 44140 22704 44192
rect 23572 44140 23624 44192
rect 27712 44183 27764 44192
rect 27712 44149 27721 44183
rect 27721 44149 27755 44183
rect 27755 44149 27764 44183
rect 27712 44140 27764 44149
rect 10982 44038 11034 44090
rect 11046 44038 11098 44090
rect 11110 44038 11162 44090
rect 11174 44038 11226 44090
rect 20982 44038 21034 44090
rect 21046 44038 21098 44090
rect 21110 44038 21162 44090
rect 21174 44038 21226 44090
rect 16488 43936 16540 43988
rect 17500 43936 17552 43988
rect 1584 43800 1636 43852
rect 7564 43800 7616 43852
rect 8576 43843 8628 43852
rect 8576 43809 8585 43843
rect 8585 43809 8619 43843
rect 8619 43809 8628 43843
rect 8576 43800 8628 43809
rect 8760 43800 8812 43852
rect 11612 43800 11664 43852
rect 12256 43868 12308 43920
rect 17592 43868 17644 43920
rect 17960 43936 18012 43988
rect 19156 43936 19208 43988
rect 19892 43936 19944 43988
rect 23848 43979 23900 43988
rect 12072 43843 12124 43852
rect 12072 43809 12081 43843
rect 12081 43809 12115 43843
rect 12115 43809 12124 43843
rect 12072 43800 12124 43809
rect 13084 43843 13136 43852
rect 13084 43809 13093 43843
rect 13093 43809 13127 43843
rect 13127 43809 13136 43843
rect 13084 43800 13136 43809
rect 16304 43843 16356 43852
rect 16304 43809 16313 43843
rect 16313 43809 16347 43843
rect 16347 43809 16356 43843
rect 16304 43800 16356 43809
rect 16488 43800 16540 43852
rect 17684 43843 17736 43852
rect 17684 43809 17693 43843
rect 17693 43809 17727 43843
rect 17727 43809 17736 43843
rect 17684 43800 17736 43809
rect 17776 43843 17828 43852
rect 17776 43809 17785 43843
rect 17785 43809 17819 43843
rect 17819 43809 17828 43843
rect 18052 43868 18104 43920
rect 18696 43868 18748 43920
rect 23848 43945 23857 43979
rect 23857 43945 23891 43979
rect 23891 43945 23900 43979
rect 23848 43936 23900 43945
rect 25412 43936 25464 43988
rect 26700 43979 26752 43988
rect 26700 43945 26709 43979
rect 26709 43945 26743 43979
rect 26743 43945 26752 43979
rect 26700 43936 26752 43945
rect 26792 43979 26844 43988
rect 26792 43945 26801 43979
rect 26801 43945 26835 43979
rect 26835 43945 26844 43979
rect 26792 43936 26844 43945
rect 21640 43868 21692 43920
rect 17776 43800 17828 43809
rect 19892 43843 19944 43852
rect 19892 43809 19901 43843
rect 19901 43809 19935 43843
rect 19935 43809 19944 43843
rect 19892 43800 19944 43809
rect 21088 43843 21140 43852
rect 21088 43809 21097 43843
rect 21097 43809 21131 43843
rect 21131 43809 21140 43843
rect 21088 43800 21140 43809
rect 23480 43868 23532 43920
rect 26516 43911 26568 43920
rect 26516 43877 26525 43911
rect 26525 43877 26559 43911
rect 26559 43877 26568 43911
rect 26516 43868 26568 43877
rect 26884 43911 26936 43920
rect 26884 43877 26893 43911
rect 26893 43877 26927 43911
rect 26927 43877 26936 43911
rect 26884 43868 26936 43877
rect 22744 43843 22796 43852
rect 22744 43809 22753 43843
rect 22753 43809 22787 43843
rect 22787 43809 22796 43843
rect 22744 43800 22796 43809
rect 23112 43800 23164 43852
rect 26792 43800 26844 43852
rect 2228 43732 2280 43784
rect 3148 43775 3200 43784
rect 3148 43741 3157 43775
rect 3157 43741 3191 43775
rect 3191 43741 3200 43775
rect 3148 43732 3200 43741
rect 7748 43775 7800 43784
rect 7748 43741 7757 43775
rect 7757 43741 7791 43775
rect 7791 43741 7800 43775
rect 7748 43732 7800 43741
rect 11336 43732 11388 43784
rect 12624 43775 12676 43784
rect 10600 43664 10652 43716
rect 12624 43741 12633 43775
rect 12633 43741 12667 43775
rect 12667 43741 12676 43775
rect 12624 43732 12676 43741
rect 13176 43732 13228 43784
rect 18420 43775 18472 43784
rect 18420 43741 18429 43775
rect 18429 43741 18463 43775
rect 18463 43741 18472 43775
rect 18420 43732 18472 43741
rect 22192 43732 22244 43784
rect 23848 43732 23900 43784
rect 24124 43732 24176 43784
rect 25872 43732 25924 43784
rect 27252 43775 27304 43784
rect 27252 43741 27261 43775
rect 27261 43741 27295 43775
rect 27295 43741 27304 43775
rect 27252 43732 27304 43741
rect 13360 43664 13412 43716
rect 15752 43664 15804 43716
rect 16120 43707 16172 43716
rect 16120 43673 16129 43707
rect 16129 43673 16163 43707
rect 16163 43673 16172 43707
rect 16120 43664 16172 43673
rect 22376 43707 22428 43716
rect 22376 43673 22385 43707
rect 22385 43673 22419 43707
rect 22419 43673 22428 43707
rect 22376 43664 22428 43673
rect 13268 43639 13320 43648
rect 13268 43605 13277 43639
rect 13277 43605 13311 43639
rect 13311 43605 13320 43639
rect 13268 43596 13320 43605
rect 18604 43596 18656 43648
rect 19984 43596 20036 43648
rect 22100 43596 22152 43648
rect 22468 43596 22520 43648
rect 24676 43596 24728 43648
rect 27528 43639 27580 43648
rect 27528 43605 27537 43639
rect 27537 43605 27571 43639
rect 27571 43605 27580 43639
rect 27528 43596 27580 43605
rect 5982 43494 6034 43546
rect 6046 43494 6098 43546
rect 6110 43494 6162 43546
rect 6174 43494 6226 43546
rect 15982 43494 16034 43546
rect 16046 43494 16098 43546
rect 16110 43494 16162 43546
rect 16174 43494 16226 43546
rect 25982 43494 26034 43546
rect 26046 43494 26098 43546
rect 26110 43494 26162 43546
rect 26174 43494 26226 43546
rect 7748 43435 7800 43444
rect 7748 43401 7757 43435
rect 7757 43401 7791 43435
rect 7791 43401 7800 43435
rect 7748 43392 7800 43401
rect 8576 43392 8628 43444
rect 8760 43324 8812 43376
rect 9680 43324 9732 43376
rect 1768 43299 1820 43308
rect 1768 43265 1777 43299
rect 1777 43265 1811 43299
rect 1811 43265 1820 43299
rect 1768 43256 1820 43265
rect 1584 43188 1636 43240
rect 3148 43231 3200 43240
rect 3148 43197 3157 43231
rect 3157 43197 3191 43231
rect 3191 43197 3200 43231
rect 3148 43188 3200 43197
rect 11520 43392 11572 43444
rect 13084 43392 13136 43444
rect 15752 43392 15804 43444
rect 16304 43392 16356 43444
rect 17408 43392 17460 43444
rect 17684 43435 17736 43444
rect 17684 43401 17693 43435
rect 17693 43401 17727 43435
rect 17727 43401 17736 43435
rect 17684 43392 17736 43401
rect 19432 43435 19484 43444
rect 19432 43401 19441 43435
rect 19441 43401 19475 43435
rect 19475 43401 19484 43435
rect 19432 43392 19484 43401
rect 21088 43392 21140 43444
rect 22928 43392 22980 43444
rect 16488 43324 16540 43376
rect 19156 43324 19208 43376
rect 20076 43367 20128 43376
rect 20076 43333 20085 43367
rect 20085 43333 20119 43367
rect 20119 43333 20128 43367
rect 20076 43324 20128 43333
rect 13820 43299 13872 43308
rect 13820 43265 13829 43299
rect 13829 43265 13863 43299
rect 13863 43265 13872 43299
rect 13820 43256 13872 43265
rect 17684 43256 17736 43308
rect 18052 43299 18104 43308
rect 18052 43265 18061 43299
rect 18061 43265 18095 43299
rect 18095 43265 18104 43299
rect 18052 43256 18104 43265
rect 20720 43256 20772 43308
rect 21272 43256 21324 43308
rect 12072 43188 12124 43240
rect 12992 43231 13044 43240
rect 12992 43197 13001 43231
rect 13001 43197 13035 43231
rect 13035 43197 13044 43231
rect 12992 43188 13044 43197
rect 13360 43231 13412 43240
rect 13360 43197 13369 43231
rect 13369 43197 13403 43231
rect 13403 43197 13412 43231
rect 13360 43188 13412 43197
rect 13728 43231 13780 43240
rect 13728 43197 13737 43231
rect 13737 43197 13771 43231
rect 13771 43197 13780 43231
rect 13728 43188 13780 43197
rect 17040 43188 17092 43240
rect 17776 43188 17828 43240
rect 18972 43188 19024 43240
rect 19984 43188 20036 43240
rect 22744 43256 22796 43308
rect 23664 43392 23716 43444
rect 24124 43392 24176 43444
rect 25780 43392 25832 43444
rect 26516 43435 26568 43444
rect 26516 43401 26525 43435
rect 26525 43401 26559 43435
rect 26559 43401 26568 43435
rect 26516 43392 26568 43401
rect 26700 43392 26752 43444
rect 27344 43435 27396 43444
rect 27344 43401 27353 43435
rect 27353 43401 27387 43435
rect 27387 43401 27396 43435
rect 27344 43392 27396 43401
rect 23480 43367 23532 43376
rect 23480 43333 23489 43367
rect 23489 43333 23523 43367
rect 23523 43333 23532 43367
rect 23480 43324 23532 43333
rect 26884 43324 26936 43376
rect 27528 43256 27580 43308
rect 19432 43120 19484 43172
rect 10600 43095 10652 43104
rect 10600 43061 10609 43095
rect 10609 43061 10643 43095
rect 10643 43061 10652 43095
rect 10600 43052 10652 43061
rect 20720 43120 20772 43172
rect 23848 43188 23900 43240
rect 24860 43231 24912 43240
rect 24860 43197 24869 43231
rect 24869 43197 24903 43231
rect 24903 43197 24912 43231
rect 24860 43188 24912 43197
rect 26332 43188 26384 43240
rect 10982 42950 11034 43002
rect 11046 42950 11098 43002
rect 11110 42950 11162 43002
rect 11174 42950 11226 43002
rect 20982 42950 21034 43002
rect 21046 42950 21098 43002
rect 21110 42950 21162 43002
rect 21174 42950 21226 43002
rect 1768 42848 1820 42900
rect 11336 42848 11388 42900
rect 17040 42891 17092 42900
rect 1584 42780 1636 42832
rect 10232 42712 10284 42764
rect 11612 42712 11664 42764
rect 12072 42755 12124 42764
rect 12072 42721 12081 42755
rect 12081 42721 12115 42755
rect 12115 42721 12124 42755
rect 12072 42712 12124 42721
rect 11980 42687 12032 42696
rect 11980 42653 11989 42687
rect 11989 42653 12023 42687
rect 12023 42653 12032 42687
rect 11980 42644 12032 42653
rect 17040 42857 17049 42891
rect 17049 42857 17083 42891
rect 17083 42857 17092 42891
rect 17040 42848 17092 42857
rect 17500 42891 17552 42900
rect 17500 42857 17509 42891
rect 17509 42857 17543 42891
rect 17543 42857 17552 42891
rect 17500 42848 17552 42857
rect 21272 42848 21324 42900
rect 26792 42848 26844 42900
rect 12440 42755 12492 42764
rect 12440 42721 12449 42755
rect 12449 42721 12483 42755
rect 12483 42721 12492 42755
rect 13820 42780 13872 42832
rect 21732 42780 21784 42832
rect 22928 42780 22980 42832
rect 23112 42780 23164 42832
rect 12440 42712 12492 42721
rect 17684 42712 17736 42764
rect 19156 42712 19208 42764
rect 19708 42712 19760 42764
rect 20076 42712 20128 42764
rect 20444 42712 20496 42764
rect 22284 42755 22336 42764
rect 22284 42721 22293 42755
rect 22293 42721 22327 42755
rect 22327 42721 22336 42755
rect 22284 42712 22336 42721
rect 22652 42755 22704 42764
rect 22652 42721 22661 42755
rect 22661 42721 22695 42755
rect 22695 42721 22704 42755
rect 22652 42712 22704 42721
rect 22744 42755 22796 42764
rect 22744 42721 22753 42755
rect 22753 42721 22787 42755
rect 22787 42721 22796 42755
rect 22744 42712 22796 42721
rect 23848 42712 23900 42764
rect 18328 42644 18380 42696
rect 22192 42644 22244 42696
rect 22468 42644 22520 42696
rect 24584 42712 24636 42764
rect 25596 42712 25648 42764
rect 26608 42755 26660 42764
rect 26608 42721 26617 42755
rect 26617 42721 26651 42755
rect 26651 42721 26660 42755
rect 26608 42712 26660 42721
rect 25780 42644 25832 42696
rect 19892 42576 19944 42628
rect 20444 42576 20496 42628
rect 2228 42508 2280 42560
rect 10232 42508 10284 42560
rect 12992 42551 13044 42560
rect 12992 42517 13001 42551
rect 13001 42517 13035 42551
rect 13035 42517 13044 42551
rect 12992 42508 13044 42517
rect 18972 42551 19024 42560
rect 18972 42517 18981 42551
rect 18981 42517 19015 42551
rect 19015 42517 19024 42551
rect 18972 42508 19024 42517
rect 22284 42508 22336 42560
rect 22560 42508 22612 42560
rect 23572 42508 23624 42560
rect 24308 42508 24360 42560
rect 25136 42508 25188 42560
rect 26792 42551 26844 42560
rect 26792 42517 26801 42551
rect 26801 42517 26835 42551
rect 26835 42517 26844 42551
rect 26792 42508 26844 42517
rect 5982 42406 6034 42458
rect 6046 42406 6098 42458
rect 6110 42406 6162 42458
rect 6174 42406 6226 42458
rect 15982 42406 16034 42458
rect 16046 42406 16098 42458
rect 16110 42406 16162 42458
rect 16174 42406 16226 42458
rect 25982 42406 26034 42458
rect 26046 42406 26098 42458
rect 26110 42406 26162 42458
rect 26174 42406 26226 42458
rect 1584 42347 1636 42356
rect 1584 42313 1593 42347
rect 1593 42313 1627 42347
rect 1627 42313 1636 42347
rect 1584 42304 1636 42313
rect 11336 42304 11388 42356
rect 8944 42143 8996 42152
rect 8944 42109 8953 42143
rect 8953 42109 8987 42143
rect 8987 42109 8996 42143
rect 8944 42100 8996 42109
rect 9220 42143 9272 42152
rect 9220 42109 9229 42143
rect 9229 42109 9263 42143
rect 9263 42109 9272 42143
rect 9220 42100 9272 42109
rect 9588 42143 9640 42152
rect 9588 42109 9597 42143
rect 9597 42109 9631 42143
rect 9631 42109 9640 42143
rect 9588 42100 9640 42109
rect 10048 42143 10100 42152
rect 10048 42109 10057 42143
rect 10057 42109 10091 42143
rect 10091 42109 10100 42143
rect 10048 42100 10100 42109
rect 10232 42143 10284 42152
rect 10232 42109 10241 42143
rect 10241 42109 10275 42143
rect 10275 42109 10284 42143
rect 10232 42100 10284 42109
rect 11980 42304 12032 42356
rect 12992 42304 13044 42356
rect 17776 42347 17828 42356
rect 17776 42313 17785 42347
rect 17785 42313 17819 42347
rect 17819 42313 17828 42347
rect 17776 42304 17828 42313
rect 18328 42347 18380 42356
rect 18328 42313 18337 42347
rect 18337 42313 18371 42347
rect 18371 42313 18380 42347
rect 18328 42304 18380 42313
rect 19708 42304 19760 42356
rect 20720 42304 20772 42356
rect 17684 42236 17736 42288
rect 18880 42279 18932 42288
rect 18880 42245 18889 42279
rect 18889 42245 18923 42279
rect 18923 42245 18932 42279
rect 18880 42236 18932 42245
rect 19892 42236 19944 42288
rect 20444 42236 20496 42288
rect 21272 42304 21324 42356
rect 21640 42304 21692 42356
rect 22192 42236 22244 42288
rect 23020 42236 23072 42288
rect 24768 42236 24820 42288
rect 9036 42032 9088 42084
rect 12440 42032 12492 42084
rect 18420 42100 18472 42152
rect 20076 42100 20128 42152
rect 15108 42075 15160 42084
rect 15108 42041 15117 42075
rect 15117 42041 15151 42075
rect 15151 42041 15160 42075
rect 15108 42032 15160 42041
rect 19340 42032 19392 42084
rect 11520 42007 11572 42016
rect 11520 41973 11529 42007
rect 11529 41973 11563 42007
rect 11563 41973 11572 42007
rect 11520 41964 11572 41973
rect 11612 41964 11664 42016
rect 12072 41964 12124 42016
rect 14004 42007 14056 42016
rect 14004 41973 14013 42007
rect 14013 41973 14047 42007
rect 14047 41973 14056 42007
rect 14004 41964 14056 41973
rect 21640 42168 21692 42220
rect 26792 42304 26844 42356
rect 25596 42279 25648 42288
rect 25596 42245 25605 42279
rect 25605 42245 25639 42279
rect 25639 42245 25648 42279
rect 25596 42236 25648 42245
rect 25964 42279 26016 42288
rect 25964 42245 25973 42279
rect 25973 42245 26007 42279
rect 26007 42245 26016 42279
rect 25964 42236 26016 42245
rect 21824 42100 21876 42152
rect 22192 42032 22244 42084
rect 22376 42143 22428 42152
rect 22376 42109 22385 42143
rect 22385 42109 22419 42143
rect 22419 42109 22428 42143
rect 25872 42168 25924 42220
rect 26332 42168 26384 42220
rect 26516 42168 26568 42220
rect 22376 42100 22428 42109
rect 24308 42143 24360 42152
rect 24308 42109 24317 42143
rect 24317 42109 24351 42143
rect 24351 42109 24360 42143
rect 24308 42100 24360 42109
rect 22652 42032 22704 42084
rect 25872 42032 25924 42084
rect 27528 42100 27580 42152
rect 22100 41964 22152 42016
rect 22468 41964 22520 42016
rect 23296 41964 23348 42016
rect 27160 41964 27212 42016
rect 10982 41862 11034 41914
rect 11046 41862 11098 41914
rect 11110 41862 11162 41914
rect 11174 41862 11226 41914
rect 20982 41862 21034 41914
rect 21046 41862 21098 41914
rect 21110 41862 21162 41914
rect 21174 41862 21226 41914
rect 10048 41760 10100 41812
rect 17408 41760 17460 41812
rect 17684 41803 17736 41812
rect 17684 41769 17693 41803
rect 17693 41769 17727 41803
rect 17727 41769 17736 41803
rect 17684 41760 17736 41769
rect 18972 41760 19024 41812
rect 19340 41760 19392 41812
rect 19892 41760 19944 41812
rect 20352 41803 20404 41812
rect 20352 41769 20361 41803
rect 20361 41769 20395 41803
rect 20395 41769 20404 41803
rect 20352 41760 20404 41769
rect 21824 41803 21876 41812
rect 21824 41769 21833 41803
rect 21833 41769 21867 41803
rect 21867 41769 21876 41803
rect 21824 41760 21876 41769
rect 22468 41760 22520 41812
rect 22744 41760 22796 41812
rect 24584 41760 24636 41812
rect 25780 41760 25832 41812
rect 26332 41760 26384 41812
rect 27528 41803 27580 41812
rect 27528 41769 27537 41803
rect 27537 41769 27571 41803
rect 27571 41769 27580 41803
rect 27528 41760 27580 41769
rect 11428 41692 11480 41744
rect 20720 41735 20772 41744
rect 20720 41701 20729 41735
rect 20729 41701 20763 41735
rect 20763 41701 20772 41735
rect 20720 41692 20772 41701
rect 22376 41692 22428 41744
rect 26516 41735 26568 41744
rect 26516 41701 26525 41735
rect 26525 41701 26559 41735
rect 26559 41701 26568 41735
rect 26516 41692 26568 41701
rect 10784 41556 10836 41608
rect 10876 41488 10928 41540
rect 19432 41624 19484 41676
rect 19984 41624 20036 41676
rect 11796 41556 11848 41608
rect 12348 41488 12400 41540
rect 19156 41488 19208 41540
rect 21272 41624 21324 41676
rect 22560 41667 22612 41676
rect 22560 41633 22569 41667
rect 22569 41633 22603 41667
rect 22603 41633 22612 41667
rect 22560 41624 22612 41633
rect 23020 41624 23072 41676
rect 24584 41624 24636 41676
rect 27160 41667 27212 41676
rect 27160 41633 27169 41667
rect 27169 41633 27203 41667
rect 27203 41633 27212 41667
rect 27160 41624 27212 41633
rect 22008 41556 22060 41608
rect 23204 41599 23256 41608
rect 23204 41565 23213 41599
rect 23213 41565 23247 41599
rect 23247 41565 23256 41599
rect 23204 41556 23256 41565
rect 22468 41488 22520 41540
rect 24400 41599 24452 41608
rect 24400 41565 24409 41599
rect 24409 41565 24443 41599
rect 24443 41565 24452 41599
rect 24400 41556 24452 41565
rect 24676 41556 24728 41608
rect 25044 41488 25096 41540
rect 9036 41463 9088 41472
rect 9036 41429 9045 41463
rect 9045 41429 9079 41463
rect 9079 41429 9088 41463
rect 9036 41420 9088 41429
rect 11336 41420 11388 41472
rect 15660 41420 15712 41472
rect 23572 41420 23624 41472
rect 5982 41318 6034 41370
rect 6046 41318 6098 41370
rect 6110 41318 6162 41370
rect 6174 41318 6226 41370
rect 15982 41318 16034 41370
rect 16046 41318 16098 41370
rect 16110 41318 16162 41370
rect 16174 41318 16226 41370
rect 25982 41318 26034 41370
rect 26046 41318 26098 41370
rect 26110 41318 26162 41370
rect 26174 41318 26226 41370
rect 11796 41259 11848 41268
rect 11796 41225 11805 41259
rect 11805 41225 11839 41259
rect 11839 41225 11848 41259
rect 11796 41216 11848 41225
rect 12532 41216 12584 41268
rect 19800 41259 19852 41268
rect 19800 41225 19809 41259
rect 19809 41225 19843 41259
rect 19843 41225 19852 41259
rect 19800 41216 19852 41225
rect 19984 41216 20036 41268
rect 22468 41259 22520 41268
rect 22468 41225 22477 41259
rect 22477 41225 22511 41259
rect 22511 41225 22520 41259
rect 22468 41216 22520 41225
rect 23020 41216 23072 41268
rect 26884 41216 26936 41268
rect 10048 41148 10100 41200
rect 16488 41148 16540 41200
rect 10692 41055 10744 41064
rect 10692 41021 10701 41055
rect 10701 41021 10735 41055
rect 10735 41021 10744 41055
rect 10692 41012 10744 41021
rect 10876 41012 10928 41064
rect 15660 41080 15712 41132
rect 11520 41012 11572 41064
rect 11704 41012 11756 41064
rect 16580 41055 16632 41064
rect 16580 41021 16589 41055
rect 16589 41021 16623 41055
rect 16623 41021 16632 41055
rect 16580 41012 16632 41021
rect 16948 41055 17000 41064
rect 16948 41021 16957 41055
rect 16957 41021 16991 41055
rect 16991 41021 17000 41055
rect 16948 41012 17000 41021
rect 19708 41148 19760 41200
rect 21640 41148 21692 41200
rect 21916 41148 21968 41200
rect 21180 41123 21232 41132
rect 21180 41089 21189 41123
rect 21189 41089 21223 41123
rect 21223 41089 21232 41123
rect 21180 41080 21232 41089
rect 27160 41148 27212 41200
rect 21548 41012 21600 41064
rect 21640 41012 21692 41064
rect 21824 41012 21876 41064
rect 23664 41012 23716 41064
rect 15752 40944 15804 40996
rect 24308 40944 24360 40996
rect 24676 40944 24728 40996
rect 10140 40919 10192 40928
rect 10140 40885 10149 40919
rect 10149 40885 10183 40919
rect 10183 40885 10192 40919
rect 10140 40876 10192 40885
rect 12072 40919 12124 40928
rect 12072 40885 12081 40919
rect 12081 40885 12115 40919
rect 12115 40885 12124 40919
rect 12072 40876 12124 40885
rect 12440 40876 12492 40928
rect 12808 40876 12860 40928
rect 13084 40919 13136 40928
rect 13084 40885 13093 40919
rect 13093 40885 13127 40919
rect 13127 40885 13136 40919
rect 13084 40876 13136 40885
rect 23940 40919 23992 40928
rect 23940 40885 23949 40919
rect 23949 40885 23983 40919
rect 23983 40885 23992 40919
rect 23940 40876 23992 40885
rect 25320 41012 25372 41064
rect 25872 40876 25924 40928
rect 10982 40774 11034 40826
rect 11046 40774 11098 40826
rect 11110 40774 11162 40826
rect 11174 40774 11226 40826
rect 20982 40774 21034 40826
rect 21046 40774 21098 40826
rect 21110 40774 21162 40826
rect 21174 40774 21226 40826
rect 10784 40672 10836 40724
rect 21272 40672 21324 40724
rect 21548 40715 21600 40724
rect 21548 40681 21557 40715
rect 21557 40681 21591 40715
rect 21591 40681 21600 40715
rect 21548 40672 21600 40681
rect 22008 40672 22060 40724
rect 23204 40672 23256 40724
rect 25044 40715 25096 40724
rect 25044 40681 25053 40715
rect 25053 40681 25087 40715
rect 25087 40681 25096 40715
rect 25044 40672 25096 40681
rect 25872 40672 25924 40724
rect 10508 40536 10560 40588
rect 12072 40579 12124 40588
rect 12072 40545 12081 40579
rect 12081 40545 12115 40579
rect 12115 40545 12124 40579
rect 12072 40536 12124 40545
rect 12348 40536 12400 40588
rect 13084 40604 13136 40656
rect 16764 40604 16816 40656
rect 22560 40647 22612 40656
rect 22560 40613 22569 40647
rect 22569 40613 22603 40647
rect 22603 40613 22612 40647
rect 22560 40604 22612 40613
rect 14188 40536 14240 40588
rect 20996 40579 21048 40588
rect 10232 40468 10284 40520
rect 11980 40511 12032 40520
rect 1492 40332 1544 40384
rect 10048 40332 10100 40384
rect 11980 40477 11989 40511
rect 11989 40477 12023 40511
rect 12023 40477 12032 40511
rect 11980 40468 12032 40477
rect 12532 40511 12584 40520
rect 12532 40477 12541 40511
rect 12541 40477 12575 40511
rect 12575 40477 12584 40511
rect 12532 40468 12584 40477
rect 20996 40545 21005 40579
rect 21005 40545 21039 40579
rect 21039 40545 21048 40579
rect 20996 40536 21048 40545
rect 21640 40536 21692 40588
rect 22192 40536 22244 40588
rect 24492 40536 24544 40588
rect 25136 40536 25188 40588
rect 17224 40468 17276 40520
rect 17408 40468 17460 40520
rect 11796 40400 11848 40452
rect 16580 40400 16632 40452
rect 23296 40468 23348 40520
rect 24584 40400 24636 40452
rect 11520 40375 11572 40384
rect 11520 40341 11529 40375
rect 11529 40341 11563 40375
rect 11563 40341 11572 40375
rect 11520 40332 11572 40341
rect 12900 40375 12952 40384
rect 12900 40341 12909 40375
rect 12909 40341 12943 40375
rect 12943 40341 12952 40375
rect 12900 40332 12952 40341
rect 12992 40332 13044 40384
rect 13912 40332 13964 40384
rect 15660 40375 15712 40384
rect 15660 40341 15669 40375
rect 15669 40341 15703 40375
rect 15703 40341 15712 40375
rect 15660 40332 15712 40341
rect 18144 40375 18196 40384
rect 18144 40341 18153 40375
rect 18153 40341 18187 40375
rect 18187 40341 18196 40375
rect 18144 40332 18196 40341
rect 24124 40332 24176 40384
rect 5982 40230 6034 40282
rect 6046 40230 6098 40282
rect 6110 40230 6162 40282
rect 6174 40230 6226 40282
rect 15982 40230 16034 40282
rect 16046 40230 16098 40282
rect 16110 40230 16162 40282
rect 16174 40230 16226 40282
rect 25982 40230 26034 40282
rect 26046 40230 26098 40282
rect 26110 40230 26162 40282
rect 26174 40230 26226 40282
rect 11704 40128 11756 40180
rect 12532 40128 12584 40180
rect 15108 40171 15160 40180
rect 15108 40137 15117 40171
rect 15117 40137 15151 40171
rect 15151 40137 15160 40171
rect 15108 40128 15160 40137
rect 16764 40128 16816 40180
rect 21640 40128 21692 40180
rect 10232 40060 10284 40112
rect 1768 40035 1820 40044
rect 1768 40001 1777 40035
rect 1777 40001 1811 40035
rect 1811 40001 1820 40035
rect 1768 39992 1820 40001
rect 9956 40035 10008 40044
rect 9956 40001 9965 40035
rect 9965 40001 9999 40035
rect 9999 40001 10008 40035
rect 9956 39992 10008 40001
rect 1492 39967 1544 39976
rect 1492 39933 1501 39967
rect 1501 39933 1535 39967
rect 1535 39933 1544 39967
rect 1492 39924 1544 39933
rect 10968 39992 11020 40044
rect 11980 40060 12032 40112
rect 23756 40060 23808 40112
rect 11704 39992 11756 40044
rect 15936 40035 15988 40044
rect 15936 40001 15945 40035
rect 15945 40001 15979 40035
rect 15979 40001 15988 40035
rect 15936 39992 15988 40001
rect 10876 39967 10928 39976
rect 3148 39899 3200 39908
rect 3148 39865 3157 39899
rect 3157 39865 3191 39899
rect 3191 39865 3200 39899
rect 3148 39856 3200 39865
rect 9680 39856 9732 39908
rect 10876 39933 10885 39967
rect 10885 39933 10919 39967
rect 10919 39933 10928 39967
rect 10876 39924 10928 39933
rect 12072 39924 12124 39976
rect 14188 39924 14240 39976
rect 17224 39924 17276 39976
rect 22008 39967 22060 39976
rect 22008 39933 22017 39967
rect 22017 39933 22051 39967
rect 22051 39933 22060 39967
rect 22008 39924 22060 39933
rect 22284 39924 22336 39976
rect 24584 39992 24636 40044
rect 25136 40035 25188 40044
rect 25136 40001 25145 40035
rect 25145 40001 25179 40035
rect 25179 40001 25188 40035
rect 25136 39992 25188 40001
rect 11980 39788 12032 39840
rect 12624 39831 12676 39840
rect 12624 39797 12633 39831
rect 12633 39797 12667 39831
rect 12667 39797 12676 39831
rect 12624 39788 12676 39797
rect 13636 39831 13688 39840
rect 13636 39797 13645 39831
rect 13645 39797 13679 39831
rect 13679 39797 13688 39831
rect 20996 39856 21048 39908
rect 22376 39856 22428 39908
rect 23480 39899 23532 39908
rect 23480 39865 23489 39899
rect 23489 39865 23523 39899
rect 23523 39865 23532 39899
rect 23480 39856 23532 39865
rect 13636 39788 13688 39797
rect 16764 39788 16816 39840
rect 21732 39788 21784 39840
rect 22560 39788 22612 39840
rect 23296 39788 23348 39840
rect 23664 39788 23716 39840
rect 24492 39856 24544 39908
rect 24584 39788 24636 39840
rect 10982 39686 11034 39738
rect 11046 39686 11098 39738
rect 11110 39686 11162 39738
rect 11174 39686 11226 39738
rect 20982 39686 21034 39738
rect 21046 39686 21098 39738
rect 21110 39686 21162 39738
rect 21174 39686 21226 39738
rect 1768 39584 1820 39636
rect 10508 39627 10560 39636
rect 10508 39593 10517 39627
rect 10517 39593 10551 39627
rect 10551 39593 10560 39627
rect 10508 39584 10560 39593
rect 16856 39584 16908 39636
rect 17316 39584 17368 39636
rect 19432 39627 19484 39636
rect 19432 39593 19441 39627
rect 19441 39593 19475 39627
rect 19475 39593 19484 39627
rect 19432 39584 19484 39593
rect 21548 39584 21600 39636
rect 22192 39584 22244 39636
rect 24492 39627 24544 39636
rect 24492 39593 24501 39627
rect 24501 39593 24535 39627
rect 24535 39593 24544 39627
rect 24492 39584 24544 39593
rect 24676 39584 24728 39636
rect 12164 39516 12216 39568
rect 21916 39516 21968 39568
rect 11520 39448 11572 39500
rect 11796 39491 11848 39500
rect 11796 39457 11805 39491
rect 11805 39457 11839 39491
rect 11839 39457 11848 39491
rect 11796 39448 11848 39457
rect 10876 39380 10928 39432
rect 12348 39380 12400 39432
rect 12992 39491 13044 39500
rect 12992 39457 13001 39491
rect 13001 39457 13035 39491
rect 13035 39457 13044 39491
rect 13544 39491 13596 39500
rect 12992 39448 13044 39457
rect 13544 39457 13553 39491
rect 13553 39457 13587 39491
rect 13587 39457 13596 39491
rect 13544 39448 13596 39457
rect 13728 39491 13780 39500
rect 13728 39457 13737 39491
rect 13737 39457 13771 39491
rect 13771 39457 13780 39491
rect 13728 39448 13780 39457
rect 15292 39491 15344 39500
rect 15292 39457 15301 39491
rect 15301 39457 15335 39491
rect 15335 39457 15344 39491
rect 15292 39448 15344 39457
rect 16764 39491 16816 39500
rect 16764 39457 16773 39491
rect 16773 39457 16807 39491
rect 16807 39457 16816 39491
rect 16764 39448 16816 39457
rect 21548 39491 21600 39500
rect 21548 39457 21557 39491
rect 21557 39457 21591 39491
rect 21591 39457 21600 39491
rect 21548 39448 21600 39457
rect 21732 39491 21784 39500
rect 21732 39457 21741 39491
rect 21741 39457 21775 39491
rect 21775 39457 21784 39491
rect 21732 39448 21784 39457
rect 23664 39448 23716 39500
rect 24584 39491 24636 39500
rect 14096 39423 14148 39432
rect 14096 39389 14105 39423
rect 14105 39389 14139 39423
rect 14139 39389 14148 39423
rect 14096 39380 14148 39389
rect 16672 39423 16724 39432
rect 16672 39389 16681 39423
rect 16681 39389 16715 39423
rect 16715 39389 16724 39423
rect 16672 39380 16724 39389
rect 17040 39380 17092 39432
rect 17224 39380 17276 39432
rect 18052 39423 18104 39432
rect 18052 39389 18061 39423
rect 18061 39389 18095 39423
rect 18095 39389 18104 39423
rect 18052 39380 18104 39389
rect 18328 39423 18380 39432
rect 18328 39389 18337 39423
rect 18337 39389 18371 39423
rect 18371 39389 18380 39423
rect 18328 39380 18380 39389
rect 13084 39312 13136 39364
rect 10048 39287 10100 39296
rect 10048 39253 10057 39287
rect 10057 39253 10091 39287
rect 10091 39253 10100 39287
rect 10048 39244 10100 39253
rect 10784 39287 10836 39296
rect 10784 39253 10793 39287
rect 10793 39253 10827 39287
rect 10827 39253 10836 39287
rect 10784 39244 10836 39253
rect 11980 39244 12032 39296
rect 12164 39244 12216 39296
rect 12808 39244 12860 39296
rect 13820 39244 13872 39296
rect 15016 39244 15068 39296
rect 15752 39287 15804 39296
rect 15752 39253 15761 39287
rect 15761 39253 15795 39287
rect 15795 39253 15804 39287
rect 15752 39244 15804 39253
rect 16396 39244 16448 39296
rect 16580 39244 16632 39296
rect 22008 39244 22060 39296
rect 23480 39244 23532 39296
rect 24584 39457 24593 39491
rect 24593 39457 24627 39491
rect 24627 39457 24636 39491
rect 24584 39448 24636 39457
rect 5982 39142 6034 39194
rect 6046 39142 6098 39194
rect 6110 39142 6162 39194
rect 6174 39142 6226 39194
rect 15982 39142 16034 39194
rect 16046 39142 16098 39194
rect 16110 39142 16162 39194
rect 16174 39142 16226 39194
rect 25982 39142 26034 39194
rect 26046 39142 26098 39194
rect 26110 39142 26162 39194
rect 26174 39142 26226 39194
rect 3332 39040 3384 39092
rect 12440 39040 12492 39092
rect 14096 39040 14148 39092
rect 16764 39040 16816 39092
rect 18328 39040 18380 39092
rect 21732 39040 21784 39092
rect 23664 39040 23716 39092
rect 24492 39040 24544 39092
rect 1492 38904 1544 38956
rect 1768 38904 1820 38956
rect 1676 38836 1728 38888
rect 8852 38836 8904 38888
rect 21548 39015 21600 39024
rect 21548 38981 21557 39015
rect 21557 38981 21591 39015
rect 21591 38981 21600 39015
rect 21548 38972 21600 38981
rect 10140 38947 10192 38956
rect 10140 38913 10149 38947
rect 10149 38913 10183 38947
rect 10183 38913 10192 38947
rect 10140 38904 10192 38913
rect 9772 38768 9824 38820
rect 9312 38700 9364 38752
rect 9496 38743 9548 38752
rect 9496 38709 9505 38743
rect 9505 38709 9539 38743
rect 9539 38709 9548 38743
rect 11336 38836 11388 38888
rect 12164 38836 12216 38888
rect 12624 38879 12676 38888
rect 12624 38845 12633 38879
rect 12633 38845 12667 38879
rect 12667 38845 12676 38879
rect 12624 38836 12676 38845
rect 12716 38879 12768 38888
rect 12716 38845 12725 38879
rect 12725 38845 12759 38879
rect 12759 38845 12768 38879
rect 12716 38836 12768 38845
rect 12900 38836 12952 38888
rect 13544 38879 13596 38888
rect 13544 38845 13553 38879
rect 13553 38845 13587 38879
rect 13587 38845 13596 38879
rect 13544 38836 13596 38845
rect 15292 38904 15344 38956
rect 15660 38904 15712 38956
rect 17776 38904 17828 38956
rect 14924 38836 14976 38888
rect 16396 38836 16448 38888
rect 18052 38879 18104 38888
rect 18052 38845 18061 38879
rect 18061 38845 18095 38879
rect 18095 38845 18104 38879
rect 18052 38836 18104 38845
rect 18420 38836 18472 38888
rect 21180 38836 21232 38888
rect 21548 38836 21600 38888
rect 21916 38836 21968 38888
rect 22376 38904 22428 38956
rect 22560 38879 22612 38888
rect 15108 38768 15160 38820
rect 15292 38768 15344 38820
rect 22560 38845 22569 38879
rect 22569 38845 22603 38879
rect 22603 38845 22612 38879
rect 22560 38836 22612 38845
rect 25780 38836 25832 38888
rect 26148 38879 26200 38888
rect 26148 38845 26157 38879
rect 26157 38845 26191 38879
rect 26191 38845 26200 38879
rect 26148 38836 26200 38845
rect 26424 38879 26476 38888
rect 26424 38845 26433 38879
rect 26433 38845 26467 38879
rect 26467 38845 26476 38879
rect 26424 38836 26476 38845
rect 9496 38700 9548 38709
rect 10048 38700 10100 38752
rect 10876 38700 10928 38752
rect 12164 38743 12216 38752
rect 12164 38709 12173 38743
rect 12173 38709 12207 38743
rect 12207 38709 12216 38743
rect 12164 38700 12216 38709
rect 14188 38700 14240 38752
rect 15476 38700 15528 38752
rect 15660 38700 15712 38752
rect 17040 38700 17092 38752
rect 23480 38700 23532 38752
rect 10982 38598 11034 38650
rect 11046 38598 11098 38650
rect 11110 38598 11162 38650
rect 11174 38598 11226 38650
rect 20982 38598 21034 38650
rect 21046 38598 21098 38650
rect 21110 38598 21162 38650
rect 21174 38598 21226 38650
rect 9312 38428 9364 38480
rect 9680 38471 9732 38480
rect 9680 38437 9689 38471
rect 9689 38437 9723 38471
rect 9723 38437 9732 38471
rect 9680 38428 9732 38437
rect 11336 38496 11388 38548
rect 16488 38539 16540 38548
rect 16488 38505 16497 38539
rect 16497 38505 16531 38539
rect 16531 38505 16540 38539
rect 16488 38496 16540 38505
rect 18328 38496 18380 38548
rect 20720 38496 20772 38548
rect 26148 38539 26200 38548
rect 26148 38505 26157 38539
rect 26157 38505 26191 38539
rect 26191 38505 26200 38539
rect 26148 38496 26200 38505
rect 12164 38428 12216 38480
rect 15108 38428 15160 38480
rect 8576 38403 8628 38412
rect 8576 38369 8585 38403
rect 8585 38369 8619 38403
rect 8619 38369 8628 38403
rect 8576 38360 8628 38369
rect 8760 38360 8812 38412
rect 9404 38360 9456 38412
rect 10232 38360 10284 38412
rect 10508 38360 10560 38412
rect 10876 38403 10928 38412
rect 10876 38369 10885 38403
rect 10885 38369 10919 38403
rect 10919 38369 10928 38403
rect 10876 38360 10928 38369
rect 12808 38360 12860 38412
rect 13544 38360 13596 38412
rect 14648 38403 14700 38412
rect 14648 38369 14657 38403
rect 14657 38369 14691 38403
rect 14691 38369 14700 38403
rect 14648 38360 14700 38369
rect 16396 38428 16448 38480
rect 9680 38292 9732 38344
rect 10600 38292 10652 38344
rect 12532 38335 12584 38344
rect 12532 38301 12541 38335
rect 12541 38301 12575 38335
rect 12575 38301 12584 38335
rect 12532 38292 12584 38301
rect 15016 38292 15068 38344
rect 16580 38360 16632 38412
rect 16488 38292 16540 38344
rect 16856 38292 16908 38344
rect 1400 38224 1452 38276
rect 1860 38224 1912 38276
rect 8300 38224 8352 38276
rect 11428 38224 11480 38276
rect 12348 38224 12400 38276
rect 14464 38224 14516 38276
rect 15108 38224 15160 38276
rect 15752 38224 15804 38276
rect 16304 38224 16356 38276
rect 1584 38199 1636 38208
rect 1584 38165 1593 38199
rect 1593 38165 1627 38199
rect 1627 38165 1636 38199
rect 1584 38156 1636 38165
rect 11520 38199 11572 38208
rect 11520 38165 11529 38199
rect 11529 38165 11563 38199
rect 11563 38165 11572 38199
rect 11520 38156 11572 38165
rect 12900 38156 12952 38208
rect 13360 38156 13412 38208
rect 14372 38199 14424 38208
rect 14372 38165 14381 38199
rect 14381 38165 14415 38199
rect 14415 38165 14424 38199
rect 14372 38156 14424 38165
rect 15016 38199 15068 38208
rect 15016 38165 15025 38199
rect 15025 38165 15059 38199
rect 15059 38165 15068 38199
rect 15016 38156 15068 38165
rect 15384 38156 15436 38208
rect 16396 38156 16448 38208
rect 16764 38199 16816 38208
rect 16764 38165 16773 38199
rect 16773 38165 16807 38199
rect 16807 38165 16816 38199
rect 16764 38156 16816 38165
rect 18052 38428 18104 38480
rect 23664 38403 23716 38412
rect 23664 38369 23673 38403
rect 23673 38369 23707 38403
rect 23707 38369 23716 38403
rect 23664 38360 23716 38369
rect 21732 38292 21784 38344
rect 22652 38292 22704 38344
rect 17408 38156 17460 38208
rect 19432 38156 19484 38208
rect 5982 38054 6034 38106
rect 6046 38054 6098 38106
rect 6110 38054 6162 38106
rect 6174 38054 6226 38106
rect 15982 38054 16034 38106
rect 16046 38054 16098 38106
rect 16110 38054 16162 38106
rect 16174 38054 16226 38106
rect 25982 38054 26034 38106
rect 26046 38054 26098 38106
rect 26110 38054 26162 38106
rect 26174 38054 26226 38106
rect 8668 37816 8720 37868
rect 8208 37748 8260 37800
rect 9036 37952 9088 38004
rect 11520 37952 11572 38004
rect 12348 37952 12400 38004
rect 13176 37952 13228 38004
rect 14648 37952 14700 38004
rect 15752 37952 15804 38004
rect 16580 37995 16632 38004
rect 16580 37961 16589 37995
rect 16589 37961 16623 37995
rect 16623 37961 16632 37995
rect 16580 37952 16632 37961
rect 18512 37952 18564 38004
rect 19524 37952 19576 38004
rect 23572 37952 23624 38004
rect 23756 37952 23808 38004
rect 23940 37952 23992 38004
rect 9404 37884 9456 37936
rect 10600 37884 10652 37936
rect 15660 37884 15712 37936
rect 16120 37884 16172 37936
rect 16396 37884 16448 37936
rect 4896 37680 4948 37732
rect 8484 37680 8536 37732
rect 7840 37612 7892 37664
rect 9496 37612 9548 37664
rect 10140 37680 10192 37732
rect 9864 37612 9916 37664
rect 11796 37816 11848 37868
rect 13176 37816 13228 37868
rect 14004 37816 14056 37868
rect 15384 37816 15436 37868
rect 16580 37816 16632 37868
rect 18512 37816 18564 37868
rect 20812 37816 20864 37868
rect 23664 37816 23716 37868
rect 10784 37791 10836 37800
rect 10784 37757 10793 37791
rect 10793 37757 10827 37791
rect 10827 37757 10836 37791
rect 10784 37748 10836 37757
rect 10876 37748 10928 37800
rect 12992 37748 13044 37800
rect 14280 37791 14332 37800
rect 14280 37757 14289 37791
rect 14289 37757 14323 37791
rect 14323 37757 14332 37791
rect 14280 37748 14332 37757
rect 15292 37748 15344 37800
rect 15660 37748 15712 37800
rect 16396 37748 16448 37800
rect 17316 37748 17368 37800
rect 20260 37791 20312 37800
rect 20260 37757 20269 37791
rect 20269 37757 20303 37791
rect 20303 37757 20312 37791
rect 20260 37748 20312 37757
rect 20720 37748 20772 37800
rect 23572 37748 23624 37800
rect 25412 37952 25464 38004
rect 12900 37680 12952 37732
rect 13176 37723 13228 37732
rect 13176 37689 13185 37723
rect 13185 37689 13219 37723
rect 13219 37689 13228 37723
rect 13176 37680 13228 37689
rect 12716 37655 12768 37664
rect 12716 37621 12725 37655
rect 12725 37621 12759 37655
rect 12759 37621 12768 37655
rect 12716 37612 12768 37621
rect 14188 37655 14240 37664
rect 14188 37621 14197 37655
rect 14197 37621 14231 37655
rect 14231 37621 14240 37655
rect 14188 37612 14240 37621
rect 14464 37680 14516 37732
rect 14924 37612 14976 37664
rect 15292 37655 15344 37664
rect 15292 37621 15301 37655
rect 15301 37621 15335 37655
rect 15335 37621 15344 37655
rect 15752 37723 15804 37732
rect 15752 37689 15761 37723
rect 15761 37689 15795 37723
rect 15795 37689 15804 37723
rect 15752 37680 15804 37689
rect 15936 37723 15988 37732
rect 15936 37689 15945 37723
rect 15945 37689 15979 37723
rect 15979 37689 15988 37723
rect 15936 37680 15988 37689
rect 16764 37680 16816 37732
rect 17500 37680 17552 37732
rect 20352 37723 20404 37732
rect 20352 37689 20361 37723
rect 20361 37689 20395 37723
rect 20395 37689 20404 37723
rect 20352 37680 20404 37689
rect 23848 37723 23900 37732
rect 23848 37689 23857 37723
rect 23857 37689 23891 37723
rect 23891 37689 23900 37723
rect 23848 37680 23900 37689
rect 24768 37748 24820 37800
rect 26240 37748 26292 37800
rect 15292 37612 15344 37621
rect 16304 37612 16356 37664
rect 17408 37612 17460 37664
rect 18880 37612 18932 37664
rect 23664 37612 23716 37664
rect 27528 37655 27580 37664
rect 27528 37621 27537 37655
rect 27537 37621 27571 37655
rect 27571 37621 27580 37655
rect 27528 37612 27580 37621
rect 10982 37510 11034 37562
rect 11046 37510 11098 37562
rect 11110 37510 11162 37562
rect 11174 37510 11226 37562
rect 20982 37510 21034 37562
rect 21046 37510 21098 37562
rect 21110 37510 21162 37562
rect 21174 37510 21226 37562
rect 7748 37408 7800 37460
rect 8944 37408 8996 37460
rect 9404 37451 9456 37460
rect 9404 37417 9413 37451
rect 9413 37417 9447 37451
rect 9447 37417 9456 37451
rect 9404 37408 9456 37417
rect 3148 37340 3200 37392
rect 8668 37383 8720 37392
rect 8668 37349 8677 37383
rect 8677 37349 8711 37383
rect 8711 37349 8720 37383
rect 8668 37340 8720 37349
rect 1676 37315 1728 37324
rect 1676 37281 1685 37315
rect 1685 37281 1719 37315
rect 1719 37281 1728 37315
rect 1676 37272 1728 37281
rect 1400 37247 1452 37256
rect 1400 37213 1409 37247
rect 1409 37213 1443 37247
rect 1443 37213 1452 37247
rect 1400 37204 1452 37213
rect 6552 37204 6604 37256
rect 9496 37272 9548 37324
rect 10784 37340 10836 37392
rect 10876 37383 10928 37392
rect 10876 37349 10885 37383
rect 10885 37349 10919 37383
rect 10919 37349 10928 37383
rect 12808 37408 12860 37460
rect 13636 37408 13688 37460
rect 14924 37408 14976 37460
rect 15384 37408 15436 37460
rect 19524 37408 19576 37460
rect 20260 37451 20312 37460
rect 20260 37417 20269 37451
rect 20269 37417 20303 37451
rect 20303 37417 20312 37451
rect 20260 37408 20312 37417
rect 10876 37340 10928 37349
rect 11796 37340 11848 37392
rect 12440 37340 12492 37392
rect 13544 37340 13596 37392
rect 13728 37340 13780 37392
rect 15016 37340 15068 37392
rect 15660 37340 15712 37392
rect 11336 37315 11388 37324
rect 7012 37247 7064 37256
rect 7012 37213 7021 37247
rect 7021 37213 7055 37247
rect 7055 37213 7064 37247
rect 7012 37204 7064 37213
rect 9220 37204 9272 37256
rect 11336 37281 11345 37315
rect 11345 37281 11379 37315
rect 11379 37281 11388 37315
rect 11336 37272 11388 37281
rect 11428 37315 11480 37324
rect 11428 37281 11437 37315
rect 11437 37281 11471 37315
rect 11471 37281 11480 37315
rect 11428 37272 11480 37281
rect 12808 37272 12860 37324
rect 12992 37272 13044 37324
rect 16764 37272 16816 37324
rect 16856 37315 16908 37324
rect 16856 37281 16865 37315
rect 16865 37281 16899 37315
rect 16899 37281 16908 37315
rect 16856 37272 16908 37281
rect 17408 37272 17460 37324
rect 10600 37204 10652 37256
rect 15660 37247 15712 37256
rect 11060 37136 11112 37188
rect 6368 37068 6420 37120
rect 9036 37111 9088 37120
rect 9036 37077 9045 37111
rect 9045 37077 9079 37111
rect 9079 37077 9088 37111
rect 9036 37068 9088 37077
rect 11244 37068 11296 37120
rect 15660 37213 15669 37247
rect 15669 37213 15703 37247
rect 15703 37213 15712 37247
rect 15660 37204 15712 37213
rect 17776 37204 17828 37256
rect 18144 37272 18196 37324
rect 18420 37315 18472 37324
rect 18420 37281 18429 37315
rect 18429 37281 18463 37315
rect 18463 37281 18472 37315
rect 18420 37272 18472 37281
rect 22100 37408 22152 37460
rect 25504 37451 25556 37460
rect 25504 37417 25513 37451
rect 25513 37417 25547 37451
rect 25547 37417 25556 37451
rect 25504 37408 25556 37417
rect 26240 37451 26292 37460
rect 26240 37417 26249 37451
rect 26249 37417 26283 37451
rect 26283 37417 26292 37451
rect 26240 37408 26292 37417
rect 22560 37272 22612 37324
rect 22744 37315 22796 37324
rect 22744 37281 22753 37315
rect 22753 37281 22787 37315
rect 22787 37281 22796 37315
rect 22744 37272 22796 37281
rect 23664 37315 23716 37324
rect 23664 37281 23673 37315
rect 23673 37281 23707 37315
rect 23707 37281 23716 37315
rect 23664 37272 23716 37281
rect 24032 37272 24084 37324
rect 22468 37204 22520 37256
rect 23480 37204 23532 37256
rect 24676 37204 24728 37256
rect 17592 37136 17644 37188
rect 17684 37136 17736 37188
rect 14740 37068 14792 37120
rect 15660 37068 15712 37120
rect 15752 37068 15804 37120
rect 16672 37068 16724 37120
rect 17224 37068 17276 37120
rect 18788 37068 18840 37120
rect 19064 37068 19116 37120
rect 19432 37068 19484 37120
rect 5982 36966 6034 37018
rect 6046 36966 6098 37018
rect 6110 36966 6162 37018
rect 6174 36966 6226 37018
rect 15982 36966 16034 37018
rect 16046 36966 16098 37018
rect 16110 36966 16162 37018
rect 16174 36966 16226 37018
rect 25982 36966 26034 37018
rect 26046 36966 26098 37018
rect 26110 36966 26162 37018
rect 26174 36966 26226 37018
rect 1676 36907 1728 36916
rect 1676 36873 1685 36907
rect 1685 36873 1719 36907
rect 1719 36873 1728 36907
rect 1676 36864 1728 36873
rect 6828 36864 6880 36916
rect 9496 36864 9548 36916
rect 9772 36864 9824 36916
rect 11060 36907 11112 36916
rect 11060 36873 11069 36907
rect 11069 36873 11103 36907
rect 11103 36873 11112 36907
rect 11060 36864 11112 36873
rect 11336 36864 11388 36916
rect 12348 36864 12400 36916
rect 12532 36864 12584 36916
rect 6552 36839 6604 36848
rect 6552 36805 6561 36839
rect 6561 36805 6595 36839
rect 6595 36805 6604 36839
rect 6552 36796 6604 36805
rect 10600 36839 10652 36848
rect 10600 36805 10609 36839
rect 10609 36805 10643 36839
rect 10643 36805 10652 36839
rect 10600 36796 10652 36805
rect 2136 36771 2188 36780
rect 2136 36737 2145 36771
rect 2145 36737 2179 36771
rect 2179 36737 2188 36771
rect 2136 36728 2188 36737
rect 7104 36771 7156 36780
rect 7104 36737 7113 36771
rect 7113 36737 7147 36771
rect 7147 36737 7156 36771
rect 7104 36728 7156 36737
rect 7932 36728 7984 36780
rect 8852 36728 8904 36780
rect 9312 36728 9364 36780
rect 9496 36728 9548 36780
rect 1400 36660 1452 36712
rect 2412 36660 2464 36712
rect 6368 36660 6420 36712
rect 6920 36660 6972 36712
rect 9404 36703 9456 36712
rect 9404 36669 9413 36703
rect 9413 36669 9447 36703
rect 9447 36669 9456 36703
rect 9404 36660 9456 36669
rect 11152 36771 11204 36780
rect 11152 36737 11161 36771
rect 11161 36737 11195 36771
rect 11195 36737 11204 36771
rect 11152 36728 11204 36737
rect 12624 36728 12676 36780
rect 13728 36864 13780 36916
rect 15660 36864 15712 36916
rect 16396 36864 16448 36916
rect 17684 36864 17736 36916
rect 18420 36864 18472 36916
rect 22100 36864 22152 36916
rect 22744 36864 22796 36916
rect 23940 36907 23992 36916
rect 23940 36873 23949 36907
rect 23949 36873 23983 36907
rect 23983 36873 23992 36907
rect 23940 36864 23992 36873
rect 24768 36864 24820 36916
rect 13360 36796 13412 36848
rect 15016 36796 15068 36848
rect 15292 36796 15344 36848
rect 16580 36796 16632 36848
rect 17224 36796 17276 36848
rect 14556 36728 14608 36780
rect 16764 36771 16816 36780
rect 6460 36592 6512 36644
rect 3240 36567 3292 36576
rect 3240 36533 3249 36567
rect 3249 36533 3283 36567
rect 3283 36533 3292 36567
rect 3240 36524 3292 36533
rect 6644 36524 6696 36576
rect 8852 36592 8904 36644
rect 9680 36660 9732 36712
rect 9220 36567 9272 36576
rect 9220 36533 9229 36567
rect 9229 36533 9263 36567
rect 9263 36533 9272 36567
rect 9220 36524 9272 36533
rect 9680 36567 9732 36576
rect 9680 36533 9689 36567
rect 9689 36533 9723 36567
rect 9723 36533 9732 36567
rect 9680 36524 9732 36533
rect 13084 36660 13136 36712
rect 13728 36660 13780 36712
rect 14188 36660 14240 36712
rect 16304 36703 16356 36712
rect 12440 36592 12492 36644
rect 14740 36635 14792 36644
rect 14740 36601 14749 36635
rect 14749 36601 14783 36635
rect 14783 36601 14792 36635
rect 14740 36592 14792 36601
rect 14280 36524 14332 36576
rect 14556 36524 14608 36576
rect 15292 36524 15344 36576
rect 16304 36669 16313 36703
rect 16313 36669 16347 36703
rect 16347 36669 16356 36703
rect 16304 36660 16356 36669
rect 16764 36737 16773 36771
rect 16773 36737 16807 36771
rect 16807 36737 16816 36771
rect 16764 36728 16816 36737
rect 16856 36728 16908 36780
rect 18052 36703 18104 36712
rect 18052 36669 18061 36703
rect 18061 36669 18095 36703
rect 18095 36669 18104 36703
rect 18052 36660 18104 36669
rect 19064 36703 19116 36712
rect 19064 36669 19073 36703
rect 19073 36669 19107 36703
rect 19107 36669 19116 36703
rect 21640 36728 21692 36780
rect 25872 36728 25924 36780
rect 19064 36660 19116 36669
rect 20720 36660 20772 36712
rect 26332 36728 26384 36780
rect 16120 36592 16172 36644
rect 16672 36592 16724 36644
rect 21548 36592 21600 36644
rect 22468 36592 22520 36644
rect 15936 36524 15988 36576
rect 16488 36524 16540 36576
rect 27712 36567 27764 36576
rect 27712 36533 27721 36567
rect 27721 36533 27755 36567
rect 27755 36533 27764 36567
rect 27712 36524 27764 36533
rect 10982 36422 11034 36474
rect 11046 36422 11098 36474
rect 11110 36422 11162 36474
rect 11174 36422 11226 36474
rect 20982 36422 21034 36474
rect 21046 36422 21098 36474
rect 21110 36422 21162 36474
rect 21174 36422 21226 36474
rect 2136 36320 2188 36372
rect 7104 36320 7156 36372
rect 7840 36320 7892 36372
rect 8300 36363 8352 36372
rect 8300 36329 8309 36363
rect 8309 36329 8343 36363
rect 8343 36329 8352 36363
rect 8300 36320 8352 36329
rect 10692 36320 10744 36372
rect 13544 36320 13596 36372
rect 15016 36320 15068 36372
rect 19616 36363 19668 36372
rect 19616 36329 19625 36363
rect 19625 36329 19659 36363
rect 19659 36329 19668 36363
rect 19616 36320 19668 36329
rect 19984 36363 20036 36372
rect 19984 36329 19993 36363
rect 19993 36329 20027 36363
rect 20027 36329 20036 36363
rect 19984 36320 20036 36329
rect 20444 36320 20496 36372
rect 20720 36363 20772 36372
rect 20720 36329 20729 36363
rect 20729 36329 20763 36363
rect 20763 36329 20772 36363
rect 20720 36320 20772 36329
rect 8576 36252 8628 36304
rect 10876 36252 10928 36304
rect 11704 36252 11756 36304
rect 13636 36252 13688 36304
rect 3700 36184 3752 36236
rect 5172 36184 5224 36236
rect 4160 36116 4212 36168
rect 2412 35980 2464 36032
rect 5356 35980 5408 36032
rect 7656 35980 7708 36032
rect 10140 36227 10192 36236
rect 10140 36193 10149 36227
rect 10149 36193 10183 36227
rect 10183 36193 10192 36227
rect 10140 36184 10192 36193
rect 10600 36227 10652 36236
rect 10600 36193 10609 36227
rect 10609 36193 10643 36227
rect 10643 36193 10652 36227
rect 10600 36184 10652 36193
rect 10692 36227 10744 36236
rect 10692 36193 10701 36227
rect 10701 36193 10735 36227
rect 10735 36193 10744 36227
rect 10692 36184 10744 36193
rect 8576 36116 8628 36168
rect 12624 36184 12676 36236
rect 12808 36184 12860 36236
rect 13360 36184 13412 36236
rect 14096 36252 14148 36304
rect 14740 36252 14792 36304
rect 16304 36252 16356 36304
rect 17592 36295 17644 36304
rect 14556 36184 14608 36236
rect 15936 36227 15988 36236
rect 15936 36193 15945 36227
rect 15945 36193 15979 36227
rect 15979 36193 15988 36227
rect 15936 36184 15988 36193
rect 17592 36261 17601 36295
rect 17601 36261 17635 36295
rect 17635 36261 17644 36295
rect 17592 36252 17644 36261
rect 21824 36295 21876 36304
rect 21824 36261 21833 36295
rect 21833 36261 21867 36295
rect 21867 36261 21876 36295
rect 21824 36252 21876 36261
rect 13636 36159 13688 36168
rect 13636 36125 13645 36159
rect 13645 36125 13679 36159
rect 13679 36125 13688 36159
rect 13636 36116 13688 36125
rect 16488 36116 16540 36168
rect 16856 36159 16908 36168
rect 16856 36125 16865 36159
rect 16865 36125 16899 36159
rect 16899 36125 16908 36159
rect 16856 36116 16908 36125
rect 7932 36048 7984 36100
rect 9128 36048 9180 36100
rect 11060 36048 11112 36100
rect 12440 36048 12492 36100
rect 15016 36048 15068 36100
rect 16120 36048 16172 36100
rect 16212 36048 16264 36100
rect 17776 36184 17828 36236
rect 19064 36184 19116 36236
rect 19432 36184 19484 36236
rect 21180 36184 21232 36236
rect 22836 36184 22888 36236
rect 17592 36116 17644 36168
rect 18236 36116 18288 36168
rect 20720 36116 20772 36168
rect 21548 36116 21600 36168
rect 21824 36116 21876 36168
rect 22008 36116 22060 36168
rect 22468 36116 22520 36168
rect 17224 36048 17276 36100
rect 20260 36091 20312 36100
rect 20260 36057 20269 36091
rect 20269 36057 20303 36091
rect 20303 36057 20312 36091
rect 20260 36048 20312 36057
rect 9036 36023 9088 36032
rect 9036 35989 9045 36023
rect 9045 35989 9079 36023
rect 9079 35989 9088 36023
rect 9036 35980 9088 35989
rect 11796 35980 11848 36032
rect 12532 36023 12584 36032
rect 12532 35989 12541 36023
rect 12541 35989 12575 36023
rect 12575 35989 12584 36023
rect 12532 35980 12584 35989
rect 13912 35980 13964 36032
rect 14832 36023 14884 36032
rect 14832 35989 14841 36023
rect 14841 35989 14875 36023
rect 14875 35989 14884 36023
rect 16396 36023 16448 36032
rect 14832 35980 14884 35989
rect 16396 35989 16405 36023
rect 16405 35989 16439 36023
rect 16439 35989 16448 36023
rect 16396 35980 16448 35989
rect 16672 35980 16724 36032
rect 17500 35980 17552 36032
rect 17960 35980 18012 36032
rect 19156 35980 19208 36032
rect 21180 36023 21232 36032
rect 21180 35989 21189 36023
rect 21189 35989 21223 36023
rect 21223 35989 21232 36023
rect 21180 35980 21232 35989
rect 23572 35980 23624 36032
rect 26332 35980 26384 36032
rect 5982 35878 6034 35930
rect 6046 35878 6098 35930
rect 6110 35878 6162 35930
rect 6174 35878 6226 35930
rect 15982 35878 16034 35930
rect 16046 35878 16098 35930
rect 16110 35878 16162 35930
rect 16174 35878 16226 35930
rect 25982 35878 26034 35930
rect 26046 35878 26098 35930
rect 26110 35878 26162 35930
rect 26174 35878 26226 35930
rect 4620 35819 4672 35828
rect 4620 35785 4629 35819
rect 4629 35785 4663 35819
rect 4663 35785 4672 35819
rect 4620 35776 4672 35785
rect 4896 35819 4948 35828
rect 4896 35785 4905 35819
rect 4905 35785 4939 35819
rect 4939 35785 4948 35819
rect 4896 35776 4948 35785
rect 5172 35819 5224 35828
rect 5172 35785 5181 35819
rect 5181 35785 5215 35819
rect 5215 35785 5224 35819
rect 5172 35776 5224 35785
rect 8576 35819 8628 35828
rect 8576 35785 8585 35819
rect 8585 35785 8619 35819
rect 8619 35785 8628 35819
rect 8576 35776 8628 35785
rect 15108 35776 15160 35828
rect 17224 35819 17276 35828
rect 1400 35436 1452 35488
rect 2412 35708 2464 35760
rect 4160 35751 4212 35760
rect 4160 35717 4169 35751
rect 4169 35717 4203 35751
rect 4203 35717 4212 35751
rect 4160 35708 4212 35717
rect 7656 35708 7708 35760
rect 12808 35708 12860 35760
rect 14280 35708 14332 35760
rect 2872 35683 2924 35692
rect 2872 35649 2881 35683
rect 2881 35649 2915 35683
rect 2915 35649 2924 35683
rect 2872 35640 2924 35649
rect 6644 35640 6696 35692
rect 7196 35640 7248 35692
rect 1860 35572 1912 35624
rect 6184 35615 6236 35624
rect 2320 35547 2372 35556
rect 2320 35513 2329 35547
rect 2329 35513 2363 35547
rect 2363 35513 2372 35547
rect 2320 35504 2372 35513
rect 4528 35504 4580 35556
rect 6184 35581 6193 35615
rect 6193 35581 6227 35615
rect 6227 35581 6236 35615
rect 6184 35572 6236 35581
rect 7840 35615 7892 35624
rect 7840 35581 7849 35615
rect 7849 35581 7883 35615
rect 7883 35581 7892 35615
rect 7840 35572 7892 35581
rect 8208 35640 8260 35692
rect 9772 35640 9824 35692
rect 11336 35640 11388 35692
rect 12440 35640 12492 35692
rect 13084 35640 13136 35692
rect 14556 35640 14608 35692
rect 15108 35640 15160 35692
rect 16304 35708 16356 35760
rect 17224 35785 17233 35819
rect 17233 35785 17267 35819
rect 17267 35785 17276 35819
rect 17224 35776 17276 35785
rect 18144 35776 18196 35828
rect 19340 35776 19392 35828
rect 17776 35708 17828 35760
rect 18236 35708 18288 35760
rect 15936 35683 15988 35692
rect 15936 35649 15945 35683
rect 15945 35649 15979 35683
rect 15979 35649 15988 35683
rect 15936 35640 15988 35649
rect 16856 35640 16908 35692
rect 18420 35640 18472 35692
rect 1676 35436 1728 35488
rect 6920 35436 6972 35488
rect 7104 35436 7156 35488
rect 7656 35436 7708 35488
rect 8484 35572 8536 35624
rect 9128 35615 9180 35624
rect 9128 35581 9137 35615
rect 9137 35581 9171 35615
rect 9171 35581 9180 35615
rect 9128 35572 9180 35581
rect 9496 35547 9548 35556
rect 9496 35513 9505 35547
rect 9505 35513 9539 35547
rect 9539 35513 9548 35547
rect 9496 35504 9548 35513
rect 10140 35572 10192 35624
rect 11704 35572 11756 35624
rect 10784 35504 10836 35556
rect 11060 35547 11112 35556
rect 11060 35513 11069 35547
rect 11069 35513 11103 35547
rect 11103 35513 11112 35547
rect 11060 35504 11112 35513
rect 11428 35547 11480 35556
rect 11428 35513 11437 35547
rect 11437 35513 11471 35547
rect 11471 35513 11480 35547
rect 11428 35504 11480 35513
rect 12164 35504 12216 35556
rect 12440 35547 12492 35556
rect 12440 35513 12449 35547
rect 12449 35513 12483 35547
rect 12483 35513 12492 35547
rect 12440 35504 12492 35513
rect 14188 35572 14240 35624
rect 13360 35504 13412 35556
rect 13820 35504 13872 35556
rect 16028 35572 16080 35624
rect 17224 35572 17276 35624
rect 18144 35572 18196 35624
rect 21640 35776 21692 35828
rect 22468 35819 22520 35828
rect 22468 35785 22477 35819
rect 22477 35785 22511 35819
rect 22511 35785 22520 35819
rect 22468 35776 22520 35785
rect 23940 35683 23992 35692
rect 23940 35649 23949 35683
rect 23949 35649 23983 35683
rect 23983 35649 23992 35683
rect 23940 35640 23992 35649
rect 26332 35640 26384 35692
rect 21640 35615 21692 35624
rect 21640 35581 21649 35615
rect 21649 35581 21683 35615
rect 21683 35581 21692 35615
rect 21640 35572 21692 35581
rect 23020 35572 23072 35624
rect 23572 35572 23624 35624
rect 27804 35640 27856 35692
rect 14740 35547 14792 35556
rect 14740 35513 14749 35547
rect 14749 35513 14783 35547
rect 14783 35513 14792 35547
rect 14740 35504 14792 35513
rect 16488 35504 16540 35556
rect 16764 35504 16816 35556
rect 19156 35504 19208 35556
rect 20536 35547 20588 35556
rect 20536 35513 20545 35547
rect 20545 35513 20579 35547
rect 20579 35513 20588 35547
rect 20536 35504 20588 35513
rect 22284 35504 22336 35556
rect 25320 35547 25372 35556
rect 25320 35513 25329 35547
rect 25329 35513 25363 35547
rect 25363 35513 25372 35547
rect 25320 35504 25372 35513
rect 27804 35547 27856 35556
rect 27804 35513 27813 35547
rect 27813 35513 27847 35547
rect 27847 35513 27856 35547
rect 27804 35504 27856 35513
rect 8300 35436 8352 35488
rect 9036 35436 9088 35488
rect 10140 35436 10192 35488
rect 11336 35436 11388 35488
rect 12532 35436 12584 35488
rect 12992 35436 13044 35488
rect 13912 35479 13964 35488
rect 13912 35445 13921 35479
rect 13921 35445 13955 35479
rect 13955 35445 13964 35479
rect 13912 35436 13964 35445
rect 14924 35436 14976 35488
rect 15476 35436 15528 35488
rect 17960 35436 18012 35488
rect 18236 35436 18288 35488
rect 20720 35436 20772 35488
rect 22836 35479 22888 35488
rect 22836 35445 22845 35479
rect 22845 35445 22879 35479
rect 22879 35445 22888 35479
rect 22836 35436 22888 35445
rect 10982 35334 11034 35386
rect 11046 35334 11098 35386
rect 11110 35334 11162 35386
rect 11174 35334 11226 35386
rect 20982 35334 21034 35386
rect 21046 35334 21098 35386
rect 21110 35334 21162 35386
rect 21174 35334 21226 35386
rect 4620 35275 4672 35284
rect 4620 35241 4629 35275
rect 4629 35241 4663 35275
rect 4663 35241 4672 35275
rect 4620 35232 4672 35241
rect 9496 35232 9548 35284
rect 10140 35232 10192 35284
rect 10600 35232 10652 35284
rect 10784 35232 10836 35284
rect 14188 35275 14240 35284
rect 14188 35241 14197 35275
rect 14197 35241 14231 35275
rect 14231 35241 14240 35275
rect 14188 35232 14240 35241
rect 14924 35232 14976 35284
rect 15936 35232 15988 35284
rect 16488 35232 16540 35284
rect 18052 35232 18104 35284
rect 18144 35275 18196 35284
rect 18144 35241 18153 35275
rect 18153 35241 18187 35275
rect 18187 35241 18196 35275
rect 18144 35232 18196 35241
rect 19340 35232 19392 35284
rect 19892 35275 19944 35284
rect 19892 35241 19901 35275
rect 19901 35241 19935 35275
rect 19935 35241 19944 35275
rect 19892 35232 19944 35241
rect 20536 35275 20588 35284
rect 20536 35241 20545 35275
rect 20545 35241 20579 35275
rect 20579 35241 20588 35275
rect 20536 35232 20588 35241
rect 22192 35232 22244 35284
rect 9128 35207 9180 35216
rect 9128 35173 9137 35207
rect 9137 35173 9171 35207
rect 9171 35173 9180 35207
rect 9128 35164 9180 35173
rect 11244 35207 11296 35216
rect 11244 35173 11253 35207
rect 11253 35173 11287 35207
rect 11287 35173 11296 35207
rect 11244 35164 11296 35173
rect 11980 35207 12032 35216
rect 11980 35173 11989 35207
rect 11989 35173 12023 35207
rect 12023 35173 12032 35207
rect 11980 35164 12032 35173
rect 12532 35207 12584 35216
rect 12532 35173 12541 35207
rect 12541 35173 12575 35207
rect 12575 35173 12584 35207
rect 12532 35164 12584 35173
rect 12716 35164 12768 35216
rect 5080 35139 5132 35148
rect 5080 35105 5089 35139
rect 5089 35105 5123 35139
rect 5123 35105 5132 35139
rect 5080 35096 5132 35105
rect 6644 35096 6696 35148
rect 7012 35096 7064 35148
rect 7840 35096 7892 35148
rect 8944 35096 8996 35148
rect 9864 35139 9916 35148
rect 9864 35105 9873 35139
rect 9873 35105 9907 35139
rect 9907 35105 9916 35139
rect 9864 35096 9916 35105
rect 3424 35028 3476 35080
rect 6000 35071 6052 35080
rect 5356 34960 5408 35012
rect 6000 35037 6009 35071
rect 6009 35037 6043 35071
rect 6043 35037 6052 35071
rect 6000 35028 6052 35037
rect 9036 35028 9088 35080
rect 9128 35028 9180 35080
rect 9404 35028 9456 35080
rect 1400 34892 1452 34944
rect 3424 34935 3476 34944
rect 3424 34901 3433 34935
rect 3433 34901 3467 34935
rect 3467 34901 3476 34935
rect 3424 34892 3476 34901
rect 4988 34935 5040 34944
rect 4988 34901 4997 34935
rect 4997 34901 5031 34935
rect 5031 34901 5040 34935
rect 4988 34892 5040 34901
rect 5264 34935 5316 34944
rect 5264 34901 5273 34935
rect 5273 34901 5307 34935
rect 5307 34901 5316 34935
rect 5264 34892 5316 34901
rect 6368 34892 6420 34944
rect 6552 34935 6604 34944
rect 6552 34901 6561 34935
rect 6561 34901 6595 34935
rect 6595 34901 6604 34935
rect 6552 34892 6604 34901
rect 6828 34892 6880 34944
rect 9864 34960 9916 35012
rect 9956 34960 10008 35012
rect 10140 35096 10192 35148
rect 12808 35139 12860 35148
rect 12808 35105 12817 35139
rect 12817 35105 12851 35139
rect 12851 35105 12860 35139
rect 12808 35096 12860 35105
rect 13268 35164 13320 35216
rect 14740 35164 14792 35216
rect 15108 35164 15160 35216
rect 10600 35028 10652 35080
rect 14556 35096 14608 35148
rect 14004 35028 14056 35080
rect 14280 35028 14332 35080
rect 16672 35164 16724 35216
rect 17224 35207 17276 35216
rect 17224 35173 17233 35207
rect 17233 35173 17267 35207
rect 17267 35173 17276 35207
rect 17224 35164 17276 35173
rect 17592 35207 17644 35216
rect 17592 35173 17601 35207
rect 17601 35173 17635 35207
rect 17635 35173 17644 35207
rect 17592 35164 17644 35173
rect 18420 35207 18472 35216
rect 18420 35173 18429 35207
rect 18429 35173 18463 35207
rect 18463 35173 18472 35207
rect 18420 35164 18472 35173
rect 20444 35164 20496 35216
rect 12072 34960 12124 35012
rect 12532 34960 12584 35012
rect 12716 34960 12768 35012
rect 16396 35096 16448 35148
rect 15660 35028 15712 35080
rect 16856 35071 16908 35080
rect 16856 35037 16865 35071
rect 16865 35037 16899 35071
rect 16899 35037 16908 35071
rect 16856 35028 16908 35037
rect 16580 34960 16632 35012
rect 16764 34960 16816 35012
rect 19432 35096 19484 35148
rect 22284 35164 22336 35216
rect 22008 35139 22060 35148
rect 22008 35105 22017 35139
rect 22017 35105 22051 35139
rect 22051 35105 22060 35139
rect 22008 35096 22060 35105
rect 23388 35139 23440 35148
rect 23388 35105 23397 35139
rect 23397 35105 23431 35139
rect 23431 35105 23440 35139
rect 23388 35096 23440 35105
rect 21640 35028 21692 35080
rect 22192 35071 22244 35080
rect 22192 35037 22201 35071
rect 22201 35037 22235 35071
rect 22235 35037 22244 35071
rect 22192 35028 22244 35037
rect 8668 34935 8720 34944
rect 8668 34901 8677 34935
rect 8677 34901 8711 34935
rect 8711 34901 8720 34935
rect 8668 34892 8720 34901
rect 8944 34892 8996 34944
rect 11428 34935 11480 34944
rect 11428 34901 11452 34935
rect 11452 34901 11480 34935
rect 11428 34892 11480 34901
rect 11704 34892 11756 34944
rect 12440 34892 12492 34944
rect 13820 34892 13872 34944
rect 15292 34892 15344 34944
rect 16672 34935 16724 34944
rect 16672 34901 16681 34935
rect 16681 34901 16715 34935
rect 16715 34901 16724 34935
rect 16672 34892 16724 34901
rect 17500 34892 17552 34944
rect 22468 34935 22520 34944
rect 22468 34901 22477 34935
rect 22477 34901 22511 34935
rect 22511 34901 22520 34935
rect 22468 34892 22520 34901
rect 23020 34935 23072 34944
rect 23020 34901 23029 34935
rect 23029 34901 23063 34935
rect 23063 34901 23072 34935
rect 23020 34892 23072 34901
rect 23480 34892 23532 34944
rect 24952 34892 25004 34944
rect 25504 34892 25556 34944
rect 26332 34892 26384 34944
rect 5982 34790 6034 34842
rect 6046 34790 6098 34842
rect 6110 34790 6162 34842
rect 6174 34790 6226 34842
rect 15982 34790 16034 34842
rect 16046 34790 16098 34842
rect 16110 34790 16162 34842
rect 16174 34790 16226 34842
rect 25982 34790 26034 34842
rect 26046 34790 26098 34842
rect 26110 34790 26162 34842
rect 26174 34790 26226 34842
rect 4528 34731 4580 34740
rect 4528 34697 4537 34731
rect 4537 34697 4571 34731
rect 4571 34697 4580 34731
rect 4528 34688 4580 34697
rect 4988 34688 5040 34740
rect 11244 34688 11296 34740
rect 12164 34731 12216 34740
rect 12164 34697 12173 34731
rect 12173 34697 12207 34731
rect 12207 34697 12216 34731
rect 12164 34688 12216 34697
rect 5080 34663 5132 34672
rect 5080 34629 5089 34663
rect 5089 34629 5123 34663
rect 5123 34629 5132 34663
rect 5080 34620 5132 34629
rect 3884 34595 3936 34604
rect 3884 34561 3893 34595
rect 3893 34561 3927 34595
rect 3927 34561 3936 34595
rect 3884 34552 3936 34561
rect 4988 34552 5040 34604
rect 5356 34595 5408 34604
rect 5356 34561 5365 34595
rect 5365 34561 5399 34595
rect 5399 34561 5408 34595
rect 5356 34552 5408 34561
rect 1400 34527 1452 34536
rect 1400 34493 1409 34527
rect 1409 34493 1443 34527
rect 1443 34493 1452 34527
rect 1400 34484 1452 34493
rect 1676 34527 1728 34536
rect 1676 34493 1685 34527
rect 1685 34493 1719 34527
rect 1719 34493 1728 34527
rect 1676 34484 1728 34493
rect 3976 34484 4028 34536
rect 5264 34484 5316 34536
rect 6644 34663 6696 34672
rect 6644 34629 6653 34663
rect 6653 34629 6687 34663
rect 6687 34629 6696 34663
rect 6644 34620 6696 34629
rect 5908 34595 5960 34604
rect 5908 34561 5917 34595
rect 5917 34561 5951 34595
rect 5951 34561 5960 34595
rect 5908 34552 5960 34561
rect 6552 34552 6604 34604
rect 10048 34620 10100 34672
rect 6920 34552 6972 34604
rect 8116 34595 8168 34604
rect 4620 34416 4672 34468
rect 6368 34484 6420 34536
rect 7656 34484 7708 34536
rect 8116 34561 8125 34595
rect 8125 34561 8159 34595
rect 8159 34561 8168 34595
rect 8116 34552 8168 34561
rect 8944 34595 8996 34604
rect 8944 34561 8953 34595
rect 8953 34561 8987 34595
rect 8987 34561 8996 34595
rect 8944 34552 8996 34561
rect 9496 34552 9548 34604
rect 10140 34552 10192 34604
rect 10324 34552 10376 34604
rect 11336 34620 11388 34672
rect 11612 34620 11664 34672
rect 11704 34620 11756 34672
rect 11888 34620 11940 34672
rect 8300 34484 8352 34536
rect 8484 34527 8536 34536
rect 8484 34493 8493 34527
rect 8493 34493 8527 34527
rect 8527 34493 8536 34527
rect 8484 34484 8536 34493
rect 8668 34527 8720 34536
rect 8668 34493 8677 34527
rect 8677 34493 8711 34527
rect 8711 34493 8720 34527
rect 8668 34484 8720 34493
rect 9036 34527 9088 34536
rect 9036 34493 9045 34527
rect 9045 34493 9079 34527
rect 9079 34493 9088 34527
rect 9036 34484 9088 34493
rect 10508 34527 10560 34536
rect 10508 34493 10517 34527
rect 10517 34493 10551 34527
rect 10551 34493 10560 34527
rect 10508 34484 10560 34493
rect 2780 34391 2832 34400
rect 2780 34357 2789 34391
rect 2789 34357 2823 34391
rect 2823 34357 2832 34391
rect 2780 34348 2832 34357
rect 5172 34348 5224 34400
rect 7104 34416 7156 34468
rect 6552 34348 6604 34400
rect 10784 34416 10836 34468
rect 14188 34688 14240 34740
rect 14556 34688 14608 34740
rect 15016 34688 15068 34740
rect 15108 34688 15160 34740
rect 16580 34688 16632 34740
rect 18420 34688 18472 34740
rect 19432 34731 19484 34740
rect 19432 34697 19441 34731
rect 19441 34697 19475 34731
rect 19475 34697 19484 34731
rect 19432 34688 19484 34697
rect 20076 34688 20128 34740
rect 22008 34688 22060 34740
rect 22192 34688 22244 34740
rect 23388 34688 23440 34740
rect 12992 34620 13044 34672
rect 17776 34620 17828 34672
rect 13268 34595 13320 34604
rect 13268 34561 13277 34595
rect 13277 34561 13311 34595
rect 13311 34561 13320 34595
rect 13268 34552 13320 34561
rect 14740 34552 14792 34604
rect 16488 34552 16540 34604
rect 18052 34552 18104 34604
rect 22284 34663 22336 34672
rect 19064 34595 19116 34604
rect 19064 34561 19073 34595
rect 19073 34561 19107 34595
rect 19107 34561 19116 34595
rect 19064 34552 19116 34561
rect 20536 34595 20588 34604
rect 20536 34561 20545 34595
rect 20545 34561 20579 34595
rect 20579 34561 20588 34595
rect 20536 34552 20588 34561
rect 12716 34527 12768 34536
rect 12716 34493 12725 34527
rect 12725 34493 12759 34527
rect 12759 34493 12768 34527
rect 12716 34484 12768 34493
rect 13084 34484 13136 34536
rect 14372 34527 14424 34536
rect 14372 34493 14381 34527
rect 14381 34493 14415 34527
rect 14415 34493 14424 34527
rect 14372 34484 14424 34493
rect 11980 34416 12032 34468
rect 12164 34416 12216 34468
rect 12348 34416 12400 34468
rect 12440 34416 12492 34468
rect 13820 34416 13872 34468
rect 14556 34459 14608 34468
rect 14556 34425 14565 34459
rect 14565 34425 14599 34459
rect 14599 34425 14608 34459
rect 14556 34416 14608 34425
rect 15108 34484 15160 34536
rect 15936 34484 15988 34536
rect 18880 34484 18932 34536
rect 20076 34484 20128 34536
rect 20260 34484 20312 34536
rect 22284 34629 22293 34663
rect 22293 34629 22327 34663
rect 22327 34629 22336 34663
rect 24952 34688 25004 34740
rect 25320 34688 25372 34740
rect 27712 34731 27764 34740
rect 22284 34620 22336 34629
rect 21548 34595 21600 34604
rect 21548 34561 21557 34595
rect 21557 34561 21591 34595
rect 21591 34561 21600 34595
rect 21548 34552 21600 34561
rect 25044 34595 25096 34604
rect 25044 34561 25053 34595
rect 25053 34561 25087 34595
rect 25087 34561 25096 34595
rect 25044 34552 25096 34561
rect 27712 34697 27721 34731
rect 27721 34697 27755 34731
rect 27755 34697 27764 34731
rect 27712 34688 27764 34697
rect 21640 34484 21692 34536
rect 23020 34484 23072 34536
rect 9128 34348 9180 34400
rect 10324 34348 10376 34400
rect 12808 34391 12860 34400
rect 12808 34357 12817 34391
rect 12817 34357 12851 34391
rect 12851 34357 12860 34391
rect 12808 34348 12860 34357
rect 14832 34348 14884 34400
rect 15016 34416 15068 34468
rect 15568 34416 15620 34468
rect 16488 34459 16540 34468
rect 16488 34425 16497 34459
rect 16497 34425 16531 34459
rect 16531 34425 16540 34459
rect 16488 34416 16540 34425
rect 17960 34416 18012 34468
rect 19616 34416 19668 34468
rect 20720 34416 20772 34468
rect 20904 34416 20956 34468
rect 16672 34348 16724 34400
rect 16948 34348 17000 34400
rect 17224 34348 17276 34400
rect 18512 34348 18564 34400
rect 21640 34348 21692 34400
rect 23756 34484 23808 34536
rect 26240 34484 26292 34536
rect 24308 34348 24360 34400
rect 10982 34246 11034 34298
rect 11046 34246 11098 34298
rect 11110 34246 11162 34298
rect 11174 34246 11226 34298
rect 20982 34246 21034 34298
rect 21046 34246 21098 34298
rect 21110 34246 21162 34298
rect 21174 34246 21226 34298
rect 1676 34187 1728 34196
rect 1676 34153 1685 34187
rect 1685 34153 1719 34187
rect 1719 34153 1728 34187
rect 1676 34144 1728 34153
rect 3424 34187 3476 34196
rect 3424 34153 3433 34187
rect 3433 34153 3467 34187
rect 3467 34153 3476 34187
rect 3424 34144 3476 34153
rect 4344 34187 4396 34196
rect 4344 34153 4353 34187
rect 4353 34153 4387 34187
rect 4387 34153 4396 34187
rect 4344 34144 4396 34153
rect 4620 34187 4672 34196
rect 4620 34153 4629 34187
rect 4629 34153 4663 34187
rect 4663 34153 4672 34187
rect 4620 34144 4672 34153
rect 5448 34144 5500 34196
rect 6368 34144 6420 34196
rect 6828 34144 6880 34196
rect 5356 34119 5408 34128
rect 5356 34085 5365 34119
rect 5365 34085 5399 34119
rect 5399 34085 5408 34119
rect 5356 34076 5408 34085
rect 5540 34076 5592 34128
rect 5816 34119 5868 34128
rect 5816 34085 5825 34119
rect 5825 34085 5859 34119
rect 5859 34085 5868 34119
rect 10232 34144 10284 34196
rect 10508 34144 10560 34196
rect 12164 34187 12216 34196
rect 12164 34153 12173 34187
rect 12173 34153 12207 34187
rect 12207 34153 12216 34187
rect 12164 34144 12216 34153
rect 13544 34144 13596 34196
rect 5816 34076 5868 34085
rect 4436 34051 4488 34060
rect 4436 34017 4445 34051
rect 4445 34017 4479 34051
rect 4479 34017 4488 34051
rect 4436 34008 4488 34017
rect 5264 34008 5316 34060
rect 6644 34008 6696 34060
rect 6828 34008 6880 34060
rect 9864 34008 9916 34060
rect 10876 34076 10928 34128
rect 11980 34076 12032 34128
rect 14372 34144 14424 34196
rect 16764 34187 16816 34196
rect 16764 34153 16773 34187
rect 16773 34153 16807 34187
rect 16807 34153 16816 34187
rect 16764 34144 16816 34153
rect 16856 34144 16908 34196
rect 18052 34187 18104 34196
rect 18052 34153 18061 34187
rect 18061 34153 18095 34187
rect 18095 34153 18104 34187
rect 18052 34144 18104 34153
rect 20812 34144 20864 34196
rect 22376 34187 22428 34196
rect 14188 34076 14240 34128
rect 14280 34076 14332 34128
rect 14740 34076 14792 34128
rect 15108 34076 15160 34128
rect 6184 33983 6236 33992
rect 6184 33949 6193 33983
rect 6193 33949 6227 33983
rect 6227 33949 6236 33983
rect 6184 33940 6236 33949
rect 7012 33983 7064 33992
rect 7012 33949 7021 33983
rect 7021 33949 7055 33983
rect 7055 33949 7064 33983
rect 7012 33940 7064 33949
rect 4988 33872 5040 33924
rect 3792 33847 3844 33856
rect 3792 33813 3801 33847
rect 3801 33813 3835 33847
rect 3835 33813 3844 33847
rect 3792 33804 3844 33813
rect 4528 33804 4580 33856
rect 6920 33847 6972 33856
rect 6920 33813 6929 33847
rect 6929 33813 6963 33847
rect 6963 33813 6972 33847
rect 6920 33804 6972 33813
rect 8116 33940 8168 33992
rect 8300 33940 8352 33992
rect 9956 33940 10008 33992
rect 11428 34008 11480 34060
rect 15292 34051 15344 34060
rect 15292 34017 15301 34051
rect 15301 34017 15335 34051
rect 15335 34017 15344 34051
rect 15292 34008 15344 34017
rect 17960 34076 18012 34128
rect 21640 34076 21692 34128
rect 22376 34153 22385 34187
rect 22385 34153 22419 34187
rect 22419 34153 22428 34187
rect 22376 34144 22428 34153
rect 23204 34076 23256 34128
rect 16672 34008 16724 34060
rect 16856 34051 16908 34060
rect 16856 34017 16865 34051
rect 16865 34017 16899 34051
rect 16899 34017 16908 34051
rect 16856 34008 16908 34017
rect 16948 34008 17000 34060
rect 19248 34008 19300 34060
rect 20720 34008 20772 34060
rect 21364 34008 21416 34060
rect 23388 34051 23440 34060
rect 23388 34017 23397 34051
rect 23397 34017 23431 34051
rect 23431 34017 23440 34051
rect 23388 34008 23440 34017
rect 25320 34008 25372 34060
rect 10968 33940 11020 33992
rect 12072 33940 12124 33992
rect 13268 33940 13320 33992
rect 12900 33872 12952 33924
rect 16488 33940 16540 33992
rect 17316 33983 17368 33992
rect 17316 33949 17325 33983
rect 17325 33949 17359 33983
rect 17359 33949 17368 33983
rect 17316 33940 17368 33949
rect 18236 33983 18288 33992
rect 18236 33949 18245 33983
rect 18245 33949 18279 33983
rect 18279 33949 18288 33983
rect 18236 33940 18288 33949
rect 20812 33940 20864 33992
rect 21640 33983 21692 33992
rect 15936 33872 15988 33924
rect 21640 33949 21649 33983
rect 21649 33949 21683 33983
rect 21683 33949 21692 33983
rect 21640 33940 21692 33949
rect 8208 33804 8260 33856
rect 8668 33804 8720 33856
rect 13084 33847 13136 33856
rect 13084 33813 13093 33847
rect 13093 33813 13127 33847
rect 13127 33813 13136 33847
rect 13084 33804 13136 33813
rect 14004 33804 14056 33856
rect 15568 33847 15620 33856
rect 15568 33813 15577 33847
rect 15577 33813 15611 33847
rect 15611 33813 15620 33847
rect 15568 33804 15620 33813
rect 15660 33804 15712 33856
rect 22836 33940 22888 33992
rect 23020 33940 23072 33992
rect 24952 33983 25004 33992
rect 24952 33949 24961 33983
rect 24961 33949 24995 33983
rect 24995 33949 25004 33983
rect 24952 33940 25004 33949
rect 25044 33940 25096 33992
rect 16488 33804 16540 33856
rect 20076 33804 20128 33856
rect 20720 33847 20772 33856
rect 20720 33813 20729 33847
rect 20729 33813 20763 33847
rect 20763 33813 20772 33847
rect 20720 33804 20772 33813
rect 23480 33804 23532 33856
rect 24308 33847 24360 33856
rect 24308 33813 24317 33847
rect 24317 33813 24351 33847
rect 24351 33813 24360 33847
rect 24308 33804 24360 33813
rect 26332 33804 26384 33856
rect 5982 33702 6034 33754
rect 6046 33702 6098 33754
rect 6110 33702 6162 33754
rect 6174 33702 6226 33754
rect 15982 33702 16034 33754
rect 16046 33702 16098 33754
rect 16110 33702 16162 33754
rect 16174 33702 16226 33754
rect 25982 33702 26034 33754
rect 26046 33702 26098 33754
rect 26110 33702 26162 33754
rect 26174 33702 26226 33754
rect 4528 33643 4580 33652
rect 4528 33609 4537 33643
rect 4537 33609 4571 33643
rect 4571 33609 4580 33643
rect 4528 33600 4580 33609
rect 5264 33532 5316 33584
rect 5816 33532 5868 33584
rect 6368 33600 6420 33652
rect 6644 33643 6696 33652
rect 6644 33609 6653 33643
rect 6653 33609 6687 33643
rect 6687 33609 6696 33643
rect 6644 33600 6696 33609
rect 7104 33643 7156 33652
rect 7104 33609 7113 33643
rect 7113 33609 7147 33643
rect 7147 33609 7156 33643
rect 7104 33600 7156 33609
rect 8116 33600 8168 33652
rect 8576 33600 8628 33652
rect 7748 33532 7800 33584
rect 4988 33464 5040 33516
rect 5356 33507 5408 33516
rect 5356 33473 5365 33507
rect 5365 33473 5399 33507
rect 5399 33473 5408 33507
rect 5356 33464 5408 33473
rect 7288 33507 7340 33516
rect 7288 33473 7297 33507
rect 7297 33473 7331 33507
rect 7331 33473 7340 33507
rect 7288 33464 7340 33473
rect 8116 33507 8168 33516
rect 8116 33473 8125 33507
rect 8125 33473 8159 33507
rect 8159 33473 8168 33507
rect 8116 33464 8168 33473
rect 4344 33439 4396 33448
rect 4344 33405 4353 33439
rect 4353 33405 4387 33439
rect 4387 33405 4396 33439
rect 4344 33396 4396 33405
rect 5448 33439 5500 33448
rect 5448 33405 5457 33439
rect 5457 33405 5491 33439
rect 5491 33405 5500 33439
rect 5448 33396 5500 33405
rect 6920 33396 6972 33448
rect 8208 33439 8260 33448
rect 8208 33405 8217 33439
rect 8217 33405 8251 33439
rect 8251 33405 8260 33439
rect 8208 33396 8260 33405
rect 10140 33532 10192 33584
rect 10876 33600 10928 33652
rect 12164 33600 12216 33652
rect 13544 33600 13596 33652
rect 15568 33600 15620 33652
rect 19248 33600 19300 33652
rect 20628 33600 20680 33652
rect 23020 33600 23072 33652
rect 23204 33643 23256 33652
rect 23204 33609 23213 33643
rect 23213 33609 23247 33643
rect 23247 33609 23256 33643
rect 23204 33600 23256 33609
rect 23572 33600 23624 33652
rect 10968 33575 11020 33584
rect 10968 33541 10977 33575
rect 10977 33541 11011 33575
rect 11011 33541 11020 33575
rect 10968 33532 11020 33541
rect 12072 33532 12124 33584
rect 12532 33532 12584 33584
rect 13084 33532 13136 33584
rect 15016 33532 15068 33584
rect 15384 33532 15436 33584
rect 9956 33439 10008 33448
rect 9956 33405 9965 33439
rect 9965 33405 9999 33439
rect 9999 33405 10008 33439
rect 9956 33396 10008 33405
rect 10232 33396 10284 33448
rect 10508 33396 10560 33448
rect 10784 33396 10836 33448
rect 12808 33464 12860 33516
rect 13544 33464 13596 33516
rect 14924 33464 14976 33516
rect 3884 33371 3936 33380
rect 3884 33337 3893 33371
rect 3893 33337 3927 33371
rect 3927 33337 3936 33371
rect 3884 33328 3936 33337
rect 4436 33328 4488 33380
rect 4988 33328 5040 33380
rect 5908 33371 5960 33380
rect 5540 33260 5592 33312
rect 5908 33337 5917 33371
rect 5917 33337 5951 33371
rect 5951 33337 5960 33371
rect 5908 33328 5960 33337
rect 7288 33328 7340 33380
rect 8760 33328 8812 33380
rect 9220 33371 9272 33380
rect 9220 33337 9229 33371
rect 9229 33337 9263 33371
rect 9263 33337 9272 33371
rect 9220 33328 9272 33337
rect 12164 33328 12216 33380
rect 13084 33396 13136 33448
rect 15108 33439 15160 33448
rect 15108 33405 15117 33439
rect 15117 33405 15151 33439
rect 15151 33405 15160 33439
rect 15108 33396 15160 33405
rect 15384 33396 15436 33448
rect 16212 33464 16264 33516
rect 15936 33396 15988 33448
rect 23112 33532 23164 33584
rect 25044 33600 25096 33652
rect 25504 33600 25556 33652
rect 24952 33532 25004 33584
rect 20352 33464 20404 33516
rect 20628 33464 20680 33516
rect 20904 33507 20956 33516
rect 20904 33473 20913 33507
rect 20913 33473 20947 33507
rect 20947 33473 20956 33507
rect 20904 33464 20956 33473
rect 22560 33507 22612 33516
rect 22560 33473 22569 33507
rect 22569 33473 22603 33507
rect 22603 33473 22612 33507
rect 22560 33464 22612 33473
rect 25320 33464 25372 33516
rect 18880 33396 18932 33448
rect 19616 33396 19668 33448
rect 20444 33396 20496 33448
rect 22284 33396 22336 33448
rect 26332 33464 26384 33516
rect 12348 33328 12400 33380
rect 16948 33371 17000 33380
rect 16948 33337 16957 33371
rect 16957 33337 16991 33371
rect 16991 33337 17000 33371
rect 18788 33371 18840 33380
rect 16948 33328 17000 33337
rect 18788 33337 18797 33371
rect 18797 33337 18831 33371
rect 18831 33337 18840 33371
rect 18788 33328 18840 33337
rect 20352 33328 20404 33380
rect 20904 33328 20956 33380
rect 22376 33328 22428 33380
rect 23296 33328 23348 33380
rect 8668 33303 8720 33312
rect 8668 33269 8677 33303
rect 8677 33269 8711 33303
rect 8711 33269 8720 33303
rect 8668 33260 8720 33269
rect 10324 33260 10376 33312
rect 11980 33303 12032 33312
rect 11980 33269 11989 33303
rect 11989 33269 12023 33303
rect 12023 33269 12032 33303
rect 11980 33260 12032 33269
rect 12900 33260 12952 33312
rect 14372 33303 14424 33312
rect 14372 33269 14381 33303
rect 14381 33269 14415 33303
rect 14415 33269 14424 33303
rect 14372 33260 14424 33269
rect 14832 33260 14884 33312
rect 15936 33260 15988 33312
rect 18052 33260 18104 33312
rect 19432 33303 19484 33312
rect 19432 33269 19441 33303
rect 19441 33269 19475 33303
rect 19475 33269 19484 33303
rect 19432 33260 19484 33269
rect 21364 33303 21416 33312
rect 21364 33269 21373 33303
rect 21373 33269 21407 33303
rect 21407 33269 21416 33303
rect 21364 33260 21416 33269
rect 21916 33260 21968 33312
rect 10982 33158 11034 33210
rect 11046 33158 11098 33210
rect 11110 33158 11162 33210
rect 11174 33158 11226 33210
rect 20982 33158 21034 33210
rect 21046 33158 21098 33210
rect 21110 33158 21162 33210
rect 21174 33158 21226 33210
rect 4620 33099 4672 33108
rect 4620 33065 4629 33099
rect 4629 33065 4663 33099
rect 4663 33065 4672 33099
rect 4620 33056 4672 33065
rect 5172 32920 5224 32972
rect 7012 32988 7064 33040
rect 7840 33056 7892 33108
rect 8116 33056 8168 33108
rect 8392 33056 8444 33108
rect 9496 33056 9548 33108
rect 8760 32988 8812 33040
rect 9128 32988 9180 33040
rect 10416 32988 10468 33040
rect 10508 32988 10560 33040
rect 8300 32963 8352 32972
rect 8300 32929 8309 32963
rect 8309 32929 8343 32963
rect 8343 32929 8352 32963
rect 8300 32920 8352 32929
rect 9312 32920 9364 32972
rect 9588 32920 9640 32972
rect 10324 32963 10376 32972
rect 10324 32929 10333 32963
rect 10333 32929 10367 32963
rect 10367 32929 10376 32963
rect 10324 32920 10376 32929
rect 12164 32988 12216 33040
rect 12716 33031 12768 33040
rect 12716 32997 12725 33031
rect 12725 32997 12759 33031
rect 12759 32997 12768 33031
rect 12716 32988 12768 32997
rect 12900 32988 12952 33040
rect 13084 32920 13136 32972
rect 3424 32852 3476 32904
rect 5724 32895 5776 32904
rect 5724 32861 5733 32895
rect 5733 32861 5767 32895
rect 5767 32861 5776 32895
rect 5724 32852 5776 32861
rect 5908 32852 5960 32904
rect 7748 32852 7800 32904
rect 7012 32784 7064 32836
rect 7656 32784 7708 32836
rect 3884 32759 3936 32768
rect 3884 32725 3893 32759
rect 3893 32725 3927 32759
rect 3927 32725 3936 32759
rect 3884 32716 3936 32725
rect 5448 32759 5500 32768
rect 5448 32725 5457 32759
rect 5457 32725 5491 32759
rect 5491 32725 5500 32759
rect 5448 32716 5500 32725
rect 6920 32716 6972 32768
rect 9128 32852 9180 32904
rect 10784 32895 10836 32904
rect 10784 32861 10793 32895
rect 10793 32861 10827 32895
rect 10827 32861 10836 32895
rect 10784 32852 10836 32861
rect 12256 32852 12308 32904
rect 12440 32852 12492 32904
rect 12992 32852 13044 32904
rect 13820 32895 13872 32904
rect 8116 32784 8168 32836
rect 13820 32861 13829 32895
rect 13829 32861 13863 32895
rect 13863 32861 13872 32895
rect 13820 32852 13872 32861
rect 14096 32988 14148 33040
rect 14280 33056 14332 33108
rect 14556 33099 14608 33108
rect 14556 33065 14565 33099
rect 14565 33065 14599 33099
rect 14599 33065 14608 33099
rect 14556 33056 14608 33065
rect 14832 33056 14884 33108
rect 15108 33056 15160 33108
rect 15476 33099 15528 33108
rect 14740 32988 14792 33040
rect 15476 33065 15485 33099
rect 15485 33065 15519 33099
rect 15519 33065 15528 33099
rect 15476 33056 15528 33065
rect 16212 33056 16264 33108
rect 16580 33056 16632 33108
rect 15384 32988 15436 33040
rect 16028 33031 16080 33040
rect 14188 32963 14240 32972
rect 14188 32929 14197 32963
rect 14197 32929 14231 32963
rect 14231 32929 14240 32963
rect 14188 32920 14240 32929
rect 15568 32963 15620 32972
rect 15568 32929 15577 32963
rect 15577 32929 15611 32963
rect 15611 32929 15620 32963
rect 15568 32920 15620 32929
rect 16028 32997 16037 33031
rect 16037 32997 16071 33031
rect 16071 32997 16080 33031
rect 16028 32988 16080 32997
rect 17500 33056 17552 33108
rect 18604 33099 18656 33108
rect 18604 33065 18613 33099
rect 18613 33065 18647 33099
rect 18647 33065 18656 33099
rect 18604 33056 18656 33065
rect 19616 33099 19668 33108
rect 19616 33065 19625 33099
rect 19625 33065 19659 33099
rect 19659 33065 19668 33099
rect 19616 33056 19668 33065
rect 20812 33056 20864 33108
rect 23388 33056 23440 33108
rect 23756 33056 23808 33108
rect 25136 33099 25188 33108
rect 25136 33065 25145 33099
rect 25145 33065 25179 33099
rect 25179 33065 25188 33099
rect 25136 33056 25188 33065
rect 23296 33031 23348 33040
rect 15936 32920 15988 32972
rect 14372 32852 14424 32904
rect 14556 32852 14608 32904
rect 14832 32852 14884 32904
rect 14924 32852 14976 32904
rect 23296 32997 23305 33031
rect 23305 32997 23339 33031
rect 23339 32997 23348 33031
rect 23296 32988 23348 32997
rect 18236 32920 18288 32972
rect 19156 32920 19208 32972
rect 16488 32852 16540 32904
rect 16856 32852 16908 32904
rect 17500 32895 17552 32904
rect 17500 32861 17509 32895
rect 17509 32861 17543 32895
rect 17543 32861 17552 32895
rect 17500 32852 17552 32861
rect 10140 32716 10192 32768
rect 11428 32716 11480 32768
rect 12164 32716 12216 32768
rect 14096 32784 14148 32836
rect 16304 32784 16356 32836
rect 16580 32716 16632 32768
rect 17960 32716 18012 32768
rect 19984 32716 20036 32768
rect 24308 32920 24360 32972
rect 21180 32895 21232 32904
rect 21180 32861 21189 32895
rect 21189 32861 21223 32895
rect 21223 32861 21232 32895
rect 21180 32852 21232 32861
rect 21640 32852 21692 32904
rect 22284 32895 22336 32904
rect 22284 32861 22293 32895
rect 22293 32861 22327 32895
rect 22327 32861 22336 32895
rect 22284 32852 22336 32861
rect 23756 32895 23808 32904
rect 23756 32861 23765 32895
rect 23765 32861 23799 32895
rect 23799 32861 23808 32895
rect 23756 32852 23808 32861
rect 24032 32895 24084 32904
rect 24032 32861 24041 32895
rect 24041 32861 24075 32895
rect 24075 32861 24084 32895
rect 24032 32852 24084 32861
rect 20536 32716 20588 32768
rect 21364 32716 21416 32768
rect 22008 32716 22060 32768
rect 26332 32716 26384 32768
rect 5982 32614 6034 32666
rect 6046 32614 6098 32666
rect 6110 32614 6162 32666
rect 6174 32614 6226 32666
rect 15982 32614 16034 32666
rect 16046 32614 16098 32666
rect 16110 32614 16162 32666
rect 16174 32614 16226 32666
rect 25982 32614 26034 32666
rect 26046 32614 26098 32666
rect 26110 32614 26162 32666
rect 26174 32614 26226 32666
rect 3424 32555 3476 32564
rect 3424 32521 3433 32555
rect 3433 32521 3467 32555
rect 3467 32521 3476 32555
rect 3424 32512 3476 32521
rect 4896 32555 4948 32564
rect 4896 32521 4905 32555
rect 4905 32521 4939 32555
rect 4939 32521 4948 32555
rect 4896 32512 4948 32521
rect 5172 32555 5224 32564
rect 5172 32521 5181 32555
rect 5181 32521 5215 32555
rect 5215 32521 5224 32555
rect 5172 32512 5224 32521
rect 5816 32512 5868 32564
rect 7932 32555 7984 32564
rect 7932 32521 7941 32555
rect 7941 32521 7975 32555
rect 7975 32521 7984 32555
rect 7932 32512 7984 32521
rect 5264 32444 5316 32496
rect 8116 32444 8168 32496
rect 8300 32376 8352 32428
rect 9404 32512 9456 32564
rect 10232 32512 10284 32564
rect 12164 32512 12216 32564
rect 5632 32283 5684 32292
rect 5632 32249 5641 32283
rect 5641 32249 5675 32283
rect 5675 32249 5684 32283
rect 5632 32240 5684 32249
rect 7656 32308 7708 32360
rect 8668 32444 8720 32496
rect 13084 32512 13136 32564
rect 8852 32376 8904 32428
rect 10140 32351 10192 32360
rect 10140 32317 10149 32351
rect 10149 32317 10183 32351
rect 10183 32317 10192 32351
rect 10140 32308 10192 32317
rect 10232 32308 10284 32360
rect 10600 32308 10652 32360
rect 11244 32351 11296 32360
rect 11244 32317 11253 32351
rect 11253 32317 11287 32351
rect 11287 32317 11296 32351
rect 13268 32376 13320 32428
rect 11244 32308 11296 32317
rect 8852 32283 8904 32292
rect 8852 32249 8861 32283
rect 8861 32249 8895 32283
rect 8895 32249 8904 32283
rect 8852 32240 8904 32249
rect 12532 32240 12584 32292
rect 3884 32215 3936 32224
rect 3884 32181 3893 32215
rect 3893 32181 3927 32215
rect 3927 32181 3936 32215
rect 3884 32172 3936 32181
rect 5448 32172 5500 32224
rect 5908 32215 5960 32224
rect 5908 32181 5917 32215
rect 5917 32181 5951 32215
rect 5951 32181 5960 32215
rect 5908 32172 5960 32181
rect 6460 32172 6512 32224
rect 8392 32172 8444 32224
rect 8760 32172 8812 32224
rect 9956 32172 10008 32224
rect 10140 32215 10192 32224
rect 10140 32181 10149 32215
rect 10149 32181 10183 32215
rect 10183 32181 10192 32215
rect 10140 32172 10192 32181
rect 12256 32215 12308 32224
rect 12256 32181 12265 32215
rect 12265 32181 12299 32215
rect 12299 32181 12308 32215
rect 14280 32283 14332 32292
rect 14280 32249 14289 32283
rect 14289 32249 14323 32283
rect 14323 32249 14332 32283
rect 14280 32240 14332 32249
rect 14740 32283 14792 32292
rect 12256 32172 12308 32181
rect 12992 32172 13044 32224
rect 14004 32172 14056 32224
rect 14740 32249 14749 32283
rect 14749 32249 14783 32283
rect 14783 32249 14792 32283
rect 14740 32240 14792 32249
rect 15108 32172 15160 32224
rect 15568 32512 15620 32564
rect 16672 32512 16724 32564
rect 21180 32555 21232 32564
rect 21180 32521 21189 32555
rect 21189 32521 21223 32555
rect 21223 32521 21232 32555
rect 21180 32512 21232 32521
rect 23480 32555 23532 32564
rect 23480 32521 23489 32555
rect 23489 32521 23523 32555
rect 23523 32521 23532 32555
rect 23480 32512 23532 32521
rect 18696 32444 18748 32496
rect 22284 32444 22336 32496
rect 22744 32444 22796 32496
rect 27528 32444 27580 32496
rect 15568 32376 15620 32428
rect 15844 32376 15896 32428
rect 19800 32376 19852 32428
rect 16856 32308 16908 32360
rect 17776 32308 17828 32360
rect 19156 32351 19208 32360
rect 17960 32240 18012 32292
rect 19156 32317 19165 32351
rect 19165 32317 19199 32351
rect 19199 32317 19208 32351
rect 19156 32308 19208 32317
rect 23112 32376 23164 32428
rect 21732 32308 21784 32360
rect 22560 32351 22612 32360
rect 22560 32317 22569 32351
rect 22569 32317 22603 32351
rect 22603 32317 22612 32351
rect 22560 32308 22612 32317
rect 23020 32308 23072 32360
rect 18144 32240 18196 32292
rect 15568 32172 15620 32224
rect 16948 32172 17000 32224
rect 17500 32172 17552 32224
rect 18236 32172 18288 32224
rect 18604 32172 18656 32224
rect 21640 32172 21692 32224
rect 24032 32172 24084 32224
rect 24676 32172 24728 32224
rect 10982 32070 11034 32122
rect 11046 32070 11098 32122
rect 11110 32070 11162 32122
rect 11174 32070 11226 32122
rect 20982 32070 21034 32122
rect 21046 32070 21098 32122
rect 21110 32070 21162 32122
rect 21174 32070 21226 32122
rect 2872 32011 2924 32020
rect 2872 31977 2881 32011
rect 2881 31977 2915 32011
rect 2915 31977 2924 32011
rect 2872 31968 2924 31977
rect 5080 31968 5132 32020
rect 5264 32011 5316 32020
rect 5264 31977 5273 32011
rect 5273 31977 5307 32011
rect 5307 31977 5316 32011
rect 5264 31968 5316 31977
rect 8300 32011 8352 32020
rect 3884 31900 3936 31952
rect 5724 31943 5776 31952
rect 5724 31909 5733 31943
rect 5733 31909 5767 31943
rect 5767 31909 5776 31943
rect 5724 31900 5776 31909
rect 8300 31977 8309 32011
rect 8309 31977 8343 32011
rect 8343 31977 8352 32011
rect 8300 31968 8352 31977
rect 8576 31968 8628 32020
rect 9128 32011 9180 32020
rect 9128 31977 9137 32011
rect 9137 31977 9171 32011
rect 9171 31977 9180 32011
rect 9128 31968 9180 31977
rect 9404 32011 9456 32020
rect 9404 31977 9413 32011
rect 9413 31977 9447 32011
rect 9447 31977 9456 32011
rect 9404 31968 9456 31977
rect 10048 32011 10100 32020
rect 10048 31977 10057 32011
rect 10057 31977 10091 32011
rect 10091 31977 10100 32011
rect 10048 31968 10100 31977
rect 10324 31968 10376 32020
rect 7656 31900 7708 31952
rect 9036 31900 9088 31952
rect 1400 31832 1452 31884
rect 5908 31832 5960 31884
rect 7932 31832 7984 31884
rect 9312 31832 9364 31884
rect 9956 31875 10008 31884
rect 9956 31841 9965 31875
rect 9965 31841 9999 31875
rect 9999 31841 10008 31875
rect 9956 31832 10008 31841
rect 10968 31900 11020 31952
rect 12624 31968 12676 32020
rect 14004 31968 14056 32020
rect 15016 31968 15068 32020
rect 17776 31968 17828 32020
rect 19524 31968 19576 32020
rect 20444 31968 20496 32020
rect 21732 32011 21784 32020
rect 21732 31977 21741 32011
rect 21741 31977 21775 32011
rect 21775 31977 21784 32011
rect 21732 31968 21784 31977
rect 22560 31968 22612 32020
rect 23480 32011 23532 32020
rect 23480 31977 23489 32011
rect 23489 31977 23523 32011
rect 23523 31977 23532 32011
rect 23480 31968 23532 31977
rect 10324 31832 10376 31884
rect 10508 31875 10560 31884
rect 10508 31841 10517 31875
rect 10517 31841 10551 31875
rect 10551 31841 10560 31875
rect 10508 31832 10560 31841
rect 11796 31875 11848 31884
rect 11796 31841 11805 31875
rect 11805 31841 11839 31875
rect 11839 31841 11848 31875
rect 11796 31832 11848 31841
rect 12164 31875 12216 31884
rect 12164 31841 12173 31875
rect 12173 31841 12207 31875
rect 12207 31841 12216 31875
rect 12164 31832 12216 31841
rect 12348 31900 12400 31952
rect 12900 31900 12952 31952
rect 13360 31900 13412 31952
rect 13544 31900 13596 31952
rect 14280 31900 14332 31952
rect 17960 31943 18012 31952
rect 17960 31909 17969 31943
rect 17969 31909 18003 31943
rect 18003 31909 18012 31943
rect 17960 31900 18012 31909
rect 19892 31900 19944 31952
rect 20720 31900 20772 31952
rect 23112 31943 23164 31952
rect 23112 31909 23121 31943
rect 23121 31909 23155 31943
rect 23155 31909 23164 31943
rect 23112 31900 23164 31909
rect 1676 31764 1728 31816
rect 1952 31764 2004 31816
rect 5724 31764 5776 31816
rect 11244 31764 11296 31816
rect 8760 31739 8812 31748
rect 8760 31705 8769 31739
rect 8769 31705 8803 31739
rect 8803 31705 8812 31739
rect 8760 31696 8812 31705
rect 12164 31696 12216 31748
rect 12716 31832 12768 31884
rect 13176 31875 13228 31884
rect 13176 31841 13185 31875
rect 13185 31841 13219 31875
rect 13219 31841 13228 31875
rect 13176 31832 13228 31841
rect 13912 31832 13964 31884
rect 14004 31832 14056 31884
rect 14648 31832 14700 31884
rect 15292 31875 15344 31884
rect 15292 31841 15301 31875
rect 15301 31841 15335 31875
rect 15335 31841 15344 31875
rect 15292 31832 15344 31841
rect 15844 31832 15896 31884
rect 12348 31764 12400 31816
rect 12808 31807 12860 31816
rect 12808 31773 12817 31807
rect 12817 31773 12851 31807
rect 12851 31773 12860 31807
rect 12808 31764 12860 31773
rect 13360 31764 13412 31816
rect 13728 31764 13780 31816
rect 14372 31764 14424 31816
rect 15476 31764 15528 31816
rect 16856 31832 16908 31884
rect 18880 31832 18932 31884
rect 19616 31832 19668 31884
rect 13084 31696 13136 31748
rect 13636 31696 13688 31748
rect 14924 31696 14976 31748
rect 15844 31696 15896 31748
rect 7196 31628 7248 31680
rect 8944 31628 8996 31680
rect 12716 31628 12768 31680
rect 15568 31628 15620 31680
rect 17500 31764 17552 31816
rect 18972 31807 19024 31816
rect 18972 31773 18981 31807
rect 18981 31773 19015 31807
rect 19015 31773 19024 31807
rect 18972 31764 19024 31773
rect 19064 31696 19116 31748
rect 19524 31764 19576 31816
rect 19984 31764 20036 31816
rect 21732 31832 21784 31884
rect 22928 31875 22980 31884
rect 22928 31841 22937 31875
rect 22937 31841 22971 31875
rect 22971 31841 22980 31875
rect 22928 31832 22980 31841
rect 23480 31832 23532 31884
rect 23664 31832 23716 31884
rect 20812 31764 20864 31816
rect 17960 31628 18012 31680
rect 21180 31671 21232 31680
rect 21180 31637 21189 31671
rect 21189 31637 21223 31671
rect 21223 31637 21232 31671
rect 21180 31628 21232 31637
rect 5982 31526 6034 31578
rect 6046 31526 6098 31578
rect 6110 31526 6162 31578
rect 6174 31526 6226 31578
rect 15982 31526 16034 31578
rect 16046 31526 16098 31578
rect 16110 31526 16162 31578
rect 16174 31526 16226 31578
rect 25982 31526 26034 31578
rect 26046 31526 26098 31578
rect 26110 31526 26162 31578
rect 26174 31526 26226 31578
rect 6644 31467 6696 31476
rect 6644 31433 6653 31467
rect 6653 31433 6687 31467
rect 6687 31433 6696 31467
rect 6644 31424 6696 31433
rect 7196 31424 7248 31476
rect 7932 31467 7984 31476
rect 7932 31433 7941 31467
rect 7941 31433 7975 31467
rect 7975 31433 7984 31467
rect 7932 31424 7984 31433
rect 8208 31424 8260 31476
rect 8484 31424 8536 31476
rect 8852 31467 8904 31476
rect 8852 31433 8861 31467
rect 8861 31433 8895 31467
rect 8895 31433 8904 31467
rect 8852 31424 8904 31433
rect 11520 31424 11572 31476
rect 11796 31424 11848 31476
rect 5540 31399 5592 31408
rect 5540 31365 5549 31399
rect 5549 31365 5583 31399
rect 5583 31365 5592 31399
rect 5540 31356 5592 31365
rect 6920 31356 6972 31408
rect 12440 31356 12492 31408
rect 13360 31424 13412 31476
rect 13912 31467 13964 31476
rect 13912 31433 13921 31467
rect 13921 31433 13955 31467
rect 13955 31433 13964 31467
rect 13912 31424 13964 31433
rect 14096 31424 14148 31476
rect 14372 31424 14424 31476
rect 15292 31424 15344 31476
rect 16396 31467 16448 31476
rect 16396 31433 16405 31467
rect 16405 31433 16439 31467
rect 16439 31433 16448 31467
rect 16396 31424 16448 31433
rect 16764 31424 16816 31476
rect 19616 31467 19668 31476
rect 19616 31433 19625 31467
rect 19625 31433 19659 31467
rect 19659 31433 19668 31467
rect 19616 31424 19668 31433
rect 21732 31467 21784 31476
rect 21732 31433 21741 31467
rect 21741 31433 21775 31467
rect 21775 31433 21784 31467
rect 21732 31424 21784 31433
rect 14188 31356 14240 31408
rect 8300 31288 8352 31340
rect 8668 31288 8720 31340
rect 8944 31288 8996 31340
rect 10600 31288 10652 31340
rect 11152 31288 11204 31340
rect 11888 31288 11940 31340
rect 12072 31288 12124 31340
rect 12624 31288 12676 31340
rect 16580 31356 16632 31408
rect 8852 31220 8904 31272
rect 10048 31263 10100 31272
rect 1952 31195 2004 31204
rect 1952 31161 1961 31195
rect 1961 31161 1995 31195
rect 1995 31161 2004 31195
rect 1952 31152 2004 31161
rect 8576 31195 8628 31204
rect 8576 31161 8585 31195
rect 8585 31161 8619 31195
rect 8619 31161 8628 31195
rect 8576 31152 8628 31161
rect 9404 31195 9456 31204
rect 9404 31161 9413 31195
rect 9413 31161 9447 31195
rect 9447 31161 9456 31195
rect 9404 31152 9456 31161
rect 10048 31229 10057 31263
rect 10057 31229 10091 31263
rect 10091 31229 10100 31263
rect 10048 31220 10100 31229
rect 10508 31220 10560 31272
rect 9956 31152 10008 31204
rect 1676 31127 1728 31136
rect 1676 31093 1685 31127
rect 1685 31093 1719 31127
rect 1719 31093 1728 31127
rect 1676 31084 1728 31093
rect 2964 31084 3016 31136
rect 4804 31127 4856 31136
rect 4804 31093 4813 31127
rect 4813 31093 4847 31127
rect 4847 31093 4856 31127
rect 4804 31084 4856 31093
rect 5448 31084 5500 31136
rect 5816 31127 5868 31136
rect 5816 31093 5825 31127
rect 5825 31093 5859 31127
rect 5859 31093 5868 31127
rect 5816 31084 5868 31093
rect 8668 31084 8720 31136
rect 9128 31084 9180 31136
rect 10968 31220 11020 31272
rect 11796 31220 11848 31272
rect 12716 31220 12768 31272
rect 13360 31220 13412 31272
rect 14188 31220 14240 31272
rect 14372 31288 14424 31340
rect 13728 31152 13780 31204
rect 14280 31152 14332 31204
rect 14832 31288 14884 31340
rect 15844 31288 15896 31340
rect 16304 31288 16356 31340
rect 17960 31288 18012 31340
rect 23940 31331 23992 31340
rect 23940 31297 23949 31331
rect 23949 31297 23983 31331
rect 23983 31297 23992 31331
rect 23940 31288 23992 31297
rect 27620 31331 27672 31340
rect 27620 31297 27629 31331
rect 27629 31297 27663 31331
rect 27663 31297 27672 31331
rect 27620 31288 27672 31297
rect 16488 31263 16540 31272
rect 16488 31229 16497 31263
rect 16497 31229 16531 31263
rect 16531 31229 16540 31263
rect 16488 31220 16540 31229
rect 16580 31220 16632 31272
rect 15108 31195 15160 31204
rect 12256 31127 12308 31136
rect 12256 31093 12265 31127
rect 12265 31093 12299 31127
rect 12299 31093 12308 31127
rect 12256 31084 12308 31093
rect 12532 31084 12584 31136
rect 13820 31084 13872 31136
rect 15108 31161 15117 31195
rect 15117 31161 15151 31195
rect 15151 31161 15160 31195
rect 15108 31152 15160 31161
rect 16856 31152 16908 31204
rect 19064 31220 19116 31272
rect 20536 31263 20588 31272
rect 20536 31229 20545 31263
rect 20545 31229 20579 31263
rect 20579 31229 20588 31263
rect 20536 31220 20588 31229
rect 20812 31220 20864 31272
rect 20904 31220 20956 31272
rect 22928 31220 22980 31272
rect 23756 31220 23808 31272
rect 24676 31220 24728 31272
rect 25780 31220 25832 31272
rect 26240 31220 26292 31272
rect 26424 31263 26476 31272
rect 26424 31229 26433 31263
rect 26433 31229 26467 31263
rect 26467 31229 26476 31263
rect 26424 31220 26476 31229
rect 15568 31084 15620 31136
rect 19984 31127 20036 31136
rect 19984 31093 19993 31127
rect 19993 31093 20027 31127
rect 20027 31093 20036 31127
rect 19984 31084 20036 31093
rect 21732 31152 21784 31204
rect 25044 31127 25096 31136
rect 25044 31093 25053 31127
rect 25053 31093 25087 31127
rect 25087 31093 25096 31127
rect 25044 31084 25096 31093
rect 10982 30982 11034 31034
rect 11046 30982 11098 31034
rect 11110 30982 11162 31034
rect 11174 30982 11226 31034
rect 20982 30982 21034 31034
rect 21046 30982 21098 31034
rect 21110 30982 21162 31034
rect 21174 30982 21226 31034
rect 6368 30880 6420 30932
rect 7196 30880 7248 30932
rect 7472 30880 7524 30932
rect 10416 30880 10468 30932
rect 10876 30880 10928 30932
rect 12624 30880 12676 30932
rect 13176 30880 13228 30932
rect 13820 30923 13872 30932
rect 13820 30889 13829 30923
rect 13829 30889 13863 30923
rect 13863 30889 13872 30923
rect 13820 30880 13872 30889
rect 16672 30923 16724 30932
rect 16672 30889 16681 30923
rect 16681 30889 16715 30923
rect 16715 30889 16724 30923
rect 16672 30880 16724 30889
rect 8760 30812 8812 30864
rect 9588 30812 9640 30864
rect 4804 30744 4856 30796
rect 5724 30744 5776 30796
rect 6644 30744 6696 30796
rect 8668 30744 8720 30796
rect 9128 30787 9180 30796
rect 9128 30753 9137 30787
rect 9137 30753 9171 30787
rect 9171 30753 9180 30787
rect 9128 30744 9180 30753
rect 9312 30744 9364 30796
rect 10048 30744 10100 30796
rect 6828 30676 6880 30728
rect 9956 30676 10008 30728
rect 10968 30812 11020 30864
rect 12256 30812 12308 30864
rect 13084 30812 13136 30864
rect 15016 30812 15068 30864
rect 11520 30744 11572 30796
rect 12440 30787 12492 30796
rect 12440 30753 12449 30787
rect 12449 30753 12483 30787
rect 12483 30753 12492 30787
rect 12440 30744 12492 30753
rect 5632 30608 5684 30660
rect 8944 30608 8996 30660
rect 10968 30676 11020 30728
rect 12164 30676 12216 30728
rect 13176 30787 13228 30796
rect 12716 30676 12768 30728
rect 13176 30753 13185 30787
rect 13185 30753 13219 30787
rect 13219 30753 13228 30787
rect 13176 30744 13228 30753
rect 14280 30744 14332 30796
rect 14464 30744 14516 30796
rect 15292 30787 15344 30796
rect 15292 30753 15301 30787
rect 15301 30753 15335 30787
rect 15335 30753 15344 30787
rect 15292 30744 15344 30753
rect 15384 30744 15436 30796
rect 17960 30880 18012 30932
rect 21916 30880 21968 30932
rect 23756 30923 23808 30932
rect 23756 30889 23765 30923
rect 23765 30889 23799 30923
rect 23799 30889 23808 30923
rect 23756 30880 23808 30889
rect 22192 30812 22244 30864
rect 19156 30744 19208 30796
rect 20904 30787 20956 30796
rect 20904 30753 20913 30787
rect 20913 30753 20947 30787
rect 20947 30753 20956 30787
rect 20904 30744 20956 30753
rect 13268 30676 13320 30728
rect 11796 30608 11848 30660
rect 12624 30608 12676 30660
rect 13452 30608 13504 30660
rect 5540 30583 5592 30592
rect 5540 30549 5549 30583
rect 5549 30549 5583 30583
rect 5583 30549 5592 30583
rect 5540 30540 5592 30549
rect 6368 30540 6420 30592
rect 7472 30583 7524 30592
rect 7472 30549 7481 30583
rect 7481 30549 7515 30583
rect 7515 30549 7524 30583
rect 7472 30540 7524 30549
rect 9312 30540 9364 30592
rect 9864 30540 9916 30592
rect 10232 30540 10284 30592
rect 11520 30540 11572 30592
rect 13360 30540 13412 30592
rect 14924 30676 14976 30728
rect 16580 30676 16632 30728
rect 16672 30676 16724 30728
rect 18144 30676 18196 30728
rect 19064 30676 19116 30728
rect 19892 30676 19944 30728
rect 22192 30719 22244 30728
rect 22192 30685 22201 30719
rect 22201 30685 22235 30719
rect 22235 30685 22244 30719
rect 22192 30676 22244 30685
rect 23388 30676 23440 30728
rect 13636 30608 13688 30660
rect 14464 30608 14516 30660
rect 16304 30608 16356 30660
rect 19340 30608 19392 30660
rect 21088 30651 21140 30660
rect 21088 30617 21097 30651
rect 21097 30617 21131 30651
rect 21131 30617 21140 30651
rect 21088 30608 21140 30617
rect 22100 30608 22152 30660
rect 14740 30540 14792 30592
rect 17960 30540 18012 30592
rect 19064 30583 19116 30592
rect 19064 30549 19073 30583
rect 19073 30549 19107 30583
rect 19107 30549 19116 30583
rect 19064 30540 19116 30549
rect 19616 30583 19668 30592
rect 19616 30549 19625 30583
rect 19625 30549 19659 30583
rect 19659 30549 19668 30583
rect 19616 30540 19668 30549
rect 25780 30540 25832 30592
rect 5982 30438 6034 30490
rect 6046 30438 6098 30490
rect 6110 30438 6162 30490
rect 6174 30438 6226 30490
rect 15982 30438 16034 30490
rect 16046 30438 16098 30490
rect 16110 30438 16162 30490
rect 16174 30438 16226 30490
rect 25982 30438 26034 30490
rect 26046 30438 26098 30490
rect 26110 30438 26162 30490
rect 26174 30438 26226 30490
rect 8668 30379 8720 30388
rect 8668 30345 8677 30379
rect 8677 30345 8711 30379
rect 8711 30345 8720 30379
rect 8668 30336 8720 30345
rect 9772 30336 9824 30388
rect 10876 30336 10928 30388
rect 5264 30311 5316 30320
rect 5264 30277 5273 30311
rect 5273 30277 5307 30311
rect 5307 30277 5316 30311
rect 5264 30268 5316 30277
rect 7472 30268 7524 30320
rect 9956 30268 10008 30320
rect 5632 30243 5684 30252
rect 5632 30209 5641 30243
rect 5641 30209 5675 30243
rect 5675 30209 5684 30243
rect 5632 30200 5684 30209
rect 7196 30200 7248 30252
rect 5540 30132 5592 30184
rect 6828 30132 6880 30184
rect 7472 30175 7524 30184
rect 7472 30141 7481 30175
rect 7481 30141 7515 30175
rect 7515 30141 7524 30175
rect 7472 30132 7524 30141
rect 8576 30200 8628 30252
rect 10508 30200 10560 30252
rect 7932 30175 7984 30184
rect 7932 30141 7941 30175
rect 7941 30141 7975 30175
rect 7975 30141 7984 30175
rect 7932 30132 7984 30141
rect 10048 30175 10100 30184
rect 7656 30064 7708 30116
rect 9588 30064 9640 30116
rect 10048 30141 10057 30175
rect 10057 30141 10091 30175
rect 10091 30141 10100 30175
rect 10048 30132 10100 30141
rect 11428 30200 11480 30252
rect 12348 30336 12400 30388
rect 12900 30336 12952 30388
rect 15384 30336 15436 30388
rect 18144 30336 18196 30388
rect 18512 30336 18564 30388
rect 20904 30379 20956 30388
rect 20904 30345 20913 30379
rect 20913 30345 20947 30379
rect 20947 30345 20956 30379
rect 20904 30336 20956 30345
rect 14280 30311 14332 30320
rect 14280 30277 14289 30311
rect 14289 30277 14323 30311
rect 14323 30277 14332 30311
rect 14280 30268 14332 30277
rect 15292 30268 15344 30320
rect 16304 30268 16356 30320
rect 17500 30268 17552 30320
rect 19248 30268 19300 30320
rect 20260 30311 20312 30320
rect 20260 30277 20269 30311
rect 20269 30277 20303 30311
rect 20303 30277 20312 30311
rect 20260 30268 20312 30277
rect 12164 30200 12216 30252
rect 13360 30200 13412 30252
rect 13820 30200 13872 30252
rect 14004 30200 14056 30252
rect 17224 30200 17276 30252
rect 18512 30243 18564 30252
rect 18512 30209 18521 30243
rect 18521 30209 18555 30243
rect 18555 30209 18564 30243
rect 18512 30200 18564 30209
rect 14740 30175 14792 30184
rect 14740 30141 14749 30175
rect 14749 30141 14783 30175
rect 14783 30141 14792 30175
rect 14740 30132 14792 30141
rect 14924 30175 14976 30184
rect 14924 30141 14933 30175
rect 14933 30141 14967 30175
rect 14967 30141 14976 30175
rect 14924 30132 14976 30141
rect 15108 30132 15160 30184
rect 15936 30175 15988 30184
rect 15936 30141 15945 30175
rect 15945 30141 15979 30175
rect 15979 30141 15988 30175
rect 15936 30132 15988 30141
rect 16488 30132 16540 30184
rect 17960 30132 18012 30184
rect 18604 30132 18656 30184
rect 19064 30175 19116 30184
rect 11428 30064 11480 30116
rect 13544 30064 13596 30116
rect 14004 30064 14056 30116
rect 14188 30064 14240 30116
rect 14280 30064 14332 30116
rect 16672 30064 16724 30116
rect 19064 30141 19073 30175
rect 19073 30141 19107 30175
rect 19107 30141 19116 30175
rect 19064 30132 19116 30141
rect 20076 30175 20128 30184
rect 18880 30064 18932 30116
rect 19248 30064 19300 30116
rect 20076 30141 20085 30175
rect 20085 30141 20119 30175
rect 20119 30141 20128 30175
rect 20076 30132 20128 30141
rect 19432 30064 19484 30116
rect 21640 30107 21692 30116
rect 21640 30073 21649 30107
rect 21649 30073 21683 30107
rect 21683 30073 21692 30107
rect 21640 30064 21692 30073
rect 4620 29996 4672 30048
rect 6644 29996 6696 30048
rect 6920 29996 6972 30048
rect 8300 29996 8352 30048
rect 8852 29996 8904 30048
rect 10140 29996 10192 30048
rect 12256 29996 12308 30048
rect 12440 29996 12492 30048
rect 15016 29996 15068 30048
rect 15384 29996 15436 30048
rect 17500 29996 17552 30048
rect 17960 29996 18012 30048
rect 19340 29996 19392 30048
rect 19616 29996 19668 30048
rect 10982 29894 11034 29946
rect 11046 29894 11098 29946
rect 11110 29894 11162 29946
rect 11174 29894 11226 29946
rect 20982 29894 21034 29946
rect 21046 29894 21098 29946
rect 21110 29894 21162 29946
rect 21174 29894 21226 29946
rect 6552 29835 6604 29844
rect 6552 29801 6561 29835
rect 6561 29801 6595 29835
rect 6595 29801 6604 29835
rect 6552 29792 6604 29801
rect 8300 29835 8352 29844
rect 8300 29801 8309 29835
rect 8309 29801 8343 29835
rect 8343 29801 8352 29835
rect 8300 29792 8352 29801
rect 8576 29792 8628 29844
rect 9312 29792 9364 29844
rect 11796 29792 11848 29844
rect 6828 29724 6880 29776
rect 7656 29724 7708 29776
rect 10048 29724 10100 29776
rect 12348 29767 12400 29776
rect 12348 29733 12357 29767
rect 12357 29733 12391 29767
rect 12391 29733 12400 29767
rect 12348 29724 12400 29733
rect 12900 29724 12952 29776
rect 13176 29792 13228 29844
rect 13360 29792 13412 29844
rect 15016 29792 15068 29844
rect 15752 29792 15804 29844
rect 14648 29724 14700 29776
rect 15108 29767 15160 29776
rect 15108 29733 15117 29767
rect 15117 29733 15151 29767
rect 15151 29733 15160 29767
rect 15108 29724 15160 29733
rect 7104 29656 7156 29708
rect 8116 29699 8168 29708
rect 8116 29665 8125 29699
rect 8125 29665 8159 29699
rect 8159 29665 8168 29699
rect 8116 29656 8168 29665
rect 6920 29588 6972 29640
rect 9220 29656 9272 29708
rect 9864 29588 9916 29640
rect 10140 29588 10192 29640
rect 10416 29588 10468 29640
rect 11428 29520 11480 29572
rect 13268 29656 13320 29708
rect 13636 29699 13688 29708
rect 13636 29665 13645 29699
rect 13645 29665 13679 29699
rect 13679 29665 13688 29699
rect 13636 29656 13688 29665
rect 13820 29699 13872 29708
rect 13820 29665 13826 29699
rect 13826 29665 13872 29699
rect 13820 29656 13872 29665
rect 15384 29724 15436 29776
rect 16212 29724 16264 29776
rect 12716 29588 12768 29640
rect 16488 29656 16540 29708
rect 16580 29656 16632 29708
rect 16856 29699 16908 29708
rect 16856 29665 16865 29699
rect 16865 29665 16899 29699
rect 16899 29665 16908 29699
rect 16856 29656 16908 29665
rect 17500 29792 17552 29844
rect 18052 29792 18104 29844
rect 17776 29724 17828 29776
rect 18880 29724 18932 29776
rect 20076 29792 20128 29844
rect 21916 29792 21968 29844
rect 14188 29588 14240 29640
rect 14924 29588 14976 29640
rect 16304 29588 16356 29640
rect 16672 29588 16724 29640
rect 17776 29588 17828 29640
rect 13360 29520 13412 29572
rect 13544 29520 13596 29572
rect 6552 29452 6604 29504
rect 9312 29452 9364 29504
rect 9680 29452 9732 29504
rect 11060 29495 11112 29504
rect 11060 29461 11069 29495
rect 11069 29461 11103 29495
rect 11103 29461 11112 29495
rect 11060 29452 11112 29461
rect 12256 29452 12308 29504
rect 12532 29452 12584 29504
rect 13912 29495 13964 29504
rect 13912 29461 13921 29495
rect 13921 29461 13955 29495
rect 13955 29461 13964 29495
rect 13912 29452 13964 29461
rect 14280 29495 14332 29504
rect 14280 29461 14289 29495
rect 14289 29461 14323 29495
rect 14323 29461 14332 29495
rect 14280 29452 14332 29461
rect 15384 29452 15436 29504
rect 15752 29495 15804 29504
rect 15752 29461 15761 29495
rect 15761 29461 15795 29495
rect 15795 29461 15804 29495
rect 15752 29452 15804 29461
rect 16764 29520 16816 29572
rect 19064 29656 19116 29708
rect 19892 29656 19944 29708
rect 19156 29588 19208 29640
rect 22192 29724 22244 29776
rect 20352 29656 20404 29708
rect 21824 29699 21876 29708
rect 21824 29665 21833 29699
rect 21833 29665 21867 29699
rect 21867 29665 21876 29699
rect 21824 29656 21876 29665
rect 18880 29452 18932 29504
rect 19340 29452 19392 29504
rect 22376 29452 22428 29504
rect 5982 29350 6034 29402
rect 6046 29350 6098 29402
rect 6110 29350 6162 29402
rect 6174 29350 6226 29402
rect 15982 29350 16034 29402
rect 16046 29350 16098 29402
rect 16110 29350 16162 29402
rect 16174 29350 16226 29402
rect 25982 29350 26034 29402
rect 26046 29350 26098 29402
rect 26110 29350 26162 29402
rect 26174 29350 26226 29402
rect 6644 29291 6696 29300
rect 6644 29257 6653 29291
rect 6653 29257 6687 29291
rect 6687 29257 6696 29291
rect 6644 29248 6696 29257
rect 7104 29291 7156 29300
rect 7104 29257 7113 29291
rect 7113 29257 7147 29291
rect 7147 29257 7156 29291
rect 7104 29248 7156 29257
rect 9128 29291 9180 29300
rect 9128 29257 9137 29291
rect 9137 29257 9171 29291
rect 9171 29257 9180 29291
rect 9128 29248 9180 29257
rect 11428 29291 11480 29300
rect 11428 29257 11437 29291
rect 11437 29257 11471 29291
rect 11471 29257 11480 29291
rect 11428 29248 11480 29257
rect 12348 29248 12400 29300
rect 9312 29180 9364 29232
rect 10508 29180 10560 29232
rect 12716 29180 12768 29232
rect 10416 29112 10468 29164
rect 11060 29112 11112 29164
rect 11428 29112 11480 29164
rect 12440 29112 12492 29164
rect 6184 29044 6236 29096
rect 6828 29044 6880 29096
rect 8208 29087 8260 29096
rect 8208 29053 8217 29087
rect 8217 29053 8251 29087
rect 8251 29053 8260 29087
rect 8208 29044 8260 29053
rect 9128 29044 9180 29096
rect 9404 29044 9456 29096
rect 1400 28976 1452 29028
rect 1952 28976 2004 29028
rect 4620 28976 4672 29028
rect 5448 28976 5500 29028
rect 5816 29019 5868 29028
rect 5816 28985 5825 29019
rect 5825 28985 5859 29019
rect 5859 28985 5868 29019
rect 5816 28976 5868 28985
rect 8116 29019 8168 29028
rect 8116 28985 8125 29019
rect 8125 28985 8159 29019
rect 8159 28985 8168 29019
rect 8116 28976 8168 28985
rect 8668 28976 8720 29028
rect 9312 28976 9364 29028
rect 8944 28908 8996 28960
rect 9496 28908 9548 28960
rect 9772 28908 9824 28960
rect 10692 29044 10744 29096
rect 10876 29044 10928 29096
rect 13176 29087 13228 29096
rect 13176 29053 13185 29087
rect 13185 29053 13219 29087
rect 13219 29053 13228 29087
rect 13176 29044 13228 29053
rect 10876 28908 10928 28960
rect 12624 28976 12676 29028
rect 15108 29248 15160 29300
rect 15292 29248 15344 29300
rect 16396 29248 16448 29300
rect 16764 29248 16816 29300
rect 16856 29248 16908 29300
rect 18052 29248 18104 29300
rect 18512 29248 18564 29300
rect 19892 29291 19944 29300
rect 19892 29257 19901 29291
rect 19901 29257 19935 29291
rect 19935 29257 19944 29291
rect 19892 29248 19944 29257
rect 20996 29291 21048 29300
rect 20996 29257 21005 29291
rect 21005 29257 21039 29291
rect 21039 29257 21048 29291
rect 20996 29248 21048 29257
rect 21824 29248 21876 29300
rect 13912 29180 13964 29232
rect 13636 29112 13688 29164
rect 13268 28908 13320 28960
rect 14832 29112 14884 29164
rect 15108 29112 15160 29164
rect 13820 29044 13872 29096
rect 13820 28908 13872 28960
rect 14648 29044 14700 29096
rect 14924 29087 14976 29096
rect 14924 29053 14933 29087
rect 14933 29053 14967 29087
rect 14967 29053 14976 29087
rect 14924 29044 14976 29053
rect 17224 29180 17276 29232
rect 15752 29044 15804 29096
rect 16580 29044 16632 29096
rect 14924 28908 14976 28960
rect 15752 28908 15804 28960
rect 16120 28951 16172 28960
rect 16120 28917 16129 28951
rect 16129 28917 16163 28951
rect 16163 28917 16172 28951
rect 16120 28908 16172 28917
rect 17040 29112 17092 29164
rect 17408 29112 17460 29164
rect 18696 29180 18748 29232
rect 18880 29223 18932 29232
rect 18880 29189 18889 29223
rect 18889 29189 18923 29223
rect 18923 29189 18932 29223
rect 18880 29180 18932 29189
rect 19064 29180 19116 29232
rect 19340 29223 19392 29232
rect 19340 29189 19349 29223
rect 19349 29189 19383 29223
rect 19383 29189 19392 29223
rect 19340 29180 19392 29189
rect 17224 29044 17276 29096
rect 18420 29112 18472 29164
rect 17776 29044 17828 29096
rect 18696 29044 18748 29096
rect 19432 29087 19484 29096
rect 19432 29053 19441 29087
rect 19441 29053 19475 29087
rect 19475 29053 19484 29087
rect 19432 29044 19484 29053
rect 17040 29019 17092 29028
rect 17040 28985 17049 29019
rect 17049 28985 17083 29019
rect 17083 28985 17092 29019
rect 17040 28976 17092 28985
rect 18880 28976 18932 29028
rect 19432 28908 19484 28960
rect 10982 28806 11034 28858
rect 11046 28806 11098 28858
rect 11110 28806 11162 28858
rect 11174 28806 11226 28858
rect 20982 28806 21034 28858
rect 21046 28806 21098 28858
rect 21110 28806 21162 28858
rect 21174 28806 21226 28858
rect 5540 28747 5592 28756
rect 5540 28713 5549 28747
rect 5549 28713 5583 28747
rect 5583 28713 5592 28747
rect 5540 28704 5592 28713
rect 6184 28747 6236 28756
rect 6184 28713 6193 28747
rect 6193 28713 6227 28747
rect 6227 28713 6236 28747
rect 6184 28704 6236 28713
rect 6552 28747 6604 28756
rect 6552 28713 6561 28747
rect 6561 28713 6595 28747
rect 6595 28713 6604 28747
rect 6552 28704 6604 28713
rect 9404 28747 9456 28756
rect 9404 28713 9413 28747
rect 9413 28713 9447 28747
rect 9447 28713 9456 28747
rect 9404 28704 9456 28713
rect 9680 28747 9732 28756
rect 9680 28713 9689 28747
rect 9689 28713 9723 28747
rect 9723 28713 9732 28747
rect 9680 28704 9732 28713
rect 11428 28704 11480 28756
rect 9128 28679 9180 28688
rect 9128 28645 9137 28679
rect 9137 28645 9171 28679
rect 9171 28645 9180 28679
rect 9128 28636 9180 28645
rect 1400 28611 1452 28620
rect 1400 28577 1409 28611
rect 1409 28577 1443 28611
rect 1443 28577 1452 28611
rect 1400 28568 1452 28577
rect 5724 28611 5776 28620
rect 5724 28577 5733 28611
rect 5733 28577 5767 28611
rect 5767 28577 5776 28611
rect 5724 28568 5776 28577
rect 8484 28568 8536 28620
rect 9220 28568 9272 28620
rect 9404 28568 9456 28620
rect 11612 28636 11664 28688
rect 11520 28568 11572 28620
rect 12532 28704 12584 28756
rect 12348 28636 12400 28688
rect 13084 28704 13136 28756
rect 13176 28704 13228 28756
rect 15384 28704 15436 28756
rect 15752 28704 15804 28756
rect 16304 28747 16356 28756
rect 16304 28713 16313 28747
rect 16313 28713 16347 28747
rect 16347 28713 16356 28747
rect 16304 28704 16356 28713
rect 16580 28704 16632 28756
rect 13268 28636 13320 28688
rect 15292 28636 15344 28688
rect 12716 28611 12768 28620
rect 12716 28577 12725 28611
rect 12725 28577 12759 28611
rect 12759 28577 12768 28611
rect 12716 28568 12768 28577
rect 13728 28568 13780 28620
rect 14556 28568 14608 28620
rect 14924 28611 14976 28620
rect 14924 28577 14933 28611
rect 14933 28577 14967 28611
rect 14967 28577 14976 28611
rect 14924 28568 14976 28577
rect 16028 28636 16080 28688
rect 1584 28500 1636 28552
rect 7840 28500 7892 28552
rect 7932 28432 7984 28484
rect 8392 28500 8444 28552
rect 11428 28543 11480 28552
rect 11428 28509 11437 28543
rect 11437 28509 11471 28543
rect 11471 28509 11480 28543
rect 11428 28500 11480 28509
rect 11612 28500 11664 28552
rect 11704 28500 11756 28552
rect 13268 28543 13320 28552
rect 13268 28509 13277 28543
rect 13277 28509 13311 28543
rect 13311 28509 13320 28543
rect 13268 28500 13320 28509
rect 13820 28500 13872 28552
rect 15384 28500 15436 28552
rect 9496 28432 9548 28484
rect 10416 28432 10468 28484
rect 13360 28432 13412 28484
rect 14372 28432 14424 28484
rect 14924 28432 14976 28484
rect 16396 28568 16448 28620
rect 15660 28500 15712 28552
rect 15936 28432 15988 28484
rect 16120 28432 16172 28484
rect 17040 28636 17092 28688
rect 17224 28636 17276 28688
rect 16856 28500 16908 28552
rect 17224 28543 17276 28552
rect 17224 28509 17233 28543
rect 17233 28509 17267 28543
rect 17267 28509 17276 28543
rect 17224 28500 17276 28509
rect 17592 28500 17644 28552
rect 18696 28704 18748 28756
rect 18880 28747 18932 28756
rect 18880 28713 18889 28747
rect 18889 28713 18923 28747
rect 18923 28713 18932 28747
rect 18880 28704 18932 28713
rect 19340 28747 19392 28756
rect 19340 28713 19349 28747
rect 19349 28713 19383 28747
rect 19383 28713 19392 28747
rect 19340 28704 19392 28713
rect 20076 28704 20128 28756
rect 20352 28747 20404 28756
rect 20352 28713 20361 28747
rect 20361 28713 20395 28747
rect 20395 28713 20404 28747
rect 20352 28704 20404 28713
rect 17960 28568 18012 28620
rect 18512 28568 18564 28620
rect 19432 28611 19484 28620
rect 19432 28577 19441 28611
rect 19441 28577 19475 28611
rect 19475 28577 19484 28611
rect 19432 28568 19484 28577
rect 4068 28364 4120 28416
rect 8208 28364 8260 28416
rect 9772 28364 9824 28416
rect 13912 28364 13964 28416
rect 16580 28364 16632 28416
rect 17040 28364 17092 28416
rect 18052 28364 18104 28416
rect 19616 28407 19668 28416
rect 19616 28373 19625 28407
rect 19625 28373 19659 28407
rect 19659 28373 19668 28407
rect 19616 28364 19668 28373
rect 22560 28364 22612 28416
rect 5982 28262 6034 28314
rect 6046 28262 6098 28314
rect 6110 28262 6162 28314
rect 6174 28262 6226 28314
rect 15982 28262 16034 28314
rect 16046 28262 16098 28314
rect 16110 28262 16162 28314
rect 16174 28262 16226 28314
rect 25982 28262 26034 28314
rect 26046 28262 26098 28314
rect 26110 28262 26162 28314
rect 26174 28262 26226 28314
rect 3148 28203 3200 28212
rect 3148 28169 3157 28203
rect 3157 28169 3191 28203
rect 3191 28169 3200 28203
rect 3148 28160 3200 28169
rect 7288 28160 7340 28212
rect 7840 28160 7892 28212
rect 8392 28160 8444 28212
rect 8944 28203 8996 28212
rect 8668 28092 8720 28144
rect 8944 28169 8953 28203
rect 8953 28169 8987 28203
rect 8987 28169 8996 28203
rect 8944 28160 8996 28169
rect 1400 28024 1452 28076
rect 6828 28024 6880 28076
rect 1860 27999 1912 28008
rect 1860 27965 1869 27999
rect 1869 27965 1903 27999
rect 1903 27965 1912 27999
rect 1860 27956 1912 27965
rect 7104 27956 7156 28008
rect 9312 27956 9364 28008
rect 9864 28092 9916 28144
rect 12532 28160 12584 28212
rect 13728 28203 13780 28212
rect 13728 28169 13737 28203
rect 13737 28169 13771 28203
rect 13771 28169 13780 28203
rect 13728 28160 13780 28169
rect 14096 28160 14148 28212
rect 14372 28160 14424 28212
rect 12440 28092 12492 28144
rect 10324 28024 10376 28076
rect 5724 27888 5776 27940
rect 6460 27888 6512 27940
rect 9220 27888 9272 27940
rect 9680 27999 9732 28008
rect 9680 27965 9689 27999
rect 9689 27965 9723 27999
rect 9723 27965 9732 27999
rect 10048 27999 10100 28008
rect 9680 27956 9732 27965
rect 10048 27965 10057 27999
rect 10057 27965 10091 27999
rect 10091 27965 10100 27999
rect 10048 27956 10100 27965
rect 10692 27956 10744 28008
rect 12440 27999 12492 28008
rect 12440 27965 12449 27999
rect 12449 27965 12483 27999
rect 12483 27965 12492 27999
rect 12440 27956 12492 27965
rect 12716 28092 12768 28144
rect 16396 28203 16448 28212
rect 16396 28169 16405 28203
rect 16405 28169 16439 28203
rect 16439 28169 16448 28203
rect 16396 28160 16448 28169
rect 16764 28203 16816 28212
rect 16764 28169 16773 28203
rect 16773 28169 16807 28203
rect 16807 28169 16816 28203
rect 16764 28160 16816 28169
rect 17224 28160 17276 28212
rect 19432 28203 19484 28212
rect 19432 28169 19441 28203
rect 19441 28169 19475 28203
rect 19475 28169 19484 28203
rect 19432 28160 19484 28169
rect 20352 28160 20404 28212
rect 21548 28203 21600 28212
rect 21548 28169 21557 28203
rect 21557 28169 21591 28203
rect 21591 28169 21600 28203
rect 21548 28160 21600 28169
rect 14924 28092 14976 28144
rect 14096 28024 14148 28076
rect 15568 28024 15620 28076
rect 13176 27999 13228 28008
rect 6828 27820 6880 27872
rect 8208 27863 8260 27872
rect 8208 27829 8217 27863
rect 8217 27829 8251 27863
rect 8251 27829 8260 27863
rect 8208 27820 8260 27829
rect 8484 27820 8536 27872
rect 9772 27888 9824 27940
rect 9864 27888 9916 27940
rect 10140 27888 10192 27940
rect 13176 27965 13185 27999
rect 13185 27965 13219 27999
rect 13219 27965 13228 27999
rect 13176 27956 13228 27965
rect 14004 27956 14056 28008
rect 13084 27888 13136 27940
rect 14372 27956 14424 28008
rect 14924 27999 14976 28008
rect 14924 27965 14933 27999
rect 14933 27965 14967 27999
rect 14967 27965 14976 27999
rect 14924 27956 14976 27965
rect 15108 27956 15160 28008
rect 15936 27956 15988 28008
rect 16212 27999 16264 28008
rect 16212 27965 16221 27999
rect 16221 27965 16255 27999
rect 16255 27965 16264 27999
rect 16212 27956 16264 27965
rect 17592 28024 17644 28076
rect 18236 28092 18288 28144
rect 20720 28135 20772 28144
rect 20720 28101 20729 28135
rect 20729 28101 20763 28135
rect 20763 28101 20772 28135
rect 20720 28092 20772 28101
rect 17960 27956 18012 28008
rect 18696 27999 18748 28008
rect 15568 27888 15620 27940
rect 9680 27820 9732 27872
rect 11704 27820 11756 27872
rect 14372 27820 14424 27872
rect 15384 27820 15436 27872
rect 16672 27888 16724 27940
rect 18696 27965 18705 27999
rect 18705 27965 18739 27999
rect 18739 27965 18748 27999
rect 18696 27956 18748 27965
rect 18788 27956 18840 28008
rect 19984 28024 20036 28076
rect 21916 28024 21968 28076
rect 23388 28024 23440 28076
rect 20720 27956 20772 28008
rect 22560 27999 22612 28008
rect 22560 27965 22569 27999
rect 22569 27965 22603 27999
rect 22603 27965 22612 27999
rect 22560 27956 22612 27965
rect 23664 27956 23716 28008
rect 19248 27888 19300 27940
rect 21824 27931 21876 27940
rect 21824 27897 21833 27931
rect 21833 27897 21867 27931
rect 21867 27897 21876 27931
rect 21824 27888 21876 27897
rect 20076 27863 20128 27872
rect 20076 27829 20085 27863
rect 20085 27829 20119 27863
rect 20119 27829 20128 27863
rect 20076 27820 20128 27829
rect 10982 27718 11034 27770
rect 11046 27718 11098 27770
rect 11110 27718 11162 27770
rect 11174 27718 11226 27770
rect 20982 27718 21034 27770
rect 21046 27718 21098 27770
rect 21110 27718 21162 27770
rect 21174 27718 21226 27770
rect 1400 27616 1452 27668
rect 7380 27659 7432 27668
rect 7380 27625 7389 27659
rect 7389 27625 7423 27659
rect 7423 27625 7432 27659
rect 7380 27616 7432 27625
rect 8208 27616 8260 27668
rect 13360 27659 13412 27668
rect 4620 27591 4672 27600
rect 4620 27557 4629 27591
rect 4629 27557 4663 27591
rect 4663 27557 4672 27591
rect 4620 27548 4672 27557
rect 8484 27548 8536 27600
rect 9588 27548 9640 27600
rect 13360 27625 13369 27659
rect 13369 27625 13403 27659
rect 13403 27625 13412 27659
rect 13360 27616 13412 27625
rect 13912 27616 13964 27668
rect 14464 27659 14516 27668
rect 14464 27625 14473 27659
rect 14473 27625 14507 27659
rect 14507 27625 14516 27659
rect 14464 27616 14516 27625
rect 15108 27616 15160 27668
rect 15292 27616 15344 27668
rect 16212 27616 16264 27668
rect 17592 27616 17644 27668
rect 18512 27659 18564 27668
rect 18512 27625 18521 27659
rect 18521 27625 18555 27659
rect 18555 27625 18564 27659
rect 18512 27616 18564 27625
rect 18788 27616 18840 27668
rect 7932 27523 7984 27532
rect 7932 27489 7941 27523
rect 7941 27489 7975 27523
rect 7975 27489 7984 27523
rect 7932 27480 7984 27489
rect 8392 27480 8444 27532
rect 10416 27523 10468 27532
rect 10416 27489 10425 27523
rect 10425 27489 10459 27523
rect 10459 27489 10468 27523
rect 10416 27480 10468 27489
rect 11060 27548 11112 27600
rect 12072 27523 12124 27532
rect 12072 27489 12081 27523
rect 12081 27489 12115 27523
rect 12115 27489 12124 27523
rect 12072 27480 12124 27489
rect 14556 27548 14608 27600
rect 15476 27548 15528 27600
rect 16304 27548 16356 27600
rect 16396 27548 16448 27600
rect 20720 27548 20772 27600
rect 20812 27548 20864 27600
rect 21916 27548 21968 27600
rect 13912 27523 13964 27532
rect 13912 27489 13921 27523
rect 13921 27489 13955 27523
rect 13955 27489 13964 27523
rect 13912 27480 13964 27489
rect 14464 27480 14516 27532
rect 14648 27480 14700 27532
rect 16672 27523 16724 27532
rect 16672 27489 16681 27523
rect 16681 27489 16715 27523
rect 16715 27489 16724 27523
rect 16672 27480 16724 27489
rect 17592 27480 17644 27532
rect 17776 27480 17828 27532
rect 18880 27523 18932 27532
rect 5080 27455 5132 27464
rect 5080 27421 5089 27455
rect 5089 27421 5123 27455
rect 5123 27421 5132 27455
rect 5080 27412 5132 27421
rect 7288 27412 7340 27464
rect 7840 27412 7892 27464
rect 9036 27412 9088 27464
rect 11428 27412 11480 27464
rect 10324 27344 10376 27396
rect 13176 27412 13228 27464
rect 18052 27412 18104 27464
rect 12440 27344 12492 27396
rect 18880 27489 18889 27523
rect 18889 27489 18923 27523
rect 18923 27489 18932 27523
rect 18880 27480 18932 27489
rect 20076 27523 20128 27532
rect 20076 27489 20085 27523
rect 20085 27489 20119 27523
rect 20119 27489 20128 27523
rect 20076 27480 20128 27489
rect 19340 27412 19392 27464
rect 1584 27319 1636 27328
rect 1584 27285 1593 27319
rect 1593 27285 1627 27319
rect 1627 27285 1636 27319
rect 1584 27276 1636 27285
rect 1860 27276 1912 27328
rect 5724 27276 5776 27328
rect 9220 27276 9272 27328
rect 9496 27276 9548 27328
rect 10968 27276 11020 27328
rect 11612 27276 11664 27328
rect 12348 27276 12400 27328
rect 13728 27319 13780 27328
rect 13728 27285 13737 27319
rect 13737 27285 13771 27319
rect 13771 27285 13780 27319
rect 13728 27276 13780 27285
rect 14924 27276 14976 27328
rect 15108 27276 15160 27328
rect 15292 27276 15344 27328
rect 16304 27319 16356 27328
rect 16304 27285 16313 27319
rect 16313 27285 16347 27319
rect 16347 27285 16356 27319
rect 16304 27276 16356 27285
rect 17040 27276 17092 27328
rect 17776 27319 17828 27328
rect 17776 27285 17785 27319
rect 17785 27285 17819 27319
rect 17819 27285 17828 27319
rect 17776 27276 17828 27285
rect 19892 27276 19944 27328
rect 20812 27412 20864 27464
rect 5982 27174 6034 27226
rect 6046 27174 6098 27226
rect 6110 27174 6162 27226
rect 6174 27174 6226 27226
rect 15982 27174 16034 27226
rect 16046 27174 16098 27226
rect 16110 27174 16162 27226
rect 16174 27174 16226 27226
rect 25982 27174 26034 27226
rect 26046 27174 26098 27226
rect 26110 27174 26162 27226
rect 26174 27174 26226 27226
rect 1400 27072 1452 27124
rect 7840 27072 7892 27124
rect 7932 27072 7984 27124
rect 8852 27072 8904 27124
rect 8392 27004 8444 27056
rect 6644 26936 6696 26988
rect 4712 26911 4764 26920
rect 4712 26877 4721 26911
rect 4721 26877 4755 26911
rect 4755 26877 4764 26911
rect 4712 26868 4764 26877
rect 5080 26868 5132 26920
rect 5356 26911 5408 26920
rect 5356 26877 5365 26911
rect 5365 26877 5399 26911
rect 5399 26877 5408 26911
rect 5356 26868 5408 26877
rect 5724 26911 5776 26920
rect 5724 26877 5733 26911
rect 5733 26877 5767 26911
rect 5767 26877 5776 26911
rect 5724 26868 5776 26877
rect 6368 26868 6420 26920
rect 6920 26911 6972 26920
rect 6920 26877 6929 26911
rect 6929 26877 6963 26911
rect 6963 26877 6972 26911
rect 6920 26868 6972 26877
rect 8852 26868 8904 26920
rect 9220 26868 9272 26920
rect 9588 26911 9640 26920
rect 9588 26877 9616 26911
rect 9616 26877 9640 26911
rect 9588 26868 9640 26877
rect 10876 27072 10928 27124
rect 12072 27072 12124 27124
rect 12808 27072 12860 27124
rect 13360 27072 13412 27124
rect 15568 27072 15620 27124
rect 15752 27072 15804 27124
rect 16396 27072 16448 27124
rect 19524 27072 19576 27124
rect 19800 27072 19852 27124
rect 20076 27115 20128 27124
rect 20076 27081 20085 27115
rect 20085 27081 20119 27115
rect 20119 27081 20128 27115
rect 20076 27072 20128 27081
rect 13912 27047 13964 27056
rect 13912 27013 13921 27047
rect 13921 27013 13955 27047
rect 13955 27013 13964 27047
rect 13912 27004 13964 27013
rect 15108 27004 15160 27056
rect 13544 26936 13596 26988
rect 16580 26936 16632 26988
rect 18420 26936 18472 26988
rect 3332 26732 3384 26784
rect 9220 26775 9272 26784
rect 9220 26741 9229 26775
rect 9229 26741 9263 26775
rect 9263 26741 9272 26775
rect 9220 26732 9272 26741
rect 9588 26732 9640 26784
rect 11060 26868 11112 26920
rect 12624 26911 12676 26920
rect 12624 26877 12633 26911
rect 12633 26877 12667 26911
rect 12667 26877 12676 26911
rect 12624 26868 12676 26877
rect 13728 26868 13780 26920
rect 14004 26868 14056 26920
rect 15016 26911 15068 26920
rect 12808 26843 12860 26852
rect 11520 26775 11572 26784
rect 11520 26741 11529 26775
rect 11529 26741 11563 26775
rect 11563 26741 11572 26775
rect 11520 26732 11572 26741
rect 11704 26732 11756 26784
rect 12256 26775 12308 26784
rect 12256 26741 12265 26775
rect 12265 26741 12299 26775
rect 12299 26741 12308 26775
rect 12808 26809 12817 26843
rect 12817 26809 12851 26843
rect 12851 26809 12860 26843
rect 12808 26800 12860 26809
rect 13544 26800 13596 26852
rect 15016 26877 15025 26911
rect 15025 26877 15059 26911
rect 15059 26877 15068 26911
rect 15016 26868 15068 26877
rect 15476 26911 15528 26920
rect 15476 26877 15485 26911
rect 15485 26877 15519 26911
rect 15519 26877 15528 26911
rect 15476 26868 15528 26877
rect 17224 26911 17276 26920
rect 15108 26800 15160 26852
rect 12716 26775 12768 26784
rect 12256 26732 12308 26741
rect 12716 26741 12725 26775
rect 12725 26741 12759 26775
rect 12759 26741 12768 26775
rect 12716 26732 12768 26741
rect 14280 26732 14332 26784
rect 17224 26877 17233 26911
rect 17233 26877 17267 26911
rect 17267 26877 17276 26911
rect 17224 26868 17276 26877
rect 18052 26911 18104 26920
rect 18052 26877 18061 26911
rect 18061 26877 18095 26911
rect 18095 26877 18104 26911
rect 18052 26868 18104 26877
rect 18696 26868 18748 26920
rect 19156 26868 19208 26920
rect 16948 26843 17000 26852
rect 16948 26809 16957 26843
rect 16957 26809 16991 26843
rect 16991 26809 17000 26843
rect 16948 26800 17000 26809
rect 10982 26630 11034 26682
rect 11046 26630 11098 26682
rect 11110 26630 11162 26682
rect 11174 26630 11226 26682
rect 20982 26630 21034 26682
rect 21046 26630 21098 26682
rect 21110 26630 21162 26682
rect 21174 26630 21226 26682
rect 6920 26528 6972 26580
rect 7104 26528 7156 26580
rect 8116 26571 8168 26580
rect 8116 26537 8125 26571
rect 8125 26537 8159 26571
rect 8159 26537 8168 26571
rect 8116 26528 8168 26537
rect 8760 26571 8812 26580
rect 8760 26537 8769 26571
rect 8769 26537 8803 26571
rect 8803 26537 8812 26571
rect 8760 26528 8812 26537
rect 9404 26528 9456 26580
rect 11520 26528 11572 26580
rect 3056 26503 3108 26512
rect 3056 26469 3065 26503
rect 3065 26469 3099 26503
rect 3099 26469 3108 26503
rect 3056 26460 3108 26469
rect 8668 26460 8720 26512
rect 9956 26460 10008 26512
rect 12716 26528 12768 26580
rect 13176 26528 13228 26580
rect 14004 26528 14056 26580
rect 14832 26571 14884 26580
rect 14832 26537 14841 26571
rect 14841 26537 14875 26571
rect 14875 26537 14884 26571
rect 14832 26528 14884 26537
rect 16488 26528 16540 26580
rect 16856 26571 16908 26580
rect 16856 26537 16865 26571
rect 16865 26537 16899 26571
rect 16899 26537 16908 26571
rect 16856 26528 16908 26537
rect 16948 26528 17000 26580
rect 18880 26571 18932 26580
rect 18880 26537 18889 26571
rect 18889 26537 18923 26571
rect 18923 26537 18932 26571
rect 18880 26528 18932 26537
rect 1400 26435 1452 26444
rect 1400 26401 1409 26435
rect 1409 26401 1443 26435
rect 1443 26401 1452 26435
rect 1400 26392 1452 26401
rect 2136 26392 2188 26444
rect 4620 26392 4672 26444
rect 5632 26392 5684 26444
rect 10324 26435 10376 26444
rect 10324 26401 10333 26435
rect 10333 26401 10367 26435
rect 10367 26401 10376 26435
rect 10324 26392 10376 26401
rect 10508 26435 10560 26444
rect 10508 26401 10517 26435
rect 10517 26401 10551 26435
rect 10551 26401 10560 26435
rect 10508 26392 10560 26401
rect 12440 26460 12492 26512
rect 12348 26392 12400 26444
rect 1676 26367 1728 26376
rect 1676 26333 1685 26367
rect 1685 26333 1719 26367
rect 1719 26333 1728 26367
rect 1676 26324 1728 26333
rect 5172 26324 5224 26376
rect 7012 26324 7064 26376
rect 8208 26324 8260 26376
rect 8668 26324 8720 26376
rect 9128 26324 9180 26376
rect 9404 26324 9456 26376
rect 10416 26324 10468 26376
rect 3332 26256 3384 26308
rect 5080 26299 5132 26308
rect 5080 26265 5089 26299
rect 5089 26265 5123 26299
rect 5123 26265 5132 26299
rect 5080 26256 5132 26265
rect 7288 26299 7340 26308
rect 7288 26265 7297 26299
rect 7297 26265 7331 26299
rect 7331 26265 7340 26299
rect 7288 26256 7340 26265
rect 10600 26324 10652 26376
rect 11244 26367 11296 26376
rect 11244 26333 11253 26367
rect 11253 26333 11287 26367
rect 11287 26333 11296 26367
rect 11244 26324 11296 26333
rect 11428 26324 11480 26376
rect 12164 26324 12216 26376
rect 12256 26324 12308 26376
rect 11612 26256 11664 26308
rect 11888 26256 11940 26308
rect 5264 26188 5316 26240
rect 5724 26188 5776 26240
rect 9220 26188 9272 26240
rect 9588 26188 9640 26240
rect 10876 26188 10928 26240
rect 12624 26392 12676 26444
rect 13360 26460 13412 26512
rect 13544 26460 13596 26512
rect 15476 26460 15528 26512
rect 17960 26460 18012 26512
rect 18144 26503 18196 26512
rect 18144 26469 18153 26503
rect 18153 26469 18187 26503
rect 18187 26469 18196 26503
rect 18144 26460 18196 26469
rect 18236 26460 18288 26512
rect 13268 26392 13320 26444
rect 15568 26392 15620 26444
rect 13360 26324 13412 26376
rect 15476 26324 15528 26376
rect 16672 26392 16724 26444
rect 17776 26392 17828 26444
rect 15844 26324 15896 26376
rect 16304 26324 16356 26376
rect 17592 26324 17644 26376
rect 16948 26256 17000 26308
rect 17500 26256 17552 26308
rect 12716 26188 12768 26240
rect 15016 26188 15068 26240
rect 16672 26188 16724 26240
rect 25136 26188 25188 26240
rect 25320 26188 25372 26240
rect 5982 26086 6034 26138
rect 6046 26086 6098 26138
rect 6110 26086 6162 26138
rect 6174 26086 6226 26138
rect 15982 26086 16034 26138
rect 16046 26086 16098 26138
rect 16110 26086 16162 26138
rect 16174 26086 16226 26138
rect 25982 26086 26034 26138
rect 26046 26086 26098 26138
rect 26110 26086 26162 26138
rect 26174 26086 26226 26138
rect 1676 26027 1728 26036
rect 1676 25993 1685 26027
rect 1685 25993 1719 26027
rect 1719 25993 1728 26027
rect 1676 25984 1728 25993
rect 2136 25984 2188 26036
rect 6644 26027 6696 26036
rect 6644 25993 6653 26027
rect 6653 25993 6687 26027
rect 6687 25993 6696 26027
rect 6644 25984 6696 25993
rect 7196 26027 7248 26036
rect 7196 25993 7205 26027
rect 7205 25993 7239 26027
rect 7239 25993 7248 26027
rect 7196 25984 7248 25993
rect 8576 25984 8628 26036
rect 10692 26027 10744 26036
rect 10692 25993 10701 26027
rect 10701 25993 10735 26027
rect 10735 25993 10744 26027
rect 10692 25984 10744 25993
rect 9128 25916 9180 25968
rect 10140 25959 10192 25968
rect 10140 25925 10149 25959
rect 10149 25925 10183 25959
rect 10183 25925 10192 25959
rect 10140 25916 10192 25925
rect 10600 25916 10652 25968
rect 11244 25984 11296 26036
rect 13544 25984 13596 26036
rect 14464 25984 14516 26036
rect 17776 26027 17828 26036
rect 11704 25916 11756 25968
rect 14740 25916 14792 25968
rect 11888 25848 11940 25900
rect 12624 25848 12676 25900
rect 13268 25891 13320 25900
rect 13268 25857 13277 25891
rect 13277 25857 13311 25891
rect 13311 25857 13320 25891
rect 13268 25848 13320 25857
rect 13636 25848 13688 25900
rect 14004 25848 14056 25900
rect 15108 25891 15160 25900
rect 15108 25857 15117 25891
rect 15117 25857 15151 25891
rect 15151 25857 15160 25891
rect 15108 25848 15160 25857
rect 17776 25993 17785 26027
rect 17785 25993 17819 26027
rect 17819 25993 17828 26027
rect 17776 25984 17828 25993
rect 18420 25984 18472 26036
rect 18696 26027 18748 26036
rect 18696 25993 18705 26027
rect 18705 25993 18739 26027
rect 18739 25993 18748 26027
rect 18696 25984 18748 25993
rect 4160 25780 4212 25832
rect 5172 25823 5224 25832
rect 5172 25789 5181 25823
rect 5181 25789 5215 25823
rect 5215 25789 5224 25823
rect 5172 25780 5224 25789
rect 5356 25823 5408 25832
rect 5356 25789 5365 25823
rect 5365 25789 5399 25823
rect 5399 25789 5408 25823
rect 5356 25780 5408 25789
rect 5724 25823 5776 25832
rect 5724 25789 5733 25823
rect 5733 25789 5767 25823
rect 5767 25789 5776 25823
rect 5724 25780 5776 25789
rect 6368 25780 6420 25832
rect 9220 25780 9272 25832
rect 10876 25712 10928 25764
rect 11152 25755 11204 25764
rect 11152 25721 11161 25755
rect 11161 25721 11195 25755
rect 11195 25721 11204 25755
rect 12256 25780 12308 25832
rect 12992 25823 13044 25832
rect 12992 25789 13001 25823
rect 13001 25789 13035 25823
rect 13035 25789 13044 25823
rect 12992 25780 13044 25789
rect 16672 25780 16724 25832
rect 16856 25780 16908 25832
rect 11152 25712 11204 25721
rect 14556 25755 14608 25764
rect 14556 25721 14565 25755
rect 14565 25721 14599 25755
rect 14599 25721 14608 25755
rect 14556 25712 14608 25721
rect 14740 25755 14792 25764
rect 14740 25721 14749 25755
rect 14749 25721 14783 25755
rect 14783 25721 14792 25755
rect 14740 25712 14792 25721
rect 16028 25712 16080 25764
rect 17776 25712 17828 25764
rect 8392 25644 8444 25696
rect 10692 25644 10744 25696
rect 11520 25644 11572 25696
rect 14832 25644 14884 25696
rect 15476 25687 15528 25696
rect 15476 25653 15485 25687
rect 15485 25653 15519 25687
rect 15519 25653 15528 25687
rect 15476 25644 15528 25653
rect 16212 25687 16264 25696
rect 16212 25653 16221 25687
rect 16221 25653 16255 25687
rect 16255 25653 16264 25687
rect 16212 25644 16264 25653
rect 16304 25644 16356 25696
rect 16764 25644 16816 25696
rect 17592 25644 17644 25696
rect 18236 25644 18288 25696
rect 10982 25542 11034 25594
rect 11046 25542 11098 25594
rect 11110 25542 11162 25594
rect 11174 25542 11226 25594
rect 20982 25542 21034 25594
rect 21046 25542 21098 25594
rect 21110 25542 21162 25594
rect 21174 25542 21226 25594
rect 1676 25483 1728 25492
rect 1676 25449 1685 25483
rect 1685 25449 1719 25483
rect 1719 25449 1728 25483
rect 1676 25440 1728 25449
rect 5632 25483 5684 25492
rect 5632 25449 5641 25483
rect 5641 25449 5675 25483
rect 5675 25449 5684 25483
rect 5632 25440 5684 25449
rect 7104 25440 7156 25492
rect 9128 25483 9180 25492
rect 9128 25449 9137 25483
rect 9137 25449 9171 25483
rect 9171 25449 9180 25483
rect 9128 25440 9180 25449
rect 9588 25440 9640 25492
rect 9956 25483 10008 25492
rect 9956 25449 9965 25483
rect 9965 25449 9999 25483
rect 9999 25449 10008 25483
rect 9956 25440 10008 25449
rect 10692 25440 10744 25492
rect 10876 25483 10928 25492
rect 10876 25449 10885 25483
rect 10885 25449 10919 25483
rect 10919 25449 10928 25483
rect 10876 25440 10928 25449
rect 11336 25440 11388 25492
rect 12256 25440 12308 25492
rect 14924 25483 14976 25492
rect 1768 25372 1820 25424
rect 1400 25347 1452 25356
rect 1400 25313 1409 25347
rect 1409 25313 1443 25347
rect 1443 25313 1452 25347
rect 1400 25304 1452 25313
rect 1952 25304 2004 25356
rect 14924 25449 14933 25483
rect 14933 25449 14967 25483
rect 14967 25449 14976 25483
rect 14924 25440 14976 25449
rect 15568 25483 15620 25492
rect 15568 25449 15577 25483
rect 15577 25449 15611 25483
rect 15611 25449 15620 25483
rect 15568 25440 15620 25449
rect 16028 25483 16080 25492
rect 16028 25449 16037 25483
rect 16037 25449 16071 25483
rect 16071 25449 16080 25483
rect 16028 25440 16080 25449
rect 9312 25304 9364 25356
rect 9588 25304 9640 25356
rect 10048 25304 10100 25356
rect 10508 25304 10560 25356
rect 10876 25304 10928 25356
rect 11704 25347 11756 25356
rect 11704 25313 11713 25347
rect 11713 25313 11747 25347
rect 11747 25313 11756 25347
rect 11704 25304 11756 25313
rect 12072 25347 12124 25356
rect 12072 25313 12081 25347
rect 12081 25313 12115 25347
rect 12115 25313 12124 25347
rect 12072 25304 12124 25313
rect 12256 25347 12308 25356
rect 12256 25313 12265 25347
rect 12265 25313 12299 25347
rect 12299 25313 12308 25347
rect 12256 25304 12308 25313
rect 12716 25304 12768 25356
rect 14004 25372 14056 25424
rect 8392 25236 8444 25288
rect 9864 25236 9916 25288
rect 13820 25279 13872 25288
rect 13820 25245 13829 25279
rect 13829 25245 13863 25279
rect 13863 25245 13872 25279
rect 13820 25236 13872 25245
rect 16764 25304 16816 25356
rect 16396 25279 16448 25288
rect 16396 25245 16405 25279
rect 16405 25245 16439 25279
rect 16439 25245 16448 25279
rect 16396 25236 16448 25245
rect 5172 25168 5224 25220
rect 8852 25168 8904 25220
rect 13268 25168 13320 25220
rect 5356 25100 5408 25152
rect 6644 25100 6696 25152
rect 8300 25100 8352 25152
rect 10600 25100 10652 25152
rect 11520 25100 11572 25152
rect 11980 25100 12032 25152
rect 13360 25143 13412 25152
rect 13360 25109 13369 25143
rect 13369 25109 13403 25143
rect 13403 25109 13412 25143
rect 13360 25100 13412 25109
rect 13544 25100 13596 25152
rect 13728 25143 13780 25152
rect 13728 25109 13737 25143
rect 13737 25109 13771 25143
rect 13771 25109 13780 25143
rect 13728 25100 13780 25109
rect 16580 25100 16632 25152
rect 16856 25100 16908 25152
rect 5982 24998 6034 25050
rect 6046 24998 6098 25050
rect 6110 24998 6162 25050
rect 6174 24998 6226 25050
rect 15982 24998 16034 25050
rect 16046 24998 16098 25050
rect 16110 24998 16162 25050
rect 16174 24998 16226 25050
rect 25982 24998 26034 25050
rect 26046 24998 26098 25050
rect 26110 24998 26162 25050
rect 26174 24998 26226 25050
rect 10508 24896 10560 24948
rect 11888 24939 11940 24948
rect 11888 24905 11897 24939
rect 11897 24905 11931 24939
rect 11931 24905 11940 24939
rect 11888 24896 11940 24905
rect 14464 24896 14516 24948
rect 16580 24939 16632 24948
rect 16580 24905 16589 24939
rect 16589 24905 16623 24939
rect 16623 24905 16632 24939
rect 16580 24896 16632 24905
rect 16764 24896 16816 24948
rect 18144 24896 18196 24948
rect 18696 24896 18748 24948
rect 9220 24828 9272 24880
rect 11980 24828 12032 24880
rect 14740 24828 14792 24880
rect 2688 24692 2740 24744
rect 8116 24803 8168 24812
rect 8116 24769 8125 24803
rect 8125 24769 8159 24803
rect 8159 24769 8168 24803
rect 8116 24760 8168 24769
rect 9772 24760 9824 24812
rect 10600 24803 10652 24812
rect 10600 24769 10609 24803
rect 10609 24769 10643 24803
rect 10643 24769 10652 24803
rect 10600 24760 10652 24769
rect 13360 24803 13412 24812
rect 13360 24769 13369 24803
rect 13369 24769 13403 24803
rect 13403 24769 13412 24803
rect 13360 24760 13412 24769
rect 8208 24692 8260 24744
rect 8392 24735 8444 24744
rect 8392 24701 8401 24735
rect 8401 24701 8435 24735
rect 8435 24701 8444 24735
rect 8392 24692 8444 24701
rect 9036 24692 9088 24744
rect 10140 24692 10192 24744
rect 12716 24692 12768 24744
rect 12900 24735 12952 24744
rect 12900 24701 12909 24735
rect 12909 24701 12943 24735
rect 12943 24701 12952 24735
rect 12900 24692 12952 24701
rect 13268 24735 13320 24744
rect 13268 24701 13277 24735
rect 13277 24701 13311 24735
rect 13311 24701 13320 24735
rect 13268 24692 13320 24701
rect 14464 24692 14516 24744
rect 15292 24692 15344 24744
rect 16396 24692 16448 24744
rect 18052 24735 18104 24744
rect 1400 24624 1452 24676
rect 2964 24624 3016 24676
rect 7288 24667 7340 24676
rect 7288 24633 7297 24667
rect 7297 24633 7331 24667
rect 7331 24633 7340 24667
rect 7288 24624 7340 24633
rect 8116 24624 8168 24676
rect 12440 24667 12492 24676
rect 12440 24633 12449 24667
rect 12449 24633 12483 24667
rect 12483 24633 12492 24667
rect 12440 24624 12492 24633
rect 18052 24701 18061 24735
rect 18061 24701 18095 24735
rect 18095 24701 18104 24735
rect 18052 24692 18104 24701
rect 1952 24599 2004 24608
rect 1952 24565 1961 24599
rect 1961 24565 1995 24599
rect 1995 24565 2004 24599
rect 1952 24556 2004 24565
rect 8392 24556 8444 24608
rect 9956 24556 10008 24608
rect 10140 24556 10192 24608
rect 10508 24556 10560 24608
rect 11612 24556 11664 24608
rect 12992 24556 13044 24608
rect 13820 24556 13872 24608
rect 15568 24556 15620 24608
rect 16856 24599 16908 24608
rect 16856 24565 16865 24599
rect 16865 24565 16899 24599
rect 16899 24565 16908 24599
rect 16856 24556 16908 24565
rect 18236 24599 18288 24608
rect 18236 24565 18245 24599
rect 18245 24565 18279 24599
rect 18279 24565 18288 24599
rect 18236 24556 18288 24565
rect 10982 24454 11034 24506
rect 11046 24454 11098 24506
rect 11110 24454 11162 24506
rect 11174 24454 11226 24506
rect 20982 24454 21034 24506
rect 21046 24454 21098 24506
rect 21110 24454 21162 24506
rect 21174 24454 21226 24506
rect 7104 24395 7156 24404
rect 7104 24361 7113 24395
rect 7113 24361 7147 24395
rect 7147 24361 7156 24395
rect 7104 24352 7156 24361
rect 8392 24352 8444 24404
rect 9772 24352 9824 24404
rect 10876 24352 10928 24404
rect 12256 24352 12308 24404
rect 12532 24395 12584 24404
rect 12532 24361 12541 24395
rect 12541 24361 12575 24395
rect 12575 24361 12584 24395
rect 12532 24352 12584 24361
rect 12716 24352 12768 24404
rect 13820 24352 13872 24404
rect 14372 24352 14424 24404
rect 14924 24395 14976 24404
rect 14924 24361 14933 24395
rect 14933 24361 14967 24395
rect 14967 24361 14976 24395
rect 14924 24352 14976 24361
rect 9036 24284 9088 24336
rect 10232 24284 10284 24336
rect 10968 24284 11020 24336
rect 12900 24284 12952 24336
rect 11428 24259 11480 24268
rect 11428 24225 11437 24259
rect 11437 24225 11471 24259
rect 11471 24225 11480 24259
rect 11428 24216 11480 24225
rect 13636 24284 13688 24336
rect 14556 24284 14608 24336
rect 15108 24284 15160 24336
rect 17500 24352 17552 24404
rect 15292 24284 15344 24336
rect 13176 24259 13228 24268
rect 13176 24225 13185 24259
rect 13185 24225 13219 24259
rect 13219 24225 13228 24259
rect 13176 24216 13228 24225
rect 13268 24216 13320 24268
rect 11336 24191 11388 24200
rect 11336 24157 11345 24191
rect 11345 24157 11379 24191
rect 11379 24157 11388 24191
rect 11336 24148 11388 24157
rect 13728 24148 13780 24200
rect 14004 24148 14056 24200
rect 16304 24216 16356 24268
rect 11796 24080 11848 24132
rect 14280 24080 14332 24132
rect 19064 24216 19116 24268
rect 16856 24080 16908 24132
rect 17960 24080 18012 24132
rect 10876 24055 10928 24064
rect 10876 24021 10885 24055
rect 10885 24021 10919 24055
rect 10919 24021 10928 24055
rect 10876 24012 10928 24021
rect 14372 24012 14424 24064
rect 14924 24012 14976 24064
rect 15476 24012 15528 24064
rect 17500 24012 17552 24064
rect 5982 23910 6034 23962
rect 6046 23910 6098 23962
rect 6110 23910 6162 23962
rect 6174 23910 6226 23962
rect 15982 23910 16034 23962
rect 16046 23910 16098 23962
rect 16110 23910 16162 23962
rect 16174 23910 16226 23962
rect 25982 23910 26034 23962
rect 26046 23910 26098 23962
rect 26110 23910 26162 23962
rect 26174 23910 26226 23962
rect 7104 23851 7156 23860
rect 7104 23817 7113 23851
rect 7113 23817 7147 23851
rect 7147 23817 7156 23851
rect 7104 23808 7156 23817
rect 8576 23851 8628 23860
rect 8576 23817 8585 23851
rect 8585 23817 8619 23851
rect 8619 23817 8628 23851
rect 8576 23808 8628 23817
rect 9680 23808 9732 23860
rect 10324 23851 10376 23860
rect 10324 23817 10333 23851
rect 10333 23817 10367 23851
rect 10367 23817 10376 23851
rect 10324 23808 10376 23817
rect 10968 23808 11020 23860
rect 11428 23808 11480 23860
rect 11704 23740 11756 23792
rect 13636 23808 13688 23860
rect 14004 23808 14056 23860
rect 12256 23740 12308 23792
rect 13176 23740 13228 23792
rect 13544 23740 13596 23792
rect 16304 23808 16356 23860
rect 16396 23808 16448 23860
rect 19064 23808 19116 23860
rect 16488 23783 16540 23792
rect 16488 23749 16497 23783
rect 16497 23749 16531 23783
rect 16531 23749 16540 23783
rect 16488 23740 16540 23749
rect 12992 23715 13044 23724
rect 12992 23681 13001 23715
rect 13001 23681 13035 23715
rect 13035 23681 13044 23715
rect 12992 23672 13044 23681
rect 15292 23672 15344 23724
rect 8576 23536 8628 23588
rect 12348 23604 12400 23656
rect 14280 23647 14332 23656
rect 14280 23613 14289 23647
rect 14289 23613 14323 23647
rect 14323 23613 14332 23647
rect 14280 23604 14332 23613
rect 14372 23604 14424 23656
rect 14832 23647 14884 23656
rect 13452 23536 13504 23588
rect 14832 23613 14841 23647
rect 14841 23613 14875 23647
rect 14875 23613 14884 23647
rect 14832 23604 14884 23613
rect 14924 23604 14976 23656
rect 15292 23536 15344 23588
rect 11704 23468 11756 23520
rect 12256 23468 12308 23520
rect 14648 23468 14700 23520
rect 16304 23647 16356 23656
rect 16304 23613 16313 23647
rect 16313 23613 16347 23647
rect 16347 23613 16356 23647
rect 16304 23604 16356 23613
rect 18236 23604 18288 23656
rect 16856 23468 16908 23520
rect 17224 23468 17276 23520
rect 10982 23366 11034 23418
rect 11046 23366 11098 23418
rect 11110 23366 11162 23418
rect 11174 23366 11226 23418
rect 20982 23366 21034 23418
rect 21046 23366 21098 23418
rect 21110 23366 21162 23418
rect 21174 23366 21226 23418
rect 8484 23264 8536 23316
rect 11336 23264 11388 23316
rect 11520 23264 11572 23316
rect 12072 23307 12124 23316
rect 10784 23196 10836 23248
rect 12072 23273 12081 23307
rect 12081 23273 12115 23307
rect 12115 23273 12124 23307
rect 12072 23264 12124 23273
rect 13912 23264 13964 23316
rect 14372 23264 14424 23316
rect 14832 23264 14884 23316
rect 15108 23307 15160 23316
rect 15108 23273 15117 23307
rect 15117 23273 15151 23307
rect 15151 23273 15160 23307
rect 15108 23264 15160 23273
rect 15292 23264 15344 23316
rect 18144 23307 18196 23316
rect 12348 23196 12400 23248
rect 14556 23196 14608 23248
rect 15660 23239 15712 23248
rect 15660 23205 15669 23239
rect 15669 23205 15703 23239
rect 15703 23205 15712 23239
rect 15660 23196 15712 23205
rect 18144 23273 18153 23307
rect 18153 23273 18187 23307
rect 18187 23273 18196 23307
rect 18144 23264 18196 23273
rect 6644 23128 6696 23180
rect 6828 23171 6880 23180
rect 6828 23137 6837 23171
rect 6837 23137 6871 23171
rect 6871 23137 6880 23171
rect 6828 23128 6880 23137
rect 7196 23171 7248 23180
rect 7196 23137 7205 23171
rect 7205 23137 7239 23171
rect 7239 23137 7248 23171
rect 7196 23128 7248 23137
rect 8576 23171 8628 23180
rect 5540 23060 5592 23112
rect 6920 23103 6972 23112
rect 6920 23069 6929 23103
rect 6929 23069 6963 23103
rect 6963 23069 6972 23103
rect 6920 23060 6972 23069
rect 7288 23060 7340 23112
rect 8576 23137 8585 23171
rect 8585 23137 8619 23171
rect 8619 23137 8628 23171
rect 8576 23128 8628 23137
rect 10968 23171 11020 23180
rect 10968 23137 10977 23171
rect 10977 23137 11011 23171
rect 11011 23137 11020 23171
rect 10968 23128 11020 23137
rect 6276 22992 6328 23044
rect 9496 23060 9548 23112
rect 9956 23060 10008 23112
rect 11520 23128 11572 23180
rect 12072 23128 12124 23180
rect 12532 23128 12584 23180
rect 13176 23128 13228 23180
rect 13544 23128 13596 23180
rect 16488 23128 16540 23180
rect 11152 23103 11204 23112
rect 11152 23069 11161 23103
rect 11161 23069 11195 23103
rect 11195 23069 11204 23103
rect 11152 23060 11204 23069
rect 14188 23060 14240 23112
rect 15292 23103 15344 23112
rect 15292 23069 15301 23103
rect 15301 23069 15335 23103
rect 15335 23069 15344 23103
rect 15292 23060 15344 23069
rect 13728 22992 13780 23044
rect 14648 22992 14700 23044
rect 7840 22924 7892 22976
rect 13268 22924 13320 22976
rect 14004 22924 14056 22976
rect 14280 22924 14332 22976
rect 15476 22924 15528 22976
rect 16304 22924 16356 22976
rect 16764 22924 16816 22976
rect 5982 22822 6034 22874
rect 6046 22822 6098 22874
rect 6110 22822 6162 22874
rect 6174 22822 6226 22874
rect 15982 22822 16034 22874
rect 16046 22822 16098 22874
rect 16110 22822 16162 22874
rect 16174 22822 16226 22874
rect 25982 22822 26034 22874
rect 26046 22822 26098 22874
rect 26110 22822 26162 22874
rect 26174 22822 26226 22874
rect 7196 22720 7248 22772
rect 9956 22720 10008 22772
rect 11152 22720 11204 22772
rect 11704 22763 11756 22772
rect 11704 22729 11713 22763
rect 11713 22729 11747 22763
rect 11747 22729 11756 22763
rect 11704 22720 11756 22729
rect 6276 22695 6328 22704
rect 6276 22661 6285 22695
rect 6285 22661 6319 22695
rect 6319 22661 6328 22695
rect 6276 22652 6328 22661
rect 6644 22695 6696 22704
rect 6644 22661 6653 22695
rect 6653 22661 6687 22695
rect 6687 22661 6696 22695
rect 6644 22652 6696 22661
rect 11520 22652 11572 22704
rect 12624 22652 12676 22704
rect 6828 22627 6880 22636
rect 6828 22593 6837 22627
rect 6837 22593 6871 22627
rect 6871 22593 6880 22627
rect 6828 22584 6880 22593
rect 7104 22627 7156 22636
rect 7104 22593 7113 22627
rect 7113 22593 7147 22627
rect 7147 22593 7156 22627
rect 7104 22584 7156 22593
rect 7288 22584 7340 22636
rect 7840 22584 7892 22636
rect 12440 22627 12492 22636
rect 12440 22593 12449 22627
rect 12449 22593 12483 22627
rect 12483 22593 12492 22627
rect 12440 22584 12492 22593
rect 12900 22584 12952 22636
rect 8576 22516 8628 22568
rect 13820 22720 13872 22772
rect 14004 22720 14056 22772
rect 15108 22720 15160 22772
rect 19616 22720 19668 22772
rect 21272 22720 21324 22772
rect 13544 22652 13596 22704
rect 13452 22584 13504 22636
rect 13636 22584 13688 22636
rect 8944 22448 8996 22500
rect 9404 22448 9456 22500
rect 10968 22448 11020 22500
rect 11336 22448 11388 22500
rect 12992 22491 13044 22500
rect 12992 22457 13001 22491
rect 13001 22457 13035 22491
rect 13035 22457 13044 22491
rect 12992 22448 13044 22457
rect 7104 22380 7156 22432
rect 9496 22423 9548 22432
rect 9496 22389 9505 22423
rect 9505 22389 9539 22423
rect 9539 22389 9548 22423
rect 9496 22380 9548 22389
rect 10048 22380 10100 22432
rect 16304 22652 16356 22704
rect 16488 22652 16540 22704
rect 14832 22584 14884 22636
rect 18420 22584 18472 22636
rect 25872 22584 25924 22636
rect 14280 22559 14332 22568
rect 14280 22525 14289 22559
rect 14289 22525 14323 22559
rect 14323 22525 14332 22559
rect 14280 22516 14332 22525
rect 14648 22559 14700 22568
rect 14648 22525 14657 22559
rect 14657 22525 14691 22559
rect 14691 22525 14700 22559
rect 14648 22516 14700 22525
rect 15292 22516 15344 22568
rect 15660 22516 15712 22568
rect 18144 22516 18196 22568
rect 26148 22559 26200 22568
rect 26148 22525 26157 22559
rect 26157 22525 26191 22559
rect 26191 22525 26200 22559
rect 26148 22516 26200 22525
rect 14924 22448 14976 22500
rect 15476 22448 15528 22500
rect 16672 22448 16724 22500
rect 15384 22380 15436 22432
rect 15844 22380 15896 22432
rect 16396 22380 16448 22432
rect 16580 22380 16632 22432
rect 19340 22380 19392 22432
rect 27712 22423 27764 22432
rect 27712 22389 27721 22423
rect 27721 22389 27755 22423
rect 27755 22389 27764 22423
rect 27712 22380 27764 22389
rect 10982 22278 11034 22330
rect 11046 22278 11098 22330
rect 11110 22278 11162 22330
rect 11174 22278 11226 22330
rect 20982 22278 21034 22330
rect 21046 22278 21098 22330
rect 21110 22278 21162 22330
rect 21174 22278 21226 22330
rect 9496 22176 9548 22228
rect 12900 22176 12952 22228
rect 14280 22176 14332 22228
rect 14924 22176 14976 22228
rect 16580 22176 16632 22228
rect 14740 22108 14792 22160
rect 18420 22176 18472 22228
rect 18880 22176 18932 22228
rect 25780 22176 25832 22228
rect 26148 22219 26200 22228
rect 26148 22185 26157 22219
rect 26157 22185 26191 22219
rect 26191 22185 26200 22219
rect 26148 22176 26200 22185
rect 6828 22040 6880 22092
rect 8576 22083 8628 22092
rect 8576 22049 8585 22083
rect 8585 22049 8619 22083
rect 8619 22049 8628 22083
rect 8576 22040 8628 22049
rect 12072 22040 12124 22092
rect 12256 22040 12308 22092
rect 6276 21972 6328 22024
rect 6368 22015 6420 22024
rect 6368 21981 6377 22015
rect 6377 21981 6411 22015
rect 6411 21981 6420 22015
rect 6368 21972 6420 21981
rect 8300 21972 8352 22024
rect 9956 22015 10008 22024
rect 9956 21981 9965 22015
rect 9965 21981 9999 22015
rect 9999 21981 10008 22015
rect 9956 21972 10008 21981
rect 13176 22015 13228 22024
rect 13176 21981 13185 22015
rect 13185 21981 13219 22015
rect 13219 21981 13228 22015
rect 13176 21972 13228 21981
rect 16580 22040 16632 22092
rect 16764 22040 16816 22092
rect 18604 22040 18656 22092
rect 19340 22083 19392 22092
rect 19340 22049 19349 22083
rect 19349 22049 19383 22083
rect 19383 22049 19392 22083
rect 19340 22040 19392 22049
rect 15016 21972 15068 22024
rect 15108 21972 15160 22024
rect 16488 21972 16540 22024
rect 17040 21972 17092 22024
rect 17500 21972 17552 22024
rect 18420 22015 18472 22024
rect 18420 21981 18429 22015
rect 18429 21981 18463 22015
rect 18463 21981 18472 22015
rect 18420 21972 18472 21981
rect 19064 22015 19116 22024
rect 19064 21981 19073 22015
rect 19073 21981 19107 22015
rect 19107 21981 19116 22015
rect 19064 21972 19116 21981
rect 19248 22015 19300 22024
rect 19248 21981 19257 22015
rect 19257 21981 19291 22015
rect 19291 21981 19300 22015
rect 19248 21972 19300 21981
rect 13820 21904 13872 21956
rect 18880 21904 18932 21956
rect 7932 21836 7984 21888
rect 8760 21879 8812 21888
rect 8760 21845 8769 21879
rect 8769 21845 8803 21879
rect 8803 21845 8812 21879
rect 8760 21836 8812 21845
rect 11704 21836 11756 21888
rect 12256 21836 12308 21888
rect 12440 21836 12492 21888
rect 12716 21879 12768 21888
rect 12716 21845 12725 21879
rect 12725 21845 12759 21879
rect 12759 21845 12768 21879
rect 12716 21836 12768 21845
rect 13452 21879 13504 21888
rect 13452 21845 13461 21879
rect 13461 21845 13495 21879
rect 13495 21845 13504 21879
rect 13452 21836 13504 21845
rect 14188 21836 14240 21888
rect 16672 21879 16724 21888
rect 16672 21845 16681 21879
rect 16681 21845 16715 21879
rect 16715 21845 16724 21879
rect 16672 21836 16724 21845
rect 18144 21879 18196 21888
rect 18144 21845 18153 21879
rect 18153 21845 18187 21879
rect 18187 21845 18196 21879
rect 18144 21836 18196 21845
rect 5982 21734 6034 21786
rect 6046 21734 6098 21786
rect 6110 21734 6162 21786
rect 6174 21734 6226 21786
rect 15982 21734 16034 21786
rect 16046 21734 16098 21786
rect 16110 21734 16162 21786
rect 16174 21734 16226 21786
rect 25982 21734 26034 21786
rect 26046 21734 26098 21786
rect 26110 21734 26162 21786
rect 26174 21734 26226 21786
rect 8576 21675 8628 21684
rect 8576 21641 8585 21675
rect 8585 21641 8619 21675
rect 8619 21641 8628 21675
rect 8576 21632 8628 21641
rect 9956 21632 10008 21684
rect 10784 21675 10836 21684
rect 10784 21641 10793 21675
rect 10793 21641 10827 21675
rect 10827 21641 10836 21675
rect 10784 21632 10836 21641
rect 12072 21632 12124 21684
rect 12624 21632 12676 21684
rect 13820 21675 13872 21684
rect 13820 21641 13829 21675
rect 13829 21641 13863 21675
rect 13863 21641 13872 21675
rect 13820 21632 13872 21641
rect 16304 21632 16356 21684
rect 16396 21632 16448 21684
rect 16764 21632 16816 21684
rect 17684 21675 17736 21684
rect 17684 21641 17693 21675
rect 17693 21641 17727 21675
rect 17727 21641 17736 21675
rect 17684 21632 17736 21641
rect 19340 21675 19392 21684
rect 19340 21641 19349 21675
rect 19349 21641 19383 21675
rect 19383 21641 19392 21675
rect 19340 21632 19392 21641
rect 6368 21564 6420 21616
rect 8852 21496 8904 21548
rect 13176 21564 13228 21616
rect 7932 21471 7984 21480
rect 7932 21437 7941 21471
rect 7941 21437 7975 21471
rect 7975 21437 7984 21471
rect 7932 21428 7984 21437
rect 6644 21360 6696 21412
rect 6920 21403 6972 21412
rect 6920 21369 6929 21403
rect 6929 21369 6963 21403
rect 6963 21369 6972 21403
rect 6920 21360 6972 21369
rect 7288 21292 7340 21344
rect 8760 21428 8812 21480
rect 8944 21471 8996 21480
rect 8944 21437 8953 21471
rect 8953 21437 8987 21471
rect 8987 21437 8996 21471
rect 8944 21428 8996 21437
rect 9496 21428 9548 21480
rect 10600 21428 10652 21480
rect 12440 21428 12492 21480
rect 13820 21496 13872 21548
rect 14004 21496 14056 21548
rect 17776 21564 17828 21616
rect 17408 21496 17460 21548
rect 17684 21496 17736 21548
rect 18788 21564 18840 21616
rect 18052 21539 18104 21548
rect 18052 21505 18061 21539
rect 18061 21505 18095 21539
rect 18095 21505 18104 21539
rect 18052 21496 18104 21505
rect 11520 21403 11572 21412
rect 11520 21369 11529 21403
rect 11529 21369 11563 21403
rect 11563 21369 11572 21403
rect 11520 21360 11572 21369
rect 12716 21428 12768 21480
rect 13176 21428 13228 21480
rect 13452 21471 13504 21480
rect 13452 21437 13461 21471
rect 13461 21437 13495 21471
rect 13495 21437 13504 21471
rect 13452 21428 13504 21437
rect 16488 21471 16540 21480
rect 14280 21360 14332 21412
rect 16488 21437 16497 21471
rect 16497 21437 16531 21471
rect 16531 21437 16540 21471
rect 16488 21428 16540 21437
rect 16672 21471 16724 21480
rect 16672 21437 16681 21471
rect 16681 21437 16715 21471
rect 16715 21437 16724 21471
rect 16672 21428 16724 21437
rect 18144 21428 18196 21480
rect 15660 21360 15712 21412
rect 16764 21360 16816 21412
rect 25044 21360 25096 21412
rect 25320 21360 25372 21412
rect 10324 21292 10376 21344
rect 10600 21292 10652 21344
rect 12256 21292 12308 21344
rect 15016 21292 15068 21344
rect 15936 21292 15988 21344
rect 16212 21292 16264 21344
rect 16488 21292 16540 21344
rect 10982 21190 11034 21242
rect 11046 21190 11098 21242
rect 11110 21190 11162 21242
rect 11174 21190 11226 21242
rect 20982 21190 21034 21242
rect 21046 21190 21098 21242
rect 21110 21190 21162 21242
rect 21174 21190 21226 21242
rect 6276 21088 6328 21140
rect 6644 21088 6696 21140
rect 7932 21088 7984 21140
rect 8944 21131 8996 21140
rect 8944 21097 8953 21131
rect 8953 21097 8987 21131
rect 8987 21097 8996 21131
rect 8944 21088 8996 21097
rect 9496 21131 9548 21140
rect 9496 21097 9505 21131
rect 9505 21097 9539 21131
rect 9539 21097 9548 21131
rect 9496 21088 9548 21097
rect 9864 21131 9916 21140
rect 9864 21097 9873 21131
rect 9873 21097 9907 21131
rect 9907 21097 9916 21131
rect 9864 21088 9916 21097
rect 11428 21088 11480 21140
rect 13084 21131 13136 21140
rect 13084 21097 13093 21131
rect 13093 21097 13127 21131
rect 13127 21097 13136 21131
rect 13084 21088 13136 21097
rect 14280 21088 14332 21140
rect 14740 21088 14792 21140
rect 16488 21088 16540 21140
rect 16672 21088 16724 21140
rect 19248 21088 19300 21140
rect 3148 21063 3200 21072
rect 3148 21029 3157 21063
rect 3157 21029 3191 21063
rect 3191 21029 3200 21063
rect 3148 21020 3200 21029
rect 12072 21020 12124 21072
rect 13452 21020 13504 21072
rect 13820 21020 13872 21072
rect 14648 21020 14700 21072
rect 18604 21020 18656 21072
rect 1584 20952 1636 21004
rect 9864 20952 9916 21004
rect 10048 20952 10100 21004
rect 11060 20995 11112 21004
rect 11060 20961 11069 20995
rect 11069 20961 11103 20995
rect 11103 20961 11112 20995
rect 11060 20952 11112 20961
rect 2136 20884 2188 20936
rect 10876 20884 10928 20936
rect 11520 20952 11572 21004
rect 12992 20995 13044 21004
rect 12992 20961 13001 20995
rect 13001 20961 13035 20995
rect 13035 20961 13044 20995
rect 12992 20952 13044 20961
rect 14188 20995 14240 21004
rect 14188 20961 14197 20995
rect 14197 20961 14231 20995
rect 14231 20961 14240 20995
rect 14188 20952 14240 20961
rect 15476 20952 15528 21004
rect 15568 20952 15620 21004
rect 15936 20952 15988 21004
rect 18972 20952 19024 21004
rect 22468 20952 22520 21004
rect 22928 20952 22980 21004
rect 11704 20884 11756 20936
rect 11980 20884 12032 20936
rect 16304 20884 16356 20936
rect 16672 20927 16724 20936
rect 16672 20893 16681 20927
rect 16681 20893 16715 20927
rect 16715 20893 16724 20927
rect 16672 20884 16724 20893
rect 10968 20816 11020 20868
rect 10048 20748 10100 20800
rect 10600 20748 10652 20800
rect 12256 20816 12308 20868
rect 11336 20791 11388 20800
rect 11336 20757 11345 20791
rect 11345 20757 11379 20791
rect 11379 20757 11388 20791
rect 11336 20748 11388 20757
rect 11980 20748 12032 20800
rect 13636 20791 13688 20800
rect 13636 20757 13645 20791
rect 13645 20757 13679 20791
rect 13679 20757 13688 20791
rect 13636 20748 13688 20757
rect 15016 20791 15068 20800
rect 15016 20757 15025 20791
rect 15025 20757 15059 20791
rect 15059 20757 15068 20791
rect 15016 20748 15068 20757
rect 15660 20748 15712 20800
rect 16672 20748 16724 20800
rect 19064 20748 19116 20800
rect 19248 20748 19300 20800
rect 23756 20791 23808 20800
rect 23756 20757 23765 20791
rect 23765 20757 23799 20791
rect 23799 20757 23808 20791
rect 23756 20748 23808 20757
rect 5982 20646 6034 20698
rect 6046 20646 6098 20698
rect 6110 20646 6162 20698
rect 6174 20646 6226 20698
rect 15982 20646 16034 20698
rect 16046 20646 16098 20698
rect 16110 20646 16162 20698
rect 16174 20646 16226 20698
rect 25982 20646 26034 20698
rect 26046 20646 26098 20698
rect 26110 20646 26162 20698
rect 26174 20646 26226 20698
rect 2136 20544 2188 20596
rect 9496 20544 9548 20596
rect 10140 20587 10192 20596
rect 10140 20553 10149 20587
rect 10149 20553 10183 20587
rect 10183 20553 10192 20587
rect 10140 20544 10192 20553
rect 10232 20544 10284 20596
rect 10876 20544 10928 20596
rect 12992 20544 13044 20596
rect 15476 20587 15528 20596
rect 15476 20553 15485 20587
rect 15485 20553 15519 20587
rect 15519 20553 15528 20587
rect 15476 20544 15528 20553
rect 12624 20476 12676 20528
rect 10692 20408 10744 20460
rect 10968 20340 11020 20392
rect 11336 20383 11388 20392
rect 11336 20349 11345 20383
rect 11345 20349 11379 20383
rect 11379 20349 11388 20383
rect 11336 20340 11388 20349
rect 10324 20315 10376 20324
rect 10324 20281 10333 20315
rect 10333 20281 10367 20315
rect 10367 20281 10376 20315
rect 10324 20272 10376 20281
rect 13728 20476 13780 20528
rect 12992 20408 13044 20460
rect 13452 20340 13504 20392
rect 13636 20383 13688 20392
rect 13636 20349 13645 20383
rect 13645 20349 13679 20383
rect 13679 20349 13688 20383
rect 13636 20340 13688 20349
rect 16212 20408 16264 20460
rect 16672 20544 16724 20596
rect 17408 20544 17460 20596
rect 17684 20544 17736 20596
rect 16488 20476 16540 20528
rect 22928 20544 22980 20596
rect 18512 20476 18564 20528
rect 14188 20383 14240 20392
rect 14188 20349 14197 20383
rect 14197 20349 14231 20383
rect 14231 20349 14240 20383
rect 14188 20340 14240 20349
rect 16580 20340 16632 20392
rect 16856 20383 16908 20392
rect 16856 20349 16865 20383
rect 16865 20349 16899 20383
rect 16899 20349 16908 20383
rect 16856 20340 16908 20349
rect 18236 20340 18288 20392
rect 18696 20383 18748 20392
rect 18696 20349 18705 20383
rect 18705 20349 18739 20383
rect 18739 20349 18748 20383
rect 18696 20340 18748 20349
rect 14832 20272 14884 20324
rect 1584 20247 1636 20256
rect 1584 20213 1593 20247
rect 1593 20213 1627 20247
rect 1627 20213 1636 20247
rect 1584 20204 1636 20213
rect 9864 20204 9916 20256
rect 14648 20204 14700 20256
rect 16764 20204 16816 20256
rect 22376 20247 22428 20256
rect 22376 20213 22385 20247
rect 22385 20213 22419 20247
rect 22419 20213 22428 20247
rect 22376 20204 22428 20213
rect 10982 20102 11034 20154
rect 11046 20102 11098 20154
rect 11110 20102 11162 20154
rect 11174 20102 11226 20154
rect 20982 20102 21034 20154
rect 21046 20102 21098 20154
rect 21110 20102 21162 20154
rect 21174 20102 21226 20154
rect 7472 20043 7524 20052
rect 7472 20009 7481 20043
rect 7481 20009 7515 20043
rect 7515 20009 7524 20043
rect 7472 20000 7524 20009
rect 10324 20000 10376 20052
rect 11336 20000 11388 20052
rect 10876 19932 10928 19984
rect 8208 19907 8260 19916
rect 8208 19873 8217 19907
rect 8217 19873 8251 19907
rect 8251 19873 8260 19907
rect 8208 19864 8260 19873
rect 8944 19864 8996 19916
rect 11520 19864 11572 19916
rect 12164 19864 12216 19916
rect 12440 19864 12492 19916
rect 14280 20000 14332 20052
rect 14740 20000 14792 20052
rect 13176 19975 13228 19984
rect 13176 19941 13185 19975
rect 13185 19941 13219 19975
rect 13219 19941 13228 19975
rect 13176 19932 13228 19941
rect 12992 19864 13044 19916
rect 14004 19907 14056 19916
rect 14004 19873 14013 19907
rect 14013 19873 14047 19907
rect 14047 19873 14056 19907
rect 16488 20000 16540 20052
rect 16580 19932 16632 19984
rect 18972 19932 19024 19984
rect 19524 19975 19576 19984
rect 14004 19864 14056 19873
rect 15752 19864 15804 19916
rect 16304 19864 16356 19916
rect 17408 19864 17460 19916
rect 19524 19941 19533 19975
rect 19533 19941 19567 19975
rect 19567 19941 19576 19975
rect 19524 19932 19576 19941
rect 11428 19796 11480 19848
rect 12624 19839 12676 19848
rect 12624 19805 12633 19839
rect 12633 19805 12667 19839
rect 12667 19805 12676 19839
rect 12624 19796 12676 19805
rect 16488 19839 16540 19848
rect 16488 19805 16497 19839
rect 16497 19805 16531 19839
rect 16531 19805 16540 19839
rect 16488 19796 16540 19805
rect 16764 19839 16816 19848
rect 16764 19805 16773 19839
rect 16773 19805 16807 19839
rect 16807 19805 16816 19839
rect 16764 19796 16816 19805
rect 18696 19796 18748 19848
rect 19248 19796 19300 19848
rect 11244 19728 11296 19780
rect 11612 19728 11664 19780
rect 12900 19728 12952 19780
rect 13176 19728 13228 19780
rect 8116 19660 8168 19712
rect 13452 19660 13504 19712
rect 14372 19660 14424 19712
rect 14740 19660 14792 19712
rect 16856 19660 16908 19712
rect 18144 19660 18196 19712
rect 5982 19558 6034 19610
rect 6046 19558 6098 19610
rect 6110 19558 6162 19610
rect 6174 19558 6226 19610
rect 15982 19558 16034 19610
rect 16046 19558 16098 19610
rect 16110 19558 16162 19610
rect 16174 19558 16226 19610
rect 25982 19558 26034 19610
rect 26046 19558 26098 19610
rect 26110 19558 26162 19610
rect 26174 19558 26226 19610
rect 8944 19499 8996 19508
rect 8944 19465 8953 19499
rect 8953 19465 8987 19499
rect 8987 19465 8996 19499
rect 8944 19456 8996 19465
rect 11520 19456 11572 19508
rect 12164 19456 12216 19508
rect 14004 19499 14056 19508
rect 14004 19465 14013 19499
rect 14013 19465 14047 19499
rect 14047 19465 14056 19499
rect 14004 19456 14056 19465
rect 15752 19456 15804 19508
rect 16856 19499 16908 19508
rect 16856 19465 16865 19499
rect 16865 19465 16899 19499
rect 16899 19465 16908 19499
rect 16856 19456 16908 19465
rect 17132 19456 17184 19508
rect 18236 19456 18288 19508
rect 18972 19499 19024 19508
rect 18972 19465 18981 19499
rect 18981 19465 19015 19499
rect 19015 19465 19024 19499
rect 18972 19456 19024 19465
rect 7472 19320 7524 19372
rect 7288 19295 7340 19304
rect 7288 19261 7297 19295
rect 7297 19261 7331 19295
rect 7331 19261 7340 19295
rect 7288 19252 7340 19261
rect 8116 19363 8168 19372
rect 8116 19329 8125 19363
rect 8125 19329 8159 19363
rect 8159 19329 8168 19363
rect 8116 19320 8168 19329
rect 9496 19320 9548 19372
rect 10324 19320 10376 19372
rect 12440 19363 12492 19372
rect 12440 19329 12449 19363
rect 12449 19329 12483 19363
rect 12483 19329 12492 19363
rect 12440 19320 12492 19329
rect 16488 19320 16540 19372
rect 16856 19320 16908 19372
rect 19248 19320 19300 19372
rect 8208 19252 8260 19304
rect 8392 19295 8444 19304
rect 8392 19261 8401 19295
rect 8401 19261 8435 19295
rect 8435 19261 8444 19295
rect 8392 19252 8444 19261
rect 6644 19159 6696 19168
rect 6644 19125 6653 19159
rect 6653 19125 6687 19159
rect 6687 19125 6696 19159
rect 6644 19116 6696 19125
rect 8024 19116 8076 19168
rect 8484 19116 8536 19168
rect 8944 19252 8996 19304
rect 9312 19295 9364 19304
rect 9312 19261 9321 19295
rect 9321 19261 9355 19295
rect 9355 19261 9364 19295
rect 9312 19252 9364 19261
rect 10232 19252 10284 19304
rect 9496 19184 9548 19236
rect 9772 19159 9824 19168
rect 9772 19125 9781 19159
rect 9781 19125 9815 19159
rect 9815 19125 9824 19159
rect 9772 19116 9824 19125
rect 9956 19184 10008 19236
rect 10048 19116 10100 19168
rect 12164 19252 12216 19304
rect 12900 19295 12952 19304
rect 11152 19184 11204 19236
rect 12256 19227 12308 19236
rect 12256 19193 12265 19227
rect 12265 19193 12299 19227
rect 12299 19193 12308 19227
rect 12256 19184 12308 19193
rect 12900 19261 12909 19295
rect 12909 19261 12943 19295
rect 12943 19261 12952 19295
rect 12900 19252 12952 19261
rect 13084 19295 13136 19304
rect 13084 19261 13093 19295
rect 13093 19261 13127 19295
rect 13127 19261 13136 19295
rect 13084 19252 13136 19261
rect 14372 19252 14424 19304
rect 15108 19252 15160 19304
rect 16212 19252 16264 19304
rect 17408 19252 17460 19304
rect 18144 19295 18196 19304
rect 18144 19261 18153 19295
rect 18153 19261 18187 19295
rect 18187 19261 18196 19295
rect 18144 19252 18196 19261
rect 19432 19252 19484 19304
rect 12164 19116 12216 19168
rect 12624 19116 12676 19168
rect 12900 19116 12952 19168
rect 14648 19159 14700 19168
rect 14648 19125 14657 19159
rect 14657 19125 14691 19159
rect 14691 19125 14700 19159
rect 14648 19116 14700 19125
rect 15568 19116 15620 19168
rect 16764 19116 16816 19168
rect 17776 19159 17828 19168
rect 17776 19125 17785 19159
rect 17785 19125 17819 19159
rect 17819 19125 17828 19159
rect 17776 19116 17828 19125
rect 10982 19014 11034 19066
rect 11046 19014 11098 19066
rect 11110 19014 11162 19066
rect 11174 19014 11226 19066
rect 20982 19014 21034 19066
rect 21046 19014 21098 19066
rect 21110 19014 21162 19066
rect 21174 19014 21226 19066
rect 6644 18912 6696 18964
rect 8392 18912 8444 18964
rect 9956 18955 10008 18964
rect 9956 18921 9965 18955
rect 9965 18921 9999 18955
rect 9999 18921 10008 18955
rect 9956 18912 10008 18921
rect 10784 18955 10836 18964
rect 10784 18921 10793 18955
rect 10793 18921 10827 18955
rect 10827 18921 10836 18955
rect 10784 18912 10836 18921
rect 12716 18912 12768 18964
rect 13084 18912 13136 18964
rect 14188 18912 14240 18964
rect 15016 18912 15068 18964
rect 15752 18955 15804 18964
rect 15752 18921 15761 18955
rect 15761 18921 15795 18955
rect 15795 18921 15804 18955
rect 15752 18912 15804 18921
rect 16212 18912 16264 18964
rect 18144 18955 18196 18964
rect 18144 18921 18153 18955
rect 18153 18921 18187 18955
rect 18187 18921 18196 18955
rect 18144 18912 18196 18921
rect 13452 18844 13504 18896
rect 7196 18776 7248 18828
rect 8116 18776 8168 18828
rect 10876 18776 10928 18828
rect 11704 18819 11756 18828
rect 11704 18785 11713 18819
rect 11713 18785 11747 18819
rect 11747 18785 11756 18819
rect 11704 18776 11756 18785
rect 12440 18776 12492 18828
rect 16304 18776 16356 18828
rect 16580 18776 16632 18828
rect 17684 18776 17736 18828
rect 7104 18751 7156 18760
rect 7104 18717 7113 18751
rect 7113 18717 7147 18751
rect 7147 18717 7156 18751
rect 7104 18708 7156 18717
rect 11428 18751 11480 18760
rect 11428 18717 11437 18751
rect 11437 18717 11471 18751
rect 11471 18717 11480 18751
rect 11428 18708 11480 18717
rect 12716 18751 12768 18760
rect 10508 18640 10560 18692
rect 12716 18717 12725 18751
rect 12725 18717 12759 18751
rect 12759 18717 12768 18751
rect 12716 18708 12768 18717
rect 13176 18708 13228 18760
rect 13728 18751 13780 18760
rect 13728 18717 13737 18751
rect 13737 18717 13771 18751
rect 13771 18717 13780 18751
rect 13728 18708 13780 18717
rect 3332 18572 3384 18624
rect 9496 18572 9548 18624
rect 10232 18615 10284 18624
rect 10232 18581 10241 18615
rect 10241 18581 10275 18615
rect 10275 18581 10284 18615
rect 10232 18572 10284 18581
rect 12440 18640 12492 18692
rect 15108 18640 15160 18692
rect 16488 18572 16540 18624
rect 16580 18572 16632 18624
rect 17132 18615 17184 18624
rect 17132 18581 17141 18615
rect 17141 18581 17175 18615
rect 17175 18581 17184 18615
rect 17132 18572 17184 18581
rect 17408 18572 17460 18624
rect 5982 18470 6034 18522
rect 6046 18470 6098 18522
rect 6110 18470 6162 18522
rect 6174 18470 6226 18522
rect 15982 18470 16034 18522
rect 16046 18470 16098 18522
rect 16110 18470 16162 18522
rect 16174 18470 16226 18522
rect 25982 18470 26034 18522
rect 26046 18470 26098 18522
rect 26110 18470 26162 18522
rect 26174 18470 26226 18522
rect 3332 18368 3384 18420
rect 7104 18368 7156 18420
rect 7840 18368 7892 18420
rect 8300 18368 8352 18420
rect 8668 18368 8720 18420
rect 7196 18343 7248 18352
rect 7196 18309 7205 18343
rect 7205 18309 7239 18343
rect 7239 18309 7248 18343
rect 7196 18300 7248 18309
rect 9956 18368 10008 18420
rect 11704 18368 11756 18420
rect 11980 18368 12032 18420
rect 13728 18368 13780 18420
rect 14372 18411 14424 18420
rect 14372 18377 14381 18411
rect 14381 18377 14415 18411
rect 14415 18377 14424 18411
rect 14372 18368 14424 18377
rect 16304 18411 16356 18420
rect 16304 18377 16313 18411
rect 16313 18377 16347 18411
rect 16347 18377 16356 18411
rect 16304 18368 16356 18377
rect 17316 18411 17368 18420
rect 17316 18377 17325 18411
rect 17325 18377 17359 18411
rect 17359 18377 17368 18411
rect 17316 18368 17368 18377
rect 17684 18411 17736 18420
rect 17684 18377 17693 18411
rect 17693 18377 17727 18411
rect 17727 18377 17736 18411
rect 17684 18368 17736 18377
rect 10692 18300 10744 18352
rect 13176 18300 13228 18352
rect 9312 18232 9364 18284
rect 9680 18232 9732 18284
rect 10232 18232 10284 18284
rect 10324 18275 10376 18284
rect 10324 18241 10333 18275
rect 10333 18241 10367 18275
rect 10367 18241 10376 18275
rect 10324 18232 10376 18241
rect 1860 18207 1912 18216
rect 1860 18173 1869 18207
rect 1869 18173 1903 18207
rect 1903 18173 1912 18207
rect 1860 18164 1912 18173
rect 1492 18028 1544 18080
rect 9588 18164 9640 18216
rect 11428 18164 11480 18216
rect 13452 18207 13504 18216
rect 11244 18096 11296 18148
rect 13452 18173 13461 18207
rect 13461 18173 13495 18207
rect 13495 18173 13504 18207
rect 13452 18164 13504 18173
rect 14648 18164 14700 18216
rect 15752 18300 15804 18352
rect 16488 18300 16540 18352
rect 15016 18275 15068 18284
rect 15016 18241 15025 18275
rect 15025 18241 15059 18275
rect 15059 18241 15068 18275
rect 15016 18232 15068 18241
rect 15108 18164 15160 18216
rect 16580 18232 16632 18284
rect 13544 18096 13596 18148
rect 11704 18028 11756 18080
rect 11980 18028 12032 18080
rect 14740 18028 14792 18080
rect 15568 18164 15620 18216
rect 17316 18164 17368 18216
rect 10982 17926 11034 17978
rect 11046 17926 11098 17978
rect 11110 17926 11162 17978
rect 11174 17926 11226 17978
rect 20982 17926 21034 17978
rect 21046 17926 21098 17978
rect 21110 17926 21162 17978
rect 21174 17926 21226 17978
rect 8300 17867 8352 17876
rect 8300 17833 8309 17867
rect 8309 17833 8343 17867
rect 8343 17833 8352 17867
rect 8300 17824 8352 17833
rect 9312 17824 9364 17876
rect 11428 17824 11480 17876
rect 12348 17824 12400 17876
rect 13544 17867 13596 17876
rect 13544 17833 13553 17867
rect 13553 17833 13587 17867
rect 13587 17833 13596 17867
rect 13544 17824 13596 17833
rect 14648 17867 14700 17876
rect 14648 17833 14657 17867
rect 14657 17833 14691 17867
rect 14691 17833 14700 17867
rect 14648 17824 14700 17833
rect 15568 17867 15620 17876
rect 15568 17833 15577 17867
rect 15577 17833 15611 17867
rect 15611 17833 15620 17867
rect 15568 17824 15620 17833
rect 16304 17824 16356 17876
rect 16488 17824 16540 17876
rect 17960 17824 18012 17876
rect 9680 17756 9732 17808
rect 10876 17756 10928 17808
rect 13728 17756 13780 17808
rect 11152 17731 11204 17740
rect 11152 17697 11161 17731
rect 11161 17697 11195 17731
rect 11195 17697 11204 17731
rect 11152 17688 11204 17697
rect 12532 17731 12584 17740
rect 12532 17697 12541 17731
rect 12541 17697 12575 17731
rect 12575 17697 12584 17731
rect 12532 17688 12584 17697
rect 12992 17688 13044 17740
rect 13268 17731 13320 17740
rect 13268 17697 13277 17731
rect 13277 17697 13311 17731
rect 13311 17697 13320 17731
rect 13268 17688 13320 17697
rect 5172 17620 5224 17672
rect 9588 17620 9640 17672
rect 10324 17620 10376 17672
rect 11336 17663 11388 17672
rect 11336 17629 11345 17663
rect 11345 17629 11379 17663
rect 11379 17629 11388 17663
rect 11336 17620 11388 17629
rect 12164 17620 12216 17672
rect 12624 17620 12676 17672
rect 15016 17620 15068 17672
rect 15752 17663 15804 17672
rect 15752 17629 15761 17663
rect 15761 17629 15795 17663
rect 15795 17629 15804 17663
rect 15752 17620 15804 17629
rect 16488 17688 16540 17740
rect 17408 17688 17460 17740
rect 10784 17552 10836 17604
rect 1952 17527 2004 17536
rect 1952 17493 1961 17527
rect 1961 17493 1995 17527
rect 1995 17493 2004 17527
rect 1952 17484 2004 17493
rect 17316 17484 17368 17536
rect 5982 17382 6034 17434
rect 6046 17382 6098 17434
rect 6110 17382 6162 17434
rect 6174 17382 6226 17434
rect 15982 17382 16034 17434
rect 16046 17382 16098 17434
rect 16110 17382 16162 17434
rect 16174 17382 16226 17434
rect 25982 17382 26034 17434
rect 26046 17382 26098 17434
rect 26110 17382 26162 17434
rect 26174 17382 26226 17434
rect 2780 17323 2832 17332
rect 2780 17289 2789 17323
rect 2789 17289 2823 17323
rect 2823 17289 2832 17323
rect 2780 17280 2832 17289
rect 9404 17280 9456 17332
rect 9956 17280 10008 17332
rect 10692 17280 10744 17332
rect 8576 17212 8628 17264
rect 1676 17187 1728 17196
rect 1676 17153 1685 17187
rect 1685 17153 1719 17187
rect 1719 17153 1728 17187
rect 1676 17144 1728 17153
rect 8300 17144 8352 17196
rect 1952 17076 2004 17128
rect 8944 17187 8996 17196
rect 8944 17153 8953 17187
rect 8953 17153 8987 17187
rect 8987 17153 8996 17187
rect 9680 17212 9732 17264
rect 10232 17212 10284 17264
rect 11152 17212 11204 17264
rect 8944 17144 8996 17153
rect 10784 17187 10836 17196
rect 10784 17153 10793 17187
rect 10793 17153 10827 17187
rect 10827 17153 10836 17187
rect 10784 17144 10836 17153
rect 11244 17187 11296 17196
rect 11244 17153 11253 17187
rect 11253 17153 11287 17187
rect 11287 17153 11296 17187
rect 11244 17144 11296 17153
rect 10140 17076 10192 17128
rect 10600 17076 10652 17128
rect 10876 17076 10928 17128
rect 12164 17280 12216 17332
rect 12992 17280 13044 17332
rect 13820 17280 13872 17332
rect 14464 17280 14516 17332
rect 15384 17280 15436 17332
rect 15568 17280 15620 17332
rect 16304 17280 16356 17332
rect 16488 17212 16540 17264
rect 14188 17187 14240 17196
rect 14188 17153 14197 17187
rect 14197 17153 14231 17187
rect 14231 17153 14240 17187
rect 14188 17144 14240 17153
rect 16580 17144 16632 17196
rect 16948 17144 17000 17196
rect 12716 17119 12768 17128
rect 12716 17085 12725 17119
rect 12725 17085 12759 17119
rect 12759 17085 12768 17119
rect 12716 17076 12768 17085
rect 14280 17119 14332 17128
rect 14280 17085 14289 17119
rect 14289 17085 14323 17119
rect 14323 17085 14332 17119
rect 14280 17076 14332 17085
rect 14464 17076 14516 17128
rect 15016 17119 15068 17128
rect 15016 17085 15025 17119
rect 15025 17085 15059 17119
rect 15059 17085 15068 17119
rect 15016 17076 15068 17085
rect 15752 17076 15804 17128
rect 17408 17119 17460 17128
rect 9680 17008 9732 17060
rect 17408 17085 17417 17119
rect 17417 17085 17451 17119
rect 17451 17085 17460 17119
rect 17408 17076 17460 17085
rect 8944 16940 8996 16992
rect 9772 16940 9824 16992
rect 10600 16983 10652 16992
rect 10600 16949 10609 16983
rect 10609 16949 10643 16983
rect 10643 16949 10652 16983
rect 10600 16940 10652 16949
rect 14280 16940 14332 16992
rect 16672 17008 16724 17060
rect 17316 16940 17368 16992
rect 18052 16940 18104 16992
rect 10982 16838 11034 16890
rect 11046 16838 11098 16890
rect 11110 16838 11162 16890
rect 11174 16838 11226 16890
rect 20982 16838 21034 16890
rect 21046 16838 21098 16890
rect 21110 16838 21162 16890
rect 21174 16838 21226 16890
rect 1676 16779 1728 16788
rect 1676 16745 1685 16779
rect 1685 16745 1719 16779
rect 1719 16745 1728 16779
rect 1676 16736 1728 16745
rect 8484 16736 8536 16788
rect 9496 16779 9548 16788
rect 9496 16745 9505 16779
rect 9505 16745 9539 16779
rect 9539 16745 9548 16779
rect 9496 16736 9548 16745
rect 10324 16779 10376 16788
rect 10324 16745 10333 16779
rect 10333 16745 10367 16779
rect 10367 16745 10376 16779
rect 10324 16736 10376 16745
rect 10784 16736 10836 16788
rect 9312 16668 9364 16720
rect 10876 16668 10928 16720
rect 5816 16600 5868 16652
rect 13268 16736 13320 16788
rect 15568 16779 15620 16788
rect 15568 16745 15577 16779
rect 15577 16745 15611 16779
rect 15611 16745 15620 16779
rect 15568 16736 15620 16745
rect 16672 16779 16724 16788
rect 16672 16745 16681 16779
rect 16681 16745 16715 16779
rect 16715 16745 16724 16779
rect 16672 16736 16724 16745
rect 23664 16779 23716 16788
rect 23664 16745 23673 16779
rect 23673 16745 23707 16779
rect 23707 16745 23716 16779
rect 23664 16736 23716 16745
rect 11704 16668 11756 16720
rect 12072 16711 12124 16720
rect 12072 16677 12081 16711
rect 12081 16677 12115 16711
rect 12115 16677 12124 16711
rect 12072 16668 12124 16677
rect 12716 16668 12768 16720
rect 15016 16711 15068 16720
rect 15016 16677 15025 16711
rect 15025 16677 15059 16711
rect 15059 16677 15068 16711
rect 15016 16668 15068 16677
rect 15108 16668 15160 16720
rect 12532 16600 12584 16652
rect 13820 16643 13872 16652
rect 13820 16609 13829 16643
rect 13829 16609 13863 16643
rect 13863 16609 13872 16643
rect 13820 16600 13872 16609
rect 14096 16643 14148 16652
rect 14096 16609 14105 16643
rect 14105 16609 14139 16643
rect 14139 16609 14148 16643
rect 14096 16600 14148 16609
rect 15476 16643 15528 16652
rect 15476 16609 15485 16643
rect 15485 16609 15519 16643
rect 15519 16609 15528 16643
rect 15476 16600 15528 16609
rect 15844 16643 15896 16652
rect 15844 16609 15853 16643
rect 15853 16609 15887 16643
rect 15887 16609 15896 16643
rect 15844 16600 15896 16609
rect 16580 16600 16632 16652
rect 16764 16600 16816 16652
rect 17316 16600 17368 16652
rect 6552 16532 6604 16584
rect 11336 16532 11388 16584
rect 11980 16532 12032 16584
rect 13452 16575 13504 16584
rect 13452 16541 13461 16575
rect 13461 16541 13495 16575
rect 13495 16541 13504 16575
rect 13452 16532 13504 16541
rect 14648 16532 14700 16584
rect 22468 16532 22520 16584
rect 22744 16532 22796 16584
rect 1952 16396 2004 16448
rect 3424 16396 3476 16448
rect 17408 16439 17460 16448
rect 17408 16405 17417 16439
rect 17417 16405 17451 16439
rect 17451 16405 17460 16439
rect 17408 16396 17460 16405
rect 5982 16294 6034 16346
rect 6046 16294 6098 16346
rect 6110 16294 6162 16346
rect 6174 16294 6226 16346
rect 15982 16294 16034 16346
rect 16046 16294 16098 16346
rect 16110 16294 16162 16346
rect 16174 16294 16226 16346
rect 25982 16294 26034 16346
rect 26046 16294 26098 16346
rect 26110 16294 26162 16346
rect 26174 16294 26226 16346
rect 5172 16192 5224 16244
rect 6644 16192 6696 16244
rect 7840 16235 7892 16244
rect 7840 16201 7849 16235
rect 7849 16201 7883 16235
rect 7883 16201 7892 16235
rect 7840 16192 7892 16201
rect 9680 16235 9732 16244
rect 9680 16201 9689 16235
rect 9689 16201 9723 16235
rect 9723 16201 9732 16235
rect 9680 16192 9732 16201
rect 10692 16192 10744 16244
rect 13820 16192 13872 16244
rect 15844 16192 15896 16244
rect 16580 16192 16632 16244
rect 17316 16235 17368 16244
rect 17316 16201 17325 16235
rect 17325 16201 17359 16235
rect 17359 16201 17368 16235
rect 17316 16192 17368 16201
rect 19708 16192 19760 16244
rect 10784 16124 10836 16176
rect 15292 16124 15344 16176
rect 3424 16031 3476 16040
rect 3424 15997 3433 16031
rect 3433 15997 3467 16031
rect 3467 15997 3476 16031
rect 3424 15988 3476 15997
rect 3700 16031 3752 16040
rect 3700 15997 3709 16031
rect 3709 15997 3743 16031
rect 3743 15997 3752 16031
rect 3700 15988 3752 15997
rect 7840 15988 7892 16040
rect 9588 15988 9640 16040
rect 10140 15988 10192 16040
rect 10784 16031 10836 16040
rect 10784 15997 10793 16031
rect 10793 15997 10827 16031
rect 10827 15997 10836 16031
rect 10784 15988 10836 15997
rect 13084 15988 13136 16040
rect 11980 15920 12032 15972
rect 13452 15920 13504 15972
rect 13820 15920 13872 15972
rect 14740 15988 14792 16040
rect 15568 16031 15620 16040
rect 15568 15997 15577 16031
rect 15577 15997 15611 16031
rect 15611 15997 15620 16031
rect 15568 15988 15620 15997
rect 15844 16031 15896 16040
rect 15844 15997 15853 16031
rect 15853 15997 15887 16031
rect 15887 15997 15896 16031
rect 15844 15988 15896 15997
rect 18052 16031 18104 16040
rect 18052 15997 18061 16031
rect 18061 15997 18095 16031
rect 18095 15997 18104 16031
rect 18052 15988 18104 15997
rect 5816 15852 5868 15904
rect 11336 15895 11388 15904
rect 11336 15861 11345 15895
rect 11345 15861 11379 15895
rect 11379 15861 11388 15895
rect 11336 15852 11388 15861
rect 17684 15852 17736 15904
rect 22468 15852 22520 15904
rect 22744 15895 22796 15904
rect 22744 15861 22753 15895
rect 22753 15861 22787 15895
rect 22787 15861 22796 15895
rect 22744 15852 22796 15861
rect 10982 15750 11034 15802
rect 11046 15750 11098 15802
rect 11110 15750 11162 15802
rect 11174 15750 11226 15802
rect 20982 15750 21034 15802
rect 21046 15750 21098 15802
rect 21110 15750 21162 15802
rect 21174 15750 21226 15802
rect 3424 15648 3476 15700
rect 6644 15691 6696 15700
rect 6644 15657 6653 15691
rect 6653 15657 6687 15691
rect 6687 15657 6696 15691
rect 6644 15648 6696 15657
rect 10048 15691 10100 15700
rect 10048 15657 10057 15691
rect 10057 15657 10091 15691
rect 10091 15657 10100 15691
rect 10048 15648 10100 15657
rect 10876 15648 10928 15700
rect 7012 15580 7064 15632
rect 8668 15623 8720 15632
rect 8668 15589 8677 15623
rect 8677 15589 8711 15623
rect 8711 15589 8720 15623
rect 8668 15580 8720 15589
rect 7288 15555 7340 15564
rect 7288 15521 7297 15555
rect 7297 15521 7331 15555
rect 7331 15521 7340 15555
rect 7288 15512 7340 15521
rect 10324 15512 10376 15564
rect 12348 15512 12400 15564
rect 12900 15512 12952 15564
rect 13360 15580 13412 15632
rect 15844 15648 15896 15700
rect 14648 15623 14700 15632
rect 14648 15589 14657 15623
rect 14657 15589 14691 15623
rect 14691 15589 14700 15623
rect 14648 15580 14700 15589
rect 15476 15623 15528 15632
rect 15476 15589 15485 15623
rect 15485 15589 15519 15623
rect 15519 15589 15528 15623
rect 15476 15580 15528 15589
rect 6644 15444 6696 15496
rect 13820 15512 13872 15564
rect 16212 15555 16264 15564
rect 16212 15521 16221 15555
rect 16221 15521 16255 15555
rect 16255 15521 16264 15555
rect 16212 15512 16264 15521
rect 15752 15444 15804 15496
rect 18052 15487 18104 15496
rect 18052 15453 18061 15487
rect 18061 15453 18095 15487
rect 18095 15453 18104 15487
rect 18052 15444 18104 15453
rect 12992 15308 13044 15360
rect 17316 15351 17368 15360
rect 17316 15317 17325 15351
rect 17325 15317 17359 15351
rect 17359 15317 17368 15351
rect 17316 15308 17368 15317
rect 5982 15206 6034 15258
rect 6046 15206 6098 15258
rect 6110 15206 6162 15258
rect 6174 15206 6226 15258
rect 15982 15206 16034 15258
rect 16046 15206 16098 15258
rect 16110 15206 16162 15258
rect 16174 15206 16226 15258
rect 25982 15206 26034 15258
rect 26046 15206 26098 15258
rect 26110 15206 26162 15258
rect 26174 15206 26226 15258
rect 6644 15147 6696 15156
rect 6644 15113 6653 15147
rect 6653 15113 6687 15147
rect 6687 15113 6696 15147
rect 6644 15104 6696 15113
rect 7288 15104 7340 15156
rect 7840 15147 7892 15156
rect 7840 15113 7849 15147
rect 7849 15113 7883 15147
rect 7883 15113 7892 15147
rect 7840 15104 7892 15113
rect 10324 15147 10376 15156
rect 10324 15113 10333 15147
rect 10333 15113 10367 15147
rect 10367 15113 10376 15147
rect 10324 15104 10376 15113
rect 12348 15104 12400 15156
rect 13360 15104 13412 15156
rect 13636 15104 13688 15156
rect 16304 15104 16356 15156
rect 14924 15036 14976 15088
rect 13268 15011 13320 15020
rect 13268 14977 13277 15011
rect 13277 14977 13311 15011
rect 13311 14977 13320 15011
rect 13268 14968 13320 14977
rect 7840 14900 7892 14952
rect 9864 14900 9916 14952
rect 12624 14943 12676 14952
rect 12624 14909 12633 14943
rect 12633 14909 12667 14943
rect 12667 14909 12676 14943
rect 12624 14900 12676 14909
rect 13268 14832 13320 14884
rect 14464 14900 14516 14952
rect 15016 14900 15068 14952
rect 14924 14832 14976 14884
rect 7012 14764 7064 14816
rect 8576 14764 8628 14816
rect 10324 14764 10376 14816
rect 11428 14764 11480 14816
rect 11888 14764 11940 14816
rect 17316 14900 17368 14952
rect 17132 14875 17184 14884
rect 17132 14841 17141 14875
rect 17141 14841 17175 14875
rect 17175 14841 17184 14875
rect 17132 14832 17184 14841
rect 17776 14764 17828 14816
rect 10982 14662 11034 14714
rect 11046 14662 11098 14714
rect 11110 14662 11162 14714
rect 11174 14662 11226 14714
rect 20982 14662 21034 14714
rect 21046 14662 21098 14714
rect 21110 14662 21162 14714
rect 21174 14662 21226 14714
rect 8576 14560 8628 14612
rect 9772 14560 9824 14612
rect 11796 14560 11848 14612
rect 14464 14603 14516 14612
rect 14464 14569 14473 14603
rect 14473 14569 14507 14603
rect 14507 14569 14516 14603
rect 14464 14560 14516 14569
rect 7564 14535 7616 14544
rect 7564 14501 7573 14535
rect 7573 14501 7607 14535
rect 7607 14501 7616 14535
rect 7564 14492 7616 14501
rect 11520 14492 11572 14544
rect 13728 14535 13780 14544
rect 8300 14424 8352 14476
rect 8576 14467 8628 14476
rect 8576 14433 8585 14467
rect 8585 14433 8619 14467
rect 8619 14433 8628 14467
rect 8576 14424 8628 14433
rect 9588 14424 9640 14476
rect 9956 14467 10008 14476
rect 9956 14433 9965 14467
rect 9965 14433 9999 14467
rect 9999 14433 10008 14467
rect 9956 14424 10008 14433
rect 10232 14424 10284 14476
rect 10692 14424 10744 14476
rect 8116 14399 8168 14408
rect 8116 14365 8125 14399
rect 8125 14365 8159 14399
rect 8159 14365 8168 14399
rect 8116 14356 8168 14365
rect 8484 14399 8536 14408
rect 8484 14365 8493 14399
rect 8493 14365 8527 14399
rect 8527 14365 8536 14399
rect 8484 14356 8536 14365
rect 13728 14501 13737 14535
rect 13737 14501 13771 14535
rect 13771 14501 13780 14535
rect 13728 14492 13780 14501
rect 13820 14492 13872 14544
rect 15016 14492 15068 14544
rect 16304 14492 16356 14544
rect 13084 14467 13136 14476
rect 12348 14356 12400 14408
rect 8760 14288 8812 14340
rect 9496 14288 9548 14340
rect 11612 14288 11664 14340
rect 13084 14433 13093 14467
rect 13093 14433 13127 14467
rect 13127 14433 13136 14467
rect 13084 14424 13136 14433
rect 14648 14424 14700 14476
rect 17132 14467 17184 14476
rect 17132 14433 17141 14467
rect 17141 14433 17175 14467
rect 17175 14433 17184 14467
rect 17132 14424 17184 14433
rect 20444 14492 20496 14544
rect 20628 14492 20680 14544
rect 17408 14424 17460 14476
rect 17592 14424 17644 14476
rect 14924 14399 14976 14408
rect 14924 14365 14933 14399
rect 14933 14365 14967 14399
rect 14967 14365 14976 14399
rect 14924 14356 14976 14365
rect 13636 14288 13688 14340
rect 17776 14288 17828 14340
rect 9128 14263 9180 14272
rect 9128 14229 9137 14263
rect 9137 14229 9171 14263
rect 9171 14229 9180 14263
rect 9128 14220 9180 14229
rect 15752 14220 15804 14272
rect 5982 14118 6034 14170
rect 6046 14118 6098 14170
rect 6110 14118 6162 14170
rect 6174 14118 6226 14170
rect 15982 14118 16034 14170
rect 16046 14118 16098 14170
rect 16110 14118 16162 14170
rect 16174 14118 16226 14170
rect 25982 14118 26034 14170
rect 26046 14118 26098 14170
rect 26110 14118 26162 14170
rect 26174 14118 26226 14170
rect 8484 14016 8536 14068
rect 9956 14059 10008 14068
rect 9956 14025 9965 14059
rect 9965 14025 9999 14059
rect 9999 14025 10008 14059
rect 9956 14016 10008 14025
rect 10692 14059 10744 14068
rect 10692 14025 10701 14059
rect 10701 14025 10735 14059
rect 10735 14025 10744 14059
rect 10692 14016 10744 14025
rect 12164 14016 12216 14068
rect 13084 14016 13136 14068
rect 13636 14016 13688 14068
rect 14280 14059 14332 14068
rect 14280 14025 14289 14059
rect 14289 14025 14323 14059
rect 14323 14025 14332 14059
rect 14280 14016 14332 14025
rect 15384 14059 15436 14068
rect 15384 14025 15393 14059
rect 15393 14025 15427 14059
rect 15427 14025 15436 14059
rect 15384 14016 15436 14025
rect 17132 14059 17184 14068
rect 17132 14025 17141 14059
rect 17141 14025 17175 14059
rect 17175 14025 17184 14059
rect 17132 14016 17184 14025
rect 17408 14059 17460 14068
rect 17408 14025 17417 14059
rect 17417 14025 17451 14059
rect 17451 14025 17460 14059
rect 17408 14016 17460 14025
rect 8116 13948 8168 14000
rect 8300 13880 8352 13932
rect 17592 13948 17644 14000
rect 8392 13855 8444 13864
rect 8392 13821 8401 13855
rect 8401 13821 8435 13855
rect 8435 13821 8444 13855
rect 8392 13812 8444 13821
rect 8760 13812 8812 13864
rect 15568 13923 15620 13932
rect 9128 13812 9180 13864
rect 12164 13855 12216 13864
rect 8944 13744 8996 13796
rect 9220 13744 9272 13796
rect 10048 13744 10100 13796
rect 12164 13821 12173 13855
rect 12173 13821 12207 13855
rect 12207 13821 12216 13855
rect 12164 13812 12216 13821
rect 12808 13855 12860 13864
rect 12808 13821 12817 13855
rect 12817 13821 12851 13855
rect 12851 13821 12860 13855
rect 12808 13812 12860 13821
rect 15568 13889 15577 13923
rect 15577 13889 15611 13923
rect 15611 13889 15620 13923
rect 15568 13880 15620 13889
rect 27620 13923 27672 13932
rect 14648 13855 14700 13864
rect 14648 13821 14657 13855
rect 14657 13821 14691 13855
rect 14691 13821 14700 13855
rect 14648 13812 14700 13821
rect 15384 13812 15436 13864
rect 27620 13889 27629 13923
rect 27629 13889 27663 13923
rect 27663 13889 27672 13923
rect 27620 13880 27672 13889
rect 26516 13812 26568 13864
rect 26240 13744 26292 13796
rect 10876 13676 10928 13728
rect 10982 13574 11034 13626
rect 11046 13574 11098 13626
rect 11110 13574 11162 13626
rect 11174 13574 11226 13626
rect 20982 13574 21034 13626
rect 21046 13574 21098 13626
rect 21110 13574 21162 13626
rect 21174 13574 21226 13626
rect 8300 13472 8352 13524
rect 12808 13472 12860 13524
rect 22560 13515 22612 13524
rect 22560 13481 22569 13515
rect 22569 13481 22603 13515
rect 22603 13481 22612 13515
rect 22560 13472 22612 13481
rect 26240 13515 26292 13524
rect 26240 13481 26249 13515
rect 26249 13481 26283 13515
rect 26283 13481 26292 13515
rect 26240 13472 26292 13481
rect 8484 13447 8536 13456
rect 8484 13413 8493 13447
rect 8493 13413 8527 13447
rect 8527 13413 8536 13447
rect 8484 13404 8536 13413
rect 7380 13336 7432 13388
rect 10692 13379 10744 13388
rect 10692 13345 10701 13379
rect 10701 13345 10735 13379
rect 10735 13345 10744 13379
rect 10692 13336 10744 13345
rect 12256 13379 12308 13388
rect 12256 13345 12265 13379
rect 12265 13345 12299 13379
rect 12299 13345 12308 13379
rect 13544 13379 13596 13388
rect 12256 13336 12308 13345
rect 13544 13345 13553 13379
rect 13553 13345 13587 13379
rect 13587 13345 13596 13379
rect 13544 13336 13596 13345
rect 20536 13336 20588 13388
rect 21548 13336 21600 13388
rect 12348 13268 12400 13320
rect 13912 13268 13964 13320
rect 21456 13311 21508 13320
rect 21456 13277 21465 13311
rect 21465 13277 21499 13311
rect 21499 13277 21508 13311
rect 21456 13268 21508 13277
rect 10784 13200 10836 13252
rect 7012 13132 7064 13184
rect 11060 13175 11112 13184
rect 11060 13141 11069 13175
rect 11069 13141 11103 13175
rect 11103 13141 11112 13175
rect 11060 13132 11112 13141
rect 12348 13132 12400 13184
rect 25044 13132 25096 13184
rect 26516 13132 26568 13184
rect 5982 13030 6034 13082
rect 6046 13030 6098 13082
rect 6110 13030 6162 13082
rect 6174 13030 6226 13082
rect 15982 13030 16034 13082
rect 16046 13030 16098 13082
rect 16110 13030 16162 13082
rect 16174 13030 16226 13082
rect 25982 13030 26034 13082
rect 26046 13030 26098 13082
rect 26110 13030 26162 13082
rect 26174 13030 26226 13082
rect 7380 12971 7432 12980
rect 7380 12937 7389 12971
rect 7389 12937 7423 12971
rect 7423 12937 7432 12971
rect 7380 12928 7432 12937
rect 10048 12971 10100 12980
rect 10048 12937 10057 12971
rect 10057 12937 10091 12971
rect 10091 12937 10100 12971
rect 10048 12928 10100 12937
rect 10692 12971 10744 12980
rect 10692 12937 10701 12971
rect 10701 12937 10735 12971
rect 10735 12937 10744 12971
rect 10692 12928 10744 12937
rect 12256 12928 12308 12980
rect 13912 12971 13964 12980
rect 13912 12937 13921 12971
rect 13921 12937 13955 12971
rect 13955 12937 13964 12971
rect 13912 12928 13964 12937
rect 21456 12928 21508 12980
rect 21640 12971 21692 12980
rect 21640 12937 21649 12971
rect 21649 12937 21683 12971
rect 21683 12937 21692 12971
rect 21640 12928 21692 12937
rect 13544 12903 13596 12912
rect 13544 12869 13553 12903
rect 13553 12869 13587 12903
rect 13587 12869 13596 12903
rect 13544 12860 13596 12869
rect 8944 12835 8996 12844
rect 8944 12801 8953 12835
rect 8953 12801 8987 12835
rect 8987 12801 8996 12835
rect 8944 12792 8996 12801
rect 8668 12767 8720 12776
rect 8668 12733 8677 12767
rect 8677 12733 8711 12767
rect 8711 12733 8720 12767
rect 8668 12724 8720 12733
rect 11060 12724 11112 12776
rect 11336 12631 11388 12640
rect 11336 12597 11345 12631
rect 11345 12597 11379 12631
rect 11379 12597 11388 12631
rect 21272 12724 21324 12776
rect 21732 12724 21784 12776
rect 12624 12631 12676 12640
rect 11336 12588 11388 12597
rect 12624 12597 12633 12631
rect 12633 12597 12667 12631
rect 12667 12597 12676 12631
rect 12624 12588 12676 12597
rect 10982 12486 11034 12538
rect 11046 12486 11098 12538
rect 11110 12486 11162 12538
rect 11174 12486 11226 12538
rect 20982 12486 21034 12538
rect 21046 12486 21098 12538
rect 21110 12486 21162 12538
rect 21174 12486 21226 12538
rect 12624 12384 12676 12436
rect 9864 12248 9916 12300
rect 12348 12316 12400 12368
rect 12992 12316 13044 12368
rect 11704 12248 11756 12300
rect 11980 12291 12032 12300
rect 10324 12180 10376 12232
rect 10600 12180 10652 12232
rect 11980 12257 11989 12291
rect 11989 12257 12023 12291
rect 12023 12257 12032 12291
rect 11980 12248 12032 12257
rect 12532 12180 12584 12232
rect 13268 12291 13320 12300
rect 13268 12257 13277 12291
rect 13277 12257 13311 12291
rect 13311 12257 13320 12291
rect 13268 12248 13320 12257
rect 16948 12248 17000 12300
rect 11428 12155 11480 12164
rect 11428 12121 11437 12155
rect 11437 12121 11471 12155
rect 11471 12121 11480 12155
rect 11428 12112 11480 12121
rect 15292 12112 15344 12164
rect 15752 12112 15804 12164
rect 7932 12044 7984 12096
rect 8668 12087 8720 12096
rect 8668 12053 8677 12087
rect 8677 12053 8711 12087
rect 8711 12053 8720 12087
rect 8668 12044 8720 12053
rect 9956 12087 10008 12096
rect 9956 12053 9965 12087
rect 9965 12053 9999 12087
rect 9999 12053 10008 12087
rect 9956 12044 10008 12053
rect 10416 12087 10468 12096
rect 10416 12053 10425 12087
rect 10425 12053 10459 12087
rect 10459 12053 10468 12087
rect 10416 12044 10468 12053
rect 14188 12087 14240 12096
rect 14188 12053 14197 12087
rect 14197 12053 14231 12087
rect 14231 12053 14240 12087
rect 14188 12044 14240 12053
rect 15568 12087 15620 12096
rect 15568 12053 15577 12087
rect 15577 12053 15611 12087
rect 15611 12053 15620 12087
rect 15568 12044 15620 12053
rect 15844 12087 15896 12096
rect 15844 12053 15853 12087
rect 15853 12053 15887 12087
rect 15887 12053 15896 12087
rect 15844 12044 15896 12053
rect 5982 11942 6034 11994
rect 6046 11942 6098 11994
rect 6110 11942 6162 11994
rect 6174 11942 6226 11994
rect 15982 11942 16034 11994
rect 16046 11942 16098 11994
rect 16110 11942 16162 11994
rect 16174 11942 16226 11994
rect 25982 11942 26034 11994
rect 26046 11942 26098 11994
rect 26110 11942 26162 11994
rect 26174 11942 26226 11994
rect 8944 11840 8996 11892
rect 9496 11883 9548 11892
rect 9496 11849 9505 11883
rect 9505 11849 9539 11883
rect 9539 11849 9548 11883
rect 9496 11840 9548 11849
rect 9864 11883 9916 11892
rect 9864 11849 9873 11883
rect 9873 11849 9907 11883
rect 9907 11849 9916 11883
rect 9864 11840 9916 11849
rect 11980 11840 12032 11892
rect 12992 11840 13044 11892
rect 14924 11883 14976 11892
rect 14924 11849 14933 11883
rect 14933 11849 14967 11883
rect 14967 11849 14976 11883
rect 14924 11840 14976 11849
rect 15384 11883 15436 11892
rect 15384 11849 15393 11883
rect 15393 11849 15427 11883
rect 15427 11849 15436 11883
rect 15384 11840 15436 11849
rect 16948 11883 17000 11892
rect 16948 11849 16957 11883
rect 16957 11849 16991 11883
rect 16991 11849 17000 11883
rect 16948 11840 17000 11849
rect 10416 11636 10468 11688
rect 10324 11611 10376 11620
rect 10324 11577 10333 11611
rect 10333 11577 10367 11611
rect 10367 11577 10376 11611
rect 10324 11568 10376 11577
rect 10876 11636 10928 11688
rect 12532 11772 12584 11824
rect 15752 11772 15804 11824
rect 12164 11747 12216 11756
rect 12164 11713 12173 11747
rect 12173 11713 12207 11747
rect 12207 11713 12216 11747
rect 15568 11747 15620 11756
rect 12164 11704 12216 11713
rect 12440 11679 12492 11688
rect 12440 11645 12449 11679
rect 12449 11645 12483 11679
rect 12483 11645 12492 11679
rect 12624 11679 12676 11688
rect 12440 11636 12492 11645
rect 12624 11645 12633 11679
rect 12633 11645 12667 11679
rect 12667 11645 12676 11679
rect 12624 11636 12676 11645
rect 15568 11713 15577 11747
rect 15577 11713 15611 11747
rect 15611 11713 15620 11747
rect 15568 11704 15620 11713
rect 11336 11568 11388 11620
rect 15936 11636 15988 11688
rect 13728 11611 13780 11620
rect 13728 11577 13737 11611
rect 13737 11577 13771 11611
rect 13771 11577 13780 11611
rect 13728 11568 13780 11577
rect 15660 11568 15712 11620
rect 10982 11398 11034 11450
rect 11046 11398 11098 11450
rect 11110 11398 11162 11450
rect 11174 11398 11226 11450
rect 20982 11398 21034 11450
rect 21046 11398 21098 11450
rect 21110 11398 21162 11450
rect 21174 11398 21226 11450
rect 10876 11296 10928 11348
rect 11704 11296 11756 11348
rect 12348 11296 12400 11348
rect 12440 11339 12492 11348
rect 12440 11305 12449 11339
rect 12449 11305 12483 11339
rect 12483 11305 12492 11339
rect 12440 11296 12492 11305
rect 12624 11296 12676 11348
rect 10784 11228 10836 11280
rect 11336 11271 11388 11280
rect 7012 11160 7064 11212
rect 7840 11160 7892 11212
rect 11336 11237 11345 11271
rect 11345 11237 11379 11271
rect 11379 11237 11388 11271
rect 11336 11228 11388 11237
rect 13268 11296 13320 11348
rect 15936 11296 15988 11348
rect 16948 11296 17000 11348
rect 18052 11296 18104 11348
rect 13360 11228 13412 11280
rect 13636 11203 13688 11212
rect 13636 11169 13645 11203
rect 13645 11169 13679 11203
rect 13679 11169 13688 11203
rect 13636 11160 13688 11169
rect 11520 11092 11572 11144
rect 12808 11092 12860 11144
rect 15660 11160 15712 11212
rect 17960 11203 18012 11212
rect 17960 11169 17969 11203
rect 17969 11169 18003 11203
rect 18003 11169 18012 11203
rect 17960 11160 18012 11169
rect 15292 11135 15344 11144
rect 15292 11101 15301 11135
rect 15301 11101 15335 11135
rect 15335 11101 15344 11135
rect 15292 11092 15344 11101
rect 7932 11024 7984 11076
rect 5982 10854 6034 10906
rect 6046 10854 6098 10906
rect 6110 10854 6162 10906
rect 6174 10854 6226 10906
rect 15982 10854 16034 10906
rect 16046 10854 16098 10906
rect 16110 10854 16162 10906
rect 16174 10854 16226 10906
rect 25982 10854 26034 10906
rect 26046 10854 26098 10906
rect 26110 10854 26162 10906
rect 26174 10854 26226 10906
rect 7840 10795 7892 10804
rect 7840 10761 7849 10795
rect 7849 10761 7883 10795
rect 7883 10761 7892 10795
rect 7840 10752 7892 10761
rect 10784 10795 10836 10804
rect 10784 10761 10793 10795
rect 10793 10761 10827 10795
rect 10827 10761 10836 10795
rect 10784 10752 10836 10761
rect 11336 10752 11388 10804
rect 11520 10752 11572 10804
rect 13452 10752 13504 10804
rect 13636 10752 13688 10804
rect 15660 10752 15712 10804
rect 17868 10795 17920 10804
rect 17868 10761 17877 10795
rect 17877 10761 17911 10795
rect 17911 10761 17920 10795
rect 17868 10752 17920 10761
rect 21364 10752 21416 10804
rect 13360 10727 13412 10736
rect 13360 10693 13369 10727
rect 13369 10693 13403 10727
rect 13403 10693 13412 10727
rect 13360 10684 13412 10693
rect 19248 10659 19300 10668
rect 19248 10625 19257 10659
rect 19257 10625 19291 10659
rect 19291 10625 19300 10659
rect 19248 10616 19300 10625
rect 20536 10616 20588 10668
rect 19064 10523 19116 10532
rect 19064 10489 19073 10523
rect 19073 10489 19107 10523
rect 19107 10489 19116 10523
rect 19064 10480 19116 10489
rect 12808 10412 12860 10464
rect 15292 10412 15344 10464
rect 10982 10310 11034 10362
rect 11046 10310 11098 10362
rect 11110 10310 11162 10362
rect 11174 10310 11226 10362
rect 20982 10310 21034 10362
rect 21046 10310 21098 10362
rect 21110 10310 21162 10362
rect 21174 10310 21226 10362
rect 17960 10208 18012 10260
rect 19248 10251 19300 10260
rect 19248 10217 19257 10251
rect 19257 10217 19291 10251
rect 19291 10217 19300 10251
rect 19248 10208 19300 10217
rect 16396 10115 16448 10124
rect 16396 10081 16405 10115
rect 16405 10081 16439 10115
rect 16439 10081 16448 10115
rect 16396 10072 16448 10081
rect 18052 10072 18104 10124
rect 18788 10072 18840 10124
rect 15752 10004 15804 10056
rect 16488 10004 16540 10056
rect 16580 9911 16632 9920
rect 16580 9877 16589 9911
rect 16589 9877 16623 9911
rect 16623 9877 16632 9911
rect 16580 9868 16632 9877
rect 5982 9766 6034 9818
rect 6046 9766 6098 9818
rect 6110 9766 6162 9818
rect 6174 9766 6226 9818
rect 15982 9766 16034 9818
rect 16046 9766 16098 9818
rect 16110 9766 16162 9818
rect 16174 9766 16226 9818
rect 25982 9766 26034 9818
rect 26046 9766 26098 9818
rect 26110 9766 26162 9818
rect 26174 9766 26226 9818
rect 12624 9664 12676 9716
rect 16396 9664 16448 9716
rect 18788 9707 18840 9716
rect 14924 9528 14976 9580
rect 15476 9571 15528 9580
rect 15476 9537 15485 9571
rect 15485 9537 15519 9571
rect 15519 9537 15528 9571
rect 15476 9528 15528 9537
rect 18788 9673 18797 9707
rect 18797 9673 18831 9707
rect 18831 9673 18840 9707
rect 18788 9664 18840 9673
rect 20536 9596 20588 9648
rect 20720 9596 20772 9648
rect 12440 9460 12492 9512
rect 14464 9503 14516 9512
rect 14464 9469 14473 9503
rect 14473 9469 14507 9503
rect 14507 9469 14516 9503
rect 14464 9460 14516 9469
rect 15292 9460 15344 9512
rect 16488 9460 16540 9512
rect 13268 9324 13320 9376
rect 10982 9222 11034 9274
rect 11046 9222 11098 9274
rect 11110 9222 11162 9274
rect 11174 9222 11226 9274
rect 20982 9222 21034 9274
rect 21046 9222 21098 9274
rect 21110 9222 21162 9274
rect 21174 9222 21226 9274
rect 3056 9095 3108 9104
rect 3056 9061 3065 9095
rect 3065 9061 3099 9095
rect 3099 9061 3108 9095
rect 3056 9052 3108 9061
rect 11612 9052 11664 9104
rect 2044 8984 2096 9036
rect 9680 9027 9732 9036
rect 9680 8993 9689 9027
rect 9689 8993 9723 9027
rect 9723 8993 9732 9027
rect 9680 8984 9732 8993
rect 10324 8984 10376 9036
rect 12624 9027 12676 9036
rect 12624 8993 12633 9027
rect 12633 8993 12667 9027
rect 12667 8993 12676 9027
rect 12624 8984 12676 8993
rect 12992 9027 13044 9036
rect 12992 8993 13001 9027
rect 13001 8993 13035 9027
rect 13035 8993 13044 9027
rect 12992 8984 13044 8993
rect 15476 9052 15528 9104
rect 16580 8984 16632 9036
rect 16948 8984 17000 9036
rect 17040 9027 17092 9036
rect 17040 8993 17049 9027
rect 17049 8993 17083 9027
rect 17083 8993 17092 9027
rect 17040 8984 17092 8993
rect 17592 8984 17644 9036
rect 1584 8916 1636 8968
rect 12164 8959 12216 8968
rect 12164 8925 12173 8959
rect 12173 8925 12207 8959
rect 12207 8925 12216 8959
rect 12164 8916 12216 8925
rect 16488 8891 16540 8900
rect 16488 8857 16497 8891
rect 16497 8857 16531 8891
rect 16531 8857 16540 8891
rect 16488 8848 16540 8857
rect 9680 8780 9732 8832
rect 14096 8780 14148 8832
rect 15476 8823 15528 8832
rect 15476 8789 15485 8823
rect 15485 8789 15519 8823
rect 15519 8789 15528 8823
rect 15476 8780 15528 8789
rect 5982 8678 6034 8730
rect 6046 8678 6098 8730
rect 6110 8678 6162 8730
rect 6174 8678 6226 8730
rect 15982 8678 16034 8730
rect 16046 8678 16098 8730
rect 16110 8678 16162 8730
rect 16174 8678 16226 8730
rect 25982 8678 26034 8730
rect 26046 8678 26098 8730
rect 26110 8678 26162 8730
rect 26174 8678 26226 8730
rect 2044 8619 2096 8628
rect 2044 8585 2053 8619
rect 2053 8585 2087 8619
rect 2087 8585 2096 8619
rect 2044 8576 2096 8585
rect 8852 8619 8904 8628
rect 8852 8585 8861 8619
rect 8861 8585 8895 8619
rect 8895 8585 8904 8619
rect 8852 8576 8904 8585
rect 10232 8576 10284 8628
rect 10324 8576 10376 8628
rect 10600 8576 10652 8628
rect 12624 8619 12676 8628
rect 9680 8415 9732 8424
rect 1584 8347 1636 8356
rect 1584 8313 1593 8347
rect 1593 8313 1627 8347
rect 1627 8313 1636 8347
rect 1584 8304 1636 8313
rect 9036 8347 9088 8356
rect 9036 8313 9045 8347
rect 9045 8313 9079 8347
rect 9079 8313 9088 8347
rect 9036 8304 9088 8313
rect 9680 8381 9689 8415
rect 9689 8381 9723 8415
rect 9723 8381 9732 8415
rect 9680 8372 9732 8381
rect 11612 8508 11664 8560
rect 12624 8585 12633 8619
rect 12633 8585 12667 8619
rect 12667 8585 12676 8619
rect 12624 8576 12676 8585
rect 14004 8576 14056 8628
rect 15568 8576 15620 8628
rect 16580 8619 16632 8628
rect 16580 8585 16589 8619
rect 16589 8585 16623 8619
rect 16623 8585 16632 8619
rect 16580 8576 16632 8585
rect 16948 8619 17000 8628
rect 16948 8585 16957 8619
rect 16957 8585 16991 8619
rect 16991 8585 17000 8619
rect 16948 8576 17000 8585
rect 12992 8508 13044 8560
rect 13268 8508 13320 8560
rect 13728 8483 13780 8492
rect 13728 8449 13737 8483
rect 13737 8449 13771 8483
rect 13771 8449 13780 8483
rect 13728 8440 13780 8449
rect 14004 8483 14056 8492
rect 14004 8449 14013 8483
rect 14013 8449 14047 8483
rect 14047 8449 14056 8483
rect 14004 8440 14056 8449
rect 17040 8508 17092 8560
rect 10232 8415 10284 8424
rect 10232 8381 10241 8415
rect 10241 8381 10275 8415
rect 10275 8381 10284 8415
rect 13268 8415 13320 8424
rect 10232 8372 10284 8381
rect 13268 8381 13277 8415
rect 13277 8381 13311 8415
rect 13311 8381 13320 8415
rect 13268 8372 13320 8381
rect 14096 8415 14148 8424
rect 14096 8381 14105 8415
rect 14105 8381 14139 8415
rect 14139 8381 14148 8415
rect 14096 8372 14148 8381
rect 9128 8236 9180 8288
rect 9864 8304 9916 8356
rect 13820 8304 13872 8356
rect 10982 8134 11034 8186
rect 11046 8134 11098 8186
rect 11110 8134 11162 8186
rect 11174 8134 11226 8186
rect 20982 8134 21034 8186
rect 21046 8134 21098 8186
rect 21110 8134 21162 8186
rect 21174 8134 21226 8186
rect 9128 8075 9180 8084
rect 9128 8041 9137 8075
rect 9137 8041 9171 8075
rect 9171 8041 9180 8075
rect 9128 8032 9180 8041
rect 9772 8032 9824 8084
rect 12440 8075 12492 8084
rect 12440 8041 12449 8075
rect 12449 8041 12483 8075
rect 12483 8041 12492 8075
rect 13820 8075 13872 8084
rect 12440 8032 12492 8041
rect 13820 8041 13829 8075
rect 13829 8041 13863 8075
rect 13863 8041 13872 8075
rect 13820 8032 13872 8041
rect 18144 8075 18196 8084
rect 18144 8041 18153 8075
rect 18153 8041 18187 8075
rect 18187 8041 18196 8075
rect 18144 8032 18196 8041
rect 13452 7964 13504 8016
rect 14004 7964 14056 8016
rect 11060 7939 11112 7948
rect 11060 7905 11069 7939
rect 11069 7905 11103 7939
rect 11103 7905 11112 7939
rect 11060 7896 11112 7905
rect 11612 7896 11664 7948
rect 16856 7939 16908 7948
rect 16856 7905 16865 7939
rect 16865 7905 16899 7939
rect 16899 7905 16908 7939
rect 16856 7896 16908 7905
rect 16948 7828 17000 7880
rect 5982 7590 6034 7642
rect 6046 7590 6098 7642
rect 6110 7590 6162 7642
rect 6174 7590 6226 7642
rect 15982 7590 16034 7642
rect 16046 7590 16098 7642
rect 16110 7590 16162 7642
rect 16174 7590 16226 7642
rect 25982 7590 26034 7642
rect 26046 7590 26098 7642
rect 26110 7590 26162 7642
rect 26174 7590 26226 7642
rect 11612 7488 11664 7540
rect 14096 7488 14148 7540
rect 16856 7488 16908 7540
rect 16948 7488 17000 7540
rect 17868 7488 17920 7540
rect 11060 7420 11112 7472
rect 13820 7352 13872 7404
rect 13084 7327 13136 7336
rect 13084 7293 13093 7327
rect 13093 7293 13127 7327
rect 13127 7293 13136 7327
rect 13084 7284 13136 7293
rect 10982 7046 11034 7098
rect 11046 7046 11098 7098
rect 11110 7046 11162 7098
rect 11174 7046 11226 7098
rect 20982 7046 21034 7098
rect 21046 7046 21098 7098
rect 21110 7046 21162 7098
rect 21174 7046 21226 7098
rect 13084 6647 13136 6656
rect 13084 6613 13093 6647
rect 13093 6613 13127 6647
rect 13127 6613 13136 6647
rect 14556 6647 14608 6656
rect 13084 6604 13136 6613
rect 14556 6613 14565 6647
rect 14565 6613 14599 6647
rect 14599 6613 14608 6647
rect 14556 6604 14608 6613
rect 5982 6502 6034 6554
rect 6046 6502 6098 6554
rect 6110 6502 6162 6554
rect 6174 6502 6226 6554
rect 15982 6502 16034 6554
rect 16046 6502 16098 6554
rect 16110 6502 16162 6554
rect 16174 6502 16226 6554
rect 25982 6502 26034 6554
rect 26046 6502 26098 6554
rect 26110 6502 26162 6554
rect 26174 6502 26226 6554
rect 14188 6400 14240 6452
rect 16304 6264 16356 6316
rect 14556 6239 14608 6248
rect 14556 6205 14565 6239
rect 14565 6205 14599 6239
rect 14599 6205 14608 6239
rect 14556 6196 14608 6205
rect 15936 6103 15988 6112
rect 15936 6069 15945 6103
rect 15945 6069 15979 6103
rect 15979 6069 15988 6103
rect 15936 6060 15988 6069
rect 10982 5958 11034 6010
rect 11046 5958 11098 6010
rect 11110 5958 11162 6010
rect 11174 5958 11226 6010
rect 20982 5958 21034 6010
rect 21046 5958 21098 6010
rect 21110 5958 21162 6010
rect 21174 5958 21226 6010
rect 13360 5788 13412 5840
rect 13820 5763 13872 5772
rect 13820 5729 13829 5763
rect 13829 5729 13863 5763
rect 13863 5729 13872 5763
rect 13820 5720 13872 5729
rect 14188 5763 14240 5772
rect 14188 5729 14197 5763
rect 14197 5729 14231 5763
rect 14231 5729 14240 5763
rect 14188 5720 14240 5729
rect 15292 5788 15344 5840
rect 15752 5788 15804 5840
rect 15936 5763 15988 5772
rect 15936 5729 15945 5763
rect 15945 5729 15979 5763
rect 15979 5729 15988 5763
rect 15936 5720 15988 5729
rect 16304 5763 16356 5772
rect 16304 5729 16313 5763
rect 16313 5729 16347 5763
rect 16347 5729 16356 5763
rect 16304 5720 16356 5729
rect 13728 5652 13780 5704
rect 14004 5652 14056 5704
rect 15660 5584 15712 5636
rect 13084 5559 13136 5568
rect 13084 5525 13093 5559
rect 13093 5525 13127 5559
rect 13127 5525 13136 5559
rect 13084 5516 13136 5525
rect 13452 5559 13504 5568
rect 13452 5525 13461 5559
rect 13461 5525 13495 5559
rect 13495 5525 13504 5559
rect 13452 5516 13504 5525
rect 15568 5559 15620 5568
rect 15568 5525 15577 5559
rect 15577 5525 15611 5559
rect 15611 5525 15620 5559
rect 15568 5516 15620 5525
rect 5982 5414 6034 5466
rect 6046 5414 6098 5466
rect 6110 5414 6162 5466
rect 6174 5414 6226 5466
rect 15982 5414 16034 5466
rect 16046 5414 16098 5466
rect 16110 5414 16162 5466
rect 16174 5414 16226 5466
rect 25982 5414 26034 5466
rect 26046 5414 26098 5466
rect 26110 5414 26162 5466
rect 26174 5414 26226 5466
rect 11428 5312 11480 5364
rect 13360 5312 13412 5364
rect 15292 5355 15344 5364
rect 15292 5321 15301 5355
rect 15301 5321 15335 5355
rect 15335 5321 15344 5355
rect 15292 5312 15344 5321
rect 15660 5355 15712 5364
rect 15660 5321 15669 5355
rect 15669 5321 15703 5355
rect 15703 5321 15712 5355
rect 15660 5312 15712 5321
rect 15844 5312 15896 5364
rect 13084 5151 13136 5160
rect 13084 5117 13093 5151
rect 13093 5117 13127 5151
rect 13127 5117 13136 5151
rect 13084 5108 13136 5117
rect 14188 5108 14240 5160
rect 13636 4972 13688 5024
rect 13820 4972 13872 5024
rect 10982 4870 11034 4922
rect 11046 4870 11098 4922
rect 11110 4870 11162 4922
rect 11174 4870 11226 4922
rect 20982 4870 21034 4922
rect 21046 4870 21098 4922
rect 21110 4870 21162 4922
rect 21174 4870 21226 4922
rect 13636 4811 13688 4820
rect 13636 4777 13645 4811
rect 13645 4777 13679 4811
rect 13679 4777 13688 4811
rect 13636 4768 13688 4777
rect 14188 4768 14240 4820
rect 16304 4768 16356 4820
rect 13544 4700 13596 4752
rect 10876 4632 10928 4684
rect 11520 4632 11572 4684
rect 13728 4632 13780 4684
rect 5982 4326 6034 4378
rect 6046 4326 6098 4378
rect 6110 4326 6162 4378
rect 6174 4326 6226 4378
rect 15982 4326 16034 4378
rect 16046 4326 16098 4378
rect 16110 4326 16162 4378
rect 16174 4326 16226 4378
rect 25982 4326 26034 4378
rect 26046 4326 26098 4378
rect 26110 4326 26162 4378
rect 26174 4326 26226 4378
rect 2780 4088 2832 4140
rect 3700 4088 3752 4140
rect 10876 4088 10928 4140
rect 13820 4088 13872 4140
rect 15108 4088 15160 4140
rect 11520 3952 11572 4004
rect 10982 3782 11034 3834
rect 11046 3782 11098 3834
rect 11110 3782 11162 3834
rect 11174 3782 11226 3834
rect 20982 3782 21034 3834
rect 21046 3782 21098 3834
rect 21110 3782 21162 3834
rect 21174 3782 21226 3834
rect 9864 3680 9916 3732
rect 10784 3680 10836 3732
rect 11796 3723 11848 3732
rect 11796 3689 11805 3723
rect 11805 3689 11839 3723
rect 11839 3689 11848 3723
rect 11796 3680 11848 3689
rect 19432 3723 19484 3732
rect 19432 3689 19441 3723
rect 19441 3689 19475 3723
rect 19475 3689 19484 3723
rect 19432 3680 19484 3689
rect 17960 3544 18012 3596
rect 10600 3476 10652 3528
rect 18144 3519 18196 3528
rect 18144 3485 18153 3519
rect 18153 3485 18187 3519
rect 18187 3485 18196 3519
rect 18144 3476 18196 3485
rect 5982 3238 6034 3290
rect 6046 3238 6098 3290
rect 6110 3238 6162 3290
rect 6174 3238 6226 3290
rect 15982 3238 16034 3290
rect 16046 3238 16098 3290
rect 16110 3238 16162 3290
rect 16174 3238 16226 3290
rect 25982 3238 26034 3290
rect 26046 3238 26098 3290
rect 26110 3238 26162 3290
rect 26174 3238 26226 3290
rect 11336 3136 11388 3188
rect 18144 3136 18196 3188
rect 18420 3136 18472 3188
rect 17960 3068 18012 3120
rect 10140 3043 10192 3052
rect 10140 3009 10149 3043
rect 10149 3009 10183 3043
rect 10183 3009 10192 3043
rect 10140 3000 10192 3009
rect 9864 2975 9916 2984
rect 9864 2941 9873 2975
rect 9873 2941 9907 2975
rect 9907 2941 9916 2975
rect 9864 2932 9916 2941
rect 10982 2694 11034 2746
rect 11046 2694 11098 2746
rect 11110 2694 11162 2746
rect 11174 2694 11226 2746
rect 20982 2694 21034 2746
rect 21046 2694 21098 2746
rect 21110 2694 21162 2746
rect 21174 2694 21226 2746
rect 10784 2635 10836 2644
rect 10784 2601 10793 2635
rect 10793 2601 10827 2635
rect 10827 2601 10836 2635
rect 10784 2592 10836 2601
rect 14004 2635 14056 2644
rect 14004 2601 14013 2635
rect 14013 2601 14047 2635
rect 14047 2601 14056 2635
rect 14004 2592 14056 2601
rect 17960 2592 18012 2644
rect 21456 2592 21508 2644
rect 12440 2456 12492 2508
rect 13084 2388 13136 2440
rect 17960 2388 18012 2440
rect 18604 2431 18656 2440
rect 18604 2397 18613 2431
rect 18613 2397 18647 2431
rect 18647 2397 18656 2431
rect 18604 2388 18656 2397
rect 21456 2431 21508 2440
rect 21456 2397 21465 2431
rect 21465 2397 21499 2431
rect 21499 2397 21508 2431
rect 21456 2388 21508 2397
rect 20260 2320 20312 2372
rect 20628 2320 20680 2372
rect 20904 2363 20956 2372
rect 20904 2329 20913 2363
rect 20913 2329 20947 2363
rect 20947 2329 20956 2363
rect 20904 2320 20956 2329
rect 10600 2252 10652 2304
rect 12440 2295 12492 2304
rect 12440 2261 12449 2295
rect 12449 2261 12483 2295
rect 12483 2261 12492 2295
rect 12440 2252 12492 2261
rect 18144 2252 18196 2304
rect 24860 2252 24912 2304
rect 5982 2150 6034 2202
rect 6046 2150 6098 2202
rect 6110 2150 6162 2202
rect 6174 2150 6226 2202
rect 15982 2150 16034 2202
rect 16046 2150 16098 2202
rect 16110 2150 16162 2202
rect 16174 2150 16226 2202
rect 25982 2150 26034 2202
rect 26046 2150 26098 2202
rect 26110 2150 26162 2202
rect 26174 2150 26226 2202
<< metal2 >>
rect 18 79200 74 80000
rect 938 79200 994 80000
rect 1858 79200 1914 80000
rect 2318 79200 2374 80000
rect 3238 79200 3294 80000
rect 4066 79656 4122 79665
rect 4066 79591 4122 79600
rect 32 76922 60 79200
rect 952 79098 980 79200
rect 952 79070 1348 79098
rect 32 76894 152 76922
rect 124 72729 152 76894
rect 110 72720 166 72729
rect 110 72655 166 72664
rect 1320 21593 1348 79070
rect 1872 75886 1900 79200
rect 1400 75880 1452 75886
rect 1400 75822 1452 75828
rect 1860 75880 1912 75886
rect 2332 75857 2360 79200
rect 1860 75822 1912 75828
rect 2318 75848 2374 75857
rect 1412 73681 1440 75822
rect 2318 75783 2374 75792
rect 2962 75576 3018 75585
rect 2962 75511 3018 75520
rect 1398 73672 1454 73681
rect 1398 73607 1454 73616
rect 1766 72176 1822 72185
rect 1766 72111 1822 72120
rect 1676 69896 1728 69902
rect 1676 69838 1728 69844
rect 1584 69420 1636 69426
rect 1584 69362 1636 69368
rect 1596 61402 1624 69362
rect 1688 69358 1716 69838
rect 1676 69352 1728 69358
rect 1674 69320 1676 69329
rect 1728 69320 1730 69329
rect 1674 69255 1730 69264
rect 1584 61396 1636 61402
rect 1584 61338 1636 61344
rect 1596 60722 1624 61338
rect 1584 60716 1636 60722
rect 1584 60658 1636 60664
rect 1676 60648 1728 60654
rect 1676 60590 1728 60596
rect 1688 59974 1716 60590
rect 1676 59968 1728 59974
rect 1676 59910 1728 59916
rect 1674 57216 1730 57225
rect 1674 57151 1730 57160
rect 1688 56914 1716 57151
rect 1676 56908 1728 56914
rect 1676 56850 1728 56856
rect 1584 56840 1636 56846
rect 1584 56782 1636 56788
rect 1596 52494 1624 56782
rect 1688 56506 1716 56850
rect 1676 56500 1728 56506
rect 1676 56442 1728 56448
rect 1674 53816 1730 53825
rect 1674 53751 1730 53760
rect 1688 52562 1716 53751
rect 1676 52556 1728 52562
rect 1676 52498 1728 52504
rect 1584 52488 1636 52494
rect 1584 52430 1636 52436
rect 1596 51814 1624 52430
rect 1688 52154 1716 52498
rect 1676 52148 1728 52154
rect 1676 52090 1728 52096
rect 1584 51808 1636 51814
rect 1584 51750 1636 51756
rect 1596 50969 1624 51750
rect 1582 50960 1638 50969
rect 1582 50895 1638 50904
rect 1596 45830 1624 50895
rect 1584 45824 1636 45830
rect 1584 45766 1636 45772
rect 1596 45490 1624 45766
rect 1780 45490 1808 72111
rect 2778 71496 2834 71505
rect 2778 71431 2834 71440
rect 2792 70106 2820 71431
rect 2780 70100 2832 70106
rect 2780 70042 2832 70048
rect 2044 69964 2096 69970
rect 2044 69906 2096 69912
rect 2056 69465 2084 69906
rect 2042 69456 2098 69465
rect 2042 69391 2044 69400
rect 2096 69391 2098 69400
rect 2044 69362 2096 69368
rect 2778 61976 2834 61985
rect 2778 61911 2834 61920
rect 2792 60858 2820 61911
rect 2780 60852 2832 60858
rect 2780 60794 2832 60800
rect 2044 59968 2096 59974
rect 2044 59910 2096 59916
rect 2870 59936 2926 59945
rect 1950 45656 2006 45665
rect 1950 45591 2006 45600
rect 1584 45484 1636 45490
rect 1584 45426 1636 45432
rect 1768 45484 1820 45490
rect 1768 45426 1820 45432
rect 1596 44742 1624 45426
rect 1780 45082 1808 45426
rect 1964 45082 1992 45591
rect 1768 45076 1820 45082
rect 1768 45018 1820 45024
rect 1952 45076 2004 45082
rect 1952 45018 2004 45024
rect 1766 44976 1822 44985
rect 1766 44911 1822 44920
rect 1584 44736 1636 44742
rect 1584 44678 1636 44684
rect 1596 44402 1624 44678
rect 1584 44396 1636 44402
rect 1584 44338 1636 44344
rect 1596 43858 1624 44338
rect 1584 43852 1636 43858
rect 1584 43794 1636 43800
rect 1596 43246 1624 43794
rect 1780 43314 1808 44911
rect 1964 44334 1992 45018
rect 1952 44328 2004 44334
rect 1952 44270 2004 44276
rect 1768 43308 1820 43314
rect 1768 43250 1820 43256
rect 1584 43240 1636 43246
rect 1584 43182 1636 43188
rect 1596 42838 1624 43182
rect 1780 42906 1808 43250
rect 1768 42900 1820 42906
rect 1768 42842 1820 42848
rect 1584 42832 1636 42838
rect 1584 42774 1636 42780
rect 1596 42362 1624 42774
rect 1584 42356 1636 42362
rect 1584 42298 1636 42304
rect 1766 41576 1822 41585
rect 1766 41511 1822 41520
rect 1492 40384 1544 40390
rect 1492 40326 1544 40332
rect 1504 39982 1532 40326
rect 1780 40050 1808 41511
rect 1768 40044 1820 40050
rect 1768 39986 1820 39992
rect 1492 39976 1544 39982
rect 1492 39918 1544 39924
rect 1504 38962 1532 39918
rect 1780 39642 1808 39986
rect 1768 39636 1820 39642
rect 1768 39578 1820 39584
rect 1492 38956 1544 38962
rect 1492 38898 1544 38904
rect 1768 38956 1820 38962
rect 1768 38898 1820 38904
rect 1676 38888 1728 38894
rect 1596 38836 1676 38842
rect 1596 38830 1728 38836
rect 1780 38842 1808 38898
rect 1596 38814 1716 38830
rect 1780 38814 1900 38842
rect 1400 38276 1452 38282
rect 1400 38218 1452 38224
rect 1412 37262 1440 38218
rect 1596 38214 1624 38814
rect 1872 38282 1900 38814
rect 1860 38276 1912 38282
rect 1860 38218 1912 38224
rect 1584 38208 1636 38214
rect 1584 38150 1636 38156
rect 1400 37256 1452 37262
rect 1400 37198 1452 37204
rect 1412 36718 1440 37198
rect 1400 36712 1452 36718
rect 1400 36654 1452 36660
rect 1400 35488 1452 35494
rect 1596 35465 1624 38150
rect 1674 37496 1730 37505
rect 1674 37431 1730 37440
rect 1688 37330 1716 37431
rect 1676 37324 1728 37330
rect 1676 37266 1728 37272
rect 1688 36922 1716 37266
rect 1676 36916 1728 36922
rect 1676 36858 1728 36864
rect 1860 35624 1912 35630
rect 1860 35566 1912 35572
rect 1676 35488 1728 35494
rect 1400 35430 1452 35436
rect 1582 35456 1638 35465
rect 1412 34950 1440 35430
rect 1676 35430 1728 35436
rect 1582 35391 1638 35400
rect 1400 34944 1452 34950
rect 1400 34886 1452 34892
rect 1412 34542 1440 34886
rect 1688 34542 1716 35430
rect 1400 34536 1452 34542
rect 1400 34478 1452 34484
rect 1676 34536 1728 34542
rect 1676 34478 1728 34484
rect 1412 31890 1440 34478
rect 1688 34202 1716 34478
rect 1676 34196 1728 34202
rect 1676 34138 1728 34144
rect 1400 31884 1452 31890
rect 1400 31826 1452 31832
rect 1676 31816 1728 31822
rect 1676 31758 1728 31764
rect 1688 31142 1716 31758
rect 1676 31136 1728 31142
rect 1872 31090 1900 35566
rect 1952 31816 2004 31822
rect 1952 31758 2004 31764
rect 1964 31210 1992 31758
rect 1952 31204 2004 31210
rect 1952 31146 2004 31152
rect 1676 31078 1728 31084
rect 1780 31062 1900 31090
rect 1400 29028 1452 29034
rect 1400 28970 1452 28976
rect 1412 28626 1440 28970
rect 1400 28620 1452 28626
rect 1400 28562 1452 28568
rect 1412 28082 1440 28562
rect 1584 28552 1636 28558
rect 1584 28494 1636 28500
rect 1400 28076 1452 28082
rect 1400 28018 1452 28024
rect 1412 27674 1440 28018
rect 1400 27668 1452 27674
rect 1400 27610 1452 27616
rect 1412 27130 1440 27610
rect 1596 27334 1624 28494
rect 1584 27328 1636 27334
rect 1584 27270 1636 27276
rect 1400 27124 1452 27130
rect 1400 27066 1452 27072
rect 1412 26450 1440 27066
rect 1596 26625 1624 27270
rect 1582 26616 1638 26625
rect 1582 26551 1638 26560
rect 1400 26444 1452 26450
rect 1400 26386 1452 26392
rect 1676 26376 1728 26382
rect 1676 26318 1728 26324
rect 1688 26042 1716 26318
rect 1676 26036 1728 26042
rect 1676 25978 1728 25984
rect 1688 25498 1716 25978
rect 1676 25492 1728 25498
rect 1676 25434 1728 25440
rect 1780 25430 1808 31062
rect 1964 29034 1992 31146
rect 1952 29028 2004 29034
rect 1952 28970 2004 28976
rect 1860 28008 1912 28014
rect 1860 27950 1912 27956
rect 1872 27334 1900 27950
rect 1860 27328 1912 27334
rect 1860 27270 1912 27276
rect 1768 25424 1820 25430
rect 1768 25366 1820 25372
rect 1400 25356 1452 25362
rect 1400 25298 1452 25304
rect 1412 24682 1440 25298
rect 1400 24676 1452 24682
rect 1400 24618 1452 24624
rect 1306 21584 1362 21593
rect 1306 21519 1362 21528
rect 1584 21004 1636 21010
rect 1584 20946 1636 20952
rect 1596 20262 1624 20946
rect 1872 20505 1900 27270
rect 1952 25356 2004 25362
rect 1952 25298 2004 25304
rect 1964 24614 1992 25298
rect 1952 24608 2004 24614
rect 1952 24550 2004 24556
rect 1964 23905 1992 24550
rect 1950 23896 2006 23905
rect 1950 23831 2006 23840
rect 1858 20496 1914 20505
rect 1858 20431 1914 20440
rect 1584 20256 1636 20262
rect 1584 20198 1636 20204
rect 1492 18080 1544 18086
rect 1492 18022 1544 18028
rect 1504 17105 1532 18022
rect 1490 17096 1546 17105
rect 1490 17031 1546 17040
rect 1596 12345 1624 20198
rect 1860 18216 1912 18222
rect 1912 18176 1992 18204
rect 1860 18158 1912 18164
rect 1964 17542 1992 18176
rect 1952 17536 2004 17542
rect 1952 17478 2004 17484
rect 1674 17232 1730 17241
rect 1674 17167 1676 17176
rect 1728 17167 1730 17176
rect 1676 17138 1728 17144
rect 1688 16794 1716 17138
rect 1964 17134 1992 17478
rect 1952 17128 2004 17134
rect 1952 17070 2004 17076
rect 1676 16788 1728 16794
rect 1676 16730 1728 16736
rect 1964 16454 1992 17070
rect 1952 16448 2004 16454
rect 1952 16390 2004 16396
rect 2056 13705 2084 59910
rect 2870 59871 2926 59880
rect 2884 58682 2912 59871
rect 2872 58676 2924 58682
rect 2872 58618 2924 58624
rect 2686 57488 2742 57497
rect 2976 57458 3004 75511
rect 3252 74905 3280 79200
rect 3330 78296 3386 78305
rect 3330 78231 3386 78240
rect 3344 77382 3372 78231
rect 4080 77489 4108 79591
rect 4158 79200 4214 80000
rect 4618 79200 4674 80000
rect 5538 79200 5594 80000
rect 6458 79200 6514 80000
rect 6918 79200 6974 80000
rect 7838 79200 7894 80000
rect 8758 79200 8814 80000
rect 9678 79200 9734 80000
rect 10138 79200 10194 80000
rect 11058 79200 11114 80000
rect 11978 79200 12034 80000
rect 12438 79200 12494 80000
rect 13358 79200 13414 80000
rect 14278 79200 14334 80000
rect 14738 79200 14794 80000
rect 15658 79200 15714 80000
rect 16578 79200 16634 80000
rect 17498 79200 17554 80000
rect 17958 79200 18014 80000
rect 18878 79200 18934 80000
rect 19798 79200 19854 80000
rect 20258 79200 20314 80000
rect 21178 79200 21234 80000
rect 22098 79200 22154 80000
rect 22558 79200 22614 80000
rect 23478 79200 23534 80000
rect 24398 79200 24454 80000
rect 24674 79656 24730 79665
rect 24674 79591 24730 79600
rect 4066 77480 4122 77489
rect 4066 77415 4122 77424
rect 3332 77376 3384 77382
rect 3332 77318 3384 77324
rect 3238 74896 3294 74905
rect 3238 74831 3294 74840
rect 4172 74798 4200 79200
rect 4160 74792 4212 74798
rect 3422 74760 3478 74769
rect 4160 74734 4212 74740
rect 3422 74695 3478 74704
rect 3238 68776 3294 68785
rect 3238 68711 3294 68720
rect 3054 58576 3110 58585
rect 3054 58511 3110 58520
rect 2686 57423 2688 57432
rect 2740 57423 2742 57432
rect 2964 57452 3016 57458
rect 2688 57394 2740 57400
rect 2964 57394 3016 57400
rect 2136 57248 2188 57254
rect 2136 57190 2188 57196
rect 2226 57216 2282 57225
rect 2148 57050 2176 57190
rect 2226 57151 2282 57160
rect 2136 57044 2188 57050
rect 2136 56986 2188 56992
rect 2136 56840 2188 56846
rect 2240 56794 2268 57151
rect 2188 56788 2268 56794
rect 2136 56782 2268 56788
rect 2148 56766 2268 56782
rect 2240 56506 2268 56766
rect 2228 56500 2280 56506
rect 2228 56442 2280 56448
rect 2962 44568 3018 44577
rect 2962 44503 2964 44512
rect 3016 44503 3018 44512
rect 2964 44474 3016 44480
rect 2228 43784 2280 43790
rect 2228 43726 2280 43732
rect 2240 42566 2268 43726
rect 2228 42560 2280 42566
rect 2228 42502 2280 42508
rect 2134 40216 2190 40225
rect 2134 40151 2190 40160
rect 2148 36786 2176 40151
rect 2136 36780 2188 36786
rect 2136 36722 2188 36728
rect 2148 36378 2176 36722
rect 2136 36372 2188 36378
rect 2136 36314 2188 36320
rect 2136 26444 2188 26450
rect 2136 26386 2188 26392
rect 2148 26042 2176 26386
rect 2136 26036 2188 26042
rect 2136 25978 2188 25984
rect 2148 20942 2176 25978
rect 2136 20936 2188 20942
rect 2136 20878 2188 20884
rect 2148 20602 2176 20878
rect 2136 20596 2188 20602
rect 2136 20538 2188 20544
rect 2042 13696 2098 13705
rect 2042 13631 2098 13640
rect 1582 12336 1638 12345
rect 1582 12271 1638 12280
rect 2042 9072 2098 9081
rect 2042 9007 2044 9016
rect 2096 9007 2098 9016
rect 2044 8978 2096 8984
rect 1584 8968 1636 8974
rect 1584 8910 1636 8916
rect 1596 8362 1624 8910
rect 2056 8634 2084 8978
rect 2044 8628 2096 8634
rect 2044 8570 2096 8576
rect 1584 8356 1636 8362
rect 1584 8298 1636 8304
rect 18 7984 74 7993
rect 18 7919 74 7928
rect 32 800 60 7919
rect 1596 7585 1624 8298
rect 1582 7576 1638 7585
rect 1582 7511 1638 7520
rect 2240 6610 2268 42502
rect 2318 41440 2374 41449
rect 2318 41375 2374 41384
rect 2332 35562 2360 41375
rect 2412 36712 2464 36718
rect 2412 36654 2464 36660
rect 2424 36038 2452 36654
rect 2412 36032 2464 36038
rect 2412 35974 2464 35980
rect 2424 35766 2452 35974
rect 2412 35760 2464 35766
rect 2412 35702 2464 35708
rect 2870 35728 2926 35737
rect 2870 35663 2872 35672
rect 2924 35663 2926 35672
rect 2872 35634 2924 35640
rect 2320 35556 2372 35562
rect 2320 35498 2372 35504
rect 2780 34400 2832 34406
rect 2780 34342 2832 34348
rect 2792 34105 2820 34342
rect 2778 34096 2834 34105
rect 2778 34031 2834 34040
rect 2870 33416 2926 33425
rect 2870 33351 2926 33360
rect 2884 32026 2912 33351
rect 2872 32020 2924 32026
rect 2872 31962 2924 31968
rect 2964 31136 3016 31142
rect 2964 31078 3016 31084
rect 2686 25256 2742 25265
rect 2686 25191 2742 25200
rect 2700 24750 2728 25191
rect 2976 24800 3004 31078
rect 3068 26518 3096 58511
rect 3148 58472 3200 58478
rect 3148 58414 3200 58420
rect 3160 57934 3188 58414
rect 3148 57928 3200 57934
rect 3148 57870 3200 57876
rect 3148 43784 3200 43790
rect 3146 43752 3148 43761
rect 3200 43752 3202 43761
rect 3146 43687 3202 43696
rect 3148 43240 3200 43246
rect 3146 43208 3148 43217
rect 3200 43208 3202 43217
rect 3146 43143 3202 43152
rect 3252 41449 3280 68711
rect 3436 62801 3464 74695
rect 4632 74662 4660 79200
rect 5354 75848 5410 75857
rect 5354 75783 5410 75792
rect 4620 74656 4672 74662
rect 4620 74598 4672 74604
rect 5368 73137 5396 75783
rect 5448 74792 5500 74798
rect 5552 74769 5580 79200
rect 5956 77276 6252 77296
rect 6012 77274 6036 77276
rect 6092 77274 6116 77276
rect 6172 77274 6196 77276
rect 6034 77222 6036 77274
rect 6098 77222 6110 77274
rect 6172 77222 6174 77274
rect 6012 77220 6036 77222
rect 6092 77220 6116 77222
rect 6172 77220 6196 77222
rect 5956 77200 6252 77220
rect 5956 76188 6252 76208
rect 6012 76186 6036 76188
rect 6092 76186 6116 76188
rect 6172 76186 6196 76188
rect 6034 76134 6036 76186
rect 6098 76134 6110 76186
rect 6172 76134 6174 76186
rect 6012 76132 6036 76134
rect 6092 76132 6116 76134
rect 6172 76132 6196 76134
rect 5956 76112 6252 76132
rect 5956 75100 6252 75120
rect 6012 75098 6036 75100
rect 6092 75098 6116 75100
rect 6172 75098 6196 75100
rect 6034 75046 6036 75098
rect 6098 75046 6110 75098
rect 6172 75046 6174 75098
rect 6012 75044 6036 75046
rect 6092 75044 6116 75046
rect 6172 75044 6196 75046
rect 5956 75024 6252 75044
rect 5630 74896 5686 74905
rect 5630 74831 5686 74840
rect 5448 74734 5500 74740
rect 5538 74760 5594 74769
rect 5354 73128 5410 73137
rect 5354 73063 5410 73072
rect 4066 66736 4122 66745
rect 4066 66671 4122 66680
rect 4080 66065 4108 66671
rect 4066 66056 4122 66065
rect 4066 65991 4122 66000
rect 4802 65240 4858 65249
rect 4802 65175 4858 65184
rect 4816 64569 4844 65175
rect 4802 64560 4858 64569
rect 4802 64495 4858 64504
rect 3790 63336 3846 63345
rect 3790 63271 3846 63280
rect 3422 62792 3478 62801
rect 3422 62727 3478 62736
rect 3332 57928 3384 57934
rect 3330 57896 3332 57905
rect 3384 57896 3386 57905
rect 3330 57831 3386 57840
rect 3608 57860 3660 57866
rect 3344 57225 3372 57831
rect 3608 57802 3660 57808
rect 3620 57390 3648 57802
rect 3608 57384 3660 57390
rect 3608 57326 3660 57332
rect 3620 57225 3648 57326
rect 3330 57216 3386 57225
rect 3330 57151 3386 57160
rect 3606 57216 3662 57225
rect 3606 57151 3662 57160
rect 3422 55856 3478 55865
rect 3422 55791 3478 55800
rect 3436 43625 3464 55791
rect 3698 49056 3754 49065
rect 3698 48991 3754 49000
rect 3514 48648 3570 48657
rect 3514 48583 3570 48592
rect 3422 43616 3478 43625
rect 3422 43551 3478 43560
rect 3330 43072 3386 43081
rect 3330 43007 3386 43016
rect 3238 41440 3294 41449
rect 3238 41375 3294 41384
rect 3148 39908 3200 39914
rect 3148 39850 3200 39856
rect 3160 39545 3188 39850
rect 3146 39536 3202 39545
rect 3146 39471 3202 39480
rect 3344 39098 3372 43007
rect 3332 39092 3384 39098
rect 3332 39034 3384 39040
rect 3146 38992 3202 39001
rect 3146 38927 3202 38936
rect 3160 37398 3188 38927
rect 3148 37392 3200 37398
rect 3148 37334 3200 37340
rect 3240 36576 3292 36582
rect 3240 36518 3292 36524
rect 3252 30569 3280 36518
rect 3424 35080 3476 35086
rect 3424 35022 3476 35028
rect 3436 34950 3464 35022
rect 3424 34944 3476 34950
rect 3424 34886 3476 34892
rect 3436 34202 3464 34886
rect 3424 34196 3476 34202
rect 3424 34138 3476 34144
rect 3424 32904 3476 32910
rect 3424 32846 3476 32852
rect 3436 32570 3464 32846
rect 3424 32564 3476 32570
rect 3424 32506 3476 32512
rect 3238 30560 3294 30569
rect 3238 30495 3294 30504
rect 3146 29200 3202 29209
rect 3146 29135 3202 29144
rect 3160 28218 3188 29135
rect 3148 28212 3200 28218
rect 3148 28154 3200 28160
rect 3332 26784 3384 26790
rect 3332 26726 3384 26732
rect 3056 26512 3108 26518
rect 3056 26454 3108 26460
rect 3344 26314 3372 26726
rect 3332 26308 3384 26314
rect 3332 26250 3384 26256
rect 2884 24772 3004 24800
rect 2688 24744 2740 24750
rect 2688 24686 2740 24692
rect 2778 21584 2834 21593
rect 2778 21519 2834 21528
rect 2792 17338 2820 21519
rect 2884 19360 2912 24772
rect 3238 24712 3294 24721
rect 2964 24676 3016 24682
rect 3238 24647 3294 24656
rect 2964 24618 3016 24624
rect 2976 19961 3004 24618
rect 3146 21584 3202 21593
rect 3146 21519 3202 21528
rect 3160 21078 3188 21519
rect 3148 21072 3200 21078
rect 3148 21014 3200 21020
rect 2962 19952 3018 19961
rect 2962 19887 3018 19896
rect 2884 19332 3004 19360
rect 2780 17332 2832 17338
rect 2780 17274 2832 17280
rect 2318 10704 2374 10713
rect 2318 10639 2374 10648
rect 1412 6582 2268 6610
rect 478 6216 534 6225
rect 478 6151 534 6160
rect 492 800 520 6151
rect 1412 800 1440 6582
rect 2332 800 2360 10639
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2792 800 2820 4082
rect 2976 921 3004 19332
rect 3252 18465 3280 24647
rect 3344 18630 3372 26250
rect 3332 18624 3384 18630
rect 3332 18566 3384 18572
rect 3238 18456 3294 18465
rect 3344 18426 3372 18566
rect 3238 18391 3294 18400
rect 3332 18420 3384 18426
rect 3332 18362 3384 18368
rect 3424 16448 3476 16454
rect 3424 16390 3476 16396
rect 3436 16046 3464 16390
rect 3424 16040 3476 16046
rect 3424 15982 3476 15988
rect 3436 15706 3464 15982
rect 3424 15700 3476 15706
rect 3424 15642 3476 15648
rect 3054 13424 3110 13433
rect 3054 13359 3110 13368
rect 3068 9110 3096 13359
rect 3330 13288 3386 13297
rect 3330 13223 3386 13232
rect 3056 9104 3108 9110
rect 3056 9046 3108 9052
rect 3344 8945 3372 13223
rect 3528 10305 3556 48583
rect 3606 48240 3662 48249
rect 3606 48175 3662 48184
rect 3620 30705 3648 48175
rect 3712 36242 3740 48991
rect 3804 48113 3832 63271
rect 5460 60761 5488 74734
rect 5538 74695 5594 74704
rect 5540 74656 5592 74662
rect 5540 74598 5592 74604
rect 5552 71097 5580 74598
rect 5538 71088 5594 71097
rect 5538 71023 5594 71032
rect 5644 69873 5672 74831
rect 6472 74662 6500 79200
rect 6932 75313 6960 79200
rect 6918 75304 6974 75313
rect 6918 75239 6974 75248
rect 7470 74760 7526 74769
rect 7470 74695 7526 74704
rect 6460 74656 6512 74662
rect 6460 74598 6512 74604
rect 6920 74656 6972 74662
rect 6920 74598 6972 74604
rect 5956 74012 6252 74032
rect 6012 74010 6036 74012
rect 6092 74010 6116 74012
rect 6172 74010 6196 74012
rect 6034 73958 6036 74010
rect 6098 73958 6110 74010
rect 6172 73958 6174 74010
rect 6012 73956 6036 73958
rect 6092 73956 6116 73958
rect 6172 73956 6196 73958
rect 5956 73936 6252 73956
rect 6932 73817 6960 74598
rect 6918 73808 6974 73817
rect 6918 73743 6974 73752
rect 5956 72924 6252 72944
rect 6012 72922 6036 72924
rect 6092 72922 6116 72924
rect 6172 72922 6196 72924
rect 6034 72870 6036 72922
rect 6098 72870 6110 72922
rect 6172 72870 6174 72922
rect 6012 72868 6036 72870
rect 6092 72868 6116 72870
rect 6172 72868 6196 72870
rect 5956 72848 6252 72868
rect 7286 72584 7342 72593
rect 7286 72519 7342 72528
rect 5956 71836 6252 71856
rect 6012 71834 6036 71836
rect 6092 71834 6116 71836
rect 6172 71834 6196 71836
rect 6034 71782 6036 71834
rect 6098 71782 6110 71834
rect 6172 71782 6174 71834
rect 6012 71780 6036 71782
rect 6092 71780 6116 71782
rect 6172 71780 6196 71782
rect 5956 71760 6252 71780
rect 5956 70748 6252 70768
rect 6012 70746 6036 70748
rect 6092 70746 6116 70748
rect 6172 70746 6196 70748
rect 6034 70694 6036 70746
rect 6098 70694 6110 70746
rect 6172 70694 6174 70746
rect 6012 70692 6036 70694
rect 6092 70692 6116 70694
rect 6172 70692 6196 70694
rect 5956 70672 6252 70692
rect 5630 69864 5686 69873
rect 5630 69799 5686 69808
rect 5956 69660 6252 69680
rect 6012 69658 6036 69660
rect 6092 69658 6116 69660
rect 6172 69658 6196 69660
rect 6034 69606 6036 69658
rect 6098 69606 6110 69658
rect 6172 69606 6174 69658
rect 6012 69604 6036 69606
rect 6092 69604 6116 69606
rect 6172 69604 6196 69606
rect 5956 69584 6252 69604
rect 5956 68572 6252 68592
rect 6012 68570 6036 68572
rect 6092 68570 6116 68572
rect 6172 68570 6196 68572
rect 6034 68518 6036 68570
rect 6098 68518 6110 68570
rect 6172 68518 6174 68570
rect 6012 68516 6036 68518
rect 6092 68516 6116 68518
rect 6172 68516 6196 68518
rect 5956 68496 6252 68516
rect 5956 67484 6252 67504
rect 6012 67482 6036 67484
rect 6092 67482 6116 67484
rect 6172 67482 6196 67484
rect 6034 67430 6036 67482
rect 6098 67430 6110 67482
rect 6172 67430 6174 67482
rect 6012 67428 6036 67430
rect 6092 67428 6116 67430
rect 6172 67428 6196 67430
rect 5956 67408 6252 67428
rect 5956 66396 6252 66416
rect 6012 66394 6036 66396
rect 6092 66394 6116 66396
rect 6172 66394 6196 66396
rect 6034 66342 6036 66394
rect 6098 66342 6110 66394
rect 6172 66342 6174 66394
rect 6012 66340 6036 66342
rect 6092 66340 6116 66342
rect 6172 66340 6196 66342
rect 5956 66320 6252 66340
rect 5956 65308 6252 65328
rect 6012 65306 6036 65308
rect 6092 65306 6116 65308
rect 6172 65306 6196 65308
rect 6034 65254 6036 65306
rect 6098 65254 6110 65306
rect 6172 65254 6174 65306
rect 6012 65252 6036 65254
rect 6092 65252 6116 65254
rect 6172 65252 6196 65254
rect 5956 65232 6252 65252
rect 5956 64220 6252 64240
rect 6012 64218 6036 64220
rect 6092 64218 6116 64220
rect 6172 64218 6196 64220
rect 6034 64166 6036 64218
rect 6098 64166 6110 64218
rect 6172 64166 6174 64218
rect 6012 64164 6036 64166
rect 6092 64164 6116 64166
rect 6172 64164 6196 64166
rect 5956 64144 6252 64164
rect 5956 63132 6252 63152
rect 6012 63130 6036 63132
rect 6092 63130 6116 63132
rect 6172 63130 6196 63132
rect 6034 63078 6036 63130
rect 6098 63078 6110 63130
rect 6172 63078 6174 63130
rect 6012 63076 6036 63078
rect 6092 63076 6116 63078
rect 6172 63076 6196 63078
rect 5956 63056 6252 63076
rect 5956 62044 6252 62064
rect 6012 62042 6036 62044
rect 6092 62042 6116 62044
rect 6172 62042 6196 62044
rect 6034 61990 6036 62042
rect 6098 61990 6110 62042
rect 6172 61990 6174 62042
rect 6012 61988 6036 61990
rect 6092 61988 6116 61990
rect 6172 61988 6196 61990
rect 5956 61968 6252 61988
rect 5956 60956 6252 60976
rect 6012 60954 6036 60956
rect 6092 60954 6116 60956
rect 6172 60954 6196 60956
rect 6034 60902 6036 60954
rect 6098 60902 6110 60954
rect 6172 60902 6174 60954
rect 6012 60900 6036 60902
rect 6092 60900 6116 60902
rect 6172 60900 6196 60902
rect 5956 60880 6252 60900
rect 5446 60752 5502 60761
rect 5446 60687 5502 60696
rect 5956 59868 6252 59888
rect 6012 59866 6036 59868
rect 6092 59866 6116 59868
rect 6172 59866 6196 59868
rect 6034 59814 6036 59866
rect 6098 59814 6110 59866
rect 6172 59814 6174 59866
rect 6012 59812 6036 59814
rect 6092 59812 6116 59814
rect 6172 59812 6196 59814
rect 5956 59792 6252 59812
rect 5956 58780 6252 58800
rect 6012 58778 6036 58780
rect 6092 58778 6116 58780
rect 6172 58778 6196 58780
rect 6034 58726 6036 58778
rect 6098 58726 6110 58778
rect 6172 58726 6174 58778
rect 6012 58724 6036 58726
rect 6092 58724 6116 58726
rect 6172 58724 6196 58726
rect 5956 58704 6252 58724
rect 5448 58404 5500 58410
rect 5448 58346 5500 58352
rect 5460 57610 5488 58346
rect 7010 57896 7066 57905
rect 7010 57831 7066 57840
rect 5956 57692 6252 57712
rect 6012 57690 6036 57692
rect 6092 57690 6116 57692
rect 6172 57690 6196 57692
rect 6034 57638 6036 57690
rect 6098 57638 6110 57690
rect 6172 57638 6174 57690
rect 6012 57636 6036 57638
rect 6092 57636 6116 57638
rect 6172 57636 6196 57638
rect 5956 57616 6252 57636
rect 5460 57594 5580 57610
rect 5460 57588 5592 57594
rect 5460 57582 5540 57588
rect 5540 57530 5592 57536
rect 7024 57390 7052 57831
rect 7012 57384 7064 57390
rect 7012 57326 7064 57332
rect 7024 57050 7052 57326
rect 7012 57044 7064 57050
rect 7012 56986 7064 56992
rect 5956 56604 6252 56624
rect 6012 56602 6036 56604
rect 6092 56602 6116 56604
rect 6172 56602 6196 56604
rect 6034 56550 6036 56602
rect 6098 56550 6110 56602
rect 6172 56550 6174 56602
rect 6012 56548 6036 56550
rect 6092 56548 6116 56550
rect 6172 56548 6196 56550
rect 5956 56528 6252 56548
rect 5956 55516 6252 55536
rect 6012 55514 6036 55516
rect 6092 55514 6116 55516
rect 6172 55514 6196 55516
rect 6034 55462 6036 55514
rect 6098 55462 6110 55514
rect 6172 55462 6174 55514
rect 6012 55460 6036 55462
rect 6092 55460 6116 55462
rect 6172 55460 6196 55462
rect 5956 55440 6252 55460
rect 5956 54428 6252 54448
rect 6012 54426 6036 54428
rect 6092 54426 6116 54428
rect 6172 54426 6196 54428
rect 6034 54374 6036 54426
rect 6098 54374 6110 54426
rect 6172 54374 6174 54426
rect 6012 54372 6036 54374
rect 6092 54372 6116 54374
rect 6172 54372 6196 54374
rect 5956 54352 6252 54372
rect 5956 53340 6252 53360
rect 6012 53338 6036 53340
rect 6092 53338 6116 53340
rect 6172 53338 6196 53340
rect 6034 53286 6036 53338
rect 6098 53286 6110 53338
rect 6172 53286 6174 53338
rect 6012 53284 6036 53286
rect 6092 53284 6116 53286
rect 6172 53284 6196 53286
rect 5956 53264 6252 53284
rect 4066 52592 4122 52601
rect 4066 52527 4068 52536
rect 4120 52527 4122 52536
rect 4068 52498 4120 52504
rect 5956 52252 6252 52272
rect 6012 52250 6036 52252
rect 6092 52250 6116 52252
rect 6172 52250 6196 52252
rect 6034 52198 6036 52250
rect 6098 52198 6110 52250
rect 6172 52198 6174 52250
rect 6012 52196 6036 52198
rect 6092 52196 6116 52198
rect 6172 52196 6196 52198
rect 5956 52176 6252 52196
rect 6276 51468 6328 51474
rect 6276 51410 6328 51416
rect 6288 51377 6316 51410
rect 6274 51368 6330 51377
rect 6274 51303 6330 51312
rect 5816 51264 5868 51270
rect 5816 51206 5868 51212
rect 5828 50969 5856 51206
rect 5956 51164 6252 51184
rect 6012 51162 6036 51164
rect 6092 51162 6116 51164
rect 6172 51162 6196 51164
rect 6034 51110 6036 51162
rect 6098 51110 6110 51162
rect 6172 51110 6174 51162
rect 6012 51108 6036 51110
rect 6092 51108 6116 51110
rect 6172 51108 6196 51110
rect 5956 51088 6252 51108
rect 6288 51066 6316 51303
rect 6276 51060 6328 51066
rect 6276 51002 6328 51008
rect 5814 50960 5870 50969
rect 5814 50895 5870 50904
rect 4066 50416 4122 50425
rect 4066 50351 4122 50360
rect 4080 49745 4108 50351
rect 5956 50076 6252 50096
rect 6012 50074 6036 50076
rect 6092 50074 6116 50076
rect 6172 50074 6196 50076
rect 6034 50022 6036 50074
rect 6098 50022 6110 50074
rect 6172 50022 6174 50074
rect 6012 50020 6036 50022
rect 6092 50020 6116 50022
rect 6172 50020 6196 50022
rect 5956 50000 6252 50020
rect 4066 49736 4122 49745
rect 4066 49671 4122 49680
rect 7196 49632 7248 49638
rect 7196 49574 7248 49580
rect 5956 48988 6252 49008
rect 6012 48986 6036 48988
rect 6092 48986 6116 48988
rect 6172 48986 6196 48988
rect 6034 48934 6036 48986
rect 6098 48934 6110 48986
rect 6172 48934 6174 48986
rect 6012 48932 6036 48934
rect 6092 48932 6116 48934
rect 6172 48932 6196 48934
rect 5956 48912 6252 48932
rect 4066 48376 4122 48385
rect 4066 48311 4122 48320
rect 3790 48104 3846 48113
rect 3790 48039 3846 48048
rect 4080 46481 4108 48311
rect 7208 48249 7236 49574
rect 7194 48240 7250 48249
rect 7194 48175 7250 48184
rect 5956 47900 6252 47920
rect 6012 47898 6036 47900
rect 6092 47898 6116 47900
rect 6172 47898 6196 47900
rect 6034 47846 6036 47898
rect 6098 47846 6110 47898
rect 6172 47846 6174 47898
rect 6012 47844 6036 47846
rect 6092 47844 6116 47846
rect 6172 47844 6196 47846
rect 5956 47824 6252 47844
rect 5956 46812 6252 46832
rect 6012 46810 6036 46812
rect 6092 46810 6116 46812
rect 6172 46810 6196 46812
rect 6034 46758 6036 46810
rect 6098 46758 6110 46810
rect 6172 46758 6174 46810
rect 6012 46756 6036 46758
rect 6092 46756 6116 46758
rect 6172 46756 6196 46758
rect 5956 46736 6252 46756
rect 4066 46472 4122 46481
rect 4066 46407 4122 46416
rect 6274 45928 6330 45937
rect 6274 45863 6330 45872
rect 5956 45724 6252 45744
rect 6012 45722 6036 45724
rect 6092 45722 6116 45724
rect 6172 45722 6196 45724
rect 6034 45670 6036 45722
rect 6098 45670 6110 45722
rect 6172 45670 6174 45722
rect 6012 45668 6036 45670
rect 6092 45668 6116 45670
rect 6172 45668 6196 45670
rect 5956 45648 6252 45668
rect 4068 45348 4120 45354
rect 4068 45290 4120 45296
rect 4080 43897 4108 45290
rect 5956 44636 6252 44656
rect 6012 44634 6036 44636
rect 6092 44634 6116 44636
rect 6172 44634 6196 44636
rect 6034 44582 6036 44634
rect 6098 44582 6110 44634
rect 6172 44582 6174 44634
rect 6012 44580 6036 44582
rect 6092 44580 6116 44582
rect 6172 44580 6196 44582
rect 5956 44560 6252 44580
rect 4066 43888 4122 43897
rect 4066 43823 4122 43832
rect 5956 43548 6252 43568
rect 6012 43546 6036 43548
rect 6092 43546 6116 43548
rect 6172 43546 6196 43548
rect 6034 43494 6036 43546
rect 6098 43494 6110 43546
rect 6172 43494 6174 43546
rect 6012 43492 6036 43494
rect 6092 43492 6116 43494
rect 6172 43492 6196 43494
rect 5956 43472 6252 43492
rect 5956 42460 6252 42480
rect 6012 42458 6036 42460
rect 6092 42458 6116 42460
rect 6172 42458 6196 42460
rect 6034 42406 6036 42458
rect 6098 42406 6110 42458
rect 6172 42406 6174 42458
rect 6012 42404 6036 42406
rect 6092 42404 6116 42406
rect 6172 42404 6196 42406
rect 5956 42384 6252 42404
rect 5956 41372 6252 41392
rect 6012 41370 6036 41372
rect 6092 41370 6116 41372
rect 6172 41370 6196 41372
rect 6034 41318 6036 41370
rect 6098 41318 6110 41370
rect 6172 41318 6174 41370
rect 6012 41316 6036 41318
rect 6092 41316 6116 41318
rect 6172 41316 6196 41318
rect 5956 41296 6252 41316
rect 5956 40284 6252 40304
rect 6012 40282 6036 40284
rect 6092 40282 6116 40284
rect 6172 40282 6196 40284
rect 6034 40230 6036 40282
rect 6098 40230 6110 40282
rect 6172 40230 6174 40282
rect 6012 40228 6036 40230
rect 6092 40228 6116 40230
rect 6172 40228 6196 40230
rect 5956 40208 6252 40228
rect 5956 39196 6252 39216
rect 6012 39194 6036 39196
rect 6092 39194 6116 39196
rect 6172 39194 6196 39196
rect 6034 39142 6036 39194
rect 6098 39142 6110 39194
rect 6172 39142 6174 39194
rect 6012 39140 6036 39142
rect 6092 39140 6116 39142
rect 6172 39140 6196 39142
rect 5956 39120 6252 39140
rect 5956 38108 6252 38128
rect 6012 38106 6036 38108
rect 6092 38106 6116 38108
rect 6172 38106 6196 38108
rect 6034 38054 6036 38106
rect 6098 38054 6110 38106
rect 6172 38054 6174 38106
rect 6012 38052 6036 38054
rect 6092 38052 6116 38054
rect 6172 38052 6196 38054
rect 5956 38032 6252 38052
rect 4896 37732 4948 37738
rect 4896 37674 4948 37680
rect 4618 36408 4674 36417
rect 4618 36343 4674 36352
rect 3700 36236 3752 36242
rect 3700 36178 3752 36184
rect 4160 36168 4212 36174
rect 4160 36110 4212 36116
rect 4172 35766 4200 36110
rect 4632 35834 4660 36343
rect 4908 35834 4936 37674
rect 5078 37224 5134 37233
rect 5078 37159 5134 37168
rect 4620 35828 4672 35834
rect 4620 35770 4672 35776
rect 4896 35828 4948 35834
rect 4896 35770 4948 35776
rect 4160 35760 4212 35766
rect 4160 35702 4212 35708
rect 4528 35556 4580 35562
rect 4528 35498 4580 35504
rect 4540 34746 4568 35498
rect 4618 35320 4674 35329
rect 4618 35255 4620 35264
rect 4672 35255 4674 35264
rect 4620 35226 4672 35232
rect 5092 35154 5120 37159
rect 5956 37020 6252 37040
rect 6012 37018 6036 37020
rect 6092 37018 6116 37020
rect 6172 37018 6196 37020
rect 6034 36966 6036 37018
rect 6098 36966 6110 37018
rect 6172 36966 6174 37018
rect 6012 36964 6036 36966
rect 6092 36964 6116 36966
rect 6172 36964 6196 36966
rect 5956 36944 6252 36964
rect 5172 36236 5224 36242
rect 5172 36178 5224 36184
rect 5184 35834 5212 36178
rect 5446 36136 5502 36145
rect 5446 36071 5502 36080
rect 5356 36032 5408 36038
rect 5356 35974 5408 35980
rect 5172 35828 5224 35834
rect 5172 35770 5224 35776
rect 5080 35148 5132 35154
rect 5080 35090 5132 35096
rect 4988 34944 5040 34950
rect 4988 34886 5040 34892
rect 5000 34746 5028 34886
rect 4528 34740 4580 34746
rect 4528 34682 4580 34688
rect 4988 34740 5040 34746
rect 4988 34682 5040 34688
rect 5092 34678 5120 35090
rect 5368 35018 5396 35974
rect 5356 35012 5408 35018
rect 5356 34954 5408 34960
rect 5264 34944 5316 34950
rect 5264 34886 5316 34892
rect 5080 34672 5132 34678
rect 3882 34640 3938 34649
rect 5080 34614 5132 34620
rect 3882 34575 3884 34584
rect 3936 34575 3938 34584
rect 4988 34604 5040 34610
rect 3884 34546 3936 34552
rect 4988 34546 5040 34552
rect 3976 34536 4028 34542
rect 3976 34478 4028 34484
rect 4342 34504 4398 34513
rect 3792 33856 3844 33862
rect 3792 33798 3844 33804
rect 3804 32756 3832 33798
rect 3882 33416 3938 33425
rect 3882 33351 3884 33360
rect 3936 33351 3938 33360
rect 3884 33322 3936 33328
rect 3884 32768 3936 32774
rect 3804 32728 3884 32756
rect 3884 32710 3936 32716
rect 3896 32473 3924 32710
rect 3882 32464 3938 32473
rect 3882 32399 3938 32408
rect 3884 32224 3936 32230
rect 3884 32166 3936 32172
rect 3896 31958 3924 32166
rect 3884 31952 3936 31958
rect 3884 31894 3936 31900
rect 3988 31249 4016 34478
rect 4342 34439 4398 34448
rect 4620 34468 4672 34474
rect 4356 34202 4384 34439
rect 4620 34410 4672 34416
rect 4632 34202 4660 34410
rect 4344 34196 4396 34202
rect 4344 34138 4396 34144
rect 4620 34196 4672 34202
rect 4620 34138 4672 34144
rect 4342 34096 4398 34105
rect 4342 34031 4398 34040
rect 4436 34060 4488 34066
rect 4356 33454 4384 34031
rect 4436 34002 4488 34008
rect 4344 33448 4396 33454
rect 4344 33390 4396 33396
rect 4448 33386 4476 34002
rect 5000 33930 5028 34546
rect 5276 34542 5304 34886
rect 5368 34610 5396 34954
rect 5356 34604 5408 34610
rect 5356 34546 5408 34552
rect 5264 34536 5316 34542
rect 5264 34478 5316 34484
rect 5172 34400 5224 34406
rect 5172 34342 5224 34348
rect 4988 33924 5040 33930
rect 4988 33866 5040 33872
rect 4528 33856 4580 33862
rect 4528 33798 4580 33804
rect 4540 33658 4568 33798
rect 4528 33652 4580 33658
rect 4528 33594 4580 33600
rect 5000 33522 5028 33866
rect 4988 33516 5040 33522
rect 5040 33476 5120 33504
rect 4988 33458 5040 33464
rect 4436 33380 4488 33386
rect 4436 33322 4488 33328
rect 4988 33380 5040 33386
rect 4988 33322 5040 33328
rect 4618 33144 4674 33153
rect 4618 33079 4620 33088
rect 4672 33079 4674 33088
rect 4620 33050 4672 33056
rect 4894 32872 4950 32881
rect 4894 32807 4950 32816
rect 4908 32570 4936 32807
rect 4896 32564 4948 32570
rect 4896 32506 4948 32512
rect 3974 31240 4030 31249
rect 3974 31175 4030 31184
rect 4804 31136 4856 31142
rect 4804 31078 4856 31084
rect 4816 30802 4844 31078
rect 4804 30796 4856 30802
rect 4804 30738 4856 30744
rect 3606 30696 3662 30705
rect 3606 30631 3662 30640
rect 4620 30048 4672 30054
rect 4620 29990 4672 29996
rect 4632 29034 4660 29990
rect 5000 29753 5028 33322
rect 5092 32026 5120 33476
rect 5184 32978 5212 34342
rect 5276 34066 5304 34478
rect 5354 34232 5410 34241
rect 5460 34202 5488 36071
rect 5956 35932 6252 35952
rect 6012 35930 6036 35932
rect 6092 35930 6116 35932
rect 6172 35930 6196 35932
rect 6034 35878 6036 35930
rect 6098 35878 6110 35930
rect 6172 35878 6174 35930
rect 6012 35876 6036 35878
rect 6092 35876 6116 35878
rect 6172 35876 6196 35878
rect 5956 35856 6252 35876
rect 6184 35624 6236 35630
rect 6182 35592 6184 35601
rect 6236 35592 6238 35601
rect 6182 35527 6238 35536
rect 6000 35080 6052 35086
rect 5998 35048 6000 35057
rect 6052 35048 6054 35057
rect 5998 34983 6054 34992
rect 5956 34844 6252 34864
rect 6012 34842 6036 34844
rect 6092 34842 6116 34844
rect 6172 34842 6196 34844
rect 6034 34790 6036 34842
rect 6098 34790 6110 34842
rect 6172 34790 6174 34842
rect 6012 34788 6036 34790
rect 6092 34788 6116 34790
rect 6172 34788 6196 34790
rect 5956 34768 6252 34788
rect 5906 34640 5962 34649
rect 5906 34575 5908 34584
rect 5960 34575 5962 34584
rect 5908 34546 5960 34552
rect 5354 34167 5410 34176
rect 5448 34196 5500 34202
rect 5368 34134 5396 34167
rect 5448 34138 5500 34144
rect 5356 34128 5408 34134
rect 5356 34070 5408 34076
rect 5540 34128 5592 34134
rect 5540 34070 5592 34076
rect 5816 34128 5868 34134
rect 5816 34070 5868 34076
rect 5264 34060 5316 34066
rect 5264 34002 5316 34008
rect 5264 33584 5316 33590
rect 5264 33526 5316 33532
rect 5354 33552 5410 33561
rect 5172 32972 5224 32978
rect 5172 32914 5224 32920
rect 5184 32570 5212 32914
rect 5172 32564 5224 32570
rect 5172 32506 5224 32512
rect 5276 32502 5304 33526
rect 5354 33487 5356 33496
rect 5408 33487 5410 33496
rect 5356 33458 5408 33464
rect 5448 33448 5500 33454
rect 5448 33390 5500 33396
rect 5460 32774 5488 33390
rect 5552 33318 5580 34070
rect 5828 33590 5856 34070
rect 6184 33992 6236 33998
rect 6182 33960 6184 33969
rect 6236 33960 6238 33969
rect 6182 33895 6238 33904
rect 5956 33756 6252 33776
rect 6012 33754 6036 33756
rect 6092 33754 6116 33756
rect 6172 33754 6196 33756
rect 6034 33702 6036 33754
rect 6098 33702 6110 33754
rect 6172 33702 6174 33754
rect 6012 33700 6036 33702
rect 6092 33700 6116 33702
rect 6172 33700 6196 33702
rect 5956 33680 6252 33700
rect 5816 33584 5868 33590
rect 5816 33526 5868 33532
rect 5908 33380 5960 33386
rect 5908 33322 5960 33328
rect 5540 33312 5592 33318
rect 5540 33254 5592 33260
rect 5448 32768 5500 32774
rect 5448 32710 5500 32716
rect 5264 32496 5316 32502
rect 5264 32438 5316 32444
rect 5460 32230 5488 32710
rect 5448 32224 5500 32230
rect 5448 32166 5500 32172
rect 5262 32056 5318 32065
rect 5080 32020 5132 32026
rect 5080 31962 5132 31968
rect 5184 32000 5262 32008
rect 5184 31980 5264 32000
rect 5184 30172 5212 31980
rect 5316 31991 5318 32000
rect 5264 31962 5316 31968
rect 5552 31498 5580 33254
rect 5920 33017 5948 33322
rect 5722 33008 5778 33017
rect 5906 33008 5962 33017
rect 5778 32966 5856 32994
rect 5722 32943 5778 32952
rect 5724 32904 5776 32910
rect 5724 32846 5776 32852
rect 5828 32892 5856 32966
rect 5906 32943 5962 32952
rect 5908 32904 5960 32910
rect 5828 32864 5908 32892
rect 5736 32450 5764 32846
rect 5828 32570 5856 32864
rect 5908 32846 5960 32852
rect 5956 32668 6252 32688
rect 6012 32666 6036 32668
rect 6092 32666 6116 32668
rect 6172 32666 6196 32668
rect 6034 32614 6036 32666
rect 6098 32614 6110 32666
rect 6172 32614 6174 32666
rect 6012 32612 6036 32614
rect 6092 32612 6116 32614
rect 6172 32612 6196 32614
rect 5956 32592 6252 32612
rect 5816 32564 5868 32570
rect 5816 32506 5868 32512
rect 5736 32422 5856 32450
rect 5630 32328 5686 32337
rect 5630 32263 5632 32272
rect 5684 32263 5686 32272
rect 5632 32234 5684 32240
rect 5724 31952 5776 31958
rect 5722 31920 5724 31929
rect 5776 31920 5778 31929
rect 5722 31855 5778 31864
rect 5724 31816 5776 31822
rect 5828 31804 5856 32422
rect 5908 32224 5960 32230
rect 5906 32192 5908 32201
rect 5960 32192 5962 32201
rect 5906 32127 5962 32136
rect 5908 31884 5960 31890
rect 5908 31826 5960 31832
rect 5776 31776 5856 31804
rect 5724 31758 5776 31764
rect 5552 31470 5672 31498
rect 5540 31408 5592 31414
rect 5538 31376 5540 31385
rect 5592 31376 5594 31385
rect 5538 31311 5594 31320
rect 5448 31136 5500 31142
rect 5448 31078 5500 31084
rect 5262 30696 5318 30705
rect 5262 30631 5318 30640
rect 5276 30326 5304 30631
rect 5264 30320 5316 30326
rect 5264 30262 5316 30268
rect 5184 30144 5304 30172
rect 4986 29744 5042 29753
rect 4986 29679 5042 29688
rect 4620 29028 4672 29034
rect 4620 28970 4672 28976
rect 4068 28416 4120 28422
rect 4068 28358 4120 28364
rect 4080 27713 4108 28358
rect 4066 27704 4122 27713
rect 4066 27639 4122 27648
rect 4632 27606 4660 28970
rect 4710 28656 4766 28665
rect 4710 28591 4766 28600
rect 4620 27600 4672 27606
rect 4620 27542 4672 27548
rect 4158 27296 4214 27305
rect 4158 27231 4214 27240
rect 4172 25838 4200 27231
rect 4632 26450 4660 27542
rect 4724 26926 4752 28591
rect 5080 27464 5132 27470
rect 5276 27452 5304 30144
rect 5460 29034 5488 31078
rect 5644 30666 5672 31470
rect 5736 30802 5764 31758
rect 5920 31736 5948 31826
rect 5828 31708 5948 31736
rect 5828 31142 5856 31708
rect 5956 31580 6252 31600
rect 6012 31578 6036 31580
rect 6092 31578 6116 31580
rect 6172 31578 6196 31580
rect 6034 31526 6036 31578
rect 6098 31526 6110 31578
rect 6172 31526 6174 31578
rect 6012 31524 6036 31526
rect 6092 31524 6116 31526
rect 6172 31524 6196 31526
rect 5956 31504 6252 31524
rect 5816 31136 5868 31142
rect 5816 31078 5868 31084
rect 5724 30796 5776 30802
rect 5724 30738 5776 30744
rect 5632 30660 5684 30666
rect 5632 30602 5684 30608
rect 5540 30592 5592 30598
rect 5540 30534 5592 30540
rect 5630 30560 5686 30569
rect 5552 30190 5580 30534
rect 5630 30495 5686 30504
rect 5644 30258 5672 30495
rect 5632 30252 5684 30258
rect 5632 30194 5684 30200
rect 5540 30184 5592 30190
rect 5540 30126 5592 30132
rect 5448 29028 5500 29034
rect 5448 28970 5500 28976
rect 5552 28762 5580 30126
rect 5828 30025 5856 31078
rect 5956 30492 6252 30512
rect 6012 30490 6036 30492
rect 6092 30490 6116 30492
rect 6172 30490 6196 30492
rect 6034 30438 6036 30490
rect 6098 30438 6110 30490
rect 6172 30438 6174 30490
rect 6012 30436 6036 30438
rect 6092 30436 6116 30438
rect 6172 30436 6196 30438
rect 5956 30416 6252 30436
rect 5814 30016 5870 30025
rect 5814 29951 5870 29960
rect 5956 29404 6252 29424
rect 6012 29402 6036 29404
rect 6092 29402 6116 29404
rect 6172 29402 6196 29404
rect 6034 29350 6036 29402
rect 6098 29350 6110 29402
rect 6172 29350 6174 29402
rect 6012 29348 6036 29350
rect 6092 29348 6116 29350
rect 6172 29348 6196 29350
rect 5956 29328 6252 29348
rect 6182 29200 6238 29209
rect 6182 29135 6238 29144
rect 6196 29102 6224 29135
rect 6184 29096 6236 29102
rect 6184 29038 6236 29044
rect 5816 29028 5868 29034
rect 5816 28970 5868 28976
rect 5540 28756 5592 28762
rect 5540 28698 5592 28704
rect 5724 28620 5776 28626
rect 5724 28562 5776 28568
rect 5736 27946 5764 28562
rect 5724 27940 5776 27946
rect 5724 27882 5776 27888
rect 5132 27424 5304 27452
rect 5080 27406 5132 27412
rect 5092 26926 5120 27406
rect 5724 27328 5776 27334
rect 5724 27270 5776 27276
rect 5736 26926 5764 27270
rect 4712 26920 4764 26926
rect 4712 26862 4764 26868
rect 5080 26920 5132 26926
rect 5080 26862 5132 26868
rect 5356 26920 5408 26926
rect 5356 26862 5408 26868
rect 5724 26920 5776 26926
rect 5724 26862 5776 26868
rect 4620 26444 4672 26450
rect 4620 26386 4672 26392
rect 5092 26314 5120 26862
rect 5172 26376 5224 26382
rect 5172 26318 5224 26324
rect 5080 26308 5132 26314
rect 5080 26250 5132 26256
rect 5184 25838 5212 26318
rect 5264 26240 5316 26246
rect 5368 26228 5396 26862
rect 5632 26444 5684 26450
rect 5632 26386 5684 26392
rect 5316 26200 5396 26228
rect 5264 26182 5316 26188
rect 5368 25838 5396 26200
rect 4160 25832 4212 25838
rect 4160 25774 4212 25780
rect 5172 25832 5224 25838
rect 5172 25774 5224 25780
rect 5356 25832 5408 25838
rect 5356 25774 5408 25780
rect 5184 25226 5212 25774
rect 5172 25220 5224 25226
rect 5172 25162 5224 25168
rect 5184 17678 5212 25162
rect 5368 25158 5396 25774
rect 5644 25498 5672 26386
rect 5724 26240 5776 26246
rect 5724 26182 5776 26188
rect 5736 25838 5764 26182
rect 5724 25832 5776 25838
rect 5724 25774 5776 25780
rect 5828 25673 5856 28970
rect 6196 28762 6224 29038
rect 6184 28756 6236 28762
rect 6184 28698 6236 28704
rect 5956 28316 6252 28336
rect 6012 28314 6036 28316
rect 6092 28314 6116 28316
rect 6172 28314 6196 28316
rect 6034 28262 6036 28314
rect 6098 28262 6110 28314
rect 6172 28262 6174 28314
rect 6012 28260 6036 28262
rect 6092 28260 6116 28262
rect 6172 28260 6196 28262
rect 5956 28240 6252 28260
rect 5956 27228 6252 27248
rect 6012 27226 6036 27228
rect 6092 27226 6116 27228
rect 6172 27226 6196 27228
rect 6034 27174 6036 27226
rect 6098 27174 6110 27226
rect 6172 27174 6174 27226
rect 6012 27172 6036 27174
rect 6092 27172 6116 27174
rect 6172 27172 6196 27174
rect 5956 27152 6252 27172
rect 5956 26140 6252 26160
rect 6012 26138 6036 26140
rect 6092 26138 6116 26140
rect 6172 26138 6196 26140
rect 6034 26086 6036 26138
rect 6098 26086 6110 26138
rect 6172 26086 6174 26138
rect 6012 26084 6036 26086
rect 6092 26084 6116 26086
rect 6172 26084 6196 26086
rect 5956 26064 6252 26084
rect 5814 25664 5870 25673
rect 5814 25599 5870 25608
rect 5632 25492 5684 25498
rect 5632 25434 5684 25440
rect 5356 25152 5408 25158
rect 5356 25094 5408 25100
rect 5956 25052 6252 25072
rect 6012 25050 6036 25052
rect 6092 25050 6116 25052
rect 6172 25050 6196 25052
rect 6034 24998 6036 25050
rect 6098 24998 6110 25050
rect 6172 24998 6174 25050
rect 6012 24996 6036 24998
rect 6092 24996 6116 24998
rect 6172 24996 6196 24998
rect 5956 24976 6252 24996
rect 6288 24721 6316 45863
rect 6734 44840 6790 44849
rect 6734 44775 6790 44784
rect 6552 37256 6604 37262
rect 6552 37198 6604 37204
rect 6368 37120 6420 37126
rect 6368 37062 6420 37068
rect 6380 36718 6408 37062
rect 6564 36854 6592 37198
rect 6552 36848 6604 36854
rect 6550 36816 6552 36825
rect 6604 36816 6606 36825
rect 6550 36751 6606 36760
rect 6368 36712 6420 36718
rect 6368 36654 6420 36660
rect 6460 36644 6512 36650
rect 6460 36586 6512 36592
rect 6368 34944 6420 34950
rect 6368 34886 6420 34892
rect 6380 34542 6408 34886
rect 6368 34536 6420 34542
rect 6368 34478 6420 34484
rect 6380 34202 6408 34478
rect 6472 34388 6500 36586
rect 6644 36576 6696 36582
rect 6644 36518 6696 36524
rect 6656 35698 6684 36518
rect 6644 35692 6696 35698
rect 6644 35634 6696 35640
rect 6642 35184 6698 35193
rect 6642 35119 6644 35128
rect 6696 35119 6698 35128
rect 6644 35090 6696 35096
rect 6552 34944 6604 34950
rect 6552 34886 6604 34892
rect 6564 34610 6592 34886
rect 6656 34678 6684 35090
rect 6644 34672 6696 34678
rect 6644 34614 6696 34620
rect 6552 34604 6604 34610
rect 6552 34546 6604 34552
rect 6552 34400 6604 34406
rect 6472 34360 6552 34388
rect 6552 34342 6604 34348
rect 6368 34196 6420 34202
rect 6368 34138 6420 34144
rect 6380 33658 6408 34138
rect 6458 34096 6514 34105
rect 6458 34031 6514 34040
rect 6472 33833 6500 34031
rect 6458 33824 6514 33833
rect 6458 33759 6514 33768
rect 6368 33652 6420 33658
rect 6368 33594 6420 33600
rect 6564 33538 6592 34342
rect 6644 34060 6696 34066
rect 6644 34002 6696 34008
rect 6656 33697 6684 34002
rect 6642 33688 6698 33697
rect 6642 33623 6644 33632
rect 6696 33623 6698 33632
rect 6644 33594 6696 33600
rect 6564 33510 6684 33538
rect 6550 33280 6606 33289
rect 6550 33215 6606 33224
rect 6564 32473 6592 33215
rect 6550 32464 6606 32473
rect 6550 32399 6606 32408
rect 6460 32224 6512 32230
rect 6460 32166 6512 32172
rect 6366 31648 6422 31657
rect 6366 31583 6422 31592
rect 6380 30938 6408 31583
rect 6368 30932 6420 30938
rect 6368 30874 6420 30880
rect 6368 30592 6420 30598
rect 6368 30534 6420 30540
rect 6380 27169 6408 30534
rect 6472 28665 6500 32166
rect 6564 29850 6592 32399
rect 6656 31793 6684 33510
rect 6642 31784 6698 31793
rect 6642 31719 6698 31728
rect 6642 31512 6698 31521
rect 6642 31447 6644 31456
rect 6696 31447 6698 31456
rect 6644 31418 6696 31424
rect 6644 30796 6696 30802
rect 6644 30738 6696 30744
rect 6656 30054 6684 30738
rect 6644 30048 6696 30054
rect 6644 29990 6696 29996
rect 6552 29844 6604 29850
rect 6552 29786 6604 29792
rect 6642 29608 6698 29617
rect 6642 29543 6698 29552
rect 6552 29504 6604 29510
rect 6552 29446 6604 29452
rect 6564 28801 6592 29446
rect 6656 29306 6684 29543
rect 6644 29300 6696 29306
rect 6644 29242 6696 29248
rect 6550 28792 6606 28801
rect 6550 28727 6552 28736
rect 6604 28727 6606 28736
rect 6552 28698 6604 28704
rect 6458 28656 6514 28665
rect 6458 28591 6514 28600
rect 6460 27940 6512 27946
rect 6460 27882 6512 27888
rect 6366 27160 6422 27169
rect 6366 27095 6422 27104
rect 6368 26920 6420 26926
rect 6368 26862 6420 26868
rect 6380 25838 6408 26862
rect 6368 25832 6420 25838
rect 6368 25774 6420 25780
rect 6274 24712 6330 24721
rect 6274 24647 6330 24656
rect 6380 24426 6408 25774
rect 6288 24398 6408 24426
rect 5956 23964 6252 23984
rect 6012 23962 6036 23964
rect 6092 23962 6116 23964
rect 6172 23962 6196 23964
rect 6034 23910 6036 23962
rect 6098 23910 6110 23962
rect 6172 23910 6174 23962
rect 6012 23908 6036 23910
rect 6092 23908 6116 23910
rect 6172 23908 6196 23910
rect 5956 23888 6252 23908
rect 5540 23112 5592 23118
rect 5540 23054 5592 23060
rect 5552 22137 5580 23054
rect 6288 23050 6316 24398
rect 6276 23044 6328 23050
rect 6276 22986 6328 22992
rect 5956 22876 6252 22896
rect 6012 22874 6036 22876
rect 6092 22874 6116 22876
rect 6172 22874 6196 22876
rect 6034 22822 6036 22874
rect 6098 22822 6110 22874
rect 6172 22822 6174 22874
rect 6012 22820 6036 22822
rect 6092 22820 6116 22822
rect 6172 22820 6196 22822
rect 5956 22800 6252 22820
rect 6288 22710 6316 22986
rect 6276 22704 6328 22710
rect 6276 22646 6328 22652
rect 5538 22128 5594 22137
rect 5538 22063 5594 22072
rect 6276 22024 6328 22030
rect 6276 21966 6328 21972
rect 6368 22024 6420 22030
rect 6368 21966 6420 21972
rect 5956 21788 6252 21808
rect 6012 21786 6036 21788
rect 6092 21786 6116 21788
rect 6172 21786 6196 21788
rect 6034 21734 6036 21786
rect 6098 21734 6110 21786
rect 6172 21734 6174 21786
rect 6012 21732 6036 21734
rect 6092 21732 6116 21734
rect 6172 21732 6196 21734
rect 5956 21712 6252 21732
rect 6288 21146 6316 21966
rect 6380 21622 6408 21966
rect 6472 21729 6500 27882
rect 6550 27704 6606 27713
rect 6550 27639 6606 27648
rect 6564 26081 6592 27639
rect 6644 26988 6696 26994
rect 6644 26930 6696 26936
rect 6550 26072 6606 26081
rect 6656 26042 6684 26930
rect 6550 26007 6606 26016
rect 6644 26036 6696 26042
rect 6644 25978 6696 25984
rect 6644 25152 6696 25158
rect 6644 25094 6696 25100
rect 6656 23186 6684 25094
rect 6644 23180 6696 23186
rect 6644 23122 6696 23128
rect 6656 22710 6684 23122
rect 6644 22704 6696 22710
rect 6644 22646 6696 22652
rect 6458 21720 6514 21729
rect 6458 21655 6514 21664
rect 6368 21616 6420 21622
rect 6366 21584 6368 21593
rect 6420 21584 6422 21593
rect 6366 21519 6422 21528
rect 6380 21493 6408 21519
rect 6656 21418 6684 22646
rect 6644 21412 6696 21418
rect 6644 21354 6696 21360
rect 6656 21146 6684 21354
rect 6276 21140 6328 21146
rect 6276 21082 6328 21088
rect 6644 21140 6696 21146
rect 6644 21082 6696 21088
rect 5956 20700 6252 20720
rect 6012 20698 6036 20700
rect 6092 20698 6116 20700
rect 6172 20698 6196 20700
rect 6034 20646 6036 20698
rect 6098 20646 6110 20698
rect 6172 20646 6174 20698
rect 6012 20644 6036 20646
rect 6092 20644 6116 20646
rect 6172 20644 6196 20646
rect 5956 20624 6252 20644
rect 5956 19612 6252 19632
rect 6012 19610 6036 19612
rect 6092 19610 6116 19612
rect 6172 19610 6196 19612
rect 6034 19558 6036 19610
rect 6098 19558 6110 19610
rect 6172 19558 6174 19610
rect 6012 19556 6036 19558
rect 6092 19556 6116 19558
rect 6172 19556 6196 19558
rect 5956 19536 6252 19556
rect 6644 19168 6696 19174
rect 6748 19145 6776 44775
rect 7012 37256 7064 37262
rect 7012 37198 7064 37204
rect 6826 36952 6882 36961
rect 6826 36887 6828 36896
rect 6880 36887 6882 36896
rect 6828 36858 6880 36864
rect 6920 36712 6972 36718
rect 7024 36700 7052 37198
rect 7104 36780 7156 36786
rect 7104 36722 7156 36728
rect 6972 36672 7052 36700
rect 6920 36654 6972 36660
rect 6920 35488 6972 35494
rect 6920 35430 6972 35436
rect 6828 34944 6880 34950
rect 6932 34921 6960 35430
rect 7024 35154 7052 36672
rect 7116 36378 7144 36722
rect 7104 36372 7156 36378
rect 7104 36314 7156 36320
rect 7196 35692 7248 35698
rect 7196 35634 7248 35640
rect 7104 35488 7156 35494
rect 7104 35430 7156 35436
rect 7012 35148 7064 35154
rect 7012 35090 7064 35096
rect 6828 34886 6880 34892
rect 6918 34912 6974 34921
rect 6840 34202 6868 34886
rect 6918 34847 6974 34856
rect 6920 34604 6972 34610
rect 6920 34546 6972 34552
rect 6828 34196 6880 34202
rect 6828 34138 6880 34144
rect 6828 34060 6880 34066
rect 6828 34002 6880 34008
rect 6840 33969 6868 34002
rect 6826 33960 6882 33969
rect 6826 33895 6882 33904
rect 6932 33862 6960 34546
rect 7024 33998 7052 35090
rect 7116 34474 7144 35430
rect 7104 34468 7156 34474
rect 7104 34410 7156 34416
rect 7102 34368 7158 34377
rect 7102 34303 7158 34312
rect 7012 33992 7064 33998
rect 7012 33934 7064 33940
rect 6920 33856 6972 33862
rect 6920 33798 6972 33804
rect 6920 33448 6972 33454
rect 6920 33390 6972 33396
rect 6932 33153 6960 33390
rect 6918 33144 6974 33153
rect 6918 33079 6974 33088
rect 7024 33046 7052 33934
rect 7116 33658 7144 34303
rect 7104 33652 7156 33658
rect 7104 33594 7156 33600
rect 7116 33561 7144 33594
rect 7102 33552 7158 33561
rect 7102 33487 7158 33496
rect 7208 33436 7236 35634
rect 7300 33522 7328 72519
rect 7378 50960 7434 50969
rect 7378 50895 7434 50904
rect 7392 49842 7420 50895
rect 7380 49836 7432 49842
rect 7380 49778 7432 49784
rect 7392 49434 7420 49778
rect 7380 49428 7432 49434
rect 7380 49370 7432 49376
rect 7378 47016 7434 47025
rect 7378 46951 7434 46960
rect 7288 33516 7340 33522
rect 7288 33458 7340 33464
rect 7116 33408 7236 33436
rect 7012 33040 7064 33046
rect 7012 32982 7064 32988
rect 7012 32836 7064 32842
rect 7012 32778 7064 32784
rect 6920 32768 6972 32774
rect 6920 32710 6972 32716
rect 6932 31414 6960 32710
rect 6920 31408 6972 31414
rect 6920 31350 6972 31356
rect 6828 30728 6880 30734
rect 6828 30670 6880 30676
rect 6840 30190 6868 30670
rect 6932 30433 6960 31350
rect 6918 30424 6974 30433
rect 6918 30359 6974 30368
rect 6828 30184 6880 30190
rect 6828 30126 6880 30132
rect 6840 29782 6868 30126
rect 6920 30048 6972 30054
rect 6920 29990 6972 29996
rect 6828 29776 6880 29782
rect 6828 29718 6880 29724
rect 6840 29345 6868 29718
rect 6932 29646 6960 29990
rect 6920 29640 6972 29646
rect 6920 29582 6972 29588
rect 6826 29336 6882 29345
rect 6826 29271 6882 29280
rect 6828 29096 6880 29102
rect 6828 29038 6880 29044
rect 6840 28082 6868 29038
rect 6828 28076 6880 28082
rect 6828 28018 6880 28024
rect 6840 27878 6868 28018
rect 6828 27872 6880 27878
rect 6828 27814 6880 27820
rect 6840 23882 6868 27814
rect 6932 26926 6960 29582
rect 6920 26920 6972 26926
rect 6920 26862 6972 26868
rect 6932 26586 6960 26862
rect 6920 26580 6972 26586
rect 6920 26522 6972 26528
rect 7024 26382 7052 32778
rect 7116 30138 7144 33408
rect 7288 33380 7340 33386
rect 7288 33322 7340 33328
rect 7196 31680 7248 31686
rect 7196 31622 7248 31628
rect 7208 31482 7236 31622
rect 7196 31476 7248 31482
rect 7196 31418 7248 31424
rect 7196 30932 7248 30938
rect 7196 30874 7248 30880
rect 7208 30258 7236 30874
rect 7196 30252 7248 30258
rect 7196 30194 7248 30200
rect 7116 30110 7236 30138
rect 7102 30016 7158 30025
rect 7102 29951 7158 29960
rect 7116 29714 7144 29951
rect 7104 29708 7156 29714
rect 7104 29650 7156 29656
rect 7116 29306 7144 29650
rect 7104 29300 7156 29306
rect 7104 29242 7156 29248
rect 7104 28008 7156 28014
rect 7102 27976 7104 27985
rect 7156 27976 7158 27985
rect 7102 27911 7158 27920
rect 7208 27554 7236 30110
rect 7300 28218 7328 33322
rect 7288 28212 7340 28218
rect 7288 28154 7340 28160
rect 7392 27674 7420 46951
rect 7484 30938 7512 74695
rect 7746 73672 7802 73681
rect 7746 73607 7802 73616
rect 7562 73128 7618 73137
rect 7562 73063 7618 73072
rect 7576 71126 7604 73063
rect 7760 71210 7788 73607
rect 7852 71346 7880 79200
rect 8772 76498 8800 79200
rect 9586 77072 9642 77081
rect 9586 77007 9642 77016
rect 8760 76492 8812 76498
rect 8760 76434 8812 76440
rect 9600 76401 9628 77007
rect 9586 76392 9642 76401
rect 9586 76327 9642 76336
rect 9692 74769 9720 79200
rect 9772 76492 9824 76498
rect 9772 76434 9824 76440
rect 9784 76090 9812 76434
rect 10048 76424 10100 76430
rect 10048 76366 10100 76372
rect 9772 76084 9824 76090
rect 9772 76026 9824 76032
rect 10060 75732 10088 76366
rect 10152 75857 10180 79200
rect 11072 78010 11100 79200
rect 11072 77982 11376 78010
rect 10956 77820 11252 77840
rect 11012 77818 11036 77820
rect 11092 77818 11116 77820
rect 11172 77818 11196 77820
rect 11034 77766 11036 77818
rect 11098 77766 11110 77818
rect 11172 77766 11174 77818
rect 11012 77764 11036 77766
rect 11092 77764 11116 77766
rect 11172 77764 11196 77766
rect 10956 77744 11252 77764
rect 10324 77376 10376 77382
rect 10324 77318 10376 77324
rect 10138 75848 10194 75857
rect 10138 75783 10194 75792
rect 10140 75744 10192 75750
rect 10060 75704 10140 75732
rect 10140 75686 10192 75692
rect 10152 75342 10180 75686
rect 10140 75336 10192 75342
rect 10140 75278 10192 75284
rect 9678 74760 9734 74769
rect 9678 74695 9734 74704
rect 7852 71318 8248 71346
rect 7760 71182 8156 71210
rect 7564 71120 7616 71126
rect 7564 71062 7616 71068
rect 8024 71120 8076 71126
rect 8024 71062 8076 71068
rect 7930 60616 7986 60625
rect 7930 60551 7986 60560
rect 7840 51808 7892 51814
rect 7840 51750 7892 51756
rect 7852 51377 7880 51750
rect 7838 51368 7894 51377
rect 7838 51303 7894 51312
rect 7838 48104 7894 48113
rect 7838 48039 7894 48048
rect 7852 47802 7880 48039
rect 7840 47796 7892 47802
rect 7840 47738 7892 47744
rect 7746 44432 7802 44441
rect 7746 44367 7802 44376
rect 7564 43852 7616 43858
rect 7564 43794 7616 43800
rect 7472 30932 7524 30938
rect 7472 30874 7524 30880
rect 7472 30592 7524 30598
rect 7472 30534 7524 30540
rect 7484 30326 7512 30534
rect 7472 30320 7524 30326
rect 7472 30262 7524 30268
rect 7472 30184 7524 30190
rect 7472 30126 7524 30132
rect 7380 27668 7432 27674
rect 7380 27610 7432 27616
rect 7208 27526 7420 27554
rect 7288 27464 7340 27470
rect 7288 27406 7340 27412
rect 7104 26580 7156 26586
rect 7104 26522 7156 26528
rect 7012 26376 7064 26382
rect 7012 26318 7064 26324
rect 7116 25498 7144 26522
rect 7300 26314 7328 27406
rect 7288 26308 7340 26314
rect 7288 26250 7340 26256
rect 7194 26208 7250 26217
rect 7194 26143 7250 26152
rect 7208 26042 7236 26143
rect 7196 26036 7248 26042
rect 7196 25978 7248 25984
rect 7104 25492 7156 25498
rect 7104 25434 7156 25440
rect 7116 24410 7144 25434
rect 7300 24682 7328 26250
rect 7392 25401 7420 27526
rect 7484 26353 7512 30126
rect 7470 26344 7526 26353
rect 7470 26279 7526 26288
rect 7378 25392 7434 25401
rect 7378 25327 7434 25336
rect 7288 24676 7340 24682
rect 7288 24618 7340 24624
rect 7104 24404 7156 24410
rect 7104 24346 7156 24352
rect 6840 23854 6960 23882
rect 7116 23866 7144 24346
rect 6826 23760 6882 23769
rect 6826 23695 6882 23704
rect 6840 23186 6868 23695
rect 6828 23180 6880 23186
rect 6828 23122 6880 23128
rect 6932 23118 6960 23854
rect 7104 23860 7156 23866
rect 7104 23802 7156 23808
rect 6920 23112 6972 23118
rect 6920 23054 6972 23060
rect 7116 22930 7144 23802
rect 7196 23180 7248 23186
rect 7196 23122 7248 23128
rect 6840 22902 7144 22930
rect 6840 22642 6868 22902
rect 7208 22778 7236 23122
rect 7288 23112 7340 23118
rect 7288 23054 7340 23060
rect 7196 22772 7248 22778
rect 7196 22714 7248 22720
rect 7300 22642 7328 23054
rect 6828 22636 6880 22642
rect 6828 22578 6880 22584
rect 7104 22636 7156 22642
rect 7104 22578 7156 22584
rect 7288 22636 7340 22642
rect 7288 22578 7340 22584
rect 6840 22098 6868 22578
rect 7116 22438 7144 22578
rect 7104 22432 7156 22438
rect 7104 22374 7156 22380
rect 6828 22092 6880 22098
rect 6828 22034 6880 22040
rect 7378 21720 7434 21729
rect 7378 21655 7434 21664
rect 6920 21412 6972 21418
rect 6920 21354 6972 21360
rect 6644 19110 6696 19116
rect 6734 19136 6790 19145
rect 6656 18970 6684 19110
rect 6734 19071 6790 19080
rect 6644 18964 6696 18970
rect 6644 18906 6696 18912
rect 5956 18524 6252 18544
rect 6012 18522 6036 18524
rect 6092 18522 6116 18524
rect 6172 18522 6196 18524
rect 6034 18470 6036 18522
rect 6098 18470 6110 18522
rect 6172 18470 6174 18522
rect 6012 18468 6036 18470
rect 6092 18468 6116 18470
rect 6172 18468 6196 18470
rect 5956 18448 6252 18468
rect 5172 17672 5224 17678
rect 5172 17614 5224 17620
rect 5184 16250 5212 17614
rect 5956 17436 6252 17456
rect 6012 17434 6036 17436
rect 6092 17434 6116 17436
rect 6172 17434 6196 17436
rect 6034 17382 6036 17434
rect 6098 17382 6110 17434
rect 6172 17382 6174 17434
rect 6012 17380 6036 17382
rect 6092 17380 6116 17382
rect 6172 17380 6196 17382
rect 5956 17360 6252 17380
rect 5816 16652 5868 16658
rect 5816 16594 5868 16600
rect 5172 16244 5224 16250
rect 5172 16186 5224 16192
rect 3700 16040 3752 16046
rect 3700 15982 3752 15988
rect 3514 10296 3570 10305
rect 3514 10231 3570 10240
rect 3330 8936 3386 8945
rect 3330 8871 3386 8880
rect 3712 4146 3740 15982
rect 5828 15910 5856 16594
rect 6552 16584 6604 16590
rect 6604 16544 6684 16572
rect 6552 16526 6604 16532
rect 5956 16348 6252 16368
rect 6012 16346 6036 16348
rect 6092 16346 6116 16348
rect 6172 16346 6196 16348
rect 6034 16294 6036 16346
rect 6098 16294 6110 16346
rect 6172 16294 6174 16346
rect 6012 16292 6036 16294
rect 6092 16292 6116 16294
rect 6172 16292 6196 16294
rect 5956 16272 6252 16292
rect 6656 16250 6684 16544
rect 6644 16244 6696 16250
rect 6644 16186 6696 16192
rect 5816 15904 5868 15910
rect 5816 15846 5868 15852
rect 3974 11248 4030 11257
rect 3974 11183 4030 11192
rect 3882 10568 3938 10577
rect 3882 10503 3938 10512
rect 3896 6905 3924 10503
rect 3882 6896 3938 6905
rect 3882 6831 3938 6840
rect 3988 4185 4016 11183
rect 5828 11121 5856 15846
rect 6656 15706 6684 16186
rect 6644 15700 6696 15706
rect 6644 15642 6696 15648
rect 6656 15502 6684 15642
rect 6644 15496 6696 15502
rect 6644 15438 6696 15444
rect 5956 15260 6252 15280
rect 6012 15258 6036 15260
rect 6092 15258 6116 15260
rect 6172 15258 6196 15260
rect 6034 15206 6036 15258
rect 6098 15206 6110 15258
rect 6172 15206 6174 15258
rect 6012 15204 6036 15206
rect 6092 15204 6116 15206
rect 6172 15204 6196 15206
rect 5956 15184 6252 15204
rect 6656 15162 6684 15438
rect 6644 15156 6696 15162
rect 6644 15098 6696 15104
rect 5956 14172 6252 14192
rect 6012 14170 6036 14172
rect 6092 14170 6116 14172
rect 6172 14170 6196 14172
rect 6034 14118 6036 14170
rect 6098 14118 6110 14170
rect 6172 14118 6174 14170
rect 6012 14116 6036 14118
rect 6092 14116 6116 14118
rect 6172 14116 6196 14118
rect 5956 14096 6252 14116
rect 5956 13084 6252 13104
rect 6012 13082 6036 13084
rect 6092 13082 6116 13084
rect 6172 13082 6196 13084
rect 6034 13030 6036 13082
rect 6098 13030 6110 13082
rect 6172 13030 6174 13082
rect 6012 13028 6036 13030
rect 6092 13028 6116 13030
rect 6172 13028 6196 13030
rect 5956 13008 6252 13028
rect 5956 11996 6252 12016
rect 6012 11994 6036 11996
rect 6092 11994 6116 11996
rect 6172 11994 6196 11996
rect 6034 11942 6036 11994
rect 6098 11942 6110 11994
rect 6172 11942 6174 11994
rect 6012 11940 6036 11942
rect 6092 11940 6116 11942
rect 6172 11940 6196 11942
rect 5956 11920 6252 11940
rect 6932 11257 6960 21354
rect 7288 21344 7340 21350
rect 7288 21286 7340 21292
rect 7300 19310 7328 21286
rect 7288 19304 7340 19310
rect 7288 19246 7340 19252
rect 7196 18828 7248 18834
rect 7196 18770 7248 18776
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 7116 18426 7144 18702
rect 7104 18420 7156 18426
rect 7104 18362 7156 18368
rect 7208 18358 7236 18770
rect 7196 18352 7248 18358
rect 7196 18294 7248 18300
rect 7286 15736 7342 15745
rect 7286 15671 7342 15680
rect 7012 15632 7064 15638
rect 7012 15574 7064 15580
rect 7024 14822 7052 15574
rect 7300 15570 7328 15671
rect 7288 15564 7340 15570
rect 7288 15506 7340 15512
rect 7300 15162 7328 15506
rect 7288 15156 7340 15162
rect 7288 15098 7340 15104
rect 7012 14816 7064 14822
rect 7012 14758 7064 14764
rect 7024 13190 7052 14758
rect 7392 13394 7420 21655
rect 7484 20058 7512 26279
rect 7472 20052 7524 20058
rect 7472 19994 7524 20000
rect 7484 19378 7512 19994
rect 7472 19372 7524 19378
rect 7472 19314 7524 19320
rect 7576 17252 7604 43794
rect 7760 43790 7788 44367
rect 7748 43784 7800 43790
rect 7748 43726 7800 43732
rect 7760 43450 7788 43726
rect 7748 43444 7800 43450
rect 7748 43386 7800 43392
rect 7840 37664 7892 37670
rect 7840 37606 7892 37612
rect 7748 37460 7800 37466
rect 7748 37402 7800 37408
rect 7656 36032 7708 36038
rect 7656 35974 7708 35980
rect 7668 35766 7696 35974
rect 7656 35760 7708 35766
rect 7656 35702 7708 35708
rect 7668 35494 7696 35702
rect 7656 35488 7708 35494
rect 7760 35465 7788 37402
rect 7852 36530 7880 37606
rect 7944 36786 7972 60551
rect 7932 36780 7984 36786
rect 7932 36722 7984 36728
rect 7852 36502 7972 36530
rect 7840 36372 7892 36378
rect 7840 36314 7892 36320
rect 7852 35630 7880 36314
rect 7944 36106 7972 36502
rect 7932 36100 7984 36106
rect 7932 36042 7984 36048
rect 7840 35624 7892 35630
rect 7840 35566 7892 35572
rect 7656 35430 7708 35436
rect 7746 35456 7802 35465
rect 7746 35391 7802 35400
rect 7656 34536 7708 34542
rect 7656 34478 7708 34484
rect 7668 34105 7696 34478
rect 7654 34096 7710 34105
rect 7654 34031 7710 34040
rect 7760 33946 7788 35391
rect 7840 35148 7892 35154
rect 7840 35090 7892 35096
rect 7852 35057 7880 35090
rect 7838 35048 7894 35057
rect 7838 34983 7894 34992
rect 7930 34776 7986 34785
rect 7930 34711 7986 34720
rect 7668 33918 7788 33946
rect 7668 32842 7696 33918
rect 7748 33584 7800 33590
rect 7748 33526 7800 33532
rect 7760 33153 7788 33526
rect 7746 33144 7802 33153
rect 7746 33079 7802 33088
rect 7840 33108 7892 33114
rect 7840 33050 7892 33056
rect 7748 32904 7800 32910
rect 7748 32846 7800 32852
rect 7656 32836 7708 32842
rect 7656 32778 7708 32784
rect 7654 32600 7710 32609
rect 7654 32535 7710 32544
rect 7668 32366 7696 32535
rect 7656 32360 7708 32366
rect 7656 32302 7708 32308
rect 7668 31958 7696 32302
rect 7656 31952 7708 31958
rect 7656 31894 7708 31900
rect 7656 30116 7708 30122
rect 7656 30058 7708 30064
rect 7668 29782 7696 30058
rect 7656 29776 7708 29782
rect 7656 29718 7708 29724
rect 7668 25265 7696 29718
rect 7654 25256 7710 25265
rect 7654 25191 7710 25200
rect 7576 17224 7696 17252
rect 7562 15056 7618 15065
rect 7562 14991 7618 15000
rect 7576 14550 7604 14991
rect 7564 14544 7616 14550
rect 7564 14486 7616 14492
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 7012 13184 7064 13190
rect 7012 13126 7064 13132
rect 6918 11248 6974 11257
rect 7024 11218 7052 13126
rect 7392 12986 7420 13330
rect 7380 12980 7432 12986
rect 7380 12922 7432 12928
rect 6918 11183 6974 11192
rect 7012 11212 7064 11218
rect 7012 11154 7064 11160
rect 4618 11112 4674 11121
rect 4618 11047 4674 11056
rect 5814 11112 5870 11121
rect 5814 11047 5870 11056
rect 4066 10976 4122 10985
rect 4066 10911 4122 10920
rect 4080 10169 4108 10911
rect 4066 10160 4122 10169
rect 4066 10095 4122 10104
rect 4066 7032 4122 7041
rect 4066 6967 4122 6976
rect 3974 4176 4030 4185
rect 3700 4140 3752 4146
rect 3974 4111 4030 4120
rect 3700 4082 3752 4088
rect 4080 3505 4108 6967
rect 4066 3496 4122 3505
rect 4066 3431 4122 3440
rect 3146 2000 3202 2009
rect 3146 1935 3202 1944
rect 2962 912 3018 921
rect 2962 847 3018 856
rect 18 0 74 800
rect 478 0 534 800
rect 1398 0 1454 800
rect 2318 0 2374 800
rect 2778 0 2834 800
rect 3160 785 3188 1935
rect 3698 912 3754 921
rect 3698 847 3754 856
rect 3712 800 3740 847
rect 4632 800 4660 11047
rect 5956 10908 6252 10928
rect 6012 10906 6036 10908
rect 6092 10906 6116 10908
rect 6172 10906 6196 10908
rect 6034 10854 6036 10906
rect 6098 10854 6110 10906
rect 6172 10854 6174 10906
rect 6012 10852 6036 10854
rect 6092 10852 6116 10854
rect 6172 10852 6196 10854
rect 5956 10832 6252 10852
rect 5956 9820 6252 9840
rect 6012 9818 6036 9820
rect 6092 9818 6116 9820
rect 6172 9818 6196 9820
rect 6034 9766 6036 9818
rect 6098 9766 6110 9818
rect 6172 9766 6174 9818
rect 6012 9764 6036 9766
rect 6092 9764 6116 9766
rect 6172 9764 6196 9766
rect 5956 9744 6252 9764
rect 5956 8732 6252 8752
rect 6012 8730 6036 8732
rect 6092 8730 6116 8732
rect 6172 8730 6196 8732
rect 6034 8678 6036 8730
rect 6098 8678 6110 8730
rect 6172 8678 6174 8730
rect 6012 8676 6036 8678
rect 6092 8676 6116 8678
rect 6172 8676 6196 8678
rect 5956 8656 6252 8676
rect 5956 7644 6252 7664
rect 6012 7642 6036 7644
rect 6092 7642 6116 7644
rect 6172 7642 6196 7644
rect 6034 7590 6036 7642
rect 6098 7590 6110 7642
rect 6172 7590 6174 7642
rect 6012 7588 6036 7590
rect 6092 7588 6116 7590
rect 6172 7588 6196 7590
rect 5956 7568 6252 7588
rect 7668 7585 7696 17224
rect 7654 7576 7710 7585
rect 7654 7511 7710 7520
rect 7760 7449 7788 32846
rect 7852 30274 7880 33050
rect 7944 32570 7972 34711
rect 7932 32564 7984 32570
rect 7932 32506 7984 32512
rect 7932 31884 7984 31890
rect 7932 31826 7984 31832
rect 7944 31482 7972 31826
rect 7932 31476 7984 31482
rect 7932 31418 7984 31424
rect 7852 30246 7972 30274
rect 7944 30190 7972 30246
rect 7932 30184 7984 30190
rect 7932 30126 7984 30132
rect 7930 28928 7986 28937
rect 7930 28863 7986 28872
rect 7840 28552 7892 28558
rect 7838 28520 7840 28529
rect 7892 28520 7894 28529
rect 7944 28490 7972 28863
rect 7838 28455 7894 28464
rect 7932 28484 7984 28490
rect 7932 28426 7984 28432
rect 7944 28393 7972 28426
rect 7930 28384 7986 28393
rect 7930 28319 7986 28328
rect 7840 28212 7892 28218
rect 7840 28154 7892 28160
rect 7852 27470 7880 28154
rect 7932 27532 7984 27538
rect 7932 27474 7984 27480
rect 7840 27464 7892 27470
rect 7840 27406 7892 27412
rect 7852 27130 7880 27406
rect 7944 27130 7972 27474
rect 7840 27124 7892 27130
rect 7840 27066 7892 27072
rect 7932 27124 7984 27130
rect 7932 27066 7984 27072
rect 7840 22976 7892 22982
rect 7840 22918 7892 22924
rect 7852 22817 7880 22918
rect 7838 22808 7894 22817
rect 7838 22743 7894 22752
rect 7852 22642 7880 22743
rect 7840 22636 7892 22642
rect 7840 22578 7892 22584
rect 7932 21888 7984 21894
rect 7932 21830 7984 21836
rect 7944 21486 7972 21830
rect 7932 21480 7984 21486
rect 7932 21422 7984 21428
rect 7944 21146 7972 21422
rect 7932 21140 7984 21146
rect 7932 21082 7984 21088
rect 8036 19174 8064 71062
rect 8128 34610 8156 71182
rect 8220 66201 8248 71318
rect 9126 69456 9182 69465
rect 9126 69391 9182 69400
rect 9140 68474 9168 69391
rect 9128 68468 9180 68474
rect 9128 68410 9180 68416
rect 8206 66192 8262 66201
rect 8206 66127 8262 66136
rect 9680 57316 9732 57322
rect 9680 57258 9732 57264
rect 8758 57216 8814 57225
rect 8758 57151 8814 57160
rect 8390 52184 8446 52193
rect 8390 52119 8392 52128
rect 8444 52119 8446 52128
rect 8392 52090 8444 52096
rect 8404 51950 8432 52090
rect 8392 51944 8444 51950
rect 8392 51886 8444 51892
rect 8206 48240 8262 48249
rect 8206 48175 8262 48184
rect 8220 47598 8248 48175
rect 8208 47592 8260 47598
rect 8208 47534 8260 47540
rect 8220 47258 8248 47534
rect 8208 47252 8260 47258
rect 8208 47194 8260 47200
rect 8298 46608 8354 46617
rect 8298 46543 8354 46552
rect 8312 38865 8340 46543
rect 8772 43897 8800 57151
rect 9692 55826 9720 57258
rect 9680 55820 9732 55826
rect 9680 55762 9732 55768
rect 8942 50280 8998 50289
rect 8942 50215 8998 50224
rect 8956 49978 8984 50215
rect 8944 49972 8996 49978
rect 8944 49914 8996 49920
rect 10336 49842 10364 77318
rect 10956 76732 11252 76752
rect 11012 76730 11036 76732
rect 11092 76730 11116 76732
rect 11172 76730 11196 76732
rect 11034 76678 11036 76730
rect 11098 76678 11110 76730
rect 11172 76678 11174 76730
rect 11012 76676 11036 76678
rect 11092 76676 11116 76678
rect 11172 76676 11196 76678
rect 10956 76656 11252 76676
rect 10956 75644 11252 75664
rect 11012 75642 11036 75644
rect 11092 75642 11116 75644
rect 11172 75642 11196 75644
rect 11034 75590 11036 75642
rect 11098 75590 11110 75642
rect 11172 75590 11174 75642
rect 11012 75588 11036 75590
rect 11092 75588 11116 75590
rect 11172 75588 11196 75590
rect 10956 75568 11252 75588
rect 11348 75410 11376 77982
rect 11612 76288 11664 76294
rect 11612 76230 11664 76236
rect 10508 75404 10560 75410
rect 10508 75346 10560 75352
rect 11336 75404 11388 75410
rect 11336 75346 11388 75352
rect 10520 75002 10548 75346
rect 10784 75336 10836 75342
rect 10784 75278 10836 75284
rect 10508 74996 10560 75002
rect 10508 74938 10560 74944
rect 10796 74662 10824 75278
rect 10784 74656 10836 74662
rect 10784 74598 10836 74604
rect 10796 69465 10824 74598
rect 10956 74556 11252 74576
rect 11012 74554 11036 74556
rect 11092 74554 11116 74556
rect 11172 74554 11196 74556
rect 11034 74502 11036 74554
rect 11098 74502 11110 74554
rect 11172 74502 11174 74554
rect 11012 74500 11036 74502
rect 11092 74500 11116 74502
rect 11172 74500 11196 74502
rect 10956 74480 11252 74500
rect 10956 73468 11252 73488
rect 11012 73466 11036 73468
rect 11092 73466 11116 73468
rect 11172 73466 11196 73468
rect 11034 73414 11036 73466
rect 11098 73414 11110 73466
rect 11172 73414 11174 73466
rect 11012 73412 11036 73414
rect 11092 73412 11116 73414
rect 11172 73412 11196 73414
rect 10956 73392 11252 73412
rect 11518 73264 11574 73273
rect 11518 73199 11574 73208
rect 10956 72380 11252 72400
rect 11012 72378 11036 72380
rect 11092 72378 11116 72380
rect 11172 72378 11196 72380
rect 11034 72326 11036 72378
rect 11098 72326 11110 72378
rect 11172 72326 11174 72378
rect 11012 72324 11036 72326
rect 11092 72324 11116 72326
rect 11172 72324 11196 72326
rect 10956 72304 11252 72324
rect 10956 71292 11252 71312
rect 11012 71290 11036 71292
rect 11092 71290 11116 71292
rect 11172 71290 11196 71292
rect 11034 71238 11036 71290
rect 11098 71238 11110 71290
rect 11172 71238 11174 71290
rect 11012 71236 11036 71238
rect 11092 71236 11116 71238
rect 11172 71236 11196 71238
rect 10956 71216 11252 71236
rect 10956 70204 11252 70224
rect 11012 70202 11036 70204
rect 11092 70202 11116 70204
rect 11172 70202 11196 70204
rect 11034 70150 11036 70202
rect 11098 70150 11110 70202
rect 11172 70150 11174 70202
rect 11012 70148 11036 70150
rect 11092 70148 11116 70150
rect 11172 70148 11196 70150
rect 10956 70128 11252 70148
rect 10782 69456 10838 69465
rect 10782 69391 10838 69400
rect 11336 69352 11388 69358
rect 11336 69294 11388 69300
rect 10956 69116 11252 69136
rect 11012 69114 11036 69116
rect 11092 69114 11116 69116
rect 11172 69114 11196 69116
rect 11034 69062 11036 69114
rect 11098 69062 11110 69114
rect 11172 69062 11174 69114
rect 11012 69060 11036 69062
rect 11092 69060 11116 69062
rect 11172 69060 11196 69062
rect 10956 69040 11252 69060
rect 11348 68474 11376 69294
rect 11532 68921 11560 73199
rect 11518 68912 11574 68921
rect 11518 68847 11574 68856
rect 10692 68468 10744 68474
rect 10692 68410 10744 68416
rect 11336 68468 11388 68474
rect 11336 68410 11388 68416
rect 10704 67386 10732 68410
rect 10956 68028 11252 68048
rect 11012 68026 11036 68028
rect 11092 68026 11116 68028
rect 11172 68026 11196 68028
rect 11034 67974 11036 68026
rect 11098 67974 11110 68026
rect 11172 67974 11174 68026
rect 11012 67972 11036 67974
rect 11092 67972 11116 67974
rect 11172 67972 11196 67974
rect 10956 67952 11252 67972
rect 11624 67697 11652 76230
rect 11992 75290 12020 79200
rect 12452 76514 12480 79200
rect 12452 76486 12572 76514
rect 12348 76424 12400 76430
rect 12348 76366 12400 76372
rect 12440 76424 12492 76430
rect 12440 76366 12492 76372
rect 12164 75880 12216 75886
rect 12162 75848 12164 75857
rect 12216 75848 12218 75857
rect 12162 75783 12218 75792
rect 12360 75750 12388 76366
rect 12452 75954 12480 76366
rect 12440 75948 12492 75954
rect 12440 75890 12492 75896
rect 12348 75744 12400 75750
rect 12348 75686 12400 75692
rect 12440 75744 12492 75750
rect 12440 75686 12492 75692
rect 11992 75262 12296 75290
rect 11980 75200 12032 75206
rect 11980 75142 12032 75148
rect 11992 74322 12020 75142
rect 11980 74316 12032 74322
rect 11980 74258 12032 74264
rect 11992 73914 12020 74258
rect 11980 73908 12032 73914
rect 11980 73850 12032 73856
rect 11242 67688 11298 67697
rect 11242 67623 11244 67632
rect 11296 67623 11298 67632
rect 11610 67688 11666 67697
rect 11610 67623 11666 67632
rect 11978 67688 12034 67697
rect 11978 67623 11980 67632
rect 11244 67594 11296 67600
rect 12032 67623 12034 67632
rect 11980 67594 12032 67600
rect 12268 67561 12296 75262
rect 12452 75206 12480 75686
rect 12440 75200 12492 75206
rect 12440 75142 12492 75148
rect 12348 74248 12400 74254
rect 12452 74202 12480 75142
rect 12544 74798 12572 76486
rect 13372 75857 13400 79200
rect 13820 77376 13872 77382
rect 13820 77318 13872 77324
rect 13832 76974 13860 77318
rect 14292 77042 14320 79200
rect 14280 77036 14332 77042
rect 14280 76978 14332 76984
rect 13820 76968 13872 76974
rect 13820 76910 13872 76916
rect 13726 76392 13782 76401
rect 13726 76327 13728 76336
rect 13780 76327 13782 76336
rect 13728 76298 13780 76304
rect 13544 75880 13596 75886
rect 13358 75848 13414 75857
rect 13832 75868 13860 76910
rect 13596 75840 13860 75868
rect 13544 75822 13596 75828
rect 13358 75783 13414 75792
rect 13360 75744 13412 75750
rect 13358 75712 13360 75721
rect 13412 75712 13414 75721
rect 13358 75647 13414 75656
rect 14752 74798 14780 79200
rect 15292 76832 15344 76838
rect 15292 76774 15344 76780
rect 15106 75848 15162 75857
rect 15106 75783 15162 75792
rect 15120 75750 15148 75783
rect 15108 75744 15160 75750
rect 15108 75686 15160 75692
rect 12532 74792 12584 74798
rect 12532 74734 12584 74740
rect 13728 74792 13780 74798
rect 13728 74734 13780 74740
rect 13820 74792 13872 74798
rect 13820 74734 13872 74740
rect 14740 74792 14792 74798
rect 14740 74734 14792 74740
rect 12400 74196 12480 74202
rect 12348 74190 12480 74196
rect 12360 74174 12480 74190
rect 12452 73574 12480 74174
rect 13084 74112 13136 74118
rect 13084 74054 13136 74060
rect 12440 73568 12492 73574
rect 12440 73510 12492 73516
rect 12452 73166 12480 73510
rect 13096 73234 13124 74054
rect 13084 73228 13136 73234
rect 13084 73170 13136 73176
rect 12440 73160 12492 73166
rect 12440 73102 12492 73108
rect 12452 72486 12480 73102
rect 13096 72826 13124 73170
rect 13084 72820 13136 72826
rect 13084 72762 13136 72768
rect 12440 72480 12492 72486
rect 12440 72422 12492 72428
rect 12348 69488 12400 69494
rect 12348 69430 12400 69436
rect 12360 69170 12388 69430
rect 12452 69170 12480 72422
rect 12622 70408 12678 70417
rect 12622 70343 12678 70352
rect 12360 69142 12480 69170
rect 12254 67552 12310 67561
rect 12254 67487 12310 67496
rect 11518 67416 11574 67425
rect 10692 67380 10744 67386
rect 11518 67351 11574 67360
rect 10692 67322 10744 67328
rect 10956 66940 11252 66960
rect 11012 66938 11036 66940
rect 11092 66938 11116 66940
rect 11172 66938 11196 66940
rect 11034 66886 11036 66938
rect 11098 66886 11110 66938
rect 11172 66886 11174 66938
rect 11012 66884 11036 66886
rect 11092 66884 11116 66886
rect 11172 66884 11196 66886
rect 10956 66864 11252 66884
rect 10956 65852 11252 65872
rect 11012 65850 11036 65852
rect 11092 65850 11116 65852
rect 11172 65850 11196 65852
rect 11034 65798 11036 65850
rect 11098 65798 11110 65850
rect 11172 65798 11174 65850
rect 11012 65796 11036 65798
rect 11092 65796 11116 65798
rect 11172 65796 11196 65798
rect 10956 65776 11252 65796
rect 10956 64764 11252 64784
rect 11012 64762 11036 64764
rect 11092 64762 11116 64764
rect 11172 64762 11196 64764
rect 11034 64710 11036 64762
rect 11098 64710 11110 64762
rect 11172 64710 11174 64762
rect 11012 64708 11036 64710
rect 11092 64708 11116 64710
rect 11172 64708 11196 64710
rect 10956 64688 11252 64708
rect 10956 63676 11252 63696
rect 11012 63674 11036 63676
rect 11092 63674 11116 63676
rect 11172 63674 11196 63676
rect 11034 63622 11036 63674
rect 11098 63622 11110 63674
rect 11172 63622 11174 63674
rect 11012 63620 11036 63622
rect 11092 63620 11116 63622
rect 11172 63620 11196 63622
rect 10956 63600 11252 63620
rect 10956 62588 11252 62608
rect 11012 62586 11036 62588
rect 11092 62586 11116 62588
rect 11172 62586 11196 62588
rect 11034 62534 11036 62586
rect 11098 62534 11110 62586
rect 11172 62534 11174 62586
rect 11012 62532 11036 62534
rect 11092 62532 11116 62534
rect 11172 62532 11196 62534
rect 10956 62512 11252 62532
rect 10956 61500 11252 61520
rect 11012 61498 11036 61500
rect 11092 61498 11116 61500
rect 11172 61498 11196 61500
rect 11034 61446 11036 61498
rect 11098 61446 11110 61498
rect 11172 61446 11174 61498
rect 11012 61444 11036 61446
rect 11092 61444 11116 61446
rect 11172 61444 11196 61446
rect 10956 61424 11252 61444
rect 10956 60412 11252 60432
rect 11012 60410 11036 60412
rect 11092 60410 11116 60412
rect 11172 60410 11196 60412
rect 11034 60358 11036 60410
rect 11098 60358 11110 60410
rect 11172 60358 11174 60410
rect 11012 60356 11036 60358
rect 11092 60356 11116 60358
rect 11172 60356 11196 60358
rect 10956 60336 11252 60356
rect 10956 59324 11252 59344
rect 11012 59322 11036 59324
rect 11092 59322 11116 59324
rect 11172 59322 11196 59324
rect 11034 59270 11036 59322
rect 11098 59270 11110 59322
rect 11172 59270 11174 59322
rect 11012 59268 11036 59270
rect 11092 59268 11116 59270
rect 11172 59268 11196 59270
rect 10956 59248 11252 59268
rect 10956 58236 11252 58256
rect 11012 58234 11036 58236
rect 11092 58234 11116 58236
rect 11172 58234 11196 58236
rect 11034 58182 11036 58234
rect 11098 58182 11110 58234
rect 11172 58182 11174 58234
rect 11012 58180 11036 58182
rect 11092 58180 11116 58182
rect 11172 58180 11196 58182
rect 10956 58160 11252 58180
rect 11532 58041 11560 67351
rect 11980 67040 12032 67046
rect 11980 66982 12032 66988
rect 11992 58138 12020 66982
rect 12452 61810 12480 69142
rect 12636 64920 12664 70343
rect 12636 64892 12756 64920
rect 12440 61804 12492 61810
rect 12440 61746 12492 61752
rect 12164 61736 12216 61742
rect 12164 61678 12216 61684
rect 11704 58132 11756 58138
rect 11704 58074 11756 58080
rect 11980 58132 12032 58138
rect 11980 58074 12032 58080
rect 11518 58032 11574 58041
rect 11518 57967 11574 57976
rect 10956 57148 11252 57168
rect 11012 57146 11036 57148
rect 11092 57146 11116 57148
rect 11172 57146 11196 57148
rect 11034 57094 11036 57146
rect 11098 57094 11110 57146
rect 11172 57094 11174 57146
rect 11012 57092 11036 57094
rect 11092 57092 11116 57094
rect 11172 57092 11196 57094
rect 10956 57072 11252 57092
rect 10956 56060 11252 56080
rect 11012 56058 11036 56060
rect 11092 56058 11116 56060
rect 11172 56058 11196 56060
rect 11034 56006 11036 56058
rect 11098 56006 11110 56058
rect 11172 56006 11174 56058
rect 11012 56004 11036 56006
rect 11092 56004 11116 56006
rect 11172 56004 11196 56006
rect 10956 55984 11252 56004
rect 10600 55820 10652 55826
rect 10600 55762 10652 55768
rect 10612 55418 10640 55762
rect 10876 55752 10928 55758
rect 10876 55694 10928 55700
rect 10888 55418 10916 55694
rect 10600 55412 10652 55418
rect 10600 55354 10652 55360
rect 10876 55412 10928 55418
rect 10876 55354 10928 55360
rect 10888 53242 10916 55354
rect 10956 54972 11252 54992
rect 11012 54970 11036 54972
rect 11092 54970 11116 54972
rect 11172 54970 11196 54972
rect 11034 54918 11036 54970
rect 11098 54918 11110 54970
rect 11172 54918 11174 54970
rect 11012 54916 11036 54918
rect 11092 54916 11116 54918
rect 11172 54916 11196 54918
rect 10956 54896 11252 54916
rect 11518 54088 11574 54097
rect 11518 54023 11574 54032
rect 11532 53990 11560 54023
rect 11520 53984 11572 53990
rect 11520 53926 11572 53932
rect 10956 53884 11252 53904
rect 11012 53882 11036 53884
rect 11092 53882 11116 53884
rect 11172 53882 11196 53884
rect 11034 53830 11036 53882
rect 11098 53830 11110 53882
rect 11172 53830 11174 53882
rect 11012 53828 11036 53830
rect 11092 53828 11116 53830
rect 11172 53828 11196 53830
rect 10956 53808 11252 53828
rect 11610 53680 11666 53689
rect 11244 53644 11296 53650
rect 11610 53615 11666 53624
rect 11244 53586 11296 53592
rect 10416 53236 10468 53242
rect 10416 53178 10468 53184
rect 10876 53236 10928 53242
rect 10876 53178 10928 53184
rect 10428 51610 10456 53178
rect 11256 52970 11284 53586
rect 11428 53440 11480 53446
rect 11426 53408 11428 53417
rect 11480 53408 11482 53417
rect 11426 53343 11482 53352
rect 11244 52964 11296 52970
rect 11244 52906 11296 52912
rect 11428 52964 11480 52970
rect 11428 52906 11480 52912
rect 10956 52796 11252 52816
rect 11012 52794 11036 52796
rect 11092 52794 11116 52796
rect 11172 52794 11196 52796
rect 11034 52742 11036 52794
rect 11098 52742 11110 52794
rect 11172 52742 11174 52794
rect 11012 52740 11036 52742
rect 11092 52740 11116 52742
rect 11172 52740 11196 52742
rect 10956 52720 11252 52740
rect 11334 52728 11390 52737
rect 10876 52692 10928 52698
rect 11334 52663 11390 52672
rect 10876 52634 10928 52640
rect 10508 51808 10560 51814
rect 10508 51750 10560 51756
rect 10416 51604 10468 51610
rect 10416 51546 10468 51552
rect 10416 51468 10468 51474
rect 10416 51410 10468 51416
rect 10428 51377 10456 51410
rect 10414 51368 10470 51377
rect 10414 51303 10470 51312
rect 10428 51066 10456 51303
rect 10416 51060 10468 51066
rect 10416 51002 10468 51008
rect 10520 49881 10548 51750
rect 10784 51604 10836 51610
rect 10784 51546 10836 51552
rect 10796 50386 10824 51546
rect 10888 51218 10916 52634
rect 11348 52426 11376 52663
rect 11440 52562 11468 52906
rect 11520 52896 11572 52902
rect 11520 52838 11572 52844
rect 11428 52556 11480 52562
rect 11428 52498 11480 52504
rect 11336 52420 11388 52426
rect 11336 52362 11388 52368
rect 10966 52320 11022 52329
rect 10966 52255 11022 52264
rect 10980 52154 11008 52255
rect 11348 52154 11376 52362
rect 10968 52148 11020 52154
rect 10968 52090 11020 52096
rect 11336 52148 11388 52154
rect 11336 52090 11388 52096
rect 10956 51708 11252 51728
rect 11012 51706 11036 51708
rect 11092 51706 11116 51708
rect 11172 51706 11196 51708
rect 11034 51654 11036 51706
rect 11098 51654 11110 51706
rect 11172 51654 11174 51706
rect 11012 51652 11036 51654
rect 11092 51652 11116 51654
rect 11172 51652 11196 51654
rect 10956 51632 11252 51652
rect 11532 51338 11560 52838
rect 11624 52465 11652 53615
rect 11610 52456 11666 52465
rect 11610 52391 11666 52400
rect 11716 52193 11744 58074
rect 12072 57996 12124 58002
rect 12072 57938 12124 57944
rect 12084 57254 12112 57938
rect 12072 57248 12124 57254
rect 12072 57190 12124 57196
rect 12084 56817 12112 57190
rect 12070 56808 12126 56817
rect 12070 56743 12126 56752
rect 12176 55865 12204 61678
rect 12452 61402 12480 61746
rect 12440 61396 12492 61402
rect 12440 61338 12492 61344
rect 12728 60704 12756 64892
rect 13360 62756 13412 62762
rect 13360 62698 13412 62704
rect 12728 60676 12940 60704
rect 12162 55856 12218 55865
rect 12162 55791 12218 55800
rect 11794 55720 11850 55729
rect 11794 55655 11850 55664
rect 11808 52698 11836 55655
rect 12072 55616 12124 55622
rect 12072 55558 12124 55564
rect 12084 55457 12112 55558
rect 12070 55448 12126 55457
rect 12070 55383 12126 55392
rect 12072 54800 12124 54806
rect 12072 54742 12124 54748
rect 11980 54596 12032 54602
rect 11980 54538 12032 54544
rect 11886 54224 11942 54233
rect 11886 54159 11888 54168
rect 11940 54159 11942 54168
rect 11888 54130 11940 54136
rect 11886 53952 11942 53961
rect 11886 53887 11942 53896
rect 11900 53242 11928 53887
rect 11992 53446 12020 54538
rect 12084 53786 12112 54742
rect 12256 54732 12308 54738
rect 12256 54674 12308 54680
rect 12268 54330 12296 54674
rect 12348 54528 12400 54534
rect 12348 54470 12400 54476
rect 12256 54324 12308 54330
rect 12256 54266 12308 54272
rect 12360 54126 12388 54470
rect 12348 54120 12400 54126
rect 12348 54062 12400 54068
rect 12072 53780 12124 53786
rect 12124 53740 12204 53768
rect 12072 53722 12124 53728
rect 12072 53644 12124 53650
rect 12072 53586 12124 53592
rect 11980 53440 12032 53446
rect 11980 53382 12032 53388
rect 11888 53236 11940 53242
rect 11888 53178 11940 53184
rect 11900 53038 11928 53178
rect 11888 53032 11940 53038
rect 11888 52974 11940 52980
rect 11888 52896 11940 52902
rect 11888 52838 11940 52844
rect 11796 52692 11848 52698
rect 11796 52634 11848 52640
rect 11900 52630 11928 52838
rect 11888 52624 11940 52630
rect 11888 52566 11940 52572
rect 11702 52184 11758 52193
rect 11702 52119 11758 52128
rect 11520 51332 11572 51338
rect 11520 51274 11572 51280
rect 10888 51190 11008 51218
rect 10980 51082 11008 51190
rect 10980 51054 11100 51082
rect 11900 51066 11928 52566
rect 11992 52358 12020 53382
rect 12084 52902 12112 53586
rect 12176 53038 12204 53740
rect 12164 53032 12216 53038
rect 12164 52974 12216 52980
rect 12072 52896 12124 52902
rect 12360 52850 12388 54062
rect 12440 53576 12492 53582
rect 12440 53518 12492 53524
rect 12452 53106 12480 53518
rect 12440 53100 12492 53106
rect 12440 53042 12492 53048
rect 12808 53100 12860 53106
rect 12808 53042 12860 53048
rect 12532 53032 12584 53038
rect 12532 52974 12584 52980
rect 12072 52838 12124 52844
rect 11980 52352 12032 52358
rect 11980 52294 12032 52300
rect 11992 52018 12020 52294
rect 11980 52012 12032 52018
rect 11980 51954 12032 51960
rect 11992 51610 12020 51954
rect 11980 51604 12032 51610
rect 11980 51546 12032 51552
rect 11980 51264 12032 51270
rect 11980 51206 12032 51212
rect 11072 50862 11100 51054
rect 11888 51060 11940 51066
rect 11888 51002 11940 51008
rect 11520 50992 11572 50998
rect 11518 50960 11520 50969
rect 11572 50960 11574 50969
rect 11518 50895 11574 50904
rect 11060 50856 11112 50862
rect 11060 50798 11112 50804
rect 10956 50620 11252 50640
rect 11012 50618 11036 50620
rect 11092 50618 11116 50620
rect 11172 50618 11196 50620
rect 11034 50566 11036 50618
rect 11098 50566 11110 50618
rect 11172 50566 11174 50618
rect 11012 50564 11036 50566
rect 11092 50564 11116 50566
rect 11172 50564 11196 50566
rect 10956 50544 11252 50564
rect 10784 50380 10836 50386
rect 10784 50322 10836 50328
rect 11428 50380 11480 50386
rect 11428 50322 11480 50328
rect 10876 50312 10928 50318
rect 10876 50254 10928 50260
rect 10888 49978 10916 50254
rect 10876 49972 10928 49978
rect 10876 49914 10928 49920
rect 10506 49872 10562 49881
rect 10324 49836 10376 49842
rect 10506 49807 10562 49816
rect 10324 49778 10376 49784
rect 10784 49768 10836 49774
rect 10784 49710 10836 49716
rect 10796 49162 10824 49710
rect 10888 49434 10916 49914
rect 11440 49638 11468 50322
rect 11796 50176 11848 50182
rect 11796 50118 11848 50124
rect 11704 49768 11756 49774
rect 11704 49710 11756 49716
rect 11428 49632 11480 49638
rect 11428 49574 11480 49580
rect 10956 49532 11252 49552
rect 11012 49530 11036 49532
rect 11092 49530 11116 49532
rect 11172 49530 11196 49532
rect 11034 49478 11036 49530
rect 11098 49478 11110 49530
rect 11172 49478 11174 49530
rect 11012 49476 11036 49478
rect 11092 49476 11116 49478
rect 11172 49476 11196 49478
rect 10956 49456 11252 49476
rect 10876 49428 10928 49434
rect 10876 49370 10928 49376
rect 11336 49224 11388 49230
rect 11336 49166 11388 49172
rect 11440 49212 11468 49574
rect 11520 49224 11572 49230
rect 11440 49184 11520 49212
rect 10784 49156 10836 49162
rect 10784 49098 10836 49104
rect 11348 48550 11376 49166
rect 11440 49094 11468 49184
rect 11520 49166 11572 49172
rect 11428 49088 11480 49094
rect 11428 49030 11480 49036
rect 11336 48544 11388 48550
rect 11336 48486 11388 48492
rect 10956 48444 11252 48464
rect 11012 48442 11036 48444
rect 11092 48442 11116 48444
rect 11172 48442 11196 48444
rect 11034 48390 11036 48442
rect 11098 48390 11110 48442
rect 11172 48390 11174 48442
rect 11012 48388 11036 48390
rect 11092 48388 11116 48390
rect 11172 48388 11196 48390
rect 10956 48368 11252 48388
rect 11440 48346 11468 49030
rect 11428 48340 11480 48346
rect 11428 48282 11480 48288
rect 11440 48249 11468 48282
rect 11426 48240 11482 48249
rect 11426 48175 11482 48184
rect 9402 48104 9458 48113
rect 9402 48039 9458 48048
rect 8574 43888 8630 43897
rect 8574 43823 8576 43832
rect 8628 43823 8630 43832
rect 8758 43888 8814 43897
rect 8758 43823 8760 43832
rect 8576 43794 8628 43800
rect 8812 43823 8814 43832
rect 8760 43794 8812 43800
rect 8588 43450 8616 43794
rect 8576 43444 8628 43450
rect 8576 43386 8628 43392
rect 8772 43382 8800 43794
rect 8760 43376 8812 43382
rect 8760 43318 8812 43324
rect 8944 42152 8996 42158
rect 9220 42152 9272 42158
rect 8944 42094 8996 42100
rect 9218 42120 9220 42129
rect 9272 42120 9274 42129
rect 8852 38888 8904 38894
rect 8298 38856 8354 38865
rect 8852 38830 8904 38836
rect 8298 38791 8354 38800
rect 8666 38448 8722 38457
rect 8576 38412 8628 38418
rect 8496 38372 8576 38400
rect 8300 38276 8352 38282
rect 8300 38218 8352 38224
rect 8208 37800 8260 37806
rect 8206 37768 8208 37777
rect 8260 37768 8262 37777
rect 8206 37703 8262 37712
rect 8312 37210 8340 38218
rect 8496 37738 8524 38372
rect 8666 38383 8722 38392
rect 8760 38412 8812 38418
rect 8576 38354 8628 38360
rect 8680 37874 8708 38383
rect 8760 38354 8812 38360
rect 8668 37868 8720 37874
rect 8668 37810 8720 37816
rect 8484 37732 8536 37738
rect 8484 37674 8536 37680
rect 8496 37448 8524 37674
rect 8220 37182 8340 37210
rect 8404 37420 8524 37448
rect 8220 36825 8248 37182
rect 8298 37088 8354 37097
rect 8298 37023 8354 37032
rect 8206 36816 8262 36825
rect 8206 36751 8262 36760
rect 8220 35698 8248 36751
rect 8312 36378 8340 37023
rect 8300 36372 8352 36378
rect 8300 36314 8352 36320
rect 8208 35692 8260 35698
rect 8208 35634 8260 35640
rect 8300 35488 8352 35494
rect 8300 35430 8352 35436
rect 8116 34604 8168 34610
rect 8116 34546 8168 34552
rect 8312 34542 8340 35430
rect 8300 34536 8352 34542
rect 8300 34478 8352 34484
rect 8116 33992 8168 33998
rect 8116 33934 8168 33940
rect 8300 33992 8352 33998
rect 8300 33934 8352 33940
rect 8128 33658 8156 33934
rect 8208 33856 8260 33862
rect 8208 33798 8260 33804
rect 8116 33652 8168 33658
rect 8116 33594 8168 33600
rect 8116 33516 8168 33522
rect 8116 33458 8168 33464
rect 8128 33114 8156 33458
rect 8220 33454 8248 33798
rect 8208 33448 8260 33454
rect 8206 33416 8208 33425
rect 8260 33416 8262 33425
rect 8206 33351 8262 33360
rect 8116 33108 8168 33114
rect 8116 33050 8168 33056
rect 8312 32978 8340 33934
rect 8404 33114 8432 37420
rect 8680 37398 8708 37810
rect 8668 37392 8720 37398
rect 8482 37360 8538 37369
rect 8668 37334 8720 37340
rect 8482 37295 8538 37304
rect 8496 36768 8524 37295
rect 8496 36740 8616 36768
rect 8588 36417 8616 36740
rect 8574 36408 8630 36417
rect 8574 36343 8630 36352
rect 8588 36310 8616 36343
rect 8576 36304 8628 36310
rect 8576 36246 8628 36252
rect 8576 36168 8628 36174
rect 8576 36110 8628 36116
rect 8588 35834 8616 36110
rect 8576 35828 8628 35834
rect 8576 35770 8628 35776
rect 8484 35624 8536 35630
rect 8484 35566 8536 35572
rect 8496 34785 8524 35566
rect 8482 34776 8538 34785
rect 8482 34711 8538 34720
rect 8484 34536 8536 34542
rect 8484 34478 8536 34484
rect 8392 33108 8444 33114
rect 8392 33050 8444 33056
rect 8300 32972 8352 32978
rect 8352 32932 8432 32960
rect 8300 32914 8352 32920
rect 8116 32836 8168 32842
rect 8116 32778 8168 32784
rect 8128 32502 8156 32778
rect 8116 32496 8168 32502
rect 8116 32438 8168 32444
rect 8298 32464 8354 32473
rect 8298 32399 8300 32408
rect 8352 32399 8354 32408
rect 8300 32370 8352 32376
rect 8404 32314 8432 32932
rect 8312 32286 8432 32314
rect 8312 32026 8340 32286
rect 8392 32224 8444 32230
rect 8392 32166 8444 32172
rect 8300 32020 8352 32026
rect 8300 31962 8352 31968
rect 8208 31476 8260 31482
rect 8208 31418 8260 31424
rect 8220 31249 8248 31418
rect 8300 31340 8352 31346
rect 8300 31282 8352 31288
rect 8206 31240 8262 31249
rect 8206 31175 8262 31184
rect 8312 30054 8340 31282
rect 8300 30048 8352 30054
rect 8300 29990 8352 29996
rect 8312 29850 8340 29990
rect 8300 29844 8352 29850
rect 8300 29786 8352 29792
rect 8128 29714 8340 29730
rect 8116 29708 8340 29714
rect 8168 29702 8340 29708
rect 8116 29650 8168 29656
rect 8206 29472 8262 29481
rect 8206 29407 8262 29416
rect 8220 29102 8248 29407
rect 8312 29209 8340 29702
rect 8298 29200 8354 29209
rect 8298 29135 8354 29144
rect 8208 29096 8260 29102
rect 8114 29064 8170 29073
rect 8208 29038 8260 29044
rect 8114 28999 8116 29008
rect 8168 28999 8170 29008
rect 8116 28970 8168 28976
rect 8404 28801 8432 32166
rect 8496 31482 8524 34478
rect 8588 33658 8616 35770
rect 8668 34944 8720 34950
rect 8668 34886 8720 34892
rect 8680 34542 8708 34886
rect 8668 34536 8720 34542
rect 8666 34504 8668 34513
rect 8720 34504 8722 34513
rect 8666 34439 8722 34448
rect 8668 33856 8720 33862
rect 8668 33798 8720 33804
rect 8576 33652 8628 33658
rect 8576 33594 8628 33600
rect 8588 32026 8616 33594
rect 8680 33318 8708 33798
rect 8772 33386 8800 38354
rect 8864 36786 8892 38830
rect 8956 37466 8984 42094
rect 9036 42084 9088 42090
rect 9218 42055 9274 42064
rect 9036 42026 9088 42032
rect 9048 41478 9076 42026
rect 9036 41472 9088 41478
rect 9034 41440 9036 41449
rect 9088 41440 9090 41449
rect 9034 41375 9090 41384
rect 9312 38752 9364 38758
rect 9312 38694 9364 38700
rect 9324 38486 9352 38694
rect 9312 38480 9364 38486
rect 9312 38422 9364 38428
rect 9034 38176 9090 38185
rect 9034 38111 9090 38120
rect 9048 38010 9076 38111
rect 9324 38026 9352 38422
rect 9416 38418 9444 48039
rect 9772 47456 9824 47462
rect 9772 47398 9824 47404
rect 9784 47025 9812 47398
rect 10956 47356 11252 47376
rect 11012 47354 11036 47356
rect 11092 47354 11116 47356
rect 11172 47354 11196 47356
rect 11034 47302 11036 47354
rect 11098 47302 11110 47354
rect 11172 47302 11174 47354
rect 11012 47300 11036 47302
rect 11092 47300 11116 47302
rect 11172 47300 11196 47302
rect 10956 47280 11252 47300
rect 9770 47016 9826 47025
rect 9770 46951 9826 46960
rect 9494 46472 9550 46481
rect 9494 46407 9550 46416
rect 9508 41970 9536 46407
rect 10956 46268 11252 46288
rect 11012 46266 11036 46268
rect 11092 46266 11116 46268
rect 11172 46266 11196 46268
rect 11034 46214 11036 46266
rect 11098 46214 11110 46266
rect 11172 46214 11174 46266
rect 11012 46212 11036 46214
rect 11092 46212 11116 46214
rect 11172 46212 11196 46214
rect 10956 46192 11252 46212
rect 11520 45280 11572 45286
rect 11520 45222 11572 45228
rect 10956 45180 11252 45200
rect 11012 45178 11036 45180
rect 11092 45178 11116 45180
rect 11172 45178 11196 45180
rect 11034 45126 11036 45178
rect 11098 45126 11110 45178
rect 11172 45126 11174 45178
rect 11012 45124 11036 45126
rect 11092 45124 11116 45126
rect 11172 45124 11196 45126
rect 10956 45104 11252 45124
rect 11532 44334 11560 45222
rect 11520 44328 11572 44334
rect 11520 44270 11572 44276
rect 10784 44192 10836 44198
rect 10784 44134 10836 44140
rect 10600 43716 10652 43722
rect 10600 43658 10652 43664
rect 9680 43376 9732 43382
rect 9680 43318 9732 43324
rect 9692 42378 9720 43318
rect 10612 43110 10640 43658
rect 10600 43104 10652 43110
rect 10598 43072 10600 43081
rect 10652 43072 10654 43081
rect 10598 43007 10654 43016
rect 10232 42764 10284 42770
rect 10232 42706 10284 42712
rect 10244 42566 10272 42706
rect 10232 42560 10284 42566
rect 10232 42502 10284 42508
rect 9600 42350 9904 42378
rect 9600 42158 9628 42350
rect 9588 42152 9640 42158
rect 9588 42094 9640 42100
rect 9508 41942 9628 41970
rect 9496 38752 9548 38758
rect 9496 38694 9548 38700
rect 9404 38412 9456 38418
rect 9404 38354 9456 38360
rect 9402 38040 9458 38049
rect 9036 38004 9088 38010
rect 9324 37998 9402 38026
rect 9402 37975 9458 37984
rect 9036 37946 9088 37952
rect 9416 37942 9444 37975
rect 9404 37936 9456 37942
rect 9404 37878 9456 37884
rect 9508 37670 9536 38694
rect 9496 37664 9548 37670
rect 9496 37606 9548 37612
rect 8944 37460 8996 37466
rect 8944 37402 8996 37408
rect 9404 37460 9456 37466
rect 9404 37402 9456 37408
rect 9220 37256 9272 37262
rect 9220 37198 9272 37204
rect 9036 37120 9088 37126
rect 9036 37062 9088 37068
rect 8852 36780 8904 36786
rect 8852 36722 8904 36728
rect 8852 36644 8904 36650
rect 8852 36586 8904 36592
rect 8864 36281 8892 36586
rect 8850 36272 8906 36281
rect 8850 36207 8906 36216
rect 8760 33380 8812 33386
rect 8760 33322 8812 33328
rect 8668 33312 8720 33318
rect 8668 33254 8720 33260
rect 8680 33028 8708 33254
rect 8760 33040 8812 33046
rect 8680 33000 8760 33028
rect 8760 32982 8812 32988
rect 8668 32496 8720 32502
rect 8668 32438 8720 32444
rect 8576 32020 8628 32026
rect 8576 31962 8628 31968
rect 8574 31784 8630 31793
rect 8574 31719 8630 31728
rect 8484 31476 8536 31482
rect 8484 31418 8536 31424
rect 8588 31362 8616 31719
rect 8496 31334 8616 31362
rect 8680 31346 8708 32438
rect 8772 32230 8800 32982
rect 8864 32434 8892 36207
rect 9048 36038 9076 37062
rect 9232 36582 9260 37198
rect 9312 36780 9364 36786
rect 9312 36722 9364 36728
rect 9220 36576 9272 36582
rect 9220 36518 9272 36524
rect 9128 36100 9180 36106
rect 9128 36042 9180 36048
rect 9036 36032 9088 36038
rect 9036 35974 9088 35980
rect 9048 35494 9076 35974
rect 9140 35737 9168 36042
rect 9126 35728 9182 35737
rect 9126 35663 9182 35672
rect 9128 35624 9180 35630
rect 9128 35566 9180 35572
rect 9036 35488 9088 35494
rect 9036 35430 9088 35436
rect 9140 35222 9168 35566
rect 9128 35216 9180 35222
rect 9128 35158 9180 35164
rect 8944 35148 8996 35154
rect 8944 35090 8996 35096
rect 8956 35057 8984 35090
rect 9036 35080 9088 35086
rect 8942 35048 8998 35057
rect 9036 35022 9088 35028
rect 9128 35080 9180 35086
rect 9128 35022 9180 35028
rect 8942 34983 8998 34992
rect 8944 34944 8996 34950
rect 8944 34886 8996 34892
rect 8956 34785 8984 34886
rect 8942 34776 8998 34785
rect 8942 34711 8998 34720
rect 8944 34604 8996 34610
rect 8944 34546 8996 34552
rect 8852 32428 8904 32434
rect 8852 32370 8904 32376
rect 8852 32292 8904 32298
rect 8852 32234 8904 32240
rect 8760 32224 8812 32230
rect 8760 32166 8812 32172
rect 8864 32065 8892 32234
rect 8850 32056 8906 32065
rect 8850 31991 8906 32000
rect 8956 31804 8984 34546
rect 9048 34542 9076 35022
rect 9140 34921 9168 35022
rect 9126 34912 9182 34921
rect 9126 34847 9182 34856
rect 9036 34536 9088 34542
rect 9036 34478 9088 34484
rect 9140 34406 9168 34847
rect 9128 34400 9180 34406
rect 9128 34342 9180 34348
rect 9232 33946 9260 36518
rect 9048 33918 9260 33946
rect 9048 32201 9076 33918
rect 9220 33380 9272 33386
rect 9220 33322 9272 33328
rect 9128 33040 9180 33046
rect 9126 33008 9128 33017
rect 9180 33008 9182 33017
rect 9126 32943 9182 32952
rect 9128 32904 9180 32910
rect 9128 32846 9180 32852
rect 9034 32192 9090 32201
rect 9034 32127 9090 32136
rect 9140 32026 9168 32846
rect 9128 32020 9180 32026
rect 9128 31962 9180 31968
rect 9036 31952 9088 31958
rect 9088 31900 9168 31906
rect 9036 31894 9168 31900
rect 9048 31878 9168 31894
rect 8850 31784 8906 31793
rect 8760 31748 8812 31754
rect 8956 31776 9076 31804
rect 8850 31719 8906 31728
rect 8760 31690 8812 31696
rect 8668 31340 8720 31346
rect 8390 28792 8446 28801
rect 8390 28727 8446 28736
rect 8404 28558 8432 28727
rect 8496 28626 8524 31334
rect 8668 31282 8720 31288
rect 8576 31204 8628 31210
rect 8576 31146 8628 31152
rect 8588 30258 8616 31146
rect 8668 31136 8720 31142
rect 8668 31078 8720 31084
rect 8680 30802 8708 31078
rect 8772 30870 8800 31690
rect 8864 31482 8892 31719
rect 8944 31680 8996 31686
rect 8942 31648 8944 31657
rect 8996 31648 8998 31657
rect 8942 31583 8998 31592
rect 8852 31476 8904 31482
rect 8852 31418 8904 31424
rect 8864 31278 8892 31418
rect 8944 31340 8996 31346
rect 8944 31282 8996 31288
rect 8852 31272 8904 31278
rect 8852 31214 8904 31220
rect 8850 31104 8906 31113
rect 8850 31039 8906 31048
rect 8760 30864 8812 30870
rect 8760 30806 8812 30812
rect 8668 30796 8720 30802
rect 8668 30738 8720 30744
rect 8680 30569 8708 30738
rect 8666 30560 8722 30569
rect 8666 30495 8722 30504
rect 8680 30394 8708 30495
rect 8668 30388 8720 30394
rect 8668 30330 8720 30336
rect 8576 30252 8628 30258
rect 8576 30194 8628 30200
rect 8588 29850 8616 30194
rect 8864 30138 8892 31039
rect 8956 30666 8984 31282
rect 8944 30660 8996 30666
rect 8944 30602 8996 30608
rect 8680 30110 8892 30138
rect 8576 29844 8628 29850
rect 8576 29786 8628 29792
rect 8680 29152 8708 30110
rect 8852 30048 8904 30054
rect 8852 29990 8904 29996
rect 8758 29744 8814 29753
rect 8758 29679 8814 29688
rect 8588 29124 8708 29152
rect 8484 28620 8536 28626
rect 8484 28562 8536 28568
rect 8392 28552 8444 28558
rect 8392 28494 8444 28500
rect 8208 28416 8260 28422
rect 8208 28358 8260 28364
rect 8220 27878 8248 28358
rect 8392 28212 8444 28218
rect 8392 28154 8444 28160
rect 8208 27872 8260 27878
rect 8208 27814 8260 27820
rect 8220 27674 8248 27814
rect 8404 27713 8432 28154
rect 8484 27872 8536 27878
rect 8484 27814 8536 27820
rect 8390 27704 8446 27713
rect 8208 27668 8260 27674
rect 8390 27639 8446 27648
rect 8208 27610 8260 27616
rect 8114 27432 8170 27441
rect 8114 27367 8170 27376
rect 8128 26586 8156 27367
rect 8116 26580 8168 26586
rect 8116 26522 8168 26528
rect 8220 26382 8248 27610
rect 8496 27606 8524 27814
rect 8484 27600 8536 27606
rect 8484 27542 8536 27548
rect 8392 27532 8444 27538
rect 8392 27474 8444 27480
rect 8404 27062 8432 27474
rect 8392 27056 8444 27062
rect 8392 26998 8444 27004
rect 8588 26568 8616 29124
rect 8668 29028 8720 29034
rect 8668 28970 8720 28976
rect 8680 28150 8708 28970
rect 8668 28144 8720 28150
rect 8668 28086 8720 28092
rect 8680 27305 8708 28086
rect 8666 27296 8722 27305
rect 8666 27231 8722 27240
rect 8772 26738 8800 29679
rect 8864 27130 8892 29990
rect 8944 28960 8996 28966
rect 8944 28902 8996 28908
rect 8956 28370 8984 28902
rect 9048 28472 9076 31776
rect 9140 31142 9168 31878
rect 9128 31136 9180 31142
rect 9128 31078 9180 31084
rect 9140 30802 9168 31078
rect 9128 30796 9180 30802
rect 9128 30738 9180 30744
rect 9140 29306 9168 30738
rect 9232 29714 9260 33322
rect 9324 32978 9352 36722
rect 9416 36718 9444 37402
rect 9496 37324 9548 37330
rect 9496 37266 9548 37272
rect 9508 36922 9536 37266
rect 9496 36916 9548 36922
rect 9496 36858 9548 36864
rect 9496 36780 9548 36786
rect 9496 36722 9548 36728
rect 9404 36712 9456 36718
rect 9404 36654 9456 36660
rect 9508 36530 9536 36722
rect 9416 36502 9536 36530
rect 9416 35086 9444 36502
rect 9496 35556 9548 35562
rect 9496 35498 9548 35504
rect 9508 35465 9536 35498
rect 9494 35456 9550 35465
rect 9494 35391 9550 35400
rect 9496 35284 9548 35290
rect 9496 35226 9548 35232
rect 9404 35080 9456 35086
rect 9404 35022 9456 35028
rect 9508 34610 9536 35226
rect 9496 34604 9548 34610
rect 9496 34546 9548 34552
rect 9600 34377 9628 41942
rect 9680 39908 9732 39914
rect 9680 39850 9732 39856
rect 9692 38486 9720 39850
rect 9772 38820 9824 38826
rect 9772 38762 9824 38768
rect 9680 38480 9732 38486
rect 9680 38422 9732 38428
rect 9680 38344 9732 38350
rect 9680 38286 9732 38292
rect 9692 36718 9720 38286
rect 9784 36922 9812 38762
rect 9876 37670 9904 42350
rect 10244 42158 10272 42502
rect 10048 42152 10100 42158
rect 10048 42094 10100 42100
rect 10232 42152 10284 42158
rect 10796 42129 10824 44134
rect 10956 44092 11252 44112
rect 11012 44090 11036 44092
rect 11092 44090 11116 44092
rect 11172 44090 11196 44092
rect 11034 44038 11036 44090
rect 11098 44038 11110 44090
rect 11172 44038 11174 44090
rect 11012 44036 11036 44038
rect 11092 44036 11116 44038
rect 11172 44036 11196 44038
rect 10956 44016 11252 44036
rect 11336 43784 11388 43790
rect 11336 43726 11388 43732
rect 10956 43004 11252 43024
rect 11012 43002 11036 43004
rect 11092 43002 11116 43004
rect 11172 43002 11196 43004
rect 11034 42950 11036 43002
rect 11098 42950 11110 43002
rect 11172 42950 11174 43002
rect 11012 42948 11036 42950
rect 11092 42948 11116 42950
rect 11172 42948 11196 42950
rect 10956 42928 11252 42948
rect 11348 42906 11376 43726
rect 11532 43450 11560 44270
rect 11612 43852 11664 43858
rect 11612 43794 11664 43800
rect 11520 43444 11572 43450
rect 11520 43386 11572 43392
rect 11336 42900 11388 42906
rect 11336 42842 11388 42848
rect 11348 42362 11376 42842
rect 11624 42770 11652 43794
rect 11612 42764 11664 42770
rect 11612 42706 11664 42712
rect 11336 42356 11388 42362
rect 11336 42298 11388 42304
rect 10232 42094 10284 42100
rect 10782 42120 10838 42129
rect 10060 41818 10088 42094
rect 10782 42055 10838 42064
rect 10048 41812 10100 41818
rect 10048 41754 10100 41760
rect 10060 41206 10088 41754
rect 10796 41614 10824 42055
rect 11520 42016 11572 42022
rect 11520 41958 11572 41964
rect 11612 42016 11664 42022
rect 11612 41958 11664 41964
rect 10956 41916 11252 41936
rect 11012 41914 11036 41916
rect 11092 41914 11116 41916
rect 11172 41914 11196 41916
rect 11034 41862 11036 41914
rect 11098 41862 11110 41914
rect 11172 41862 11174 41914
rect 11012 41860 11036 41862
rect 11092 41860 11116 41862
rect 11172 41860 11196 41862
rect 10956 41840 11252 41860
rect 11428 41744 11480 41750
rect 11428 41686 11480 41692
rect 10784 41608 10836 41614
rect 10784 41550 10836 41556
rect 10414 41440 10470 41449
rect 10414 41375 10470 41384
rect 10048 41200 10100 41206
rect 10048 41142 10100 41148
rect 10140 40928 10192 40934
rect 10140 40870 10192 40876
rect 10048 40384 10100 40390
rect 10048 40326 10100 40332
rect 9954 40080 10010 40089
rect 9954 40015 9956 40024
rect 10008 40015 10010 40024
rect 9956 39986 10008 39992
rect 10060 39930 10088 40326
rect 9968 39902 10088 39930
rect 9864 37664 9916 37670
rect 9862 37632 9864 37641
rect 9916 37632 9918 37641
rect 9862 37567 9918 37576
rect 9772 36916 9824 36922
rect 9772 36858 9824 36864
rect 9680 36712 9732 36718
rect 9680 36654 9732 36660
rect 9680 36576 9732 36582
rect 9680 36518 9732 36524
rect 9692 36009 9720 36518
rect 9678 36000 9734 36009
rect 9678 35935 9734 35944
rect 9784 35698 9812 36858
rect 9772 35692 9824 35698
rect 9772 35634 9824 35640
rect 9968 35465 9996 39902
rect 10048 39296 10100 39302
rect 10048 39238 10100 39244
rect 10060 38758 10088 39238
rect 10152 38962 10180 40870
rect 10232 40520 10284 40526
rect 10232 40462 10284 40468
rect 10244 40118 10272 40462
rect 10232 40112 10284 40118
rect 10232 40054 10284 40060
rect 10140 38956 10192 38962
rect 10140 38898 10192 38904
rect 10048 38752 10100 38758
rect 10048 38694 10100 38700
rect 9954 35456 10010 35465
rect 9954 35391 10010 35400
rect 10060 35272 10088 38694
rect 10232 38412 10284 38418
rect 10232 38354 10284 38360
rect 10244 37777 10272 38354
rect 10230 37768 10286 37777
rect 10140 37732 10192 37738
rect 10230 37703 10286 37712
rect 10140 37674 10192 37680
rect 10152 36242 10180 37674
rect 10140 36236 10192 36242
rect 10140 36178 10192 36184
rect 10152 35630 10180 36178
rect 10140 35624 10192 35630
rect 10140 35566 10192 35572
rect 10140 35488 10192 35494
rect 10140 35430 10192 35436
rect 10152 35290 10180 35430
rect 9692 35244 10088 35272
rect 10140 35284 10192 35290
rect 9692 34898 9720 35244
rect 10140 35226 10192 35232
rect 9864 35148 9916 35154
rect 10140 35148 10192 35154
rect 9916 35108 10088 35136
rect 9864 35090 9916 35096
rect 9864 35012 9916 35018
rect 9956 35012 10008 35018
rect 9916 34972 9956 35000
rect 9864 34954 9916 34960
rect 9956 34954 10008 34960
rect 9692 34870 9812 34898
rect 9678 34776 9734 34785
rect 9678 34711 9734 34720
rect 9586 34368 9642 34377
rect 9586 34303 9642 34312
rect 9496 33108 9548 33114
rect 9496 33050 9548 33056
rect 9312 32972 9364 32978
rect 9508 32960 9536 33050
rect 9312 32914 9364 32920
rect 9416 32932 9536 32960
rect 9586 33008 9642 33017
rect 9586 32943 9588 32952
rect 9416 32570 9444 32932
rect 9640 32943 9642 32952
rect 9588 32914 9640 32920
rect 9404 32564 9456 32570
rect 9404 32506 9456 32512
rect 9310 32056 9366 32065
rect 9416 32026 9444 32506
rect 9310 31991 9366 32000
rect 9404 32020 9456 32026
rect 9324 31890 9352 31991
rect 9404 31962 9456 31968
rect 9312 31884 9364 31890
rect 9312 31826 9364 31832
rect 9494 31648 9550 31657
rect 9494 31583 9550 31592
rect 9404 31204 9456 31210
rect 9404 31146 9456 31152
rect 9312 30796 9364 30802
rect 9312 30738 9364 30744
rect 9324 30598 9352 30738
rect 9312 30592 9364 30598
rect 9312 30534 9364 30540
rect 9324 29850 9352 30534
rect 9312 29844 9364 29850
rect 9312 29786 9364 29792
rect 9220 29708 9272 29714
rect 9220 29650 9272 29656
rect 9312 29504 9364 29510
rect 9312 29446 9364 29452
rect 9128 29300 9180 29306
rect 9128 29242 9180 29248
rect 9140 29102 9168 29242
rect 9324 29238 9352 29446
rect 9312 29232 9364 29238
rect 9312 29174 9364 29180
rect 9128 29096 9180 29102
rect 9128 29038 9180 29044
rect 9324 29034 9352 29174
rect 9416 29102 9444 31146
rect 9404 29096 9456 29102
rect 9404 29038 9456 29044
rect 9312 29028 9364 29034
rect 9312 28970 9364 28976
rect 9128 28688 9180 28694
rect 9126 28656 9128 28665
rect 9180 28656 9182 28665
rect 9126 28591 9182 28600
rect 9220 28620 9272 28626
rect 9220 28562 9272 28568
rect 9048 28444 9168 28472
rect 8956 28342 9076 28370
rect 8942 28248 8998 28257
rect 8942 28183 8944 28192
rect 8996 28183 8998 28192
rect 8944 28154 8996 28160
rect 9048 27554 9076 28342
rect 8956 27526 9076 27554
rect 8852 27124 8904 27130
rect 8852 27066 8904 27072
rect 8852 26920 8904 26926
rect 8852 26862 8904 26868
rect 8496 26540 8616 26568
rect 8680 26710 8800 26738
rect 8208 26376 8260 26382
rect 8208 26318 8260 26324
rect 8392 25696 8444 25702
rect 8392 25638 8444 25644
rect 8404 25294 8432 25638
rect 8392 25288 8444 25294
rect 8392 25230 8444 25236
rect 8300 25152 8352 25158
rect 8300 25094 8352 25100
rect 8116 24812 8168 24818
rect 8116 24754 8168 24760
rect 8128 24682 8156 24754
rect 8208 24744 8260 24750
rect 8312 24732 8340 25094
rect 8404 24750 8432 25230
rect 8496 25129 8524 26540
rect 8680 26518 8708 26710
rect 8760 26580 8812 26586
rect 8760 26522 8812 26528
rect 8668 26512 8720 26518
rect 8588 26472 8668 26500
rect 8588 26042 8616 26472
rect 8668 26454 8720 26460
rect 8668 26376 8720 26382
rect 8772 26353 8800 26522
rect 8668 26318 8720 26324
rect 8758 26344 8814 26353
rect 8576 26036 8628 26042
rect 8576 25978 8628 25984
rect 8482 25120 8538 25129
rect 8482 25055 8538 25064
rect 8260 24704 8340 24732
rect 8392 24744 8444 24750
rect 8208 24686 8260 24692
rect 8392 24686 8444 24692
rect 8116 24676 8168 24682
rect 8116 24618 8168 24624
rect 8128 21457 8156 24618
rect 8404 24614 8432 24686
rect 8392 24608 8444 24614
rect 8392 24550 8444 24556
rect 8404 24410 8432 24550
rect 8392 24404 8444 24410
rect 8392 24346 8444 24352
rect 8496 23322 8524 25055
rect 8588 24177 8616 25978
rect 8574 24168 8630 24177
rect 8574 24103 8630 24112
rect 8588 23866 8616 24103
rect 8576 23860 8628 23866
rect 8576 23802 8628 23808
rect 8576 23588 8628 23594
rect 8576 23530 8628 23536
rect 8484 23316 8536 23322
rect 8484 23258 8536 23264
rect 8588 23186 8616 23530
rect 8576 23180 8628 23186
rect 8576 23122 8628 23128
rect 8588 22574 8616 23122
rect 8576 22568 8628 22574
rect 8576 22510 8628 22516
rect 8588 22098 8616 22510
rect 8576 22092 8628 22098
rect 8576 22034 8628 22040
rect 8300 22024 8352 22030
rect 8300 21966 8352 21972
rect 8114 21448 8170 21457
rect 8114 21383 8170 21392
rect 8206 20360 8262 20369
rect 8206 20295 8262 20304
rect 8220 19922 8248 20295
rect 8208 19916 8260 19922
rect 8208 19858 8260 19864
rect 8116 19712 8168 19718
rect 8116 19654 8168 19660
rect 8128 19378 8156 19654
rect 8116 19372 8168 19378
rect 8116 19314 8168 19320
rect 8024 19168 8076 19174
rect 8024 19110 8076 19116
rect 8128 18834 8156 19314
rect 8208 19304 8260 19310
rect 8208 19246 8260 19252
rect 8116 18828 8168 18834
rect 8116 18770 8168 18776
rect 7840 18420 7892 18426
rect 7840 18362 7892 18368
rect 7852 16250 7880 18362
rect 8220 17898 8248 19246
rect 8312 18426 8340 21966
rect 8588 21690 8616 22034
rect 8576 21684 8628 21690
rect 8576 21626 8628 21632
rect 8392 19304 8444 19310
rect 8392 19246 8444 19252
rect 8404 18970 8432 19246
rect 8484 19168 8536 19174
rect 8484 19110 8536 19116
rect 8392 18964 8444 18970
rect 8392 18906 8444 18912
rect 8300 18420 8352 18426
rect 8300 18362 8352 18368
rect 8220 17882 8340 17898
rect 8220 17876 8352 17882
rect 8220 17870 8300 17876
rect 8300 17818 8352 17824
rect 8312 17202 8340 17818
rect 8496 17252 8524 19110
rect 8680 18426 8708 26318
rect 8758 26279 8814 26288
rect 8864 25226 8892 26862
rect 8852 25220 8904 25226
rect 8852 25162 8904 25168
rect 8760 21888 8812 21894
rect 8760 21830 8812 21836
rect 8772 21486 8800 21830
rect 8864 21554 8892 25162
rect 8956 22506 8984 27526
rect 9036 27464 9088 27470
rect 9036 27406 9088 27412
rect 9048 24750 9076 27406
rect 9140 26382 9168 28444
rect 9232 27946 9260 28562
rect 9324 28014 9352 28970
rect 9416 28762 9444 29038
rect 9508 28966 9536 31583
rect 9586 31240 9642 31249
rect 9586 31175 9642 31184
rect 9600 30870 9628 31175
rect 9588 30864 9640 30870
rect 9588 30806 9640 30812
rect 9588 30116 9640 30122
rect 9588 30058 9640 30064
rect 9496 28960 9548 28966
rect 9496 28902 9548 28908
rect 9404 28756 9456 28762
rect 9404 28698 9456 28704
rect 9404 28620 9456 28626
rect 9404 28562 9456 28568
rect 9312 28008 9364 28014
rect 9312 27950 9364 27956
rect 9220 27940 9272 27946
rect 9220 27882 9272 27888
rect 9232 27554 9260 27882
rect 9232 27526 9352 27554
rect 9220 27328 9272 27334
rect 9220 27270 9272 27276
rect 9232 26926 9260 27270
rect 9220 26920 9272 26926
rect 9220 26862 9272 26868
rect 9220 26784 9272 26790
rect 9220 26726 9272 26732
rect 9128 26376 9180 26382
rect 9128 26318 9180 26324
rect 9232 26246 9260 26726
rect 9220 26240 9272 26246
rect 9220 26182 9272 26188
rect 9128 25968 9180 25974
rect 9128 25910 9180 25916
rect 9140 25809 9168 25910
rect 9232 25838 9260 26182
rect 9220 25832 9272 25838
rect 9126 25800 9182 25809
rect 9220 25774 9272 25780
rect 9126 25735 9182 25744
rect 9140 25498 9168 25735
rect 9128 25492 9180 25498
rect 9128 25434 9180 25440
rect 9232 24886 9260 25774
rect 9324 25362 9352 27526
rect 9416 26586 9444 28562
rect 9496 28484 9548 28490
rect 9496 28426 9548 28432
rect 9508 27334 9536 28426
rect 9600 27606 9628 30058
rect 9692 29510 9720 34711
rect 9784 30394 9812 34870
rect 9876 34066 9904 34954
rect 10060 34678 10088 35108
rect 10140 35090 10192 35096
rect 10048 34672 10100 34678
rect 10048 34614 10100 34620
rect 10152 34610 10180 35090
rect 10140 34604 10192 34610
rect 10140 34546 10192 34552
rect 10138 34368 10194 34377
rect 10138 34303 10194 34312
rect 9864 34060 9916 34066
rect 9864 34002 9916 34008
rect 9876 30598 9904 34002
rect 9956 33992 10008 33998
rect 9956 33934 10008 33940
rect 9968 33454 9996 33934
rect 10152 33590 10180 34303
rect 10244 34202 10272 37703
rect 10322 35320 10378 35329
rect 10322 35255 10378 35264
rect 10336 34610 10364 35255
rect 10324 34604 10376 34610
rect 10324 34546 10376 34552
rect 10324 34400 10376 34406
rect 10324 34342 10376 34348
rect 10232 34196 10284 34202
rect 10232 34138 10284 34144
rect 10140 33584 10192 33590
rect 10140 33526 10192 33532
rect 9956 33448 10008 33454
rect 9956 33390 10008 33396
rect 10232 33448 10284 33454
rect 10232 33390 10284 33396
rect 9968 32230 9996 33390
rect 10140 32768 10192 32774
rect 10140 32710 10192 32716
rect 10152 32366 10180 32710
rect 10244 32570 10272 33390
rect 10336 33318 10364 34342
rect 10324 33312 10376 33318
rect 10324 33254 10376 33260
rect 10428 33046 10456 41375
rect 10692 41064 10744 41070
rect 10692 41006 10744 41012
rect 10508 40588 10560 40594
rect 10508 40530 10560 40536
rect 10520 39642 10548 40530
rect 10508 39636 10560 39642
rect 10508 39578 10560 39584
rect 10508 38412 10560 38418
rect 10508 38354 10560 38360
rect 10520 34728 10548 38354
rect 10600 38344 10652 38350
rect 10600 38286 10652 38292
rect 10612 37942 10640 38286
rect 10600 37936 10652 37942
rect 10600 37878 10652 37884
rect 10600 37256 10652 37262
rect 10600 37198 10652 37204
rect 10612 36854 10640 37198
rect 10600 36848 10652 36854
rect 10600 36790 10652 36796
rect 10704 36378 10732 41006
rect 10796 40730 10824 41550
rect 10876 41540 10928 41546
rect 10876 41482 10928 41488
rect 10888 41070 10916 41482
rect 11336 41472 11388 41478
rect 11336 41414 11388 41420
rect 10876 41064 10928 41070
rect 10876 41006 10928 41012
rect 10956 40828 11252 40848
rect 11012 40826 11036 40828
rect 11092 40826 11116 40828
rect 11172 40826 11196 40828
rect 11034 40774 11036 40826
rect 11098 40774 11110 40826
rect 11172 40774 11174 40826
rect 11012 40772 11036 40774
rect 11092 40772 11116 40774
rect 11172 40772 11196 40774
rect 10956 40752 11252 40772
rect 10784 40724 10836 40730
rect 10784 40666 10836 40672
rect 11348 40066 11376 41414
rect 10980 40050 11376 40066
rect 10968 40044 11376 40050
rect 11020 40038 11376 40044
rect 10968 39986 11020 39992
rect 10876 39976 10928 39982
rect 10876 39918 10928 39924
rect 10888 39438 10916 39918
rect 10956 39740 11252 39760
rect 11012 39738 11036 39740
rect 11092 39738 11116 39740
rect 11172 39738 11196 39740
rect 11034 39686 11036 39738
rect 11098 39686 11110 39738
rect 11172 39686 11174 39738
rect 11012 39684 11036 39686
rect 11092 39684 11116 39686
rect 11172 39684 11196 39686
rect 10956 39664 11252 39684
rect 11440 39681 11468 41686
rect 11532 41070 11560 41958
rect 11520 41064 11572 41070
rect 11520 41006 11572 41012
rect 11520 40384 11572 40390
rect 11520 40326 11572 40332
rect 11426 39672 11482 39681
rect 11426 39607 11482 39616
rect 11532 39506 11560 40326
rect 11520 39500 11572 39506
rect 11520 39442 11572 39448
rect 10876 39432 10928 39438
rect 10876 39374 10928 39380
rect 10784 39296 10836 39302
rect 10784 39238 10836 39244
rect 10796 37806 10824 39238
rect 10888 38758 10916 39374
rect 11336 38888 11388 38894
rect 11336 38830 11388 38836
rect 10876 38752 10928 38758
rect 10876 38694 10928 38700
rect 10956 38652 11252 38672
rect 11012 38650 11036 38652
rect 11092 38650 11116 38652
rect 11172 38650 11196 38652
rect 11034 38598 11036 38650
rect 11098 38598 11110 38650
rect 11172 38598 11174 38650
rect 11012 38596 11036 38598
rect 11092 38596 11116 38598
rect 11172 38596 11196 38598
rect 10956 38576 11252 38596
rect 11348 38554 11376 38830
rect 11336 38548 11388 38554
rect 11336 38490 11388 38496
rect 10874 38448 10930 38457
rect 10874 38383 10876 38392
rect 10928 38383 10930 38392
rect 10876 38354 10928 38360
rect 11348 38049 11376 38490
rect 11428 38276 11480 38282
rect 11428 38218 11480 38224
rect 11334 38040 11390 38049
rect 11334 37975 11390 37984
rect 11440 37890 11468 38218
rect 11520 38208 11572 38214
rect 11520 38150 11572 38156
rect 11532 38010 11560 38150
rect 11520 38004 11572 38010
rect 11520 37946 11572 37952
rect 11440 37862 11560 37890
rect 10784 37800 10836 37806
rect 10784 37742 10836 37748
rect 10876 37800 10928 37806
rect 10876 37742 10928 37748
rect 10796 37398 10824 37742
rect 10888 37398 10916 37742
rect 10956 37564 11252 37584
rect 11012 37562 11036 37564
rect 11092 37562 11116 37564
rect 11172 37562 11196 37564
rect 11034 37510 11036 37562
rect 11098 37510 11110 37562
rect 11172 37510 11174 37562
rect 11012 37508 11036 37510
rect 11092 37508 11116 37510
rect 11172 37508 11196 37510
rect 10956 37488 11252 37508
rect 10784 37392 10836 37398
rect 10876 37392 10928 37398
rect 10784 37334 10836 37340
rect 10874 37360 10876 37369
rect 10928 37360 10930 37369
rect 10874 37295 10930 37304
rect 11336 37324 11388 37330
rect 11336 37266 11388 37272
rect 11428 37324 11480 37330
rect 11428 37266 11480 37272
rect 11242 37224 11298 37233
rect 11060 37188 11112 37194
rect 11242 37159 11298 37168
rect 11060 37130 11112 37136
rect 11072 36961 11100 37130
rect 11256 37126 11284 37159
rect 11244 37120 11296 37126
rect 11244 37062 11296 37068
rect 11058 36952 11114 36961
rect 11348 36922 11376 37266
rect 11058 36887 11060 36896
rect 11112 36887 11114 36896
rect 11336 36916 11388 36922
rect 11060 36858 11112 36864
rect 11336 36858 11388 36864
rect 11150 36816 11206 36825
rect 11150 36751 11152 36760
rect 11204 36751 11206 36760
rect 11152 36722 11204 36728
rect 10956 36476 11252 36496
rect 11012 36474 11036 36476
rect 11092 36474 11116 36476
rect 11172 36474 11196 36476
rect 11034 36422 11036 36474
rect 11098 36422 11110 36474
rect 11172 36422 11174 36474
rect 11012 36420 11036 36422
rect 11092 36420 11116 36422
rect 11172 36420 11196 36422
rect 10956 36400 11252 36420
rect 10692 36372 10744 36378
rect 10692 36314 10744 36320
rect 10876 36304 10928 36310
rect 10876 36246 10928 36252
rect 10600 36236 10652 36242
rect 10600 36178 10652 36184
rect 10692 36236 10744 36242
rect 10692 36178 10744 36184
rect 10612 35290 10640 36178
rect 10600 35284 10652 35290
rect 10600 35226 10652 35232
rect 10600 35080 10652 35086
rect 10598 35048 10600 35057
rect 10652 35048 10654 35057
rect 10598 34983 10654 34992
rect 10704 34921 10732 36178
rect 10784 35556 10836 35562
rect 10784 35498 10836 35504
rect 10796 35290 10824 35498
rect 10784 35284 10836 35290
rect 10784 35226 10836 35232
rect 10690 34912 10746 34921
rect 10690 34847 10746 34856
rect 10520 34700 10640 34728
rect 10506 34640 10562 34649
rect 10506 34575 10562 34584
rect 10520 34542 10548 34575
rect 10508 34536 10560 34542
rect 10508 34478 10560 34484
rect 10506 34232 10562 34241
rect 10506 34167 10508 34176
rect 10560 34167 10562 34176
rect 10508 34138 10560 34144
rect 10508 33448 10560 33454
rect 10508 33390 10560 33396
rect 10520 33046 10548 33390
rect 10416 33040 10468 33046
rect 10322 33008 10378 33017
rect 10416 32982 10468 32988
rect 10508 33040 10560 33046
rect 10508 32982 10560 32988
rect 10322 32943 10324 32952
rect 10376 32943 10378 32952
rect 10324 32914 10376 32920
rect 10232 32564 10284 32570
rect 10232 32506 10284 32512
rect 10140 32360 10192 32366
rect 10140 32302 10192 32308
rect 10232 32360 10284 32366
rect 10232 32302 10284 32308
rect 9956 32224 10008 32230
rect 9956 32166 10008 32172
rect 10140 32224 10192 32230
rect 10140 32166 10192 32172
rect 9968 31890 9996 32166
rect 10046 32056 10102 32065
rect 10046 31991 10048 32000
rect 10100 31991 10102 32000
rect 10048 31962 10100 31968
rect 9956 31884 10008 31890
rect 10008 31844 10088 31872
rect 9956 31826 10008 31832
rect 10060 31278 10088 31844
rect 10048 31272 10100 31278
rect 10048 31214 10100 31220
rect 9956 31204 10008 31210
rect 9956 31146 10008 31152
rect 9968 31113 9996 31146
rect 9954 31104 10010 31113
rect 9954 31039 10010 31048
rect 9954 30832 10010 30841
rect 10060 30802 10088 31214
rect 9954 30767 10010 30776
rect 10048 30796 10100 30802
rect 9968 30734 9996 30767
rect 10048 30738 10100 30744
rect 9956 30728 10008 30734
rect 9956 30670 10008 30676
rect 9864 30592 9916 30598
rect 9864 30534 9916 30540
rect 9968 30410 9996 30670
rect 10152 30410 10180 32166
rect 10244 31521 10272 32302
rect 10336 32026 10364 32914
rect 10612 32450 10640 34700
rect 10428 32422 10640 32450
rect 10704 32450 10732 34847
rect 10784 34468 10836 34474
rect 10784 34410 10836 34416
rect 10796 33454 10824 34410
rect 10888 34134 10916 36246
rect 11060 36100 11112 36106
rect 11060 36042 11112 36048
rect 11072 35562 11100 36042
rect 11440 35986 11468 37266
rect 11348 35958 11468 35986
rect 11348 35698 11376 35958
rect 11426 35864 11482 35873
rect 11426 35799 11482 35808
rect 11336 35692 11388 35698
rect 11336 35634 11388 35640
rect 11060 35556 11112 35562
rect 11060 35498 11112 35504
rect 11348 35494 11376 35634
rect 11440 35562 11468 35799
rect 11428 35556 11480 35562
rect 11428 35498 11480 35504
rect 11336 35488 11388 35494
rect 11336 35430 11388 35436
rect 10956 35388 11252 35408
rect 11012 35386 11036 35388
rect 11092 35386 11116 35388
rect 11172 35386 11196 35388
rect 11034 35334 11036 35386
rect 11098 35334 11110 35386
rect 11172 35334 11174 35386
rect 11012 35332 11036 35334
rect 11092 35332 11116 35334
rect 11172 35332 11196 35334
rect 10956 35312 11252 35332
rect 11244 35216 11296 35222
rect 11244 35158 11296 35164
rect 11256 34746 11284 35158
rect 11348 34762 11376 35430
rect 11440 34950 11468 35498
rect 11428 34944 11480 34950
rect 11428 34886 11480 34892
rect 11244 34740 11296 34746
rect 11348 34734 11468 34762
rect 11244 34682 11296 34688
rect 11336 34672 11388 34678
rect 11336 34614 11388 34620
rect 10956 34300 11252 34320
rect 11012 34298 11036 34300
rect 11092 34298 11116 34300
rect 11172 34298 11196 34300
rect 11034 34246 11036 34298
rect 11098 34246 11110 34298
rect 11172 34246 11174 34298
rect 11012 34244 11036 34246
rect 11092 34244 11116 34246
rect 11172 34244 11196 34246
rect 10956 34224 11252 34244
rect 10876 34128 10928 34134
rect 10876 34070 10928 34076
rect 10968 33992 11020 33998
rect 10968 33934 11020 33940
rect 10876 33652 10928 33658
rect 10876 33594 10928 33600
rect 10784 33448 10836 33454
rect 10784 33390 10836 33396
rect 10796 33289 10824 33390
rect 10782 33280 10838 33289
rect 10782 33215 10838 33224
rect 10784 32904 10836 32910
rect 10784 32846 10836 32852
rect 10796 32609 10824 32846
rect 10782 32600 10838 32609
rect 10782 32535 10838 32544
rect 10704 32422 10824 32450
rect 10324 32020 10376 32026
rect 10324 31962 10376 31968
rect 10324 31884 10376 31890
rect 10324 31826 10376 31832
rect 10336 31634 10364 31826
rect 10428 31736 10456 32422
rect 10600 32360 10652 32366
rect 10600 32302 10652 32308
rect 10506 31920 10562 31929
rect 10612 31906 10640 32302
rect 10562 31878 10640 31906
rect 10506 31855 10508 31864
rect 10560 31855 10562 31864
rect 10508 31826 10560 31832
rect 10428 31708 10640 31736
rect 10336 31606 10456 31634
rect 10230 31512 10286 31521
rect 10286 31470 10364 31498
rect 10230 31447 10286 31456
rect 10336 30841 10364 31470
rect 10428 30938 10456 31606
rect 10612 31464 10640 31708
rect 10612 31436 10732 31464
rect 10600 31340 10652 31346
rect 10600 31282 10652 31288
rect 10508 31272 10560 31278
rect 10506 31240 10508 31249
rect 10560 31240 10562 31249
rect 10506 31175 10562 31184
rect 10416 30932 10468 30938
rect 10416 30874 10468 30880
rect 10322 30832 10378 30841
rect 10322 30767 10378 30776
rect 10232 30592 10284 30598
rect 10232 30534 10284 30540
rect 9772 30388 9824 30394
rect 9772 30330 9824 30336
rect 9876 30382 9996 30410
rect 10060 30382 10180 30410
rect 9876 30274 9904 30382
rect 9784 30246 9904 30274
rect 9956 30320 10008 30326
rect 9956 30262 10008 30268
rect 9680 29504 9732 29510
rect 9680 29446 9732 29452
rect 9784 29322 9812 30246
rect 9864 29640 9916 29646
rect 9864 29582 9916 29588
rect 9692 29294 9812 29322
rect 9692 28762 9720 29294
rect 9772 28960 9824 28966
rect 9772 28902 9824 28908
rect 9680 28756 9732 28762
rect 9680 28698 9732 28704
rect 9678 28520 9734 28529
rect 9678 28455 9734 28464
rect 9692 28014 9720 28455
rect 9784 28422 9812 28902
rect 9772 28416 9824 28422
rect 9772 28358 9824 28364
rect 9680 28008 9732 28014
rect 9680 27950 9732 27956
rect 9784 27946 9812 28358
rect 9876 28150 9904 29582
rect 9864 28144 9916 28150
rect 9864 28086 9916 28092
rect 9772 27940 9824 27946
rect 9772 27882 9824 27888
rect 9864 27940 9916 27946
rect 9864 27882 9916 27888
rect 9680 27872 9732 27878
rect 9680 27814 9732 27820
rect 9770 27840 9826 27849
rect 9588 27600 9640 27606
rect 9588 27542 9640 27548
rect 9496 27328 9548 27334
rect 9496 27270 9548 27276
rect 9588 26920 9640 26926
rect 9588 26862 9640 26868
rect 9600 26790 9628 26862
rect 9588 26784 9640 26790
rect 9588 26726 9640 26732
rect 9404 26580 9456 26586
rect 9404 26522 9456 26528
rect 9404 26376 9456 26382
rect 9404 26318 9456 26324
rect 9312 25356 9364 25362
rect 9312 25298 9364 25304
rect 9416 24970 9444 26318
rect 9588 26240 9640 26246
rect 9588 26182 9640 26188
rect 9600 25498 9628 26182
rect 9588 25492 9640 25498
rect 9588 25434 9640 25440
rect 9588 25356 9640 25362
rect 9588 25298 9640 25304
rect 9324 24942 9444 24970
rect 9220 24880 9272 24886
rect 9220 24822 9272 24828
rect 9036 24744 9088 24750
rect 9036 24686 9088 24692
rect 9048 24342 9076 24686
rect 9036 24336 9088 24342
rect 9036 24278 9088 24284
rect 8944 22500 8996 22506
rect 8944 22442 8996 22448
rect 8942 21584 8998 21593
rect 8852 21548 8904 21554
rect 8942 21519 8998 21528
rect 8852 21490 8904 21496
rect 8956 21486 8984 21519
rect 8760 21480 8812 21486
rect 8760 21422 8812 21428
rect 8944 21480 8996 21486
rect 8944 21422 8996 21428
rect 8956 21146 8984 21422
rect 8944 21140 8996 21146
rect 8944 21082 8996 21088
rect 9048 21026 9076 24278
rect 9324 23338 9352 24942
rect 8864 20998 9076 21026
rect 9140 23310 9352 23338
rect 8668 18420 8720 18426
rect 8668 18362 8720 18368
rect 8576 17264 8628 17270
rect 8496 17224 8576 17252
rect 8300 17196 8352 17202
rect 8300 17138 8352 17144
rect 7840 16244 7892 16250
rect 7840 16186 7892 16192
rect 7852 16046 7880 16186
rect 7840 16040 7892 16046
rect 7840 15982 7892 15988
rect 7852 15162 7880 15982
rect 8114 15600 8170 15609
rect 8114 15535 8170 15544
rect 7840 15156 7892 15162
rect 7840 15098 7892 15104
rect 7852 14958 7880 15098
rect 7840 14952 7892 14958
rect 7840 14894 7892 14900
rect 8128 14414 8156 15535
rect 8312 14482 8340 17138
rect 8496 16794 8524 17224
rect 8576 17206 8628 17212
rect 8484 16788 8536 16794
rect 8484 16730 8536 16736
rect 8300 14476 8352 14482
rect 8300 14418 8352 14424
rect 8116 14408 8168 14414
rect 8116 14350 8168 14356
rect 8128 14006 8156 14350
rect 8116 14000 8168 14006
rect 8116 13942 8168 13948
rect 8312 13938 8340 14418
rect 8496 14414 8524 16730
rect 8666 16008 8722 16017
rect 8666 15943 8722 15952
rect 8680 15638 8708 15943
rect 8668 15632 8720 15638
rect 8668 15574 8720 15580
rect 8576 14816 8628 14822
rect 8576 14758 8628 14764
rect 8588 14618 8616 14758
rect 8576 14612 8628 14618
rect 8576 14554 8628 14560
rect 8588 14482 8616 14554
rect 8576 14476 8628 14482
rect 8576 14418 8628 14424
rect 8484 14408 8536 14414
rect 8484 14350 8536 14356
rect 8496 14074 8524 14350
rect 8760 14340 8812 14346
rect 8760 14282 8812 14288
rect 8484 14068 8536 14074
rect 8484 14010 8536 14016
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8312 13530 8340 13874
rect 8392 13864 8444 13870
rect 8392 13806 8444 13812
rect 8300 13524 8352 13530
rect 8300 13466 8352 13472
rect 8404 13297 8432 13806
rect 8496 13462 8524 14010
rect 8772 13870 8800 14282
rect 8760 13864 8812 13870
rect 8760 13806 8812 13812
rect 8484 13456 8536 13462
rect 8484 13398 8536 13404
rect 8390 13288 8446 13297
rect 8390 13223 8446 13232
rect 8668 12776 8720 12782
rect 8668 12718 8720 12724
rect 8680 12102 8708 12718
rect 7932 12096 7984 12102
rect 7932 12038 7984 12044
rect 8668 12096 8720 12102
rect 8668 12038 8720 12044
rect 7840 11212 7892 11218
rect 7840 11154 7892 11160
rect 7852 10810 7880 11154
rect 7944 11082 7972 12038
rect 7932 11076 7984 11082
rect 7932 11018 7984 11024
rect 7840 10804 7892 10810
rect 7840 10746 7892 10752
rect 7944 9081 7972 11018
rect 7930 9072 7986 9081
rect 7930 9007 7986 9016
rect 8864 8634 8892 20998
rect 8944 19916 8996 19922
rect 8944 19858 8996 19864
rect 8956 19553 8984 19858
rect 8942 19544 8998 19553
rect 8942 19479 8944 19488
rect 8996 19479 8998 19488
rect 8944 19450 8996 19456
rect 8944 19304 8996 19310
rect 8944 19246 8996 19252
rect 9034 19272 9090 19281
rect 8956 17202 8984 19246
rect 9140 19258 9168 23310
rect 9218 23216 9274 23225
rect 9218 23151 9274 23160
rect 9090 19230 9168 19258
rect 9034 19207 9090 19216
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 8956 16998 8984 17138
rect 8944 16992 8996 16998
rect 8944 16934 8996 16940
rect 9128 14272 9180 14278
rect 9128 14214 9180 14220
rect 9140 13870 9168 14214
rect 9128 13864 9180 13870
rect 9128 13806 9180 13812
rect 9232 13802 9260 23151
rect 9496 23112 9548 23118
rect 9496 23054 9548 23060
rect 9404 22500 9456 22506
rect 9404 22442 9456 22448
rect 9310 20360 9366 20369
rect 9310 20295 9366 20304
rect 9324 19310 9352 20295
rect 9312 19304 9364 19310
rect 9312 19246 9364 19252
rect 9312 18284 9364 18290
rect 9312 18226 9364 18232
rect 9324 17882 9352 18226
rect 9312 17876 9364 17882
rect 9312 17818 9364 17824
rect 9324 16726 9352 17818
rect 9416 17338 9444 22442
rect 9508 22438 9536 23054
rect 9496 22432 9548 22438
rect 9496 22374 9548 22380
rect 9508 22234 9536 22374
rect 9496 22228 9548 22234
rect 9496 22170 9548 22176
rect 9496 21480 9548 21486
rect 9496 21422 9548 21428
rect 9508 21146 9536 21422
rect 9496 21140 9548 21146
rect 9496 21082 9548 21088
rect 9494 20632 9550 20641
rect 9494 20567 9496 20576
rect 9548 20567 9550 20576
rect 9496 20538 9548 20544
rect 9508 19378 9536 20538
rect 9496 19372 9548 19378
rect 9496 19314 9548 19320
rect 9496 19236 9548 19242
rect 9496 19178 9548 19184
rect 9508 18630 9536 19178
rect 9496 18624 9548 18630
rect 9496 18566 9548 18572
rect 9600 18306 9628 25298
rect 9692 24290 9720 27814
rect 9770 27775 9826 27784
rect 9784 24818 9812 27775
rect 9876 25378 9904 27882
rect 9968 26518 9996 30262
rect 10060 30190 10088 30382
rect 10048 30184 10100 30190
rect 10048 30126 10100 30132
rect 10060 29782 10088 30126
rect 10140 30048 10192 30054
rect 10138 30016 10140 30025
rect 10192 30016 10194 30025
rect 10138 29951 10194 29960
rect 10048 29776 10100 29782
rect 10048 29718 10100 29724
rect 10138 29744 10194 29753
rect 10138 29679 10194 29688
rect 10152 29646 10180 29679
rect 10140 29640 10192 29646
rect 10140 29582 10192 29588
rect 10152 29073 10180 29582
rect 10138 29064 10194 29073
rect 10138 28999 10194 29008
rect 10046 28384 10102 28393
rect 10046 28319 10102 28328
rect 10060 28014 10088 28319
rect 10048 28008 10100 28014
rect 10048 27950 10100 27956
rect 10060 27554 10088 27950
rect 10152 27946 10180 28999
rect 10140 27940 10192 27946
rect 10140 27882 10192 27888
rect 10060 27526 10180 27554
rect 10152 26772 10180 27526
rect 10060 26744 10180 26772
rect 9956 26512 10008 26518
rect 9956 26454 10008 26460
rect 9968 25498 9996 26454
rect 9956 25492 10008 25498
rect 9956 25434 10008 25440
rect 9876 25350 9996 25378
rect 10060 25362 10088 26744
rect 10140 25968 10192 25974
rect 10140 25910 10192 25916
rect 9864 25288 9916 25294
rect 9864 25230 9916 25236
rect 9772 24812 9824 24818
rect 9772 24754 9824 24760
rect 9784 24410 9812 24754
rect 9772 24404 9824 24410
rect 9772 24346 9824 24352
rect 9692 24262 9812 24290
rect 9680 23860 9732 23866
rect 9680 23802 9732 23808
rect 9692 20505 9720 23802
rect 9784 22953 9812 24262
rect 9770 22944 9826 22953
rect 9770 22879 9826 22888
rect 9876 21570 9904 25230
rect 9968 24614 9996 25350
rect 10048 25356 10100 25362
rect 10048 25298 10100 25304
rect 10046 25256 10102 25265
rect 10046 25191 10102 25200
rect 9956 24608 10008 24614
rect 9956 24550 10008 24556
rect 9956 23112 10008 23118
rect 9956 23054 10008 23060
rect 9968 22778 9996 23054
rect 9956 22772 10008 22778
rect 9956 22714 10008 22720
rect 10060 22438 10088 25191
rect 10152 24750 10180 25910
rect 10140 24744 10192 24750
rect 10140 24686 10192 24692
rect 10140 24608 10192 24614
rect 10140 24550 10192 24556
rect 10048 22432 10100 22438
rect 10048 22374 10100 22380
rect 9956 22024 10008 22030
rect 9954 21992 9956 22001
rect 10008 21992 10010 22001
rect 9954 21927 10010 21936
rect 9968 21690 9996 21927
rect 9956 21684 10008 21690
rect 9956 21626 10008 21632
rect 9876 21542 9996 21570
rect 9862 21448 9918 21457
rect 9862 21383 9918 21392
rect 9876 21146 9904 21383
rect 9864 21140 9916 21146
rect 9864 21082 9916 21088
rect 9864 21004 9916 21010
rect 9864 20946 9916 20952
rect 9678 20496 9734 20505
rect 9678 20431 9734 20440
rect 9876 20262 9904 20946
rect 9864 20256 9916 20262
rect 9678 20224 9734 20233
rect 9864 20198 9916 20204
rect 9678 20159 9734 20168
rect 9508 18278 9628 18306
rect 9692 18290 9720 20159
rect 9770 19272 9826 19281
rect 9770 19207 9826 19216
rect 9784 19174 9812 19207
rect 9772 19168 9824 19174
rect 9772 19110 9824 19116
rect 9680 18284 9732 18290
rect 9404 17332 9456 17338
rect 9404 17274 9456 17280
rect 9508 17252 9536 18278
rect 9680 18226 9732 18232
rect 9588 18216 9640 18222
rect 9640 18164 9720 18170
rect 9588 18158 9720 18164
rect 9600 18142 9720 18158
rect 9692 17814 9720 18142
rect 9680 17808 9732 17814
rect 9586 17776 9642 17785
rect 9680 17750 9732 17756
rect 9586 17711 9642 17720
rect 9600 17678 9628 17711
rect 9588 17672 9640 17678
rect 9588 17614 9640 17620
rect 9680 17264 9732 17270
rect 9508 17224 9680 17252
rect 9680 17206 9732 17212
rect 9494 17096 9550 17105
rect 9494 17031 9550 17040
rect 9680 17060 9732 17066
rect 9508 16794 9536 17031
rect 9680 17002 9732 17008
rect 9496 16788 9548 16794
rect 9496 16730 9548 16736
rect 9312 16720 9364 16726
rect 9312 16662 9364 16668
rect 9692 16250 9720 17002
rect 9772 16992 9824 16998
rect 9772 16934 9824 16940
rect 9680 16244 9732 16250
rect 9680 16186 9732 16192
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 9600 14482 9628 15982
rect 9784 14618 9812 16934
rect 9876 14958 9904 20198
rect 9968 19242 9996 21542
rect 10060 21010 10088 22374
rect 10048 21004 10100 21010
rect 10048 20946 10100 20952
rect 10048 20800 10100 20806
rect 10048 20742 10100 20748
rect 9956 19236 10008 19242
rect 9956 19178 10008 19184
rect 9968 18970 9996 19178
rect 10060 19174 10088 20742
rect 10152 20602 10180 24550
rect 10244 24342 10272 30534
rect 10428 29866 10456 30874
rect 10520 30258 10548 31175
rect 10508 30252 10560 30258
rect 10508 30194 10560 30200
rect 10336 29838 10456 29866
rect 10336 28082 10364 29838
rect 10416 29640 10468 29646
rect 10416 29582 10468 29588
rect 10428 29170 10456 29582
rect 10508 29232 10560 29238
rect 10508 29174 10560 29180
rect 10416 29164 10468 29170
rect 10416 29106 10468 29112
rect 10416 28484 10468 28490
rect 10416 28426 10468 28432
rect 10324 28076 10376 28082
rect 10324 28018 10376 28024
rect 10428 27538 10456 28426
rect 10416 27532 10468 27538
rect 10416 27474 10468 27480
rect 10428 27441 10456 27474
rect 10414 27432 10470 27441
rect 10324 27396 10376 27402
rect 10414 27367 10470 27376
rect 10324 27338 10376 27344
rect 10336 26450 10364 27338
rect 10520 26450 10548 29174
rect 10324 26444 10376 26450
rect 10324 26386 10376 26392
rect 10508 26444 10560 26450
rect 10508 26386 10560 26392
rect 10336 26217 10364 26386
rect 10612 26382 10640 31282
rect 10704 29102 10732 31436
rect 10692 29096 10744 29102
rect 10692 29038 10744 29044
rect 10690 28792 10746 28801
rect 10690 28727 10746 28736
rect 10704 28529 10732 28727
rect 10690 28520 10746 28529
rect 10690 28455 10746 28464
rect 10692 28008 10744 28014
rect 10692 27950 10744 27956
rect 10416 26376 10468 26382
rect 10416 26318 10468 26324
rect 10600 26376 10652 26382
rect 10600 26318 10652 26324
rect 10322 26208 10378 26217
rect 10322 26143 10378 26152
rect 10322 25936 10378 25945
rect 10322 25871 10378 25880
rect 10232 24336 10284 24342
rect 10232 24278 10284 24284
rect 10336 23866 10364 25871
rect 10324 23860 10376 23866
rect 10324 23802 10376 23808
rect 10322 21720 10378 21729
rect 10322 21655 10378 21664
rect 10336 21350 10364 21655
rect 10324 21344 10376 21350
rect 10324 21286 10376 21292
rect 10140 20596 10192 20602
rect 10140 20538 10192 20544
rect 10232 20596 10284 20602
rect 10232 20538 10284 20544
rect 10244 19553 10272 20538
rect 10324 20324 10376 20330
rect 10324 20266 10376 20272
rect 10336 20058 10364 20266
rect 10324 20052 10376 20058
rect 10324 19994 10376 20000
rect 10230 19544 10286 19553
rect 10230 19479 10286 19488
rect 10336 19378 10364 19994
rect 10324 19372 10376 19378
rect 10324 19314 10376 19320
rect 10232 19304 10284 19310
rect 10232 19246 10284 19252
rect 10048 19168 10100 19174
rect 10048 19110 10100 19116
rect 9956 18964 10008 18970
rect 9956 18906 10008 18912
rect 9968 18426 9996 18906
rect 10244 18630 10272 19246
rect 10232 18624 10284 18630
rect 10232 18566 10284 18572
rect 9956 18420 10008 18426
rect 9956 18362 10008 18368
rect 9968 17338 9996 18362
rect 10244 18290 10272 18566
rect 10232 18284 10284 18290
rect 10232 18226 10284 18232
rect 10324 18284 10376 18290
rect 10324 18226 10376 18232
rect 10336 17678 10364 18226
rect 10324 17672 10376 17678
rect 10324 17614 10376 17620
rect 9956 17332 10008 17338
rect 9956 17274 10008 17280
rect 10232 17264 10284 17270
rect 10232 17206 10284 17212
rect 10140 17128 10192 17134
rect 10140 17070 10192 17076
rect 10152 16046 10180 17070
rect 10140 16040 10192 16046
rect 10140 15982 10192 15988
rect 10048 15700 10100 15706
rect 10048 15642 10100 15648
rect 10060 15609 10088 15642
rect 10046 15600 10102 15609
rect 10046 15535 10102 15544
rect 9864 14952 9916 14958
rect 9864 14894 9916 14900
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9588 14476 9640 14482
rect 9588 14418 9640 14424
rect 9496 14340 9548 14346
rect 9496 14282 9548 14288
rect 8944 13796 8996 13802
rect 8944 13738 8996 13744
rect 9220 13796 9272 13802
rect 9220 13738 9272 13744
rect 8956 12850 8984 13738
rect 8944 12844 8996 12850
rect 8944 12786 8996 12792
rect 8956 11898 8984 12786
rect 9508 11898 9536 14282
rect 9784 13297 9812 14554
rect 9770 13288 9826 13297
rect 9770 13223 9826 13232
rect 9876 12306 9904 14894
rect 10244 14482 10272 17206
rect 10336 16794 10364 17614
rect 10324 16788 10376 16794
rect 10324 16730 10376 16736
rect 10428 16130 10456 26318
rect 10612 25974 10640 26318
rect 10704 26042 10732 27950
rect 10692 26036 10744 26042
rect 10692 25978 10744 25984
rect 10600 25968 10652 25974
rect 10600 25910 10652 25916
rect 10692 25696 10744 25702
rect 10690 25664 10692 25673
rect 10744 25664 10746 25673
rect 10690 25599 10746 25608
rect 10692 25492 10744 25498
rect 10692 25434 10744 25440
rect 10508 25356 10560 25362
rect 10508 25298 10560 25304
rect 10520 24954 10548 25298
rect 10600 25152 10652 25158
rect 10600 25094 10652 25100
rect 10508 24948 10560 24954
rect 10508 24890 10560 24896
rect 10612 24818 10640 25094
rect 10600 24812 10652 24818
rect 10600 24754 10652 24760
rect 10508 24608 10560 24614
rect 10508 24550 10560 24556
rect 10520 18873 10548 24550
rect 10598 22536 10654 22545
rect 10598 22471 10654 22480
rect 10612 21486 10640 22471
rect 10600 21480 10652 21486
rect 10600 21422 10652 21428
rect 10600 21344 10652 21350
rect 10600 21286 10652 21292
rect 10612 20806 10640 21286
rect 10600 20800 10652 20806
rect 10600 20742 10652 20748
rect 10704 20618 10732 25434
rect 10796 23254 10824 32422
rect 10888 30938 10916 33594
rect 10980 33590 11008 33934
rect 10968 33584 11020 33590
rect 10968 33526 11020 33532
rect 10956 33212 11252 33232
rect 11012 33210 11036 33212
rect 11092 33210 11116 33212
rect 11172 33210 11196 33212
rect 11034 33158 11036 33210
rect 11098 33158 11110 33210
rect 11172 33158 11174 33210
rect 11012 33156 11036 33158
rect 11092 33156 11116 33158
rect 11172 33156 11196 33158
rect 10956 33136 11252 33156
rect 11242 32464 11298 32473
rect 11242 32399 11298 32408
rect 11256 32366 11284 32399
rect 11244 32360 11296 32366
rect 11244 32302 11296 32308
rect 10956 32124 11252 32144
rect 11012 32122 11036 32124
rect 11092 32122 11116 32124
rect 11172 32122 11196 32124
rect 11034 32070 11036 32122
rect 11098 32070 11110 32122
rect 11172 32070 11174 32122
rect 11012 32068 11036 32070
rect 11092 32068 11116 32070
rect 11172 32068 11196 32070
rect 10956 32048 11252 32068
rect 10968 31952 11020 31958
rect 10968 31894 11020 31900
rect 11150 31920 11206 31929
rect 10980 31278 11008 31894
rect 11150 31855 11206 31864
rect 11164 31346 11192 31855
rect 11244 31816 11296 31822
rect 11244 31758 11296 31764
rect 11152 31340 11204 31346
rect 11152 31282 11204 31288
rect 10968 31272 11020 31278
rect 11256 31249 11284 31758
rect 10968 31214 11020 31220
rect 11242 31240 11298 31249
rect 11242 31175 11298 31184
rect 10956 31036 11252 31056
rect 11012 31034 11036 31036
rect 11092 31034 11116 31036
rect 11172 31034 11196 31036
rect 11034 30982 11036 31034
rect 11098 30982 11110 31034
rect 11172 30982 11174 31034
rect 11012 30980 11036 30982
rect 11092 30980 11116 30982
rect 11172 30980 11196 30982
rect 10956 30960 11252 30980
rect 10876 30932 10928 30938
rect 10876 30874 10928 30880
rect 10888 30394 10916 30874
rect 10968 30864 11020 30870
rect 10966 30832 10968 30841
rect 11020 30832 11022 30841
rect 10966 30767 11022 30776
rect 10968 30728 11020 30734
rect 10968 30670 11020 30676
rect 10876 30388 10928 30394
rect 10876 30330 10928 30336
rect 10980 30274 11008 30670
rect 10888 30246 11008 30274
rect 10888 29492 10916 30246
rect 10956 29948 11252 29968
rect 11012 29946 11036 29948
rect 11092 29946 11116 29948
rect 11172 29946 11196 29948
rect 11034 29894 11036 29946
rect 11098 29894 11110 29946
rect 11172 29894 11174 29946
rect 11012 29892 11036 29894
rect 11092 29892 11116 29894
rect 11172 29892 11196 29894
rect 10956 29872 11252 29892
rect 11060 29504 11112 29510
rect 10888 29464 11060 29492
rect 11060 29446 11112 29452
rect 10874 29200 10930 29209
rect 11072 29170 11100 29446
rect 10874 29135 10930 29144
rect 11060 29164 11112 29170
rect 10888 29102 10916 29135
rect 11060 29106 11112 29112
rect 10876 29096 10928 29102
rect 10876 29038 10928 29044
rect 10876 28960 10928 28966
rect 10876 28902 10928 28908
rect 10888 28121 10916 28902
rect 10956 28860 11252 28880
rect 11012 28858 11036 28860
rect 11092 28858 11116 28860
rect 11172 28858 11196 28860
rect 11034 28806 11036 28858
rect 11098 28806 11110 28858
rect 11172 28806 11174 28858
rect 11012 28804 11036 28806
rect 11092 28804 11116 28806
rect 11172 28804 11196 28806
rect 10956 28784 11252 28804
rect 10874 28112 10930 28121
rect 10874 28047 10930 28056
rect 10874 27976 10930 27985
rect 10874 27911 10930 27920
rect 10888 27316 10916 27911
rect 10956 27772 11252 27792
rect 11012 27770 11036 27772
rect 11092 27770 11116 27772
rect 11172 27770 11196 27772
rect 11034 27718 11036 27770
rect 11098 27718 11110 27770
rect 11172 27718 11174 27770
rect 11012 27716 11036 27718
rect 11092 27716 11116 27718
rect 11172 27716 11196 27718
rect 10956 27696 11252 27716
rect 11060 27600 11112 27606
rect 11060 27542 11112 27548
rect 10968 27328 11020 27334
rect 10888 27288 10968 27316
rect 10888 27130 10916 27288
rect 10968 27270 11020 27276
rect 10876 27124 10928 27130
rect 10876 27066 10928 27072
rect 11072 26926 11100 27542
rect 11060 26920 11112 26926
rect 11060 26862 11112 26868
rect 10956 26684 11252 26704
rect 11012 26682 11036 26684
rect 11092 26682 11116 26684
rect 11172 26682 11196 26684
rect 11034 26630 11036 26682
rect 11098 26630 11110 26682
rect 11172 26630 11174 26682
rect 11012 26628 11036 26630
rect 11092 26628 11116 26630
rect 11172 26628 11196 26630
rect 10956 26608 11252 26628
rect 11244 26376 11296 26382
rect 11242 26344 11244 26353
rect 11296 26344 11298 26353
rect 11242 26279 11298 26288
rect 10876 26240 10928 26246
rect 10876 26182 10928 26188
rect 10888 25770 10916 26182
rect 11244 26036 11296 26042
rect 11244 25978 11296 25984
rect 11150 25936 11206 25945
rect 11150 25871 11206 25880
rect 11164 25770 11192 25871
rect 11256 25809 11284 25978
rect 11242 25800 11298 25809
rect 10876 25764 10928 25770
rect 10876 25706 10928 25712
rect 11152 25764 11204 25770
rect 11242 25735 11298 25744
rect 11152 25706 11204 25712
rect 10888 25498 10916 25706
rect 10956 25596 11252 25616
rect 11012 25594 11036 25596
rect 11092 25594 11116 25596
rect 11172 25594 11196 25596
rect 11034 25542 11036 25594
rect 11098 25542 11110 25594
rect 11172 25542 11174 25594
rect 11012 25540 11036 25542
rect 11092 25540 11116 25542
rect 11172 25540 11196 25542
rect 10956 25520 11252 25540
rect 11348 25498 11376 34614
rect 11440 34066 11468 34734
rect 11428 34060 11480 34066
rect 11428 34002 11480 34008
rect 11428 32768 11480 32774
rect 11428 32710 11480 32716
rect 11440 31521 11468 32710
rect 11532 31657 11560 37862
rect 11624 34678 11652 41958
rect 11716 41313 11744 49710
rect 11808 49298 11836 50118
rect 11992 49609 12020 51206
rect 11978 49600 12034 49609
rect 11978 49535 12034 49544
rect 11796 49292 11848 49298
rect 11796 49234 11848 49240
rect 11808 48890 11836 49234
rect 11796 48884 11848 48890
rect 11796 48826 11848 48832
rect 12084 48657 12112 52838
rect 12268 52822 12388 52850
rect 12268 52714 12296 52822
rect 12176 52686 12296 52714
rect 12176 52034 12204 52686
rect 12254 52592 12310 52601
rect 12254 52527 12256 52536
rect 12308 52527 12310 52536
rect 12256 52498 12308 52504
rect 12268 52154 12296 52498
rect 12440 52488 12492 52494
rect 12544 52476 12572 52974
rect 12624 52556 12676 52562
rect 12624 52498 12676 52504
rect 12492 52448 12572 52476
rect 12440 52430 12492 52436
rect 12256 52148 12308 52154
rect 12256 52090 12308 52096
rect 12176 52006 12296 52034
rect 12268 51474 12296 52006
rect 12348 51808 12400 51814
rect 12348 51750 12400 51756
rect 12256 51468 12308 51474
rect 12256 51410 12308 51416
rect 12268 51066 12296 51410
rect 12256 51060 12308 51066
rect 12256 51002 12308 51008
rect 12254 50688 12310 50697
rect 12254 50623 12310 50632
rect 12268 49978 12296 50623
rect 12360 50454 12388 51750
rect 12452 51513 12480 52430
rect 12636 52329 12664 52498
rect 12622 52320 12678 52329
rect 12678 52278 12756 52306
rect 12622 52255 12678 52264
rect 12624 51808 12676 51814
rect 12624 51750 12676 51756
rect 12438 51504 12494 51513
rect 12438 51439 12494 51448
rect 12348 50448 12400 50454
rect 12348 50390 12400 50396
rect 12256 49972 12308 49978
rect 12256 49914 12308 49920
rect 12164 49836 12216 49842
rect 12164 49778 12216 49784
rect 12070 48648 12126 48657
rect 12070 48583 12126 48592
rect 11978 47560 12034 47569
rect 11978 47495 12034 47504
rect 11992 47462 12020 47495
rect 11980 47456 12032 47462
rect 11980 47398 12032 47404
rect 11888 46368 11940 46374
rect 11888 46310 11940 46316
rect 11900 46170 11928 46310
rect 11888 46164 11940 46170
rect 11888 46106 11940 46112
rect 11992 46050 12020 47398
rect 11900 46022 12020 46050
rect 11796 44940 11848 44946
rect 11796 44882 11848 44888
rect 11808 44538 11836 44882
rect 11796 44532 11848 44538
rect 11796 44474 11848 44480
rect 11808 44198 11836 44474
rect 11796 44192 11848 44198
rect 11796 44134 11848 44140
rect 11808 41614 11836 44134
rect 11796 41608 11848 41614
rect 11796 41550 11848 41556
rect 11702 41304 11758 41313
rect 11808 41274 11836 41550
rect 11702 41239 11758 41248
rect 11796 41268 11848 41274
rect 11796 41210 11848 41216
rect 11900 41177 11928 46022
rect 11980 44872 12032 44878
rect 11980 44814 12032 44820
rect 11992 42702 12020 44814
rect 12072 43852 12124 43858
rect 12072 43794 12124 43800
rect 12084 43246 12112 43794
rect 12072 43240 12124 43246
rect 12072 43182 12124 43188
rect 12072 42764 12124 42770
rect 12072 42706 12124 42712
rect 11980 42696 12032 42702
rect 11980 42638 12032 42644
rect 11992 42362 12020 42638
rect 11980 42356 12032 42362
rect 11980 42298 12032 42304
rect 12084 42022 12112 42706
rect 12072 42016 12124 42022
rect 12072 41958 12124 41964
rect 11886 41168 11942 41177
rect 11886 41103 11942 41112
rect 11704 41064 11756 41070
rect 11704 41006 11756 41012
rect 11716 40186 11744 41006
rect 11796 40452 11848 40458
rect 11796 40394 11848 40400
rect 11704 40180 11756 40186
rect 11704 40122 11756 40128
rect 11704 40044 11756 40050
rect 11704 39986 11756 39992
rect 11716 36310 11744 39986
rect 11808 39506 11836 40394
rect 11796 39500 11848 39506
rect 11796 39442 11848 39448
rect 11808 37874 11836 39442
rect 11796 37868 11848 37874
rect 11796 37810 11848 37816
rect 11796 37392 11848 37398
rect 11796 37334 11848 37340
rect 11704 36304 11756 36310
rect 11704 36246 11756 36252
rect 11808 36038 11836 37334
rect 11796 36032 11848 36038
rect 11796 35974 11848 35980
rect 11704 35624 11756 35630
rect 11704 35566 11756 35572
rect 11716 34950 11744 35566
rect 11704 34944 11756 34950
rect 11704 34886 11756 34892
rect 11612 34672 11664 34678
rect 11612 34614 11664 34620
rect 11704 34672 11756 34678
rect 11704 34614 11756 34620
rect 11716 34354 11744 34614
rect 11624 34326 11744 34354
rect 11518 31648 11574 31657
rect 11518 31583 11574 31592
rect 11426 31512 11482 31521
rect 11426 31447 11482 31456
rect 11520 31476 11572 31482
rect 11520 31418 11572 31424
rect 11532 31260 11560 31418
rect 11440 31232 11560 31260
rect 11440 30258 11468 31232
rect 11624 31192 11652 34326
rect 11702 34232 11758 34241
rect 11702 34167 11758 34176
rect 11716 33969 11744 34167
rect 11808 34116 11836 35974
rect 11900 34678 11928 41103
rect 12072 40928 12124 40934
rect 12072 40870 12124 40876
rect 12084 40594 12112 40870
rect 12072 40588 12124 40594
rect 12072 40530 12124 40536
rect 11980 40520 12032 40526
rect 11980 40462 12032 40468
rect 11992 40118 12020 40462
rect 11980 40112 12032 40118
rect 11980 40054 12032 40060
rect 12072 39976 12124 39982
rect 12072 39918 12124 39924
rect 11980 39840 12032 39846
rect 11980 39782 12032 39788
rect 11992 39302 12020 39782
rect 11980 39296 12032 39302
rect 11980 39238 12032 39244
rect 11978 38584 12034 38593
rect 11978 38519 12034 38528
rect 11992 35222 12020 38519
rect 11980 35216 12032 35222
rect 11980 35158 12032 35164
rect 12084 35018 12112 39918
rect 12176 39574 12204 49778
rect 12636 49745 12664 51750
rect 12728 51610 12756 52278
rect 12820 51950 12848 53042
rect 12808 51944 12860 51950
rect 12808 51886 12860 51892
rect 12716 51604 12768 51610
rect 12716 51546 12768 51552
rect 12714 51504 12770 51513
rect 12714 51439 12716 51448
rect 12768 51439 12770 51448
rect 12716 51410 12768 51416
rect 12728 50522 12756 51410
rect 12716 50516 12768 50522
rect 12716 50458 12768 50464
rect 12820 49842 12848 51886
rect 12808 49836 12860 49842
rect 12728 49796 12808 49824
rect 12622 49736 12678 49745
rect 12622 49671 12678 49680
rect 12256 49292 12308 49298
rect 12256 49234 12308 49240
rect 12268 48890 12296 49234
rect 12728 49230 12756 49796
rect 12808 49778 12860 49784
rect 12716 49224 12768 49230
rect 12716 49166 12768 49172
rect 12912 48890 12940 60676
rect 13268 56908 13320 56914
rect 13268 56850 13320 56856
rect 13280 56166 13308 56850
rect 13268 56160 13320 56166
rect 13266 56128 13268 56137
rect 13320 56128 13322 56137
rect 13266 56063 13322 56072
rect 13176 55820 13228 55826
rect 13176 55762 13228 55768
rect 13084 55616 13136 55622
rect 13084 55558 13136 55564
rect 13096 54602 13124 55558
rect 13188 55418 13216 55762
rect 13176 55412 13228 55418
rect 13176 55354 13228 55360
rect 13268 55072 13320 55078
rect 13268 55014 13320 55020
rect 13174 54632 13230 54641
rect 13084 54596 13136 54602
rect 13174 54567 13230 54576
rect 13084 54538 13136 54544
rect 13188 54097 13216 54567
rect 13174 54088 13230 54097
rect 13174 54023 13230 54032
rect 12992 52352 13044 52358
rect 12992 52294 13044 52300
rect 13004 51474 13032 52294
rect 13280 51542 13308 55014
rect 13268 51536 13320 51542
rect 13268 51478 13320 51484
rect 12992 51468 13044 51474
rect 12992 51410 13044 51416
rect 13084 51264 13136 51270
rect 13084 51206 13136 51212
rect 12992 51060 13044 51066
rect 12992 51002 13044 51008
rect 13004 50522 13032 51002
rect 13096 50697 13124 51206
rect 13082 50688 13138 50697
rect 13082 50623 13138 50632
rect 12992 50516 13044 50522
rect 12992 50458 13044 50464
rect 13096 50425 13124 50623
rect 13082 50416 13138 50425
rect 13082 50351 13138 50360
rect 13268 49836 13320 49842
rect 13268 49778 13320 49784
rect 13280 49434 13308 49778
rect 13268 49428 13320 49434
rect 13268 49370 13320 49376
rect 12256 48884 12308 48890
rect 12256 48826 12308 48832
rect 12900 48884 12952 48890
rect 12900 48826 12952 48832
rect 12912 48686 12940 48826
rect 12900 48680 12952 48686
rect 12900 48622 12952 48628
rect 13174 48648 13230 48657
rect 12808 48544 12860 48550
rect 12806 48512 12808 48521
rect 12860 48512 12862 48521
rect 12806 48447 12862 48456
rect 12912 48113 12940 48622
rect 13174 48583 13230 48592
rect 13188 48278 13216 48583
rect 13176 48272 13228 48278
rect 13176 48214 13228 48220
rect 12898 48104 12954 48113
rect 12898 48039 12954 48048
rect 13082 48104 13138 48113
rect 13082 48039 13138 48048
rect 13096 47802 13124 48039
rect 13084 47796 13136 47802
rect 13084 47738 13136 47744
rect 12532 47116 12584 47122
rect 12532 47058 12584 47064
rect 12544 46646 12572 47058
rect 12624 47048 12676 47054
rect 12624 46990 12676 46996
rect 12532 46640 12584 46646
rect 12532 46582 12584 46588
rect 12440 46504 12492 46510
rect 12440 46446 12492 46452
rect 12348 46368 12400 46374
rect 12348 46310 12400 46316
rect 12256 45620 12308 45626
rect 12256 45562 12308 45568
rect 12268 43926 12296 45562
rect 12360 45558 12388 46310
rect 12452 46034 12480 46446
rect 12440 46028 12492 46034
rect 12440 45970 12492 45976
rect 12348 45552 12400 45558
rect 12348 45494 12400 45500
rect 12452 45422 12480 45970
rect 12636 45898 12664 46990
rect 12716 46504 12768 46510
rect 12716 46446 12768 46452
rect 12728 46034 12756 46446
rect 13280 46102 13308 49370
rect 13372 48278 13400 62698
rect 13740 62354 13768 74734
rect 13728 62348 13780 62354
rect 13728 62290 13780 62296
rect 13832 61946 13860 74734
rect 14372 73296 14424 73302
rect 14370 73264 14372 73273
rect 14424 73264 14426 73273
rect 14370 73199 14426 73208
rect 15198 68912 15254 68921
rect 15198 68847 15254 68856
rect 15106 66192 15162 66201
rect 15106 66127 15162 66136
rect 14372 65612 14424 65618
rect 14372 65554 14424 65560
rect 14384 65074 14412 65554
rect 14372 65068 14424 65074
rect 14372 65010 14424 65016
rect 14096 62824 14148 62830
rect 14096 62766 14148 62772
rect 13820 61940 13872 61946
rect 13820 61882 13872 61888
rect 13452 57928 13504 57934
rect 13452 57870 13504 57876
rect 13464 57594 13492 57870
rect 13728 57860 13780 57866
rect 13728 57802 13780 57808
rect 13544 57792 13596 57798
rect 13544 57734 13596 57740
rect 13452 57588 13504 57594
rect 13452 57530 13504 57536
rect 13452 57452 13504 57458
rect 13452 57394 13504 57400
rect 13464 57050 13492 57394
rect 13556 57390 13584 57734
rect 13544 57384 13596 57390
rect 13544 57326 13596 57332
rect 13452 57044 13504 57050
rect 13452 56986 13504 56992
rect 13556 56273 13584 57326
rect 13740 57050 13768 57802
rect 14004 57248 14056 57254
rect 14004 57190 14056 57196
rect 13728 57044 13780 57050
rect 13728 56986 13780 56992
rect 13728 56432 13780 56438
rect 13726 56400 13728 56409
rect 13780 56400 13782 56409
rect 13726 56335 13782 56344
rect 13542 56264 13598 56273
rect 13542 56199 13598 56208
rect 14016 55962 14044 57190
rect 14004 55956 14056 55962
rect 14004 55898 14056 55904
rect 14004 55820 14056 55826
rect 14004 55762 14056 55768
rect 14016 55078 14044 55762
rect 14004 55072 14056 55078
rect 14004 55014 14056 55020
rect 13820 54732 13872 54738
rect 13820 54674 13872 54680
rect 13832 54330 13860 54674
rect 13912 54528 13964 54534
rect 13912 54470 13964 54476
rect 13820 54324 13872 54330
rect 13820 54266 13872 54272
rect 13452 54120 13504 54126
rect 13450 54088 13452 54097
rect 13504 54088 13506 54097
rect 13450 54023 13506 54032
rect 13832 53990 13860 54266
rect 13924 54126 13952 54470
rect 13912 54120 13964 54126
rect 13912 54062 13964 54068
rect 13820 53984 13872 53990
rect 13820 53926 13872 53932
rect 13832 53428 13860 53926
rect 13924 53718 13952 54062
rect 14016 54058 14044 55014
rect 14004 54052 14056 54058
rect 14004 53994 14056 54000
rect 14016 53961 14044 53994
rect 14002 53952 14058 53961
rect 14002 53887 14058 53896
rect 13912 53712 13964 53718
rect 13912 53654 13964 53660
rect 14004 53440 14056 53446
rect 13832 53400 14004 53428
rect 14004 53382 14056 53388
rect 14016 53038 14044 53382
rect 14004 53032 14056 53038
rect 14004 52974 14056 52980
rect 14016 52902 14044 52974
rect 14004 52896 14056 52902
rect 14004 52838 14056 52844
rect 14016 52737 14044 52838
rect 14002 52728 14058 52737
rect 13820 52692 13872 52698
rect 14002 52663 14058 52672
rect 13820 52634 13872 52640
rect 13728 52420 13780 52426
rect 13728 52362 13780 52368
rect 13542 52048 13598 52057
rect 13542 51983 13598 51992
rect 13556 51610 13584 51983
rect 13544 51604 13596 51610
rect 13544 51546 13596 51552
rect 13452 51332 13504 51338
rect 13452 51274 13504 51280
rect 13464 50930 13492 51274
rect 13452 50924 13504 50930
rect 13452 50866 13504 50872
rect 13556 50862 13584 51546
rect 13544 50856 13596 50862
rect 13544 50798 13596 50804
rect 13556 50522 13584 50798
rect 13544 50516 13596 50522
rect 13544 50458 13596 50464
rect 13452 49972 13504 49978
rect 13452 49914 13504 49920
rect 13360 48272 13412 48278
rect 13360 48214 13412 48220
rect 13464 48074 13492 49914
rect 13740 49842 13768 52362
rect 13832 50969 13860 52634
rect 13912 52556 13964 52562
rect 13912 52498 13964 52504
rect 13924 52086 13952 52498
rect 13912 52080 13964 52086
rect 13912 52022 13964 52028
rect 13912 51536 13964 51542
rect 13912 51478 13964 51484
rect 13818 50960 13874 50969
rect 13818 50895 13874 50904
rect 13924 50862 13952 51478
rect 14004 51400 14056 51406
rect 14004 51342 14056 51348
rect 14016 51066 14044 51342
rect 14004 51060 14056 51066
rect 14004 51002 14056 51008
rect 13912 50856 13964 50862
rect 13912 50798 13964 50804
rect 14002 50824 14058 50833
rect 14002 50759 14058 50768
rect 14016 50386 14044 50759
rect 14004 50380 14056 50386
rect 14004 50322 14056 50328
rect 14016 49978 14044 50322
rect 14004 49972 14056 49978
rect 14004 49914 14056 49920
rect 13728 49836 13780 49842
rect 13912 49836 13964 49842
rect 13728 49778 13780 49784
rect 13832 49796 13912 49824
rect 13728 49292 13780 49298
rect 13832 49280 13860 49796
rect 13912 49778 13964 49784
rect 13780 49252 13860 49280
rect 13728 49234 13780 49240
rect 13542 49192 13598 49201
rect 13542 49127 13598 49136
rect 13556 48890 13584 49127
rect 13912 49088 13964 49094
rect 13912 49030 13964 49036
rect 13634 48920 13690 48929
rect 13544 48884 13596 48890
rect 13634 48855 13690 48864
rect 13544 48826 13596 48832
rect 13648 48686 13676 48855
rect 13636 48680 13688 48686
rect 13636 48622 13688 48628
rect 13648 48346 13676 48622
rect 13820 48544 13872 48550
rect 13820 48486 13872 48492
rect 13636 48340 13688 48346
rect 13636 48282 13688 48288
rect 13728 48136 13780 48142
rect 13728 48078 13780 48084
rect 13452 48068 13504 48074
rect 13452 48010 13504 48016
rect 13464 47802 13492 48010
rect 13452 47796 13504 47802
rect 13452 47738 13504 47744
rect 13740 47734 13768 48078
rect 13832 47802 13860 48486
rect 13820 47796 13872 47802
rect 13820 47738 13872 47744
rect 13728 47728 13780 47734
rect 13728 47670 13780 47676
rect 13740 47258 13768 47670
rect 13728 47252 13780 47258
rect 13728 47194 13780 47200
rect 13924 47138 13952 49030
rect 14002 47288 14058 47297
rect 14108 47258 14136 62766
rect 14384 59129 14412 65010
rect 15120 63306 15148 66127
rect 15212 65482 15240 68847
rect 15200 65476 15252 65482
rect 15200 65418 15252 65424
rect 15108 63300 15160 63306
rect 15108 63242 15160 63248
rect 14556 59424 14608 59430
rect 14462 59392 14518 59401
rect 14556 59366 14608 59372
rect 14462 59327 14518 59336
rect 14370 59120 14426 59129
rect 14370 59055 14426 59064
rect 14384 58138 14412 59055
rect 14476 58682 14504 59327
rect 14464 58676 14516 58682
rect 14464 58618 14516 58624
rect 14372 58132 14424 58138
rect 14372 58074 14424 58080
rect 14372 57928 14424 57934
rect 14372 57870 14424 57876
rect 14384 57254 14412 57870
rect 14372 57248 14424 57254
rect 14372 57190 14424 57196
rect 14384 57050 14412 57190
rect 14372 57044 14424 57050
rect 14372 56986 14424 56992
rect 14568 56930 14596 59366
rect 14740 59084 14792 59090
rect 14740 59026 14792 59032
rect 14648 58880 14700 58886
rect 14648 58822 14700 58828
rect 14660 58585 14688 58822
rect 14646 58576 14702 58585
rect 14646 58511 14702 58520
rect 14752 58410 14780 59026
rect 14740 58404 14792 58410
rect 14740 58346 14792 58352
rect 14752 57798 14780 58346
rect 14832 58336 14884 58342
rect 14830 58304 14832 58313
rect 14884 58304 14886 58313
rect 14830 58239 14886 58248
rect 15108 57996 15160 58002
rect 15108 57938 15160 57944
rect 15120 57882 15148 57938
rect 15120 57854 15240 57882
rect 14740 57792 14792 57798
rect 14740 57734 14792 57740
rect 14648 57452 14700 57458
rect 14648 57394 14700 57400
rect 14660 57089 14688 57394
rect 14752 57390 14780 57734
rect 14740 57384 14792 57390
rect 14740 57326 14792 57332
rect 14646 57080 14702 57089
rect 14646 57015 14702 57024
rect 14188 56908 14240 56914
rect 14188 56850 14240 56856
rect 14384 56902 14596 56930
rect 14752 56914 14780 57326
rect 14740 56908 14792 56914
rect 14200 56409 14228 56850
rect 14186 56400 14242 56409
rect 14186 56335 14242 56344
rect 14280 56364 14332 56370
rect 14280 56306 14332 56312
rect 14186 56264 14242 56273
rect 14186 56199 14242 56208
rect 14200 52476 14228 56199
rect 14292 56166 14320 56306
rect 14280 56160 14332 56166
rect 14280 56102 14332 56108
rect 14292 55962 14320 56102
rect 14280 55956 14332 55962
rect 14280 55898 14332 55904
rect 14292 55865 14320 55898
rect 14278 55856 14334 55865
rect 14278 55791 14334 55800
rect 14384 55690 14412 56902
rect 14740 56850 14792 56856
rect 14924 56840 14976 56846
rect 14924 56782 14976 56788
rect 14832 55888 14884 55894
rect 14832 55830 14884 55836
rect 14372 55684 14424 55690
rect 14372 55626 14424 55632
rect 14278 52864 14334 52873
rect 14278 52799 14334 52808
rect 14292 52630 14320 52799
rect 14280 52624 14332 52630
rect 14280 52566 14332 52572
rect 14384 52494 14412 55626
rect 14554 55448 14610 55457
rect 14554 55383 14610 55392
rect 14464 55208 14516 55214
rect 14464 55150 14516 55156
rect 14476 54874 14504 55150
rect 14464 54868 14516 54874
rect 14464 54810 14516 54816
rect 14462 53544 14518 53553
rect 14462 53479 14518 53488
rect 14476 53242 14504 53479
rect 14464 53236 14516 53242
rect 14464 53178 14516 53184
rect 14476 52630 14504 53178
rect 14464 52624 14516 52630
rect 14464 52566 14516 52572
rect 14372 52488 14424 52494
rect 14200 52448 14320 52476
rect 14292 52170 14320 52448
rect 14372 52430 14424 52436
rect 14292 52142 14412 52170
rect 14188 51400 14240 51406
rect 14188 51342 14240 51348
rect 14200 50425 14228 51342
rect 14280 51264 14332 51270
rect 14280 51206 14332 51212
rect 14186 50416 14242 50425
rect 14186 50351 14188 50360
rect 14240 50351 14242 50360
rect 14188 50322 14240 50328
rect 14292 49201 14320 51206
rect 14278 49192 14334 49201
rect 14278 49127 14334 49136
rect 14188 48204 14240 48210
rect 14188 48146 14240 48152
rect 14200 47666 14228 48146
rect 14188 47660 14240 47666
rect 14188 47602 14240 47608
rect 14002 47223 14004 47232
rect 14056 47223 14058 47232
rect 14096 47252 14148 47258
rect 14004 47194 14056 47200
rect 14096 47194 14148 47200
rect 13740 47122 14044 47138
rect 13728 47116 14044 47122
rect 13780 47110 14044 47116
rect 13728 47058 13780 47064
rect 13740 46714 13768 47058
rect 13728 46708 13780 46714
rect 13728 46650 13780 46656
rect 13268 46096 13320 46102
rect 13268 46038 13320 46044
rect 12716 46028 12768 46034
rect 12716 45970 12768 45976
rect 13452 46028 13504 46034
rect 13452 45970 13504 45976
rect 12624 45892 12676 45898
rect 12624 45834 12676 45840
rect 12636 45422 12664 45834
rect 13464 45422 13492 45970
rect 13820 45960 13872 45966
rect 13820 45902 13872 45908
rect 13636 45484 13688 45490
rect 13636 45426 13688 45432
rect 12440 45416 12492 45422
rect 12440 45358 12492 45364
rect 12624 45416 12676 45422
rect 12624 45358 12676 45364
rect 13452 45416 13504 45422
rect 13452 45358 13504 45364
rect 12636 45082 12664 45358
rect 12624 45076 12676 45082
rect 12624 45018 12676 45024
rect 12636 44470 12664 45018
rect 13648 45014 13676 45426
rect 13636 45008 13688 45014
rect 13636 44950 13688 44956
rect 13452 44940 13504 44946
rect 13452 44882 13504 44888
rect 12624 44464 12676 44470
rect 12624 44406 12676 44412
rect 12624 44328 12676 44334
rect 12624 44270 12676 44276
rect 12256 43920 12308 43926
rect 12256 43862 12308 43868
rect 12164 39568 12216 39574
rect 12164 39510 12216 39516
rect 12164 39296 12216 39302
rect 12164 39238 12216 39244
rect 12176 38894 12204 39238
rect 12164 38888 12216 38894
rect 12164 38830 12216 38836
rect 12176 38758 12204 38830
rect 12164 38752 12216 38758
rect 12164 38694 12216 38700
rect 12176 38486 12204 38694
rect 12164 38480 12216 38486
rect 12164 38422 12216 38428
rect 12176 35873 12204 38422
rect 12162 35864 12218 35873
rect 12162 35799 12218 35808
rect 12164 35556 12216 35562
rect 12164 35498 12216 35504
rect 12072 35012 12124 35018
rect 12072 34954 12124 34960
rect 12070 34912 12126 34921
rect 12070 34847 12126 34856
rect 11888 34672 11940 34678
rect 11888 34614 11940 34620
rect 11980 34468 12032 34474
rect 11980 34410 12032 34416
rect 11992 34377 12020 34410
rect 11978 34368 12034 34377
rect 11978 34303 12034 34312
rect 11980 34128 12032 34134
rect 11808 34088 11928 34116
rect 11702 33960 11758 33969
rect 11702 33895 11758 33904
rect 11794 33824 11850 33833
rect 11794 33759 11850 33768
rect 11808 31890 11836 33759
rect 11796 31884 11848 31890
rect 11796 31826 11848 31832
rect 11702 31648 11758 31657
rect 11702 31583 11758 31592
rect 11532 31164 11652 31192
rect 11532 30802 11560 31164
rect 11610 31104 11666 31113
rect 11610 31039 11666 31048
rect 11520 30796 11572 30802
rect 11520 30738 11572 30744
rect 11532 30705 11560 30738
rect 11518 30696 11574 30705
rect 11518 30631 11574 30640
rect 11520 30592 11572 30598
rect 11520 30534 11572 30540
rect 11428 30252 11480 30258
rect 11428 30194 11480 30200
rect 11428 30116 11480 30122
rect 11428 30058 11480 30064
rect 11440 29578 11468 30058
rect 11532 29753 11560 30534
rect 11518 29744 11574 29753
rect 11518 29679 11574 29688
rect 11428 29572 11480 29578
rect 11428 29514 11480 29520
rect 11440 29306 11468 29514
rect 11518 29472 11574 29481
rect 11518 29407 11574 29416
rect 11428 29300 11480 29306
rect 11428 29242 11480 29248
rect 11428 29164 11480 29170
rect 11428 29106 11480 29112
rect 11440 28762 11468 29106
rect 11428 28756 11480 28762
rect 11428 28698 11480 28704
rect 11532 28626 11560 29407
rect 11624 28694 11652 31039
rect 11612 28688 11664 28694
rect 11612 28630 11664 28636
rect 11520 28620 11572 28626
rect 11520 28562 11572 28568
rect 11428 28552 11480 28558
rect 11428 28494 11480 28500
rect 11440 27470 11468 28494
rect 11532 28257 11560 28562
rect 11716 28558 11744 31583
rect 11808 31482 11836 31826
rect 11900 31804 11928 34088
rect 11980 34070 12032 34076
rect 11992 33318 12020 34070
rect 12084 33998 12112 34847
rect 12176 34746 12204 35498
rect 12164 34740 12216 34746
rect 12164 34682 12216 34688
rect 12164 34468 12216 34474
rect 12164 34410 12216 34416
rect 12176 34202 12204 34410
rect 12164 34196 12216 34202
rect 12164 34138 12216 34144
rect 12072 33992 12124 33998
rect 12072 33934 12124 33940
rect 12084 33697 12112 33934
rect 12070 33688 12126 33697
rect 12176 33658 12204 34138
rect 12070 33623 12126 33632
rect 12164 33652 12216 33658
rect 12164 33594 12216 33600
rect 12072 33584 12124 33590
rect 12072 33526 12124 33532
rect 11980 33312 12032 33318
rect 11980 33254 12032 33260
rect 11992 32473 12020 33254
rect 11978 32464 12034 32473
rect 11978 32399 12034 32408
rect 11992 31929 12020 32399
rect 11978 31920 12034 31929
rect 11978 31855 12034 31864
rect 11900 31776 12020 31804
rect 11796 31476 11848 31482
rect 11796 31418 11848 31424
rect 11888 31340 11940 31346
rect 11888 31282 11940 31288
rect 11796 31272 11848 31278
rect 11796 31214 11848 31220
rect 11808 30666 11836 31214
rect 11796 30660 11848 30666
rect 11796 30602 11848 30608
rect 11796 29844 11848 29850
rect 11796 29786 11848 29792
rect 11612 28552 11664 28558
rect 11612 28494 11664 28500
rect 11704 28552 11756 28558
rect 11704 28494 11756 28500
rect 11518 28248 11574 28257
rect 11518 28183 11574 28192
rect 11428 27464 11480 27470
rect 11428 27406 11480 27412
rect 11624 27418 11652 28494
rect 11716 28121 11744 28494
rect 11702 28112 11758 28121
rect 11702 28047 11758 28056
rect 11716 27878 11744 28047
rect 11704 27872 11756 27878
rect 11704 27814 11756 27820
rect 11624 27390 11744 27418
rect 11612 27328 11664 27334
rect 11612 27270 11664 27276
rect 11520 26784 11572 26790
rect 11520 26726 11572 26732
rect 11532 26586 11560 26726
rect 11520 26580 11572 26586
rect 11520 26522 11572 26528
rect 11624 26432 11652 27270
rect 11716 26790 11744 27390
rect 11704 26784 11756 26790
rect 11704 26726 11756 26732
rect 11532 26404 11652 26432
rect 11428 26376 11480 26382
rect 11428 26318 11480 26324
rect 10876 25492 10928 25498
rect 10876 25434 10928 25440
rect 11336 25492 11388 25498
rect 11336 25434 11388 25440
rect 10876 25356 10928 25362
rect 10876 25298 10928 25304
rect 10888 24410 10916 25298
rect 10956 24508 11252 24528
rect 11012 24506 11036 24508
rect 11092 24506 11116 24508
rect 11172 24506 11196 24508
rect 11034 24454 11036 24506
rect 11098 24454 11110 24506
rect 11172 24454 11174 24506
rect 11012 24452 11036 24454
rect 11092 24452 11116 24454
rect 11172 24452 11196 24454
rect 10956 24432 11252 24452
rect 10876 24404 10928 24410
rect 11440 24392 11468 26318
rect 11532 25702 11560 26404
rect 11612 26308 11664 26314
rect 11612 26250 11664 26256
rect 11520 25696 11572 25702
rect 11520 25638 11572 25644
rect 11520 25152 11572 25158
rect 11520 25094 11572 25100
rect 10876 24346 10928 24352
rect 11164 24364 11468 24392
rect 10968 24336 11020 24342
rect 10968 24278 11020 24284
rect 10876 24064 10928 24070
rect 10874 24032 10876 24041
rect 10928 24032 10930 24041
rect 10874 23967 10930 23976
rect 10980 23866 11008 24278
rect 10968 23860 11020 23866
rect 10968 23802 11020 23808
rect 11164 23508 11192 24364
rect 11428 24268 11480 24274
rect 11428 24210 11480 24216
rect 11336 24200 11388 24206
rect 11336 24142 11388 24148
rect 10888 23480 11192 23508
rect 10784 23248 10836 23254
rect 10784 23190 10836 23196
rect 10782 21720 10838 21729
rect 10782 21655 10784 21664
rect 10836 21655 10838 21664
rect 10784 21626 10836 21632
rect 10888 20942 10916 23480
rect 10956 23420 11252 23440
rect 11012 23418 11036 23420
rect 11092 23418 11116 23420
rect 11172 23418 11196 23420
rect 11034 23366 11036 23418
rect 11098 23366 11110 23418
rect 11172 23366 11174 23418
rect 11012 23364 11036 23366
rect 11092 23364 11116 23366
rect 11172 23364 11196 23366
rect 10956 23344 11252 23364
rect 11348 23322 11376 24142
rect 11440 23866 11468 24210
rect 11428 23860 11480 23866
rect 11428 23802 11480 23808
rect 11426 23624 11482 23633
rect 11426 23559 11482 23568
rect 11336 23316 11388 23322
rect 11336 23258 11388 23264
rect 10968 23180 11020 23186
rect 10968 23122 11020 23128
rect 10980 22506 11008 23122
rect 11152 23112 11204 23118
rect 11152 23054 11204 23060
rect 11164 22778 11192 23054
rect 11152 22772 11204 22778
rect 11152 22714 11204 22720
rect 11348 22681 11376 23258
rect 11334 22672 11390 22681
rect 11334 22607 11390 22616
rect 10968 22500 11020 22506
rect 10968 22442 11020 22448
rect 11336 22500 11388 22506
rect 11336 22442 11388 22448
rect 10956 22332 11252 22352
rect 11012 22330 11036 22332
rect 11092 22330 11116 22332
rect 11172 22330 11196 22332
rect 11034 22278 11036 22330
rect 11098 22278 11110 22330
rect 11172 22278 11174 22330
rect 11012 22276 11036 22278
rect 11092 22276 11116 22278
rect 11172 22276 11196 22278
rect 10956 22256 11252 22276
rect 10956 21244 11252 21264
rect 11012 21242 11036 21244
rect 11092 21242 11116 21244
rect 11172 21242 11196 21244
rect 11034 21190 11036 21242
rect 11098 21190 11110 21242
rect 11172 21190 11174 21242
rect 11012 21188 11036 21190
rect 11092 21188 11116 21190
rect 11172 21188 11196 21190
rect 10956 21168 11252 21188
rect 11060 21004 11112 21010
rect 11060 20946 11112 20952
rect 10876 20936 10928 20942
rect 10876 20878 10928 20884
rect 10782 20768 10838 20777
rect 10782 20703 10838 20712
rect 10612 20590 10732 20618
rect 10506 18864 10562 18873
rect 10506 18799 10562 18808
rect 10508 18692 10560 18698
rect 10508 18634 10560 18640
rect 10520 17785 10548 18634
rect 10506 17776 10562 17785
rect 10506 17711 10562 17720
rect 10612 17134 10640 20590
rect 10692 20460 10744 20466
rect 10692 20402 10744 20408
rect 10704 18358 10732 20402
rect 10796 18970 10824 20703
rect 10888 20602 10916 20878
rect 10968 20868 11020 20874
rect 10968 20810 11020 20816
rect 10876 20596 10928 20602
rect 10876 20538 10928 20544
rect 10980 20398 11008 20810
rect 11072 20641 11100 20946
rect 11348 20806 11376 22442
rect 11440 21146 11468 23559
rect 11532 23322 11560 25094
rect 11624 24614 11652 26250
rect 11704 25968 11756 25974
rect 11704 25910 11756 25916
rect 11716 25362 11744 25910
rect 11704 25356 11756 25362
rect 11704 25298 11756 25304
rect 11612 24608 11664 24614
rect 11612 24550 11664 24556
rect 11520 23316 11572 23322
rect 11520 23258 11572 23264
rect 11520 23180 11572 23186
rect 11520 23122 11572 23128
rect 11532 22710 11560 23122
rect 11520 22704 11572 22710
rect 11520 22646 11572 22652
rect 11520 21412 11572 21418
rect 11520 21354 11572 21360
rect 11428 21140 11480 21146
rect 11428 21082 11480 21088
rect 11336 20800 11388 20806
rect 11336 20742 11388 20748
rect 11058 20632 11114 20641
rect 11058 20567 11114 20576
rect 10968 20392 11020 20398
rect 10888 20352 10968 20380
rect 10888 19990 10916 20352
rect 10968 20334 11020 20340
rect 11336 20392 11388 20398
rect 11336 20334 11388 20340
rect 10956 20156 11252 20176
rect 11012 20154 11036 20156
rect 11092 20154 11116 20156
rect 11172 20154 11196 20156
rect 11034 20102 11036 20154
rect 11098 20102 11110 20154
rect 11172 20102 11174 20154
rect 11012 20100 11036 20102
rect 11092 20100 11116 20102
rect 11172 20100 11196 20102
rect 10956 20080 11252 20100
rect 11348 20058 11376 20334
rect 11336 20052 11388 20058
rect 11336 19994 11388 20000
rect 10876 19984 10928 19990
rect 10876 19926 10928 19932
rect 11440 19854 11468 21082
rect 11532 21010 11560 21354
rect 11520 21004 11572 21010
rect 11520 20946 11572 20952
rect 11532 19922 11560 20946
rect 11520 19916 11572 19922
rect 11520 19858 11572 19864
rect 11428 19848 11480 19854
rect 11150 19816 11206 19825
rect 11428 19790 11480 19796
rect 11150 19751 11206 19760
rect 11244 19780 11296 19786
rect 11164 19242 11192 19751
rect 11244 19722 11296 19728
rect 11152 19236 11204 19242
rect 11152 19178 11204 19184
rect 11256 19156 11284 19722
rect 11256 19128 11376 19156
rect 10956 19068 11252 19088
rect 11012 19066 11036 19068
rect 11092 19066 11116 19068
rect 11172 19066 11196 19068
rect 11034 19014 11036 19066
rect 11098 19014 11110 19066
rect 11172 19014 11174 19066
rect 11012 19012 11036 19014
rect 11092 19012 11116 19014
rect 11172 19012 11196 19014
rect 10956 18992 11252 19012
rect 10784 18964 10836 18970
rect 11348 18952 11376 19128
rect 10784 18906 10836 18912
rect 11256 18924 11376 18952
rect 10876 18828 10928 18834
rect 10876 18770 10928 18776
rect 10692 18352 10744 18358
rect 10692 18294 10744 18300
rect 10782 18184 10838 18193
rect 10782 18119 10838 18128
rect 10796 17610 10824 18119
rect 10888 17814 10916 18770
rect 11256 18154 11284 18924
rect 11440 18850 11468 19790
rect 11532 19514 11560 19858
rect 11624 19786 11652 24550
rect 11716 23798 11744 25298
rect 11808 24834 11836 29786
rect 11900 26314 11928 31282
rect 11888 26308 11940 26314
rect 11888 26250 11940 26256
rect 11888 25900 11940 25906
rect 11888 25842 11940 25848
rect 11900 24954 11928 25842
rect 11992 25158 12020 31776
rect 12084 31346 12112 33526
rect 12164 33380 12216 33386
rect 12164 33322 12216 33328
rect 12176 33046 12204 33322
rect 12164 33040 12216 33046
rect 12164 32982 12216 32988
rect 12268 32994 12296 43862
rect 12636 43790 12664 44270
rect 13464 44198 13492 44882
rect 13832 44334 13860 45902
rect 13912 45552 13964 45558
rect 13912 45494 13964 45500
rect 13820 44328 13872 44334
rect 13820 44270 13872 44276
rect 13084 44192 13136 44198
rect 13084 44134 13136 44140
rect 13452 44192 13504 44198
rect 13452 44134 13504 44140
rect 13096 43858 13124 44134
rect 13084 43852 13136 43858
rect 13084 43794 13136 43800
rect 12624 43784 12676 43790
rect 12624 43726 12676 43732
rect 13096 43450 13124 43794
rect 13176 43784 13228 43790
rect 13176 43726 13228 43732
rect 13084 43444 13136 43450
rect 13084 43386 13136 43392
rect 12992 43240 13044 43246
rect 12992 43182 13044 43188
rect 12440 42764 12492 42770
rect 12440 42706 12492 42712
rect 12452 42090 12480 42706
rect 13004 42566 13032 43182
rect 12992 42560 13044 42566
rect 12992 42502 13044 42508
rect 13004 42362 13032 42502
rect 12992 42356 13044 42362
rect 12992 42298 13044 42304
rect 12440 42084 12492 42090
rect 12440 42026 12492 42032
rect 12348 41540 12400 41546
rect 12348 41482 12400 41488
rect 12360 41426 12388 41482
rect 12360 41398 12480 41426
rect 12452 40934 12480 41398
rect 12532 41268 12584 41274
rect 12532 41210 12584 41216
rect 12440 40928 12492 40934
rect 12440 40870 12492 40876
rect 12348 40588 12400 40594
rect 12348 40530 12400 40536
rect 12360 40474 12388 40530
rect 12544 40526 12572 41210
rect 12808 40928 12860 40934
rect 13084 40928 13136 40934
rect 12808 40870 12860 40876
rect 13082 40896 13084 40905
rect 13136 40896 13138 40905
rect 12532 40520 12584 40526
rect 12360 40446 12480 40474
rect 12532 40462 12584 40468
rect 12348 39432 12400 39438
rect 12348 39374 12400 39380
rect 12360 38282 12388 39374
rect 12452 39098 12480 40446
rect 12544 40186 12572 40462
rect 12532 40180 12584 40186
rect 12532 40122 12584 40128
rect 12624 39840 12676 39846
rect 12624 39782 12676 39788
rect 12440 39092 12492 39098
rect 12440 39034 12492 39040
rect 12636 38894 12664 39782
rect 12820 39302 12848 40870
rect 13082 40831 13138 40840
rect 13096 40662 13124 40831
rect 13084 40656 13136 40662
rect 13084 40598 13136 40604
rect 12900 40384 12952 40390
rect 12900 40326 12952 40332
rect 12992 40384 13044 40390
rect 12992 40326 13044 40332
rect 12808 39296 12860 39302
rect 12808 39238 12860 39244
rect 12912 38894 12940 40326
rect 13004 39506 13032 40326
rect 12992 39500 13044 39506
rect 12992 39442 13044 39448
rect 12624 38888 12676 38894
rect 12624 38830 12676 38836
rect 12716 38888 12768 38894
rect 12716 38830 12768 38836
rect 12900 38888 12952 38894
rect 12900 38830 12952 38836
rect 12532 38344 12584 38350
rect 12532 38286 12584 38292
rect 12348 38276 12400 38282
rect 12348 38218 12400 38224
rect 12544 38185 12572 38286
rect 12530 38176 12586 38185
rect 12530 38111 12586 38120
rect 12348 38004 12400 38010
rect 12348 37946 12400 37952
rect 12360 36922 12388 37946
rect 12440 37392 12492 37398
rect 12440 37334 12492 37340
rect 12348 36916 12400 36922
rect 12348 36858 12400 36864
rect 12360 34474 12388 36858
rect 12452 36650 12480 37334
rect 12544 36922 12572 38111
rect 12728 37754 12756 38830
rect 13004 38593 13032 39442
rect 13084 39364 13136 39370
rect 13084 39306 13136 39312
rect 12990 38584 13046 38593
rect 12990 38519 13046 38528
rect 12808 38412 12860 38418
rect 12808 38354 12860 38360
rect 12636 37726 12756 37754
rect 12532 36916 12584 36922
rect 12532 36858 12584 36864
rect 12636 36786 12664 37726
rect 12716 37664 12768 37670
rect 12716 37606 12768 37612
rect 12624 36780 12676 36786
rect 12624 36722 12676 36728
rect 12440 36644 12492 36650
rect 12440 36586 12492 36592
rect 12452 36106 12480 36586
rect 12624 36236 12676 36242
rect 12624 36178 12676 36184
rect 12440 36100 12492 36106
rect 12440 36042 12492 36048
rect 12452 35698 12480 36042
rect 12532 36032 12584 36038
rect 12532 35974 12584 35980
rect 12440 35692 12492 35698
rect 12440 35634 12492 35640
rect 12438 35592 12494 35601
rect 12438 35527 12440 35536
rect 12492 35527 12494 35536
rect 12440 35498 12492 35504
rect 12544 35494 12572 35974
rect 12532 35488 12584 35494
rect 12532 35430 12584 35436
rect 12544 35222 12572 35430
rect 12532 35216 12584 35222
rect 12530 35184 12532 35193
rect 12584 35184 12586 35193
rect 12530 35119 12586 35128
rect 12532 35012 12584 35018
rect 12532 34954 12584 34960
rect 12440 34944 12492 34950
rect 12440 34886 12492 34892
rect 12452 34474 12480 34886
rect 12348 34468 12400 34474
rect 12348 34410 12400 34416
rect 12440 34468 12492 34474
rect 12440 34410 12492 34416
rect 12348 33380 12400 33386
rect 12348 33322 12400 33328
rect 12360 33289 12388 33322
rect 12346 33280 12402 33289
rect 12346 33215 12402 33224
rect 12268 32966 12388 32994
rect 12256 32904 12308 32910
rect 12256 32846 12308 32852
rect 12164 32768 12216 32774
rect 12164 32710 12216 32716
rect 12176 32570 12204 32710
rect 12164 32564 12216 32570
rect 12164 32506 12216 32512
rect 12268 32230 12296 32846
rect 12256 32224 12308 32230
rect 12256 32166 12308 32172
rect 12162 32056 12218 32065
rect 12162 31991 12218 32000
rect 12176 31890 12204 31991
rect 12268 31929 12296 32166
rect 12360 31958 12388 32966
rect 12452 32910 12480 34410
rect 12544 33590 12572 34954
rect 12532 33584 12584 33590
rect 12532 33526 12584 33532
rect 12530 33280 12586 33289
rect 12530 33215 12586 33224
rect 12440 32904 12492 32910
rect 12440 32846 12492 32852
rect 12544 32298 12572 33215
rect 12532 32292 12584 32298
rect 12532 32234 12584 32240
rect 12348 31952 12400 31958
rect 12254 31920 12310 31929
rect 12164 31884 12216 31890
rect 12348 31894 12400 31900
rect 12254 31855 12310 31864
rect 12164 31826 12216 31832
rect 12348 31816 12400 31822
rect 12348 31758 12400 31764
rect 12164 31748 12216 31754
rect 12164 31690 12216 31696
rect 12072 31340 12124 31346
rect 12072 31282 12124 31288
rect 12176 30954 12204 31690
rect 12256 31136 12308 31142
rect 12254 31104 12256 31113
rect 12308 31104 12310 31113
rect 12254 31039 12310 31048
rect 12084 30926 12204 30954
rect 12084 27538 12112 30926
rect 12256 30864 12308 30870
rect 12256 30806 12308 30812
rect 12164 30728 12216 30734
rect 12164 30670 12216 30676
rect 12176 30258 12204 30670
rect 12164 30252 12216 30258
rect 12164 30194 12216 30200
rect 12268 30054 12296 30806
rect 12360 30394 12388 31758
rect 12440 31408 12492 31414
rect 12440 31350 12492 31356
rect 12452 30802 12480 31350
rect 12544 31249 12572 32234
rect 12636 32026 12664 36178
rect 12728 36009 12756 37606
rect 12820 37466 12848 38354
rect 12900 38208 12952 38214
rect 12900 38150 12952 38156
rect 12912 37738 12940 38150
rect 12992 37800 13044 37806
rect 13096 37777 13124 39306
rect 13188 38010 13216 43726
rect 13360 43716 13412 43722
rect 13360 43658 13412 43664
rect 13268 43648 13320 43654
rect 13268 43590 13320 43596
rect 13280 42945 13308 43590
rect 13372 43246 13400 43658
rect 13360 43240 13412 43246
rect 13360 43182 13412 43188
rect 13266 42936 13322 42945
rect 13266 42871 13322 42880
rect 13372 41834 13400 43182
rect 13280 41806 13400 41834
rect 13176 38004 13228 38010
rect 13176 37946 13228 37952
rect 13174 37904 13230 37913
rect 13174 37839 13176 37848
rect 13228 37839 13230 37848
rect 13176 37810 13228 37816
rect 12992 37742 13044 37748
rect 13082 37768 13138 37777
rect 12900 37732 12952 37738
rect 12900 37674 12952 37680
rect 12808 37460 12860 37466
rect 12808 37402 12860 37408
rect 12808 37324 12860 37330
rect 12808 37266 12860 37272
rect 12820 36242 12848 37266
rect 12808 36236 12860 36242
rect 12808 36178 12860 36184
rect 12714 36000 12770 36009
rect 12714 35935 12770 35944
rect 12820 35766 12848 36178
rect 12808 35760 12860 35766
rect 12808 35702 12860 35708
rect 12716 35216 12768 35222
rect 12716 35158 12768 35164
rect 12728 35018 12756 35158
rect 12808 35148 12860 35154
rect 12808 35090 12860 35096
rect 12820 35057 12848 35090
rect 12806 35048 12862 35057
rect 12716 35012 12768 35018
rect 12806 34983 12862 34992
rect 12716 34954 12768 34960
rect 12728 34542 12756 34954
rect 12716 34536 12768 34542
rect 12912 34513 12940 37674
rect 13004 37330 13032 37742
rect 13082 37703 13138 37712
rect 13176 37732 13228 37738
rect 13176 37674 13228 37680
rect 12992 37324 13044 37330
rect 12992 37266 13044 37272
rect 12990 36816 13046 36825
rect 12990 36751 13046 36760
rect 13004 35494 13032 36751
rect 13084 36712 13136 36718
rect 13084 36654 13136 36660
rect 13096 35698 13124 36654
rect 13084 35692 13136 35698
rect 13084 35634 13136 35640
rect 12992 35488 13044 35494
rect 12992 35430 13044 35436
rect 13004 35193 13032 35430
rect 12990 35184 13046 35193
rect 12990 35119 13046 35128
rect 12992 34672 13044 34678
rect 12992 34614 13044 34620
rect 12716 34478 12768 34484
rect 12898 34504 12954 34513
rect 12898 34439 12954 34448
rect 12808 34400 12860 34406
rect 12808 34342 12860 34348
rect 12820 33522 12848 34342
rect 12898 33960 12954 33969
rect 12898 33895 12900 33904
rect 12952 33895 12954 33904
rect 12900 33866 12952 33872
rect 12808 33516 12860 33522
rect 12808 33458 12860 33464
rect 13004 33402 13032 34614
rect 13084 34536 13136 34542
rect 13084 34478 13136 34484
rect 13096 34377 13124 34478
rect 13082 34368 13138 34377
rect 13082 34303 13138 34312
rect 13082 34096 13138 34105
rect 13082 34031 13138 34040
rect 13096 33862 13124 34031
rect 13084 33856 13136 33862
rect 13084 33798 13136 33804
rect 13096 33590 13124 33798
rect 13084 33584 13136 33590
rect 13084 33526 13136 33532
rect 12820 33374 13032 33402
rect 13084 33448 13136 33454
rect 13084 33390 13136 33396
rect 12714 33144 12770 33153
rect 12714 33079 12770 33088
rect 12728 33046 12756 33079
rect 12716 33040 12768 33046
rect 12716 32982 12768 32988
rect 12820 32416 12848 33374
rect 12900 33312 12952 33318
rect 13096 33289 13124 33390
rect 12900 33254 12952 33260
rect 13082 33280 13138 33289
rect 12912 33046 12940 33254
rect 13082 33215 13138 33224
rect 12900 33040 12952 33046
rect 12900 32982 12952 32988
rect 12728 32388 12848 32416
rect 12624 32020 12676 32026
rect 12624 31962 12676 31968
rect 12728 31890 12756 32388
rect 12912 32314 12940 32982
rect 13084 32972 13136 32978
rect 13084 32914 13136 32920
rect 12992 32904 13044 32910
rect 12992 32846 13044 32852
rect 12820 32286 12940 32314
rect 12716 31884 12768 31890
rect 12716 31826 12768 31832
rect 12820 31822 12848 32286
rect 13004 32230 13032 32846
rect 13096 32570 13124 32914
rect 13084 32564 13136 32570
rect 13084 32506 13136 32512
rect 13082 32328 13138 32337
rect 13082 32263 13138 32272
rect 12992 32224 13044 32230
rect 12992 32166 13044 32172
rect 12900 31952 12952 31958
rect 12900 31894 12952 31900
rect 12808 31816 12860 31822
rect 12806 31784 12808 31793
rect 12860 31784 12862 31793
rect 12806 31719 12862 31728
rect 12716 31680 12768 31686
rect 12716 31622 12768 31628
rect 12624 31340 12676 31346
rect 12624 31282 12676 31288
rect 12530 31240 12586 31249
rect 12530 31175 12586 31184
rect 12532 31136 12584 31142
rect 12532 31078 12584 31084
rect 12440 30796 12492 30802
rect 12440 30738 12492 30744
rect 12348 30388 12400 30394
rect 12348 30330 12400 30336
rect 12256 30048 12308 30054
rect 12176 30008 12256 30036
rect 12072 27532 12124 27538
rect 12072 27474 12124 27480
rect 12084 27130 12112 27474
rect 12072 27124 12124 27130
rect 12072 27066 12124 27072
rect 12084 26194 12112 27066
rect 12176 26382 12204 30008
rect 12440 30048 12492 30054
rect 12256 29990 12308 29996
rect 12346 30016 12402 30025
rect 12440 29990 12492 29996
rect 12346 29951 12402 29960
rect 12360 29782 12388 29951
rect 12348 29776 12400 29782
rect 12348 29718 12400 29724
rect 12256 29504 12308 29510
rect 12256 29446 12308 29452
rect 12268 27849 12296 29446
rect 12360 29306 12388 29718
rect 12452 29322 12480 29990
rect 12544 29510 12572 31078
rect 12636 30938 12664 31282
rect 12728 31278 12756 31622
rect 12806 31376 12862 31385
rect 12806 31311 12862 31320
rect 12716 31272 12768 31278
rect 12716 31214 12768 31220
rect 12624 30932 12676 30938
rect 12624 30874 12676 30880
rect 12716 30728 12768 30734
rect 12716 30670 12768 30676
rect 12624 30660 12676 30666
rect 12624 30602 12676 30608
rect 12532 29504 12584 29510
rect 12532 29446 12584 29452
rect 12348 29300 12400 29306
rect 12452 29294 12572 29322
rect 12348 29242 12400 29248
rect 12440 29164 12492 29170
rect 12440 29106 12492 29112
rect 12348 28688 12400 28694
rect 12348 28630 12400 28636
rect 12254 27840 12310 27849
rect 12254 27775 12310 27784
rect 12360 27334 12388 28630
rect 12452 28150 12480 29106
rect 12544 28914 12572 29294
rect 12636 29034 12664 30602
rect 12728 29646 12756 30670
rect 12716 29640 12768 29646
rect 12716 29582 12768 29588
rect 12728 29238 12756 29582
rect 12716 29232 12768 29238
rect 12716 29174 12768 29180
rect 12624 29028 12676 29034
rect 12624 28970 12676 28976
rect 12544 28886 12664 28914
rect 12532 28756 12584 28762
rect 12532 28698 12584 28704
rect 12544 28218 12572 28698
rect 12636 28529 12664 28886
rect 12716 28620 12768 28626
rect 12716 28562 12768 28568
rect 12622 28520 12678 28529
rect 12622 28455 12678 28464
rect 12532 28212 12584 28218
rect 12532 28154 12584 28160
rect 12440 28144 12492 28150
rect 12440 28086 12492 28092
rect 12440 28008 12492 28014
rect 12440 27950 12492 27956
rect 12452 27402 12480 27950
rect 12440 27396 12492 27402
rect 12440 27338 12492 27344
rect 12348 27328 12400 27334
rect 12348 27270 12400 27276
rect 12256 26784 12308 26790
rect 12256 26726 12308 26732
rect 12268 26382 12296 26726
rect 12440 26512 12492 26518
rect 12440 26454 12492 26460
rect 12348 26444 12400 26450
rect 12348 26386 12400 26392
rect 12164 26376 12216 26382
rect 12164 26318 12216 26324
rect 12256 26376 12308 26382
rect 12256 26318 12308 26324
rect 12084 26166 12296 26194
rect 12162 26072 12218 26081
rect 12162 26007 12218 26016
rect 12072 25356 12124 25362
rect 12072 25298 12124 25304
rect 11980 25152 12032 25158
rect 11980 25094 12032 25100
rect 11888 24948 11940 24954
rect 11888 24890 11940 24896
rect 11980 24880 12032 24886
rect 11808 24806 11928 24834
rect 11980 24822 12032 24828
rect 11794 24576 11850 24585
rect 11794 24511 11850 24520
rect 11808 24138 11836 24511
rect 11796 24132 11848 24138
rect 11796 24074 11848 24080
rect 11704 23792 11756 23798
rect 11704 23734 11756 23740
rect 11704 23520 11756 23526
rect 11704 23462 11756 23468
rect 11716 22778 11744 23462
rect 11704 22772 11756 22778
rect 11704 22714 11756 22720
rect 11704 21888 11756 21894
rect 11704 21830 11756 21836
rect 11716 21049 11744 21830
rect 11702 21040 11758 21049
rect 11702 20975 11758 20984
rect 11704 20936 11756 20942
rect 11704 20878 11756 20884
rect 11612 19780 11664 19786
rect 11612 19722 11664 19728
rect 11520 19508 11572 19514
rect 11520 19450 11572 19456
rect 11716 18986 11744 20878
rect 11624 18958 11744 18986
rect 11440 18822 11560 18850
rect 11428 18760 11480 18766
rect 11428 18702 11480 18708
rect 11334 18320 11390 18329
rect 11334 18255 11390 18264
rect 11244 18148 11296 18154
rect 11244 18090 11296 18096
rect 10956 17980 11252 18000
rect 11012 17978 11036 17980
rect 11092 17978 11116 17980
rect 11172 17978 11196 17980
rect 11034 17926 11036 17978
rect 11098 17926 11110 17978
rect 11172 17926 11174 17978
rect 11012 17924 11036 17926
rect 11092 17924 11116 17926
rect 11172 17924 11196 17926
rect 10956 17904 11252 17924
rect 10876 17808 10928 17814
rect 10876 17750 10928 17756
rect 11152 17740 11204 17746
rect 11152 17682 11204 17688
rect 10784 17604 10836 17610
rect 10784 17546 10836 17552
rect 10692 17332 10744 17338
rect 10692 17274 10744 17280
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10600 16992 10652 16998
rect 10600 16934 10652 16940
rect 10612 16153 10640 16934
rect 10704 16250 10732 17274
rect 10796 17202 10824 17546
rect 11164 17270 11192 17682
rect 11348 17678 11376 18255
rect 11440 18222 11468 18702
rect 11428 18216 11480 18222
rect 11428 18158 11480 18164
rect 11440 17882 11468 18158
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 11336 17672 11388 17678
rect 11336 17614 11388 17620
rect 11152 17264 11204 17270
rect 11152 17206 11204 17212
rect 10784 17196 10836 17202
rect 10784 17138 10836 17144
rect 11244 17196 11296 17202
rect 11244 17138 11296 17144
rect 10876 17128 10928 17134
rect 11256 17105 11284 17138
rect 10876 17070 10928 17076
rect 11242 17096 11298 17105
rect 10784 16788 10836 16794
rect 10784 16730 10836 16736
rect 10692 16244 10744 16250
rect 10692 16186 10744 16192
rect 10796 16182 10824 16730
rect 10888 16726 10916 17070
rect 11242 17031 11298 17040
rect 10956 16892 11252 16912
rect 11012 16890 11036 16892
rect 11092 16890 11116 16892
rect 11172 16890 11196 16892
rect 11034 16838 11036 16890
rect 11098 16838 11110 16890
rect 11172 16838 11174 16890
rect 11012 16836 11036 16838
rect 11092 16836 11116 16838
rect 11172 16836 11196 16838
rect 10956 16816 11252 16836
rect 10876 16720 10928 16726
rect 11348 16708 11376 17614
rect 11426 17232 11482 17241
rect 11426 17167 11482 17176
rect 10876 16662 10928 16668
rect 10980 16680 11376 16708
rect 10980 16538 11008 16680
rect 10888 16510 11008 16538
rect 11336 16584 11388 16590
rect 11336 16526 11388 16532
rect 10784 16176 10836 16182
rect 10598 16144 10654 16153
rect 10428 16102 10548 16130
rect 10324 15564 10376 15570
rect 10324 15506 10376 15512
rect 10336 15337 10364 15506
rect 10322 15328 10378 15337
rect 10322 15263 10378 15272
rect 10336 15162 10364 15263
rect 10324 15156 10376 15162
rect 10324 15098 10376 15104
rect 10324 14816 10376 14822
rect 10324 14758 10376 14764
rect 9956 14476 10008 14482
rect 9956 14418 10008 14424
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 9968 14385 9996 14418
rect 9954 14376 10010 14385
rect 9954 14311 10010 14320
rect 9968 14074 9996 14311
rect 9956 14068 10008 14074
rect 9956 14010 10008 14016
rect 10048 13796 10100 13802
rect 10048 13738 10100 13744
rect 10060 12986 10088 13738
rect 10048 12980 10100 12986
rect 10048 12922 10100 12928
rect 9864 12300 9916 12306
rect 9864 12242 9916 12248
rect 9876 11898 9904 12242
rect 10336 12238 10364 14758
rect 10324 12232 10376 12238
rect 10324 12174 10376 12180
rect 9956 12096 10008 12102
rect 9956 12038 10008 12044
rect 10416 12096 10468 12102
rect 10416 12038 10468 12044
rect 8944 11892 8996 11898
rect 8944 11834 8996 11840
rect 9496 11892 9548 11898
rect 9496 11834 9548 11840
rect 9864 11892 9916 11898
rect 9864 11834 9916 11840
rect 9678 9072 9734 9081
rect 9968 9058 9996 12038
rect 10428 11694 10456 12038
rect 10416 11688 10468 11694
rect 10416 11630 10468 11636
rect 10324 11620 10376 11626
rect 10324 11562 10376 11568
rect 9876 9030 9996 9058
rect 10336 9042 10364 11562
rect 10520 9761 10548 16102
rect 10784 16118 10836 16124
rect 10598 16079 10654 16088
rect 10784 16040 10836 16046
rect 10784 15982 10836 15988
rect 10692 14476 10744 14482
rect 10692 14418 10744 14424
rect 10704 14074 10732 14418
rect 10692 14068 10744 14074
rect 10692 14010 10744 14016
rect 10692 13388 10744 13394
rect 10692 13330 10744 13336
rect 10704 12986 10732 13330
rect 10796 13258 10824 15982
rect 10888 15706 10916 16510
rect 11348 15910 11376 16526
rect 11336 15904 11388 15910
rect 11336 15846 11388 15852
rect 10956 15804 11252 15824
rect 11012 15802 11036 15804
rect 11092 15802 11116 15804
rect 11172 15802 11196 15804
rect 11034 15750 11036 15802
rect 11098 15750 11110 15802
rect 11172 15750 11174 15802
rect 11012 15748 11036 15750
rect 11092 15748 11116 15750
rect 11172 15748 11196 15750
rect 10956 15728 11252 15748
rect 10876 15700 10928 15706
rect 10876 15642 10928 15648
rect 10956 14716 11252 14736
rect 11012 14714 11036 14716
rect 11092 14714 11116 14716
rect 11172 14714 11196 14716
rect 11034 14662 11036 14714
rect 11098 14662 11110 14714
rect 11172 14662 11174 14714
rect 11012 14660 11036 14662
rect 11092 14660 11116 14662
rect 11172 14660 11196 14662
rect 10956 14640 11252 14660
rect 10876 13728 10928 13734
rect 10876 13670 10928 13676
rect 10888 13274 10916 13670
rect 10956 13628 11252 13648
rect 11012 13626 11036 13628
rect 11092 13626 11116 13628
rect 11172 13626 11196 13628
rect 11034 13574 11036 13626
rect 11098 13574 11110 13626
rect 11172 13574 11174 13626
rect 11012 13572 11036 13574
rect 11092 13572 11116 13574
rect 11172 13572 11196 13574
rect 10956 13552 11252 13572
rect 10784 13252 10836 13258
rect 10888 13246 11100 13274
rect 10784 13194 10836 13200
rect 10692 12980 10744 12986
rect 10692 12922 10744 12928
rect 10600 12232 10652 12238
rect 10600 12174 10652 12180
rect 10506 9752 10562 9761
rect 10506 9687 10562 9696
rect 10324 9036 10376 9042
rect 9734 9016 9812 9024
rect 9678 9007 9680 9016
rect 9732 8996 9812 9016
rect 9680 8978 9732 8984
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 8852 8628 8904 8634
rect 8852 8570 8904 8576
rect 9692 8430 9720 8774
rect 9680 8424 9732 8430
rect 9680 8366 9732 8372
rect 9036 8356 9088 8362
rect 9036 8298 9088 8304
rect 8298 7576 8354 7585
rect 8298 7511 8354 7520
rect 6274 7440 6330 7449
rect 6274 7375 6330 7384
rect 7746 7440 7802 7449
rect 7746 7375 7802 7384
rect 5956 6556 6252 6576
rect 6012 6554 6036 6556
rect 6092 6554 6116 6556
rect 6172 6554 6196 6556
rect 6034 6502 6036 6554
rect 6098 6502 6110 6554
rect 6172 6502 6174 6554
rect 6012 6500 6036 6502
rect 6092 6500 6116 6502
rect 6172 6500 6196 6502
rect 5956 6480 6252 6500
rect 5956 5468 6252 5488
rect 6012 5466 6036 5468
rect 6092 5466 6116 5468
rect 6172 5466 6196 5468
rect 6034 5414 6036 5466
rect 6098 5414 6110 5466
rect 6172 5414 6174 5466
rect 6012 5412 6036 5414
rect 6092 5412 6116 5414
rect 6172 5412 6196 5414
rect 5956 5392 6252 5412
rect 5956 4380 6252 4400
rect 6012 4378 6036 4380
rect 6092 4378 6116 4380
rect 6172 4378 6196 4380
rect 6034 4326 6036 4378
rect 6098 4326 6110 4378
rect 6172 4326 6174 4378
rect 6012 4324 6036 4326
rect 6092 4324 6116 4326
rect 6172 4324 6196 4326
rect 5956 4304 6252 4324
rect 5078 3632 5134 3641
rect 5078 3567 5134 3576
rect 5092 800 5120 3567
rect 5956 3292 6252 3312
rect 6012 3290 6036 3292
rect 6092 3290 6116 3292
rect 6172 3290 6196 3292
rect 6034 3238 6036 3290
rect 6098 3238 6110 3290
rect 6172 3238 6174 3290
rect 6012 3236 6036 3238
rect 6092 3236 6116 3238
rect 6172 3236 6196 3238
rect 5956 3216 6252 3236
rect 5956 2204 6252 2224
rect 6012 2202 6036 2204
rect 6092 2202 6116 2204
rect 6172 2202 6196 2204
rect 6034 2150 6036 2202
rect 6098 2150 6110 2202
rect 6172 2150 6174 2202
rect 6012 2148 6036 2150
rect 6092 2148 6116 2150
rect 6172 2148 6196 2150
rect 5956 2128 6252 2148
rect 6288 1986 6316 7375
rect 6918 3360 6974 3369
rect 6918 3295 6974 3304
rect 6012 1958 6316 1986
rect 6012 800 6040 1958
rect 6932 800 6960 3295
rect 7378 3224 7434 3233
rect 7378 3159 7434 3168
rect 7392 800 7420 3159
rect 8312 800 8340 7511
rect 9048 7041 9076 8298
rect 9128 8288 9180 8294
rect 9128 8230 9180 8236
rect 9140 8090 9168 8230
rect 9784 8090 9812 8996
rect 9876 8362 9904 9030
rect 10324 8978 10376 8984
rect 10336 8634 10364 8978
rect 10612 8634 10640 12174
rect 10796 11286 10824 13194
rect 11072 13190 11100 13246
rect 11060 13184 11112 13190
rect 11060 13126 11112 13132
rect 11072 12782 11100 13126
rect 11060 12776 11112 12782
rect 11060 12718 11112 12724
rect 11348 12646 11376 15846
rect 11440 15473 11468 17167
rect 11426 15464 11482 15473
rect 11426 15399 11482 15408
rect 11428 14816 11480 14822
rect 11428 14758 11480 14764
rect 11336 12640 11388 12646
rect 11336 12582 11388 12588
rect 10956 12540 11252 12560
rect 11012 12538 11036 12540
rect 11092 12538 11116 12540
rect 11172 12538 11196 12540
rect 11034 12486 11036 12538
rect 11098 12486 11110 12538
rect 11172 12486 11174 12538
rect 11012 12484 11036 12486
rect 11092 12484 11116 12486
rect 11172 12484 11196 12486
rect 10956 12464 11252 12484
rect 11440 12288 11468 14758
rect 11532 14550 11560 18822
rect 11520 14544 11572 14550
rect 11520 14486 11572 14492
rect 11624 14346 11652 18958
rect 11704 18828 11756 18834
rect 11704 18770 11756 18776
rect 11716 18426 11744 18770
rect 11704 18420 11756 18426
rect 11704 18362 11756 18368
rect 11704 18080 11756 18086
rect 11704 18022 11756 18028
rect 11716 16726 11744 18022
rect 11704 16720 11756 16726
rect 11704 16662 11756 16668
rect 11808 14618 11836 24074
rect 11900 14822 11928 24806
rect 11992 23225 12020 24822
rect 12084 24041 12112 25298
rect 12070 24032 12126 24041
rect 12070 23967 12126 23976
rect 12084 23322 12112 23967
rect 12072 23316 12124 23322
rect 12072 23258 12124 23264
rect 11978 23216 12034 23225
rect 11978 23151 12034 23160
rect 12072 23180 12124 23186
rect 12072 23122 12124 23128
rect 12084 23032 12112 23122
rect 11992 23004 12112 23032
rect 11992 20942 12020 23004
rect 12070 22944 12126 22953
rect 12176 22930 12204 26007
rect 12268 25838 12296 26166
rect 12256 25832 12308 25838
rect 12256 25774 12308 25780
rect 12268 25498 12296 25774
rect 12256 25492 12308 25498
rect 12256 25434 12308 25440
rect 12256 25356 12308 25362
rect 12360 25344 12388 26386
rect 12452 25378 12480 26454
rect 12544 26081 12572 28154
rect 12728 28150 12756 28562
rect 12716 28144 12768 28150
rect 12716 28086 12768 28092
rect 12714 27840 12770 27849
rect 12714 27775 12770 27784
rect 12622 27296 12678 27305
rect 12622 27231 12678 27240
rect 12636 26926 12664 27231
rect 12624 26920 12676 26926
rect 12624 26862 12676 26868
rect 12728 26790 12756 27775
rect 12820 27130 12848 31311
rect 12912 30569 12940 31894
rect 12898 30560 12954 30569
rect 12898 30495 12954 30504
rect 12912 30394 12940 30495
rect 12900 30388 12952 30394
rect 12900 30330 12952 30336
rect 12898 30288 12954 30297
rect 12898 30223 12954 30232
rect 12912 29782 12940 30223
rect 12900 29776 12952 29782
rect 12900 29718 12952 29724
rect 12912 29617 12940 29718
rect 12898 29608 12954 29617
rect 12898 29543 12954 29552
rect 12808 27124 12860 27130
rect 12808 27066 12860 27072
rect 12806 27024 12862 27033
rect 12806 26959 12862 26968
rect 12820 26858 12848 26959
rect 12808 26852 12860 26858
rect 12808 26794 12860 26800
rect 12716 26784 12768 26790
rect 12912 26738 12940 29543
rect 12716 26726 12768 26732
rect 12728 26586 12756 26726
rect 12820 26710 12940 26738
rect 12716 26580 12768 26586
rect 12716 26522 12768 26528
rect 12624 26444 12676 26450
rect 12624 26386 12676 26392
rect 12530 26072 12586 26081
rect 12530 26007 12586 26016
rect 12636 25906 12664 26386
rect 12716 26240 12768 26246
rect 12716 26182 12768 26188
rect 12624 25900 12676 25906
rect 12624 25842 12676 25848
rect 12728 25786 12756 26182
rect 12636 25758 12756 25786
rect 12452 25350 12572 25378
rect 12308 25316 12388 25344
rect 12256 25298 12308 25304
rect 12268 24410 12296 25298
rect 12438 24712 12494 24721
rect 12438 24647 12440 24656
rect 12492 24647 12494 24656
rect 12440 24618 12492 24624
rect 12544 24410 12572 25350
rect 12256 24404 12308 24410
rect 12256 24346 12308 24352
rect 12532 24404 12584 24410
rect 12532 24346 12584 24352
rect 12256 23792 12308 23798
rect 12256 23734 12308 23740
rect 12268 23526 12296 23734
rect 12348 23656 12400 23662
rect 12348 23598 12400 23604
rect 12256 23520 12308 23526
rect 12256 23462 12308 23468
rect 12360 23254 12388 23598
rect 12348 23248 12400 23254
rect 12348 23190 12400 23196
rect 12532 23180 12584 23186
rect 12532 23122 12584 23128
rect 12176 22902 12388 22930
rect 12070 22879 12126 22888
rect 12084 22794 12112 22879
rect 12084 22766 12204 22794
rect 12072 22092 12124 22098
rect 12072 22034 12124 22040
rect 12084 21690 12112 22034
rect 12072 21684 12124 21690
rect 12072 21626 12124 21632
rect 12072 21072 12124 21078
rect 12072 21014 12124 21020
rect 11980 20936 12032 20942
rect 11980 20878 12032 20884
rect 11980 20800 12032 20806
rect 11980 20742 12032 20748
rect 11992 18426 12020 20742
rect 11980 18420 12032 18426
rect 11980 18362 12032 18368
rect 11980 18080 12032 18086
rect 11980 18022 12032 18028
rect 11992 16590 12020 18022
rect 12084 16726 12112 21014
rect 12176 19922 12204 22766
rect 12254 22536 12310 22545
rect 12254 22471 12310 22480
rect 12268 22098 12296 22471
rect 12360 22273 12388 22902
rect 12438 22672 12494 22681
rect 12438 22607 12440 22616
rect 12492 22607 12494 22616
rect 12440 22578 12492 22584
rect 12346 22264 12402 22273
rect 12544 22250 12572 23122
rect 12636 22710 12664 25758
rect 12716 25356 12768 25362
rect 12716 25298 12768 25304
rect 12728 24750 12756 25298
rect 12716 24744 12768 24750
rect 12716 24686 12768 24692
rect 12728 24410 12756 24686
rect 12716 24404 12768 24410
rect 12716 24346 12768 24352
rect 12624 22704 12676 22710
rect 12624 22646 12676 22652
rect 12346 22199 12402 22208
rect 12452 22222 12572 22250
rect 12256 22092 12308 22098
rect 12256 22034 12308 22040
rect 12452 21894 12480 22222
rect 12256 21888 12308 21894
rect 12256 21830 12308 21836
rect 12440 21888 12492 21894
rect 12440 21830 12492 21836
rect 12716 21888 12768 21894
rect 12716 21830 12768 21836
rect 12268 21350 12296 21830
rect 12624 21684 12676 21690
rect 12624 21626 12676 21632
rect 12440 21480 12492 21486
rect 12440 21422 12492 21428
rect 12256 21344 12308 21350
rect 12256 21286 12308 21292
rect 12254 20904 12310 20913
rect 12254 20839 12256 20848
rect 12308 20839 12310 20848
rect 12256 20810 12308 20816
rect 12452 19922 12480 21422
rect 12636 20534 12664 21626
rect 12728 21486 12756 21830
rect 12716 21480 12768 21486
rect 12716 21422 12768 21428
rect 12624 20528 12676 20534
rect 12624 20470 12676 20476
rect 12164 19916 12216 19922
rect 12440 19916 12492 19922
rect 12164 19858 12216 19864
rect 12268 19876 12440 19904
rect 12176 19514 12204 19858
rect 12164 19508 12216 19514
rect 12164 19450 12216 19456
rect 12176 19310 12204 19450
rect 12164 19304 12216 19310
rect 12164 19246 12216 19252
rect 12268 19242 12296 19876
rect 12440 19858 12492 19864
rect 12624 19848 12676 19854
rect 12624 19790 12676 19796
rect 12440 19372 12492 19378
rect 12440 19314 12492 19320
rect 12256 19236 12308 19242
rect 12256 19178 12308 19184
rect 12164 19168 12216 19174
rect 12452 19156 12480 19314
rect 12636 19292 12664 19790
rect 12636 19264 12756 19292
rect 12164 19110 12216 19116
rect 12360 19128 12480 19156
rect 12624 19168 12676 19174
rect 12176 18986 12204 19110
rect 12176 18958 12296 18986
rect 12164 17672 12216 17678
rect 12164 17614 12216 17620
rect 12176 17338 12204 17614
rect 12164 17332 12216 17338
rect 12164 17274 12216 17280
rect 12072 16720 12124 16726
rect 12072 16662 12124 16668
rect 11980 16584 12032 16590
rect 11980 16526 12032 16532
rect 11992 15978 12020 16526
rect 11980 15972 12032 15978
rect 11980 15914 12032 15920
rect 11888 14816 11940 14822
rect 11888 14758 11940 14764
rect 11796 14612 11848 14618
rect 11796 14554 11848 14560
rect 11808 14498 11836 14554
rect 11716 14470 11836 14498
rect 11612 14340 11664 14346
rect 11612 14282 11664 14288
rect 11716 12306 11744 14470
rect 11992 14260 12020 15914
rect 12268 15609 12296 18958
rect 12360 18816 12388 19128
rect 12624 19110 12676 19116
rect 12440 18828 12492 18834
rect 12360 18788 12440 18816
rect 12360 17882 12388 18788
rect 12440 18770 12492 18776
rect 12440 18692 12492 18698
rect 12440 18634 12492 18640
rect 12348 17876 12400 17882
rect 12348 17818 12400 17824
rect 12452 17105 12480 18634
rect 12532 17740 12584 17746
rect 12532 17682 12584 17688
rect 12438 17096 12494 17105
rect 12438 17031 12494 17040
rect 12544 16658 12572 17682
rect 12636 17678 12664 19110
rect 12728 18970 12756 19264
rect 12716 18964 12768 18970
rect 12716 18906 12768 18912
rect 12716 18760 12768 18766
rect 12716 18702 12768 18708
rect 12728 18193 12756 18702
rect 12714 18184 12770 18193
rect 12714 18119 12770 18128
rect 12624 17672 12676 17678
rect 12624 17614 12676 17620
rect 12716 17128 12768 17134
rect 12716 17070 12768 17076
rect 12728 16726 12756 17070
rect 12716 16720 12768 16726
rect 12716 16662 12768 16668
rect 12532 16652 12584 16658
rect 12532 16594 12584 16600
rect 12544 16017 12572 16594
rect 12530 16008 12586 16017
rect 12530 15943 12586 15952
rect 12254 15600 12310 15609
rect 12438 15600 12494 15609
rect 12254 15535 12310 15544
rect 12348 15564 12400 15570
rect 12438 15535 12494 15544
rect 12348 15506 12400 15512
rect 12360 15162 12388 15506
rect 12348 15156 12400 15162
rect 12348 15098 12400 15104
rect 12348 14408 12400 14414
rect 12348 14350 12400 14356
rect 11808 14232 12020 14260
rect 11704 12300 11756 12306
rect 11440 12260 11560 12288
rect 11428 12164 11480 12170
rect 11428 12106 11480 12112
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10888 11354 10916 11630
rect 11336 11620 11388 11626
rect 11336 11562 11388 11568
rect 10956 11452 11252 11472
rect 11012 11450 11036 11452
rect 11092 11450 11116 11452
rect 11172 11450 11196 11452
rect 11034 11398 11036 11450
rect 11098 11398 11110 11450
rect 11172 11398 11174 11450
rect 11012 11396 11036 11398
rect 11092 11396 11116 11398
rect 11172 11396 11196 11398
rect 10956 11376 11252 11396
rect 10876 11348 10928 11354
rect 10876 11290 10928 11296
rect 11348 11286 11376 11562
rect 10784 11280 10836 11286
rect 10784 11222 10836 11228
rect 11336 11280 11388 11286
rect 11336 11222 11388 11228
rect 10796 10810 10824 11222
rect 10784 10804 10836 10810
rect 10784 10746 10836 10752
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 10956 10364 11252 10384
rect 11012 10362 11036 10364
rect 11092 10362 11116 10364
rect 11172 10362 11196 10364
rect 11034 10310 11036 10362
rect 11098 10310 11110 10362
rect 11172 10310 11174 10362
rect 11012 10308 11036 10310
rect 11092 10308 11116 10310
rect 11172 10308 11196 10310
rect 10956 10288 11252 10308
rect 10956 9276 11252 9296
rect 11012 9274 11036 9276
rect 11092 9274 11116 9276
rect 11172 9274 11196 9276
rect 11034 9222 11036 9274
rect 11098 9222 11110 9274
rect 11172 9222 11174 9274
rect 11012 9220 11036 9222
rect 11092 9220 11116 9222
rect 11172 9220 11196 9222
rect 10956 9200 11252 9220
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10600 8628 10652 8634
rect 10600 8570 10652 8576
rect 10244 8430 10272 8570
rect 10232 8424 10284 8430
rect 10232 8366 10284 8372
rect 9864 8356 9916 8362
rect 9864 8298 9916 8304
rect 9128 8084 9180 8090
rect 9128 8026 9180 8032
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9876 7993 9904 8298
rect 10956 8188 11252 8208
rect 11012 8186 11036 8188
rect 11092 8186 11116 8188
rect 11172 8186 11196 8188
rect 11034 8134 11036 8186
rect 11098 8134 11110 8186
rect 11172 8134 11174 8186
rect 11012 8132 11036 8134
rect 11092 8132 11116 8134
rect 11172 8132 11196 8134
rect 10956 8112 11252 8132
rect 9862 7984 9918 7993
rect 9862 7919 9918 7928
rect 11060 7948 11112 7954
rect 11060 7890 11112 7896
rect 11072 7478 11100 7890
rect 11060 7472 11112 7478
rect 11060 7414 11112 7420
rect 11072 7290 11100 7414
rect 10888 7262 11100 7290
rect 9034 7032 9090 7041
rect 9034 6967 9090 6976
rect 9218 5536 9274 5545
rect 9218 5471 9274 5480
rect 9232 800 9260 5471
rect 10888 4690 10916 7262
rect 10956 7100 11252 7120
rect 11012 7098 11036 7100
rect 11092 7098 11116 7100
rect 11172 7098 11196 7100
rect 11034 7046 11036 7098
rect 11098 7046 11110 7098
rect 11172 7046 11174 7098
rect 11012 7044 11036 7046
rect 11092 7044 11116 7046
rect 11172 7044 11196 7046
rect 10956 7024 11252 7044
rect 10956 6012 11252 6032
rect 11012 6010 11036 6012
rect 11092 6010 11116 6012
rect 11172 6010 11196 6012
rect 11034 5958 11036 6010
rect 11098 5958 11110 6010
rect 11172 5958 11174 6010
rect 11012 5956 11036 5958
rect 11092 5956 11116 5958
rect 11172 5956 11196 5958
rect 10956 5936 11252 5956
rect 10956 4924 11252 4944
rect 11012 4922 11036 4924
rect 11092 4922 11116 4924
rect 11172 4922 11196 4924
rect 11034 4870 11036 4922
rect 11098 4870 11110 4922
rect 11172 4870 11174 4922
rect 11012 4868 11036 4870
rect 11092 4868 11116 4870
rect 11172 4868 11196 4870
rect 10956 4848 11252 4868
rect 10876 4684 10928 4690
rect 10876 4626 10928 4632
rect 10888 4146 10916 4626
rect 10876 4140 10928 4146
rect 10876 4082 10928 4088
rect 10888 3754 10916 4082
rect 10956 3836 11252 3856
rect 11012 3834 11036 3836
rect 11092 3834 11116 3836
rect 11172 3834 11196 3836
rect 11034 3782 11036 3834
rect 11098 3782 11110 3834
rect 11172 3782 11174 3834
rect 11012 3780 11036 3782
rect 11092 3780 11116 3782
rect 11172 3780 11196 3782
rect 10956 3760 11252 3780
rect 10796 3738 10916 3754
rect 9864 3732 9916 3738
rect 9864 3674 9916 3680
rect 10784 3732 10916 3738
rect 10836 3726 10916 3732
rect 10784 3674 10836 3680
rect 9876 2990 9904 3674
rect 10600 3528 10652 3534
rect 10600 3470 10652 3476
rect 10140 3052 10192 3058
rect 10140 2994 10192 3000
rect 9864 2984 9916 2990
rect 9864 2926 9916 2932
rect 10152 800 10180 2994
rect 10612 2310 10640 3470
rect 10796 2650 10824 3674
rect 11348 3194 11376 10746
rect 11440 5370 11468 12106
rect 11532 11150 11560 12260
rect 11704 12242 11756 12248
rect 11716 11354 11744 12242
rect 11704 11348 11756 11354
rect 11704 11290 11756 11296
rect 11520 11144 11572 11150
rect 11520 11086 11572 11092
rect 11532 10810 11560 11086
rect 11610 10840 11666 10849
rect 11520 10804 11572 10810
rect 11610 10775 11666 10784
rect 11520 10746 11572 10752
rect 11624 9110 11652 10775
rect 11612 9104 11664 9110
rect 11612 9046 11664 9052
rect 11624 8566 11652 9046
rect 11612 8560 11664 8566
rect 11612 8502 11664 8508
rect 11624 7954 11652 8502
rect 11612 7948 11664 7954
rect 11612 7890 11664 7896
rect 11624 7546 11652 7890
rect 11612 7540 11664 7546
rect 11612 7482 11664 7488
rect 11428 5364 11480 5370
rect 11428 5306 11480 5312
rect 11520 4684 11572 4690
rect 11520 4626 11572 4632
rect 11532 4010 11560 4626
rect 11520 4004 11572 4010
rect 11520 3946 11572 3952
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 10956 2748 11252 2768
rect 11012 2746 11036 2748
rect 11092 2746 11116 2748
rect 11172 2746 11196 2748
rect 11034 2694 11036 2746
rect 11098 2694 11110 2746
rect 11172 2694 11174 2746
rect 11012 2692 11036 2694
rect 11092 2692 11116 2694
rect 11172 2692 11196 2694
rect 10956 2672 11252 2692
rect 10784 2644 10836 2650
rect 10784 2586 10836 2592
rect 10600 2304 10652 2310
rect 10600 2246 10652 2252
rect 10612 800 10640 2246
rect 11532 800 11560 3946
rect 11808 3738 11836 14232
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 12176 13870 12204 14010
rect 12164 13864 12216 13870
rect 12164 13806 12216 13812
rect 11978 13288 12034 13297
rect 11978 13223 12034 13232
rect 11992 12306 12020 13223
rect 11980 12300 12032 12306
rect 11980 12242 12032 12248
rect 11992 11898 12020 12242
rect 11980 11892 12032 11898
rect 11980 11834 12032 11840
rect 12176 11762 12204 13806
rect 12256 13388 12308 13394
rect 12256 13330 12308 13336
rect 12268 12986 12296 13330
rect 12360 13326 12388 14350
rect 12348 13320 12400 13326
rect 12348 13262 12400 13268
rect 12348 13184 12400 13190
rect 12348 13126 12400 13132
rect 12256 12980 12308 12986
rect 12256 12922 12308 12928
rect 12360 12374 12388 13126
rect 12348 12368 12400 12374
rect 12348 12310 12400 12316
rect 12164 11756 12216 11762
rect 12164 11698 12216 11704
rect 12360 11354 12388 12310
rect 12452 11694 12480 15535
rect 12622 15056 12678 15065
rect 12622 14991 12678 15000
rect 12636 14958 12664 14991
rect 12624 14952 12676 14958
rect 12624 14894 12676 14900
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12636 12442 12664 12582
rect 12624 12436 12676 12442
rect 12624 12378 12676 12384
rect 12532 12232 12584 12238
rect 12532 12174 12584 12180
rect 12544 11830 12572 12174
rect 12532 11824 12584 11830
rect 12532 11766 12584 11772
rect 12636 11694 12664 12378
rect 12440 11688 12492 11694
rect 12440 11630 12492 11636
rect 12624 11688 12676 11694
rect 12624 11630 12676 11636
rect 12452 11354 12480 11630
rect 12636 11354 12664 11630
rect 12348 11348 12400 11354
rect 12348 11290 12400 11296
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12624 11348 12676 11354
rect 12624 11290 12676 11296
rect 12728 11234 12756 16662
rect 12820 13870 12848 26710
rect 13004 25838 13032 32166
rect 13096 31754 13124 32263
rect 13188 31890 13216 37674
rect 13280 36961 13308 41806
rect 13464 39953 13492 44134
rect 13924 43908 13952 45494
rect 14016 45354 14044 47110
rect 14108 46170 14136 47194
rect 14384 47138 14412 52142
rect 14462 50960 14518 50969
rect 14462 50895 14518 50904
rect 14476 50726 14504 50895
rect 14464 50720 14516 50726
rect 14464 50662 14516 50668
rect 14464 47796 14516 47802
rect 14464 47738 14516 47744
rect 14200 47122 14412 47138
rect 14476 47122 14504 47738
rect 14188 47116 14412 47122
rect 14240 47110 14412 47116
rect 14464 47116 14516 47122
rect 14188 47058 14240 47064
rect 14464 47058 14516 47064
rect 14200 46374 14228 47058
rect 14476 46714 14504 47058
rect 14464 46708 14516 46714
rect 14464 46650 14516 46656
rect 14188 46368 14240 46374
rect 14188 46310 14240 46316
rect 14096 46164 14148 46170
rect 14096 46106 14148 46112
rect 14200 45966 14228 46310
rect 14568 46186 14596 55383
rect 14740 55344 14792 55350
rect 14740 55286 14792 55292
rect 14648 55276 14700 55282
rect 14648 55218 14700 55224
rect 14660 54806 14688 55218
rect 14648 54800 14700 54806
rect 14648 54742 14700 54748
rect 14752 54670 14780 55286
rect 14844 55282 14872 55830
rect 14936 55622 14964 56782
rect 15108 56704 15160 56710
rect 15108 56646 15160 56652
rect 15120 56438 15148 56646
rect 15212 56506 15240 57854
rect 15200 56500 15252 56506
rect 15200 56442 15252 56448
rect 15016 56432 15068 56438
rect 15016 56374 15068 56380
rect 15108 56432 15160 56438
rect 15108 56374 15160 56380
rect 15028 56166 15056 56374
rect 15120 56234 15148 56374
rect 15200 56364 15252 56370
rect 15200 56306 15252 56312
rect 15108 56228 15160 56234
rect 15108 56170 15160 56176
rect 15016 56160 15068 56166
rect 15016 56102 15068 56108
rect 14924 55616 14976 55622
rect 14924 55558 14976 55564
rect 15028 55418 15056 56102
rect 15108 55616 15160 55622
rect 15108 55558 15160 55564
rect 15016 55412 15068 55418
rect 15016 55354 15068 55360
rect 15120 55321 15148 55558
rect 15212 55350 15240 56306
rect 15200 55344 15252 55350
rect 15106 55312 15162 55321
rect 14832 55276 14884 55282
rect 15200 55286 15252 55292
rect 15106 55247 15162 55256
rect 14832 55218 14884 55224
rect 15108 55072 15160 55078
rect 15108 55014 15160 55020
rect 14922 54904 14978 54913
rect 14922 54839 14978 54848
rect 14832 54732 14884 54738
rect 14832 54674 14884 54680
rect 14740 54664 14792 54670
rect 14740 54606 14792 54612
rect 14844 54126 14872 54674
rect 14936 54602 14964 54839
rect 15016 54800 15068 54806
rect 15016 54742 15068 54748
rect 14924 54596 14976 54602
rect 14924 54538 14976 54544
rect 14832 54120 14884 54126
rect 14832 54062 14884 54068
rect 15028 54058 15056 54742
rect 15120 54534 15148 55014
rect 15304 54874 15332 76774
rect 15672 74798 15700 79200
rect 15956 77276 16252 77296
rect 16012 77274 16036 77276
rect 16092 77274 16116 77276
rect 16172 77274 16196 77276
rect 16034 77222 16036 77274
rect 16098 77222 16110 77274
rect 16172 77222 16174 77274
rect 16012 77220 16036 77222
rect 16092 77220 16116 77222
rect 16172 77220 16196 77222
rect 15956 77200 16252 77220
rect 15956 76188 16252 76208
rect 16012 76186 16036 76188
rect 16092 76186 16116 76188
rect 16172 76186 16196 76188
rect 16034 76134 16036 76186
rect 16098 76134 16110 76186
rect 16172 76134 16174 76186
rect 16012 76132 16036 76134
rect 16092 76132 16116 76134
rect 16172 76132 16196 76134
rect 15956 76112 16252 76132
rect 16592 75857 16620 79200
rect 17512 77178 17540 79200
rect 17500 77172 17552 77178
rect 17500 77114 17552 77120
rect 16578 75848 16634 75857
rect 16578 75783 16634 75792
rect 15956 75100 16252 75120
rect 16012 75098 16036 75100
rect 16092 75098 16116 75100
rect 16172 75098 16196 75100
rect 16034 75046 16036 75098
rect 16098 75046 16110 75098
rect 16172 75046 16174 75098
rect 16012 75044 16036 75046
rect 16092 75044 16116 75046
rect 16172 75044 16196 75046
rect 15956 75024 16252 75044
rect 17972 75002 18000 79200
rect 18602 75304 18658 75313
rect 18602 75239 18658 75248
rect 17960 74996 18012 75002
rect 17960 74938 18012 74944
rect 15660 74792 15712 74798
rect 15660 74734 15712 74740
rect 16488 74792 16540 74798
rect 16488 74734 16540 74740
rect 15956 74012 16252 74032
rect 16012 74010 16036 74012
rect 16092 74010 16116 74012
rect 16172 74010 16196 74012
rect 16034 73958 16036 74010
rect 16098 73958 16110 74010
rect 16172 73958 16174 74010
rect 16012 73956 16036 73958
rect 16092 73956 16116 73958
rect 16172 73956 16196 73958
rect 15956 73936 16252 73956
rect 15956 72924 16252 72944
rect 16012 72922 16036 72924
rect 16092 72922 16116 72924
rect 16172 72922 16196 72924
rect 16034 72870 16036 72922
rect 16098 72870 16110 72922
rect 16172 72870 16174 72922
rect 16012 72868 16036 72870
rect 16092 72868 16116 72870
rect 16172 72868 16196 72870
rect 15956 72848 16252 72868
rect 15956 71836 16252 71856
rect 16012 71834 16036 71836
rect 16092 71834 16116 71836
rect 16172 71834 16196 71836
rect 16034 71782 16036 71834
rect 16098 71782 16110 71834
rect 16172 71782 16174 71834
rect 16012 71780 16036 71782
rect 16092 71780 16116 71782
rect 16172 71780 16196 71782
rect 15956 71760 16252 71780
rect 15956 70748 16252 70768
rect 16012 70746 16036 70748
rect 16092 70746 16116 70748
rect 16172 70746 16196 70748
rect 16034 70694 16036 70746
rect 16098 70694 16110 70746
rect 16172 70694 16174 70746
rect 16012 70692 16036 70694
rect 16092 70692 16116 70694
rect 16172 70692 16196 70694
rect 15956 70672 16252 70692
rect 15956 69660 16252 69680
rect 16012 69658 16036 69660
rect 16092 69658 16116 69660
rect 16172 69658 16196 69660
rect 16034 69606 16036 69658
rect 16098 69606 16110 69658
rect 16172 69606 16174 69658
rect 16012 69604 16036 69606
rect 16092 69604 16116 69606
rect 16172 69604 16196 69606
rect 15956 69584 16252 69604
rect 15956 68572 16252 68592
rect 16012 68570 16036 68572
rect 16092 68570 16116 68572
rect 16172 68570 16196 68572
rect 16034 68518 16036 68570
rect 16098 68518 16110 68570
rect 16172 68518 16174 68570
rect 16012 68516 16036 68518
rect 16092 68516 16116 68518
rect 16172 68516 16196 68518
rect 15956 68496 16252 68516
rect 16396 67652 16448 67658
rect 16396 67594 16448 67600
rect 15382 67552 15438 67561
rect 15382 67487 15438 67496
rect 15396 65142 15424 67487
rect 15956 67484 16252 67504
rect 16012 67482 16036 67484
rect 16092 67482 16116 67484
rect 16172 67482 16196 67484
rect 16034 67430 16036 67482
rect 16098 67430 16110 67482
rect 16172 67430 16174 67482
rect 16012 67428 16036 67430
rect 16092 67428 16116 67430
rect 16172 67428 16196 67430
rect 15956 67408 16252 67428
rect 15956 66396 16252 66416
rect 16012 66394 16036 66396
rect 16092 66394 16116 66396
rect 16172 66394 16196 66396
rect 16034 66342 16036 66394
rect 16098 66342 16110 66394
rect 16172 66342 16174 66394
rect 16012 66340 16036 66342
rect 16092 66340 16116 66342
rect 16172 66340 16196 66342
rect 15956 66320 16252 66340
rect 15476 65952 15528 65958
rect 15476 65894 15528 65900
rect 15384 65136 15436 65142
rect 15384 65078 15436 65084
rect 15488 64977 15516 65894
rect 15660 65612 15712 65618
rect 15660 65554 15712 65560
rect 15844 65612 15896 65618
rect 15844 65554 15896 65560
rect 15474 64968 15530 64977
rect 15672 64938 15700 65554
rect 15856 65006 15884 65554
rect 15956 65308 16252 65328
rect 16012 65306 16036 65308
rect 16092 65306 16116 65308
rect 16172 65306 16196 65308
rect 16034 65254 16036 65306
rect 16098 65254 16110 65306
rect 16172 65254 16174 65306
rect 16012 65252 16036 65254
rect 16092 65252 16116 65254
rect 16172 65252 16196 65254
rect 15956 65232 16252 65252
rect 15844 65000 15896 65006
rect 15844 64942 15896 64948
rect 15474 64903 15530 64912
rect 15660 64932 15712 64938
rect 15488 62490 15516 64903
rect 15660 64874 15712 64880
rect 15672 64326 15700 64874
rect 15856 64394 15884 64942
rect 15844 64388 15896 64394
rect 15844 64330 15896 64336
rect 15660 64320 15712 64326
rect 15660 64262 15712 64268
rect 15672 63986 15700 64262
rect 15660 63980 15712 63986
rect 15660 63922 15712 63928
rect 15672 63442 15700 63922
rect 15752 63776 15804 63782
rect 15752 63718 15804 63724
rect 15764 63442 15792 63718
rect 15660 63436 15712 63442
rect 15660 63378 15712 63384
rect 15752 63436 15804 63442
rect 15752 63378 15804 63384
rect 15568 63368 15620 63374
rect 15568 63310 15620 63316
rect 15580 62694 15608 63310
rect 15672 62830 15700 63378
rect 15660 62824 15712 62830
rect 15660 62766 15712 62772
rect 15764 62762 15792 63378
rect 15752 62756 15804 62762
rect 15752 62698 15804 62704
rect 15568 62688 15620 62694
rect 15568 62630 15620 62636
rect 15476 62484 15528 62490
rect 15476 62426 15528 62432
rect 15476 62348 15528 62354
rect 15476 62290 15528 62296
rect 15384 57928 15436 57934
rect 15382 57896 15384 57905
rect 15436 57896 15438 57905
rect 15382 57831 15438 57840
rect 15384 57792 15436 57798
rect 15384 57734 15436 57740
rect 15292 54868 15344 54874
rect 15292 54810 15344 54816
rect 15292 54732 15344 54738
rect 15292 54674 15344 54680
rect 15200 54664 15252 54670
rect 15200 54606 15252 54612
rect 15108 54528 15160 54534
rect 15108 54470 15160 54476
rect 15120 54262 15148 54470
rect 15108 54256 15160 54262
rect 15108 54198 15160 54204
rect 15212 54097 15240 54606
rect 15198 54088 15254 54097
rect 15016 54052 15068 54058
rect 14936 54012 15016 54040
rect 14738 53680 14794 53689
rect 14738 53615 14794 53624
rect 14752 53446 14780 53615
rect 14740 53440 14792 53446
rect 14646 53408 14702 53417
rect 14740 53382 14792 53388
rect 14646 53343 14702 53352
rect 14660 50998 14688 53343
rect 14752 52630 14780 53382
rect 14830 53000 14886 53009
rect 14830 52935 14886 52944
rect 14740 52624 14792 52630
rect 14740 52566 14792 52572
rect 14740 52488 14792 52494
rect 14740 52430 14792 52436
rect 14648 50992 14700 50998
rect 14648 50934 14700 50940
rect 14660 50522 14688 50934
rect 14648 50516 14700 50522
rect 14648 50458 14700 50464
rect 14648 49768 14700 49774
rect 14648 49710 14700 49716
rect 14660 48686 14688 49710
rect 14752 48686 14780 52430
rect 14844 52358 14872 52935
rect 14832 52352 14884 52358
rect 14832 52294 14884 52300
rect 14844 52154 14872 52294
rect 14832 52148 14884 52154
rect 14832 52090 14884 52096
rect 14936 52034 14964 54012
rect 15198 54023 15200 54032
rect 15016 53994 15068 54000
rect 15252 54023 15254 54032
rect 15200 53994 15252 54000
rect 15212 53582 15240 53994
rect 15200 53576 15252 53582
rect 15200 53518 15252 53524
rect 15108 53440 15160 53446
rect 15106 53408 15108 53417
rect 15160 53408 15162 53417
rect 15106 53343 15162 53352
rect 15212 53242 15240 53518
rect 15304 53514 15332 54674
rect 15292 53508 15344 53514
rect 15292 53450 15344 53456
rect 15200 53236 15252 53242
rect 15200 53178 15252 53184
rect 15016 52896 15068 52902
rect 15016 52838 15068 52844
rect 15200 52896 15252 52902
rect 15200 52838 15252 52844
rect 15028 52737 15056 52838
rect 15014 52728 15070 52737
rect 15014 52663 15070 52672
rect 15108 52692 15160 52698
rect 15028 52630 15056 52663
rect 15108 52634 15160 52640
rect 15016 52624 15068 52630
rect 15016 52566 15068 52572
rect 14844 52006 14964 52034
rect 14844 51610 14872 52006
rect 14832 51604 14884 51610
rect 14832 51546 14884 51552
rect 14924 51536 14976 51542
rect 14924 51478 14976 51484
rect 14832 51264 14884 51270
rect 14832 51206 14884 51212
rect 14844 49094 14872 51206
rect 14936 51066 14964 51478
rect 15028 51105 15056 52566
rect 15120 52154 15148 52634
rect 15212 52601 15240 52838
rect 15198 52592 15254 52601
rect 15198 52527 15254 52536
rect 15200 52488 15252 52494
rect 15304 52476 15332 53450
rect 15252 52448 15332 52476
rect 15200 52430 15252 52436
rect 15108 52148 15160 52154
rect 15108 52090 15160 52096
rect 15212 51270 15240 52430
rect 15290 52048 15346 52057
rect 15290 51983 15292 51992
rect 15344 51983 15346 51992
rect 15292 51954 15344 51960
rect 15292 51808 15344 51814
rect 15292 51750 15344 51756
rect 15200 51264 15252 51270
rect 15120 51224 15200 51252
rect 15014 51096 15070 51105
rect 14924 51060 14976 51066
rect 15014 51031 15070 51040
rect 14924 51002 14976 51008
rect 15120 50862 15148 51224
rect 15200 51206 15252 51212
rect 15198 51096 15254 51105
rect 15198 51031 15254 51040
rect 15108 50856 15160 50862
rect 15108 50798 15160 50804
rect 15212 50454 15240 51031
rect 15304 50794 15332 51750
rect 15292 50788 15344 50794
rect 15292 50730 15344 50736
rect 15292 50516 15344 50522
rect 15292 50458 15344 50464
rect 14924 50448 14976 50454
rect 14924 50390 14976 50396
rect 15200 50448 15252 50454
rect 15200 50390 15252 50396
rect 14936 49366 14964 50390
rect 15108 50312 15160 50318
rect 15108 50254 15160 50260
rect 15016 49700 15068 49706
rect 15016 49642 15068 49648
rect 14924 49360 14976 49366
rect 14924 49302 14976 49308
rect 14832 49088 14884 49094
rect 14832 49030 14884 49036
rect 14648 48680 14700 48686
rect 14648 48622 14700 48628
rect 14740 48680 14792 48686
rect 14740 48622 14792 48628
rect 14752 48346 14780 48622
rect 14740 48340 14792 48346
rect 14740 48282 14792 48288
rect 14832 48204 14884 48210
rect 14832 48146 14884 48152
rect 14648 48068 14700 48074
rect 14648 48010 14700 48016
rect 14660 47802 14688 48010
rect 14648 47796 14700 47802
rect 14648 47738 14700 47744
rect 14738 47424 14794 47433
rect 14738 47359 14794 47368
rect 14752 47258 14780 47359
rect 14740 47252 14792 47258
rect 14740 47194 14792 47200
rect 14568 46158 14688 46186
rect 14188 45960 14240 45966
rect 14188 45902 14240 45908
rect 14464 45824 14516 45830
rect 14464 45766 14516 45772
rect 14476 45422 14504 45766
rect 14096 45416 14148 45422
rect 14096 45358 14148 45364
rect 14464 45416 14516 45422
rect 14464 45358 14516 45364
rect 14004 45348 14056 45354
rect 14004 45290 14056 45296
rect 14108 45234 14136 45358
rect 14556 45348 14608 45354
rect 14556 45290 14608 45296
rect 14016 45206 14136 45234
rect 14016 44198 14044 45206
rect 14568 45082 14596 45290
rect 14556 45076 14608 45082
rect 14556 45018 14608 45024
rect 14004 44192 14056 44198
rect 14004 44134 14056 44140
rect 14016 44033 14044 44134
rect 14002 44024 14058 44033
rect 14002 43959 14058 43968
rect 13740 43880 13952 43908
rect 13740 43246 13768 43880
rect 13820 43308 13872 43314
rect 13820 43250 13872 43256
rect 13728 43240 13780 43246
rect 13728 43182 13780 43188
rect 13832 42838 13860 43250
rect 13820 42832 13872 42838
rect 14660 42809 14688 46158
rect 13820 42774 13872 42780
rect 14646 42800 14702 42809
rect 14646 42735 14702 42744
rect 14844 42265 14872 48146
rect 15028 48074 15056 49642
rect 15120 48872 15148 50254
rect 15304 49978 15332 50458
rect 15292 49972 15344 49978
rect 15292 49914 15344 49920
rect 15292 49768 15344 49774
rect 15290 49736 15292 49745
rect 15344 49736 15346 49745
rect 15290 49671 15346 49680
rect 15292 49292 15344 49298
rect 15292 49234 15344 49240
rect 15304 49201 15332 49234
rect 15290 49192 15346 49201
rect 15290 49127 15346 49136
rect 15292 49088 15344 49094
rect 15292 49030 15344 49036
rect 15200 48884 15252 48890
rect 15120 48844 15200 48872
rect 15200 48826 15252 48832
rect 15108 48612 15160 48618
rect 15108 48554 15160 48560
rect 15120 48260 15148 48554
rect 15120 48232 15240 48260
rect 15016 48068 15068 48074
rect 15016 48010 15068 48016
rect 15108 48068 15160 48074
rect 15108 48010 15160 48016
rect 15016 47456 15068 47462
rect 15016 47398 15068 47404
rect 14924 47184 14976 47190
rect 15028 47161 15056 47398
rect 14924 47126 14976 47132
rect 15014 47152 15070 47161
rect 14936 46714 14964 47126
rect 15014 47087 15070 47096
rect 15028 46714 15056 47087
rect 14924 46708 14976 46714
rect 14924 46650 14976 46656
rect 15016 46708 15068 46714
rect 15016 46650 15068 46656
rect 15120 42276 15148 48010
rect 15212 47802 15240 48232
rect 15304 48074 15332 49030
rect 15292 48068 15344 48074
rect 15292 48010 15344 48016
rect 15200 47796 15252 47802
rect 15200 47738 15252 47744
rect 15212 47054 15240 47738
rect 15200 47048 15252 47054
rect 15200 46990 15252 46996
rect 15212 46578 15240 46990
rect 15200 46572 15252 46578
rect 15200 46514 15252 46520
rect 15396 44180 15424 57734
rect 15488 56545 15516 62290
rect 15580 59430 15608 62630
rect 15660 62484 15712 62490
rect 15660 62426 15712 62432
rect 15672 60722 15700 62426
rect 15856 62422 15884 64330
rect 15956 64220 16252 64240
rect 16012 64218 16036 64220
rect 16092 64218 16116 64220
rect 16172 64218 16196 64220
rect 16034 64166 16036 64218
rect 16098 64166 16110 64218
rect 16172 64166 16174 64218
rect 16012 64164 16036 64166
rect 16092 64164 16116 64166
rect 16172 64164 16196 64166
rect 15956 64144 16252 64164
rect 16212 63912 16264 63918
rect 16264 63860 16344 63866
rect 16212 63854 16344 63860
rect 16224 63838 16344 63854
rect 15956 63132 16252 63152
rect 16012 63130 16036 63132
rect 16092 63130 16116 63132
rect 16172 63130 16196 63132
rect 16034 63078 16036 63130
rect 16098 63078 16110 63130
rect 16172 63078 16174 63130
rect 16012 63076 16036 63078
rect 16092 63076 16116 63078
rect 16172 63076 16196 63078
rect 15956 63056 16252 63076
rect 15844 62416 15896 62422
rect 15844 62358 15896 62364
rect 16316 62354 16344 63838
rect 16304 62348 16356 62354
rect 16304 62290 16356 62296
rect 15956 62044 16252 62064
rect 16012 62042 16036 62044
rect 16092 62042 16116 62044
rect 16172 62042 16196 62044
rect 16034 61990 16036 62042
rect 16098 61990 16110 62042
rect 16172 61990 16174 62042
rect 16012 61988 16036 61990
rect 16092 61988 16116 61990
rect 16172 61988 16196 61990
rect 15956 61968 16252 61988
rect 16316 61606 16344 62290
rect 15844 61600 15896 61606
rect 15844 61542 15896 61548
rect 16304 61600 16356 61606
rect 16304 61542 16356 61548
rect 15660 60716 15712 60722
rect 15660 60658 15712 60664
rect 15660 60308 15712 60314
rect 15660 60250 15712 60256
rect 15568 59424 15620 59430
rect 15568 59366 15620 59372
rect 15672 59208 15700 60250
rect 15752 59492 15804 59498
rect 15752 59434 15804 59440
rect 15580 59180 15700 59208
rect 15580 59022 15608 59180
rect 15660 59084 15712 59090
rect 15660 59026 15712 59032
rect 15568 59016 15620 59022
rect 15568 58958 15620 58964
rect 15580 58682 15608 58958
rect 15568 58676 15620 58682
rect 15568 58618 15620 58624
rect 15672 58478 15700 59026
rect 15660 58472 15712 58478
rect 15660 58414 15712 58420
rect 15568 58336 15620 58342
rect 15568 58278 15620 58284
rect 15474 56536 15530 56545
rect 15474 56471 15530 56480
rect 15580 56386 15608 58278
rect 15672 58070 15700 58414
rect 15764 58138 15792 59434
rect 15752 58132 15804 58138
rect 15752 58074 15804 58080
rect 15660 58064 15712 58070
rect 15660 58006 15712 58012
rect 15764 57866 15792 58074
rect 15752 57860 15804 57866
rect 15752 57802 15804 57808
rect 15764 57390 15792 57802
rect 15752 57384 15804 57390
rect 15752 57326 15804 57332
rect 15660 57316 15712 57322
rect 15660 57258 15712 57264
rect 15488 56358 15608 56386
rect 15488 51406 15516 56358
rect 15568 56160 15620 56166
rect 15568 56102 15620 56108
rect 15580 55622 15608 56102
rect 15568 55616 15620 55622
rect 15568 55558 15620 55564
rect 15568 54868 15620 54874
rect 15568 54810 15620 54816
rect 15580 52426 15608 54810
rect 15568 52420 15620 52426
rect 15568 52362 15620 52368
rect 15568 52148 15620 52154
rect 15568 52090 15620 52096
rect 15476 51400 15528 51406
rect 15476 51342 15528 51348
rect 15476 50720 15528 50726
rect 15580 50697 15608 52090
rect 15476 50662 15528 50668
rect 15566 50688 15622 50697
rect 15488 48929 15516 50662
rect 15566 50623 15622 50632
rect 15568 49904 15620 49910
rect 15568 49846 15620 49852
rect 15474 48920 15530 48929
rect 15474 48855 15530 48864
rect 15476 48816 15528 48822
rect 15476 48758 15528 48764
rect 15488 48385 15516 48758
rect 15474 48376 15530 48385
rect 15474 48311 15530 48320
rect 15476 48068 15528 48074
rect 15476 48010 15528 48016
rect 15488 47122 15516 48010
rect 15476 47116 15528 47122
rect 15476 47058 15528 47064
rect 15488 46034 15516 47058
rect 15580 46458 15608 49846
rect 15672 49178 15700 57258
rect 15752 56772 15804 56778
rect 15752 56714 15804 56720
rect 15764 56681 15792 56714
rect 15750 56672 15806 56681
rect 15750 56607 15806 56616
rect 15750 56536 15806 56545
rect 15750 56471 15806 56480
rect 15764 51252 15792 56471
rect 15856 51377 15884 61542
rect 15956 60956 16252 60976
rect 16012 60954 16036 60956
rect 16092 60954 16116 60956
rect 16172 60954 16196 60956
rect 16034 60902 16036 60954
rect 16098 60902 16110 60954
rect 16172 60902 16174 60954
rect 16012 60900 16036 60902
rect 16092 60900 16116 60902
rect 16172 60900 16196 60902
rect 15956 60880 16252 60900
rect 16212 60580 16264 60586
rect 16212 60522 16264 60528
rect 16224 60314 16252 60522
rect 16212 60308 16264 60314
rect 16212 60250 16264 60256
rect 15956 59868 16252 59888
rect 16012 59866 16036 59868
rect 16092 59866 16116 59868
rect 16172 59866 16196 59868
rect 16034 59814 16036 59866
rect 16098 59814 16110 59866
rect 16172 59814 16174 59866
rect 16012 59812 16036 59814
rect 16092 59812 16116 59814
rect 16172 59812 16196 59814
rect 15956 59792 16252 59812
rect 16212 59560 16264 59566
rect 16210 59528 16212 59537
rect 16264 59528 16266 59537
rect 16210 59463 16266 59472
rect 15956 58780 16252 58800
rect 16012 58778 16036 58780
rect 16092 58778 16116 58780
rect 16172 58778 16196 58780
rect 16034 58726 16036 58778
rect 16098 58726 16110 58778
rect 16172 58726 16174 58778
rect 16012 58724 16036 58726
rect 16092 58724 16116 58726
rect 16172 58724 16196 58726
rect 15956 58704 16252 58724
rect 16210 58576 16266 58585
rect 16210 58511 16266 58520
rect 16224 58478 16252 58511
rect 16212 58472 16264 58478
rect 16212 58414 16264 58420
rect 15956 57692 16252 57712
rect 16012 57690 16036 57692
rect 16092 57690 16116 57692
rect 16172 57690 16196 57692
rect 16034 57638 16036 57690
rect 16098 57638 16110 57690
rect 16172 57638 16174 57690
rect 16012 57636 16036 57638
rect 16092 57636 16116 57638
rect 16172 57636 16196 57638
rect 15956 57616 16252 57636
rect 16212 57248 16264 57254
rect 16212 57190 16264 57196
rect 16224 56778 16252 57190
rect 16212 56772 16264 56778
rect 16212 56714 16264 56720
rect 15956 56604 16252 56624
rect 16012 56602 16036 56604
rect 16092 56602 16116 56604
rect 16172 56602 16196 56604
rect 16034 56550 16036 56602
rect 16098 56550 16110 56602
rect 16172 56550 16174 56602
rect 16012 56548 16036 56550
rect 16092 56548 16116 56550
rect 16172 56548 16196 56550
rect 15956 56528 16252 56548
rect 16120 56364 16172 56370
rect 16120 56306 16172 56312
rect 16132 55962 16160 56306
rect 16212 56160 16264 56166
rect 16212 56102 16264 56108
rect 16120 55956 16172 55962
rect 16120 55898 16172 55904
rect 16224 55894 16252 56102
rect 16212 55888 16264 55894
rect 16212 55830 16264 55836
rect 15956 55516 16252 55536
rect 16012 55514 16036 55516
rect 16092 55514 16116 55516
rect 16172 55514 16196 55516
rect 16034 55462 16036 55514
rect 16098 55462 16110 55514
rect 16172 55462 16174 55514
rect 16012 55460 16036 55462
rect 16092 55460 16116 55462
rect 16172 55460 16196 55462
rect 15956 55440 16252 55460
rect 15936 55344 15988 55350
rect 15936 55286 15988 55292
rect 15948 55078 15976 55286
rect 15936 55072 15988 55078
rect 15936 55014 15988 55020
rect 15948 54602 15976 55014
rect 16316 54670 16344 61542
rect 16304 54664 16356 54670
rect 16304 54606 16356 54612
rect 15936 54596 15988 54602
rect 15936 54538 15988 54544
rect 16304 54528 16356 54534
rect 16304 54470 16356 54476
rect 15956 54428 16252 54448
rect 16012 54426 16036 54428
rect 16092 54426 16116 54428
rect 16172 54426 16196 54428
rect 16034 54374 16036 54426
rect 16098 54374 16110 54426
rect 16172 54374 16174 54426
rect 16012 54372 16036 54374
rect 16092 54372 16116 54374
rect 16172 54372 16196 54374
rect 15956 54352 16252 54372
rect 16028 54256 16080 54262
rect 16026 54224 16028 54233
rect 16080 54224 16082 54233
rect 16026 54159 16082 54168
rect 16120 54120 16172 54126
rect 16120 54062 16172 54068
rect 16132 53514 16160 54062
rect 16212 54052 16264 54058
rect 16212 53994 16264 54000
rect 16224 53650 16252 53994
rect 16212 53644 16264 53650
rect 16212 53586 16264 53592
rect 16120 53508 16172 53514
rect 16120 53450 16172 53456
rect 15956 53340 16252 53360
rect 16012 53338 16036 53340
rect 16092 53338 16116 53340
rect 16172 53338 16196 53340
rect 16034 53286 16036 53338
rect 16098 53286 16110 53338
rect 16172 53286 16174 53338
rect 16012 53284 16036 53286
rect 16092 53284 16116 53286
rect 16172 53284 16196 53286
rect 15956 53264 16252 53284
rect 16316 53038 16344 54470
rect 16304 53032 16356 53038
rect 16304 52974 16356 52980
rect 16316 52698 16344 52974
rect 16304 52692 16356 52698
rect 16304 52634 16356 52640
rect 16304 52556 16356 52562
rect 16304 52498 16356 52504
rect 15956 52252 16252 52272
rect 16012 52250 16036 52252
rect 16092 52250 16116 52252
rect 16172 52250 16196 52252
rect 16034 52198 16036 52250
rect 16098 52198 16110 52250
rect 16172 52198 16174 52250
rect 16012 52196 16036 52198
rect 16092 52196 16116 52198
rect 16172 52196 16196 52198
rect 15956 52176 16252 52196
rect 16120 52012 16172 52018
rect 16120 51954 16172 51960
rect 16028 51876 16080 51882
rect 16028 51818 16080 51824
rect 16040 51474 16068 51818
rect 16132 51474 16160 51954
rect 16316 51814 16344 52498
rect 16304 51808 16356 51814
rect 16304 51750 16356 51756
rect 16028 51468 16080 51474
rect 16028 51410 16080 51416
rect 16120 51468 16172 51474
rect 16120 51410 16172 51416
rect 16304 51400 16356 51406
rect 15842 51368 15898 51377
rect 16304 51342 16356 51348
rect 15842 51303 15898 51312
rect 15764 51224 15884 51252
rect 15752 50516 15804 50522
rect 15752 50458 15804 50464
rect 15764 50386 15792 50458
rect 15752 50380 15804 50386
rect 15752 50322 15804 50328
rect 15752 50176 15804 50182
rect 15752 50118 15804 50124
rect 15764 49609 15792 50118
rect 15750 49600 15806 49609
rect 15750 49535 15806 49544
rect 15764 49366 15792 49535
rect 15752 49360 15804 49366
rect 15752 49302 15804 49308
rect 15672 49150 15792 49178
rect 15660 49088 15712 49094
rect 15660 49030 15712 49036
rect 15672 48346 15700 49030
rect 15660 48340 15712 48346
rect 15660 48282 15712 48288
rect 15672 47598 15700 48282
rect 15764 48278 15792 49150
rect 15752 48272 15804 48278
rect 15752 48214 15804 48220
rect 15752 48136 15804 48142
rect 15752 48078 15804 48084
rect 15660 47592 15712 47598
rect 15660 47534 15712 47540
rect 15580 46430 15700 46458
rect 15764 46442 15792 48078
rect 15568 46368 15620 46374
rect 15566 46336 15568 46345
rect 15620 46336 15622 46345
rect 15566 46271 15622 46280
rect 15568 46096 15620 46102
rect 15568 46038 15620 46044
rect 15476 46028 15528 46034
rect 15476 45970 15528 45976
rect 15488 45626 15516 45970
rect 15476 45620 15528 45626
rect 15476 45562 15528 45568
rect 15580 44538 15608 46038
rect 15672 44849 15700 46430
rect 15752 46436 15804 46442
rect 15752 46378 15804 46384
rect 15764 46034 15792 46378
rect 15752 46028 15804 46034
rect 15752 45970 15804 45976
rect 15764 45082 15792 45970
rect 15752 45076 15804 45082
rect 15752 45018 15804 45024
rect 15658 44840 15714 44849
rect 15658 44775 15714 44784
rect 15568 44532 15620 44538
rect 15568 44474 15620 44480
rect 15396 44152 15516 44180
rect 14830 42256 14886 42265
rect 15120 42248 15240 42276
rect 14830 42191 14886 42200
rect 15106 42120 15162 42129
rect 15106 42055 15108 42064
rect 15160 42055 15162 42064
rect 15108 42026 15160 42032
rect 14004 42016 14056 42022
rect 14004 41958 14056 41964
rect 14016 41857 14044 41958
rect 14002 41848 14058 41857
rect 14002 41783 14058 41792
rect 15106 41168 15162 41177
rect 15106 41103 15162 41112
rect 14188 40588 14240 40594
rect 14188 40530 14240 40536
rect 13912 40384 13964 40390
rect 13912 40326 13964 40332
rect 13450 39944 13506 39953
rect 13450 39879 13506 39888
rect 13636 39840 13688 39846
rect 13634 39808 13636 39817
rect 13688 39808 13690 39817
rect 13634 39743 13690 39752
rect 13544 39500 13596 39506
rect 13544 39442 13596 39448
rect 13728 39500 13780 39506
rect 13728 39442 13780 39448
rect 13556 38894 13584 39442
rect 13544 38888 13596 38894
rect 13542 38856 13544 38865
rect 13596 38856 13598 38865
rect 13542 38791 13598 38800
rect 13556 38418 13584 38791
rect 13740 38457 13768 39442
rect 13820 39296 13872 39302
rect 13820 39238 13872 39244
rect 13726 38448 13782 38457
rect 13544 38412 13596 38418
rect 13726 38383 13782 38392
rect 13544 38354 13596 38360
rect 13360 38208 13412 38214
rect 13360 38150 13412 38156
rect 13266 36952 13322 36961
rect 13266 36887 13322 36896
rect 13372 36854 13400 38150
rect 13542 37768 13598 37777
rect 13542 37703 13598 37712
rect 13556 37398 13584 37703
rect 13636 37460 13688 37466
rect 13636 37402 13688 37408
rect 13544 37392 13596 37398
rect 13544 37334 13596 37340
rect 13450 37224 13506 37233
rect 13450 37159 13506 37168
rect 13360 36848 13412 36854
rect 13360 36790 13412 36796
rect 13372 36417 13400 36790
rect 13358 36408 13414 36417
rect 13358 36343 13414 36352
rect 13360 36236 13412 36242
rect 13360 36178 13412 36184
rect 13372 35562 13400 36178
rect 13360 35556 13412 35562
rect 13360 35498 13412 35504
rect 13268 35216 13320 35222
rect 13268 35158 13320 35164
rect 13280 34649 13308 35158
rect 13266 34640 13322 34649
rect 13266 34575 13268 34584
rect 13320 34575 13322 34584
rect 13268 34546 13320 34552
rect 13268 33992 13320 33998
rect 13268 33934 13320 33940
rect 13280 32434 13308 33934
rect 13268 32428 13320 32434
rect 13268 32370 13320 32376
rect 13280 32065 13308 32370
rect 13266 32056 13322 32065
rect 13266 31991 13322 32000
rect 13372 31958 13400 35498
rect 13360 31952 13412 31958
rect 13360 31894 13412 31900
rect 13176 31884 13228 31890
rect 13176 31826 13228 31832
rect 13084 31748 13136 31754
rect 13084 31690 13136 31696
rect 13082 31648 13138 31657
rect 13082 31583 13138 31592
rect 13096 30870 13124 31583
rect 13188 30938 13216 31826
rect 13360 31816 13412 31822
rect 13360 31758 13412 31764
rect 13372 31482 13400 31758
rect 13360 31476 13412 31482
rect 13360 31418 13412 31424
rect 13360 31272 13412 31278
rect 13360 31214 13412 31220
rect 13176 30932 13228 30938
rect 13176 30874 13228 30880
rect 13084 30864 13136 30870
rect 13084 30806 13136 30812
rect 13174 30832 13230 30841
rect 13174 30767 13176 30776
rect 13228 30767 13230 30776
rect 13176 30738 13228 30744
rect 13268 30728 13320 30734
rect 13372 30705 13400 31214
rect 13268 30670 13320 30676
rect 13358 30696 13414 30705
rect 13082 30560 13138 30569
rect 13082 30495 13138 30504
rect 13096 28762 13124 30495
rect 13176 29844 13228 29850
rect 13176 29786 13228 29792
rect 13188 29102 13216 29786
rect 13280 29714 13308 30670
rect 13464 30666 13492 37159
rect 13544 36372 13596 36378
rect 13544 36314 13596 36320
rect 13556 35068 13584 36314
rect 13648 36310 13676 37402
rect 13728 37392 13780 37398
rect 13728 37334 13780 37340
rect 13740 36922 13768 37334
rect 13728 36916 13780 36922
rect 13728 36858 13780 36864
rect 13728 36712 13780 36718
rect 13832 36700 13860 39238
rect 13780 36672 13860 36700
rect 13728 36654 13780 36660
rect 13636 36304 13688 36310
rect 13636 36246 13688 36252
rect 13818 36272 13874 36281
rect 13818 36207 13874 36216
rect 13636 36168 13688 36174
rect 13636 36110 13688 36116
rect 13648 35193 13676 36110
rect 13832 35562 13860 36207
rect 13924 36038 13952 40326
rect 14200 39982 14228 40530
rect 15120 40186 15148 41103
rect 15108 40180 15160 40186
rect 15108 40122 15160 40128
rect 14188 39976 14240 39982
rect 14188 39918 14240 39924
rect 14096 39432 14148 39438
rect 14096 39374 14148 39380
rect 14108 39098 14136 39374
rect 14096 39092 14148 39098
rect 14096 39034 14148 39040
rect 14200 38758 14228 39918
rect 15016 39296 15068 39302
rect 15016 39238 15068 39244
rect 14924 38888 14976 38894
rect 14924 38830 14976 38836
rect 14188 38752 14240 38758
rect 14188 38694 14240 38700
rect 14004 37868 14056 37874
rect 14004 37810 14056 37816
rect 13912 36032 13964 36038
rect 13912 35974 13964 35980
rect 13820 35556 13872 35562
rect 13820 35498 13872 35504
rect 13832 35465 13860 35498
rect 13912 35488 13964 35494
rect 13818 35456 13874 35465
rect 13912 35430 13964 35436
rect 13818 35391 13874 35400
rect 13726 35320 13782 35329
rect 13726 35255 13782 35264
rect 13634 35184 13690 35193
rect 13634 35119 13690 35128
rect 13556 35040 13676 35068
rect 13648 34592 13676 35040
rect 13556 34564 13676 34592
rect 13556 34202 13584 34564
rect 13634 34504 13690 34513
rect 13634 34439 13690 34448
rect 13544 34196 13596 34202
rect 13544 34138 13596 34144
rect 13556 33658 13584 34138
rect 13544 33652 13596 33658
rect 13544 33594 13596 33600
rect 13544 33516 13596 33522
rect 13544 33458 13596 33464
rect 13556 32881 13584 33458
rect 13542 32872 13598 32881
rect 13542 32807 13598 32816
rect 13556 31958 13584 32807
rect 13544 31952 13596 31958
rect 13648 31929 13676 34439
rect 13544 31894 13596 31900
rect 13634 31920 13690 31929
rect 13634 31855 13690 31864
rect 13740 31822 13768 35255
rect 13820 34944 13872 34950
rect 13820 34886 13872 34892
rect 13832 34785 13860 34886
rect 13818 34776 13874 34785
rect 13818 34711 13874 34720
rect 13820 34468 13872 34474
rect 13820 34410 13872 34416
rect 13832 33674 13860 34410
rect 13924 33844 13952 35430
rect 14016 35086 14044 37810
rect 14200 37670 14228 38694
rect 14648 38412 14700 38418
rect 14648 38354 14700 38360
rect 14464 38276 14516 38282
rect 14464 38218 14516 38224
rect 14372 38208 14424 38214
rect 14372 38150 14424 38156
rect 14280 37800 14332 37806
rect 14280 37742 14332 37748
rect 14188 37664 14240 37670
rect 14292 37641 14320 37742
rect 14188 37606 14240 37612
rect 14278 37632 14334 37641
rect 14200 36718 14228 37606
rect 14278 37567 14334 37576
rect 14188 36712 14240 36718
rect 14188 36654 14240 36660
rect 14280 36576 14332 36582
rect 14280 36518 14332 36524
rect 14096 36304 14148 36310
rect 14096 36246 14148 36252
rect 14004 35080 14056 35086
rect 14004 35022 14056 35028
rect 14016 34105 14044 35022
rect 14002 34096 14058 34105
rect 14002 34031 14058 34040
rect 14004 33856 14056 33862
rect 13924 33816 14004 33844
rect 14004 33798 14056 33804
rect 13832 33646 13952 33674
rect 13820 32904 13872 32910
rect 13924 32881 13952 33646
rect 13820 32846 13872 32852
rect 13910 32872 13966 32881
rect 13728 31816 13780 31822
rect 13542 31784 13598 31793
rect 13728 31758 13780 31764
rect 13542 31719 13598 31728
rect 13636 31748 13688 31754
rect 13358 30631 13414 30640
rect 13452 30660 13504 30666
rect 13452 30602 13504 30608
rect 13360 30592 13412 30598
rect 13412 30540 13492 30546
rect 13360 30534 13492 30540
rect 13372 30518 13492 30534
rect 13360 30252 13412 30258
rect 13360 30194 13412 30200
rect 13372 29850 13400 30194
rect 13360 29844 13412 29850
rect 13360 29786 13412 29792
rect 13268 29708 13320 29714
rect 13268 29650 13320 29656
rect 13176 29096 13228 29102
rect 13174 29064 13176 29073
rect 13228 29064 13230 29073
rect 13174 28999 13230 29008
rect 13280 28966 13308 29650
rect 13360 29572 13412 29578
rect 13360 29514 13412 29520
rect 13268 28960 13320 28966
rect 13268 28902 13320 28908
rect 13084 28756 13136 28762
rect 13084 28698 13136 28704
rect 13176 28756 13228 28762
rect 13176 28698 13228 28704
rect 13188 28014 13216 28698
rect 13280 28694 13308 28902
rect 13268 28688 13320 28694
rect 13268 28630 13320 28636
rect 13268 28552 13320 28558
rect 13266 28520 13268 28529
rect 13320 28520 13322 28529
rect 13372 28490 13400 29514
rect 13266 28455 13322 28464
rect 13360 28484 13412 28490
rect 13360 28426 13412 28432
rect 13358 28112 13414 28121
rect 13358 28047 13414 28056
rect 13176 28008 13228 28014
rect 13176 27950 13228 27956
rect 13084 27940 13136 27946
rect 13084 27882 13136 27888
rect 12992 25832 13044 25838
rect 12992 25774 13044 25780
rect 12900 24744 12952 24750
rect 12900 24686 12952 24692
rect 12912 24342 12940 24686
rect 12992 24608 13044 24614
rect 12992 24550 13044 24556
rect 12900 24336 12952 24342
rect 12900 24278 12952 24284
rect 13004 23730 13032 24550
rect 12992 23724 13044 23730
rect 12992 23666 13044 23672
rect 12900 22636 12952 22642
rect 12900 22578 12952 22584
rect 12912 22234 12940 22578
rect 12992 22500 13044 22506
rect 12992 22442 13044 22448
rect 12900 22228 12952 22234
rect 12900 22170 12952 22176
rect 13004 21010 13032 22442
rect 13096 21146 13124 27882
rect 13372 27674 13400 28047
rect 13360 27668 13412 27674
rect 13360 27610 13412 27616
rect 13176 27464 13228 27470
rect 13176 27406 13228 27412
rect 13188 26761 13216 27406
rect 13360 27124 13412 27130
rect 13360 27066 13412 27072
rect 13174 26752 13230 26761
rect 13230 26710 13308 26738
rect 13174 26687 13230 26696
rect 13176 26580 13228 26586
rect 13176 26522 13228 26528
rect 13188 24274 13216 26522
rect 13280 26450 13308 26710
rect 13372 26518 13400 27066
rect 13360 26512 13412 26518
rect 13360 26454 13412 26460
rect 13268 26444 13320 26450
rect 13268 26386 13320 26392
rect 13280 25906 13308 26386
rect 13360 26376 13412 26382
rect 13360 26318 13412 26324
rect 13268 25900 13320 25906
rect 13268 25842 13320 25848
rect 13268 25220 13320 25226
rect 13268 25162 13320 25168
rect 13280 24750 13308 25162
rect 13372 25158 13400 26318
rect 13360 25152 13412 25158
rect 13360 25094 13412 25100
rect 13372 24818 13400 25094
rect 13360 24812 13412 24818
rect 13360 24754 13412 24760
rect 13268 24744 13320 24750
rect 13268 24686 13320 24692
rect 13176 24268 13228 24274
rect 13176 24210 13228 24216
rect 13268 24268 13320 24274
rect 13268 24210 13320 24216
rect 13188 23798 13216 24210
rect 13176 23792 13228 23798
rect 13176 23734 13228 23740
rect 13188 23186 13216 23734
rect 13176 23180 13228 23186
rect 13176 23122 13228 23128
rect 13280 22982 13308 24210
rect 13464 23594 13492 30518
rect 13556 30122 13584 31719
rect 13636 31690 13688 31696
rect 13648 30666 13676 31690
rect 13832 31226 13860 32846
rect 13910 32807 13966 32816
rect 13910 32736 13966 32745
rect 13910 32671 13966 32680
rect 13924 31890 13952 32671
rect 14016 32230 14044 33798
rect 14108 33046 14136 36246
rect 14292 35766 14320 36518
rect 14280 35760 14332 35766
rect 14280 35702 14332 35708
rect 14188 35624 14240 35630
rect 14188 35566 14240 35572
rect 14200 35290 14228 35566
rect 14188 35284 14240 35290
rect 14188 35226 14240 35232
rect 14292 35170 14320 35702
rect 14200 35142 14320 35170
rect 14200 34746 14228 35142
rect 14280 35080 14332 35086
rect 14280 35022 14332 35028
rect 14188 34740 14240 34746
rect 14188 34682 14240 34688
rect 14292 34626 14320 35022
rect 14200 34598 14320 34626
rect 14200 34134 14228 34598
rect 14384 34542 14412 38150
rect 14476 37738 14504 38218
rect 14660 38010 14688 38354
rect 14648 38004 14700 38010
rect 14648 37946 14700 37952
rect 14464 37732 14516 37738
rect 14464 37674 14516 37680
rect 14476 37641 14504 37674
rect 14936 37670 14964 38830
rect 15028 38350 15056 39238
rect 15108 38820 15160 38826
rect 15108 38762 15160 38768
rect 15120 38486 15148 38762
rect 15108 38480 15160 38486
rect 15108 38422 15160 38428
rect 15016 38344 15068 38350
rect 15016 38286 15068 38292
rect 15108 38276 15160 38282
rect 15108 38218 15160 38224
rect 15016 38208 15068 38214
rect 15016 38150 15068 38156
rect 14924 37664 14976 37670
rect 14462 37632 14518 37641
rect 14924 37606 14976 37612
rect 14462 37567 14518 37576
rect 14922 37496 14978 37505
rect 14922 37431 14924 37440
rect 14976 37431 14978 37440
rect 14924 37402 14976 37408
rect 15028 37398 15056 38150
rect 15016 37392 15068 37398
rect 14646 37360 14702 37369
rect 15016 37334 15068 37340
rect 14646 37295 14702 37304
rect 14556 36780 14608 36786
rect 14476 36740 14556 36768
rect 14372 34536 14424 34542
rect 14292 34496 14372 34524
rect 14292 34134 14320 34496
rect 14372 34478 14424 34484
rect 14372 34196 14424 34202
rect 14372 34138 14424 34144
rect 14188 34128 14240 34134
rect 14188 34070 14240 34076
rect 14280 34128 14332 34134
rect 14280 34070 14332 34076
rect 14200 33289 14228 34070
rect 14384 33318 14412 34138
rect 14372 33312 14424 33318
rect 14186 33280 14242 33289
rect 14372 33254 14424 33260
rect 14186 33215 14242 33224
rect 14280 33108 14332 33114
rect 14280 33050 14332 33056
rect 14096 33040 14148 33046
rect 14096 32982 14148 32988
rect 14188 32972 14240 32978
rect 14188 32914 14240 32920
rect 14096 32836 14148 32842
rect 14096 32778 14148 32784
rect 14004 32224 14056 32230
rect 14004 32166 14056 32172
rect 14016 32026 14044 32166
rect 14004 32020 14056 32026
rect 14004 31962 14056 31968
rect 13912 31884 13964 31890
rect 13912 31826 13964 31832
rect 14004 31884 14056 31890
rect 14004 31826 14056 31832
rect 13924 31482 13952 31826
rect 13912 31476 13964 31482
rect 13912 31418 13964 31424
rect 13728 31204 13780 31210
rect 13832 31198 13952 31226
rect 13728 31146 13780 31152
rect 13636 30660 13688 30666
rect 13636 30602 13688 30608
rect 13544 30116 13596 30122
rect 13544 30058 13596 30064
rect 13636 29708 13688 29714
rect 13636 29650 13688 29656
rect 13544 29572 13596 29578
rect 13544 29514 13596 29520
rect 13556 26994 13584 29514
rect 13648 29170 13676 29650
rect 13740 29345 13768 31146
rect 13820 31136 13872 31142
rect 13820 31078 13872 31084
rect 13832 30938 13860 31078
rect 13924 30977 13952 31198
rect 13910 30968 13966 30977
rect 13820 30932 13872 30938
rect 13910 30903 13966 30912
rect 13820 30874 13872 30880
rect 13832 30784 13860 30874
rect 13832 30756 13952 30784
rect 13818 30696 13874 30705
rect 13818 30631 13874 30640
rect 13832 30258 13860 30631
rect 13820 30252 13872 30258
rect 13820 30194 13872 30200
rect 13832 29714 13860 30194
rect 13820 29708 13872 29714
rect 13820 29650 13872 29656
rect 13924 29594 13952 30756
rect 14016 30258 14044 31826
rect 14108 31482 14136 32778
rect 14096 31476 14148 31482
rect 14096 31418 14148 31424
rect 14200 31414 14228 32914
rect 14292 32298 14320 33050
rect 14384 33017 14412 33254
rect 14370 33008 14426 33017
rect 14370 32943 14426 32952
rect 14372 32904 14424 32910
rect 14372 32846 14424 32852
rect 14280 32292 14332 32298
rect 14280 32234 14332 32240
rect 14280 31952 14332 31958
rect 14280 31894 14332 31900
rect 14188 31408 14240 31414
rect 14188 31350 14240 31356
rect 14188 31272 14240 31278
rect 14188 31214 14240 31220
rect 14004 30252 14056 30258
rect 14004 30194 14056 30200
rect 14200 30122 14228 31214
rect 14292 31210 14320 31894
rect 14384 31822 14412 32846
rect 14372 31816 14424 31822
rect 14372 31758 14424 31764
rect 14372 31476 14424 31482
rect 14372 31418 14424 31424
rect 14384 31346 14412 31418
rect 14372 31340 14424 31346
rect 14372 31282 14424 31288
rect 14280 31204 14332 31210
rect 14280 31146 14332 31152
rect 14292 31113 14320 31146
rect 14278 31104 14334 31113
rect 14278 31039 14334 31048
rect 14280 30796 14332 30802
rect 14280 30738 14332 30744
rect 14292 30326 14320 30738
rect 14280 30320 14332 30326
rect 14280 30262 14332 30268
rect 14292 30122 14320 30262
rect 14004 30116 14056 30122
rect 14004 30058 14056 30064
rect 14188 30116 14240 30122
rect 14188 30058 14240 30064
rect 14280 30116 14332 30122
rect 14280 30058 14332 30064
rect 13832 29566 13952 29594
rect 13726 29336 13782 29345
rect 13726 29271 13782 29280
rect 13636 29164 13688 29170
rect 13636 29106 13688 29112
rect 13648 28665 13676 29106
rect 13832 29102 13860 29566
rect 13912 29504 13964 29510
rect 13912 29446 13964 29452
rect 13924 29238 13952 29446
rect 13912 29232 13964 29238
rect 13912 29174 13964 29180
rect 13820 29096 13872 29102
rect 13726 29064 13782 29073
rect 13820 29038 13872 29044
rect 13726 28999 13782 29008
rect 13740 28744 13768 28999
rect 13820 28960 13872 28966
rect 13872 28920 13952 28948
rect 13820 28902 13872 28908
rect 13924 28801 13952 28920
rect 13910 28792 13966 28801
rect 13740 28716 13860 28744
rect 13910 28727 13966 28736
rect 13634 28656 13690 28665
rect 13634 28591 13690 28600
rect 13728 28620 13780 28626
rect 13728 28562 13780 28568
rect 13740 28218 13768 28562
rect 13832 28558 13860 28716
rect 13820 28552 13872 28558
rect 13820 28494 13872 28500
rect 13728 28212 13780 28218
rect 13728 28154 13780 28160
rect 13832 27418 13860 28494
rect 13912 28416 13964 28422
rect 13910 28384 13912 28393
rect 13964 28384 13966 28393
rect 13910 28319 13966 28328
rect 13924 27674 13952 28319
rect 14016 28014 14044 30058
rect 14094 29744 14150 29753
rect 14094 29679 14150 29688
rect 14108 28218 14136 29679
rect 14188 29640 14240 29646
rect 14188 29582 14240 29588
rect 14096 28212 14148 28218
rect 14096 28154 14148 28160
rect 14096 28076 14148 28082
rect 14096 28018 14148 28024
rect 14004 28008 14056 28014
rect 14004 27950 14056 27956
rect 14002 27704 14058 27713
rect 13912 27668 13964 27674
rect 14002 27639 14058 27648
rect 13912 27610 13964 27616
rect 13912 27532 13964 27538
rect 13912 27474 13964 27480
rect 13648 27390 13860 27418
rect 13544 26988 13596 26994
rect 13544 26930 13596 26936
rect 13544 26852 13596 26858
rect 13544 26794 13596 26800
rect 13556 26625 13584 26794
rect 13542 26616 13598 26625
rect 13542 26551 13598 26560
rect 13544 26512 13596 26518
rect 13544 26454 13596 26460
rect 13556 26042 13584 26454
rect 13544 26036 13596 26042
rect 13544 25978 13596 25984
rect 13648 25906 13676 27390
rect 13728 27328 13780 27334
rect 13728 27270 13780 27276
rect 13740 26926 13768 27270
rect 13924 27169 13952 27474
rect 13910 27160 13966 27169
rect 13910 27095 13966 27104
rect 13924 27062 13952 27095
rect 13912 27056 13964 27062
rect 13832 27016 13912 27044
rect 13728 26920 13780 26926
rect 13728 26862 13780 26868
rect 13636 25900 13688 25906
rect 13636 25842 13688 25848
rect 13832 25378 13860 27016
rect 13912 26998 13964 27004
rect 14016 26926 14044 27639
rect 14004 26920 14056 26926
rect 13910 26888 13966 26897
rect 14004 26862 14056 26868
rect 13910 26823 13966 26832
rect 13648 25350 13860 25378
rect 13544 25152 13596 25158
rect 13544 25094 13596 25100
rect 13556 24993 13584 25094
rect 13542 24984 13598 24993
rect 13542 24919 13598 24928
rect 13648 24342 13676 25350
rect 13820 25288 13872 25294
rect 13820 25230 13872 25236
rect 13728 25152 13780 25158
rect 13726 25120 13728 25129
rect 13780 25120 13782 25129
rect 13726 25055 13782 25064
rect 13832 24614 13860 25230
rect 13820 24608 13872 24614
rect 13820 24550 13872 24556
rect 13820 24404 13872 24410
rect 13820 24346 13872 24352
rect 13636 24336 13688 24342
rect 13636 24278 13688 24284
rect 13648 23866 13676 24278
rect 13728 24200 13780 24206
rect 13728 24142 13780 24148
rect 13636 23860 13688 23866
rect 13636 23802 13688 23808
rect 13544 23792 13596 23798
rect 13544 23734 13596 23740
rect 13452 23588 13504 23594
rect 13452 23530 13504 23536
rect 13268 22976 13320 22982
rect 13268 22918 13320 22924
rect 13176 22024 13228 22030
rect 13176 21966 13228 21972
rect 13188 21622 13216 21966
rect 13176 21616 13228 21622
rect 13176 21558 13228 21564
rect 13176 21480 13228 21486
rect 13176 21422 13228 21428
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 12992 21004 13044 21010
rect 12992 20946 13044 20952
rect 13004 20602 13032 20946
rect 12992 20596 13044 20602
rect 12992 20538 13044 20544
rect 13004 20466 13032 20538
rect 13082 20496 13138 20505
rect 12992 20460 13044 20466
rect 13082 20431 13138 20440
rect 12992 20402 13044 20408
rect 13004 19922 13032 20402
rect 12992 19916 13044 19922
rect 12992 19858 13044 19864
rect 12900 19780 12952 19786
rect 12900 19722 12952 19728
rect 12912 19310 12940 19722
rect 13096 19310 13124 20431
rect 13188 19990 13216 21422
rect 13176 19984 13228 19990
rect 13176 19926 13228 19932
rect 13188 19786 13216 19926
rect 13176 19780 13228 19786
rect 13176 19722 13228 19728
rect 12900 19304 12952 19310
rect 12900 19246 12952 19252
rect 13084 19304 13136 19310
rect 13084 19246 13136 19252
rect 12900 19168 12952 19174
rect 12900 19110 12952 19116
rect 12912 15570 12940 19110
rect 13096 18970 13124 19246
rect 13084 18964 13136 18970
rect 13084 18906 13136 18912
rect 12992 17740 13044 17746
rect 12992 17682 13044 17688
rect 13004 17377 13032 17682
rect 12990 17368 13046 17377
rect 12990 17303 12992 17312
rect 13044 17303 13046 17312
rect 12992 17274 13044 17280
rect 13004 17243 13032 17274
rect 13096 16046 13124 18906
rect 13176 18760 13228 18766
rect 13176 18702 13228 18708
rect 13188 18358 13216 18702
rect 13176 18352 13228 18358
rect 13176 18294 13228 18300
rect 13280 17921 13308 22918
rect 13464 22642 13492 23530
rect 13556 23186 13584 23734
rect 13740 23225 13768 24142
rect 13726 23216 13782 23225
rect 13544 23180 13596 23186
rect 13726 23151 13782 23160
rect 13544 23122 13596 23128
rect 13556 22710 13584 23122
rect 13728 23044 13780 23050
rect 13728 22986 13780 22992
rect 13544 22704 13596 22710
rect 13544 22646 13596 22652
rect 13452 22636 13504 22642
rect 13452 22578 13504 22584
rect 13636 22636 13688 22642
rect 13636 22578 13688 22584
rect 13358 22264 13414 22273
rect 13358 22199 13414 22208
rect 13266 17912 13322 17921
rect 13266 17847 13322 17856
rect 13372 17762 13400 22199
rect 13648 22012 13676 22578
rect 13556 21984 13676 22012
rect 13452 21888 13504 21894
rect 13452 21830 13504 21836
rect 13464 21486 13492 21830
rect 13452 21480 13504 21486
rect 13452 21422 13504 21428
rect 13464 21078 13492 21422
rect 13452 21072 13504 21078
rect 13452 21014 13504 21020
rect 13452 20392 13504 20398
rect 13452 20334 13504 20340
rect 13464 19718 13492 20334
rect 13452 19712 13504 19718
rect 13452 19654 13504 19660
rect 13464 19417 13492 19654
rect 13450 19408 13506 19417
rect 13450 19343 13506 19352
rect 13464 18902 13492 19343
rect 13452 18896 13504 18902
rect 13452 18838 13504 18844
rect 13464 18222 13492 18838
rect 13556 18306 13584 21984
rect 13636 20800 13688 20806
rect 13636 20742 13688 20748
rect 13648 20398 13676 20742
rect 13740 20534 13768 22986
rect 13832 22778 13860 24346
rect 13924 23322 13952 26823
rect 14016 26586 14044 26862
rect 14004 26580 14056 26586
rect 14004 26522 14056 26528
rect 14004 25900 14056 25906
rect 14004 25842 14056 25848
rect 14016 25430 14044 25842
rect 14004 25424 14056 25430
rect 14004 25366 14056 25372
rect 14016 24206 14044 25366
rect 14004 24200 14056 24206
rect 14004 24142 14056 24148
rect 14004 23860 14056 23866
rect 14004 23802 14056 23808
rect 13912 23316 13964 23322
rect 13912 23258 13964 23264
rect 14016 22982 14044 23802
rect 14004 22976 14056 22982
rect 14004 22918 14056 22924
rect 13820 22772 13872 22778
rect 13820 22714 13872 22720
rect 14004 22772 14056 22778
rect 14004 22714 14056 22720
rect 13820 21956 13872 21962
rect 13820 21898 13872 21904
rect 13832 21690 13860 21898
rect 13820 21684 13872 21690
rect 13820 21626 13872 21632
rect 14016 21554 14044 22714
rect 13820 21548 13872 21554
rect 13820 21490 13872 21496
rect 14004 21548 14056 21554
rect 14004 21490 14056 21496
rect 13832 21078 13860 21490
rect 13820 21072 13872 21078
rect 13820 21014 13872 21020
rect 13728 20528 13780 20534
rect 13728 20470 13780 20476
rect 13636 20392 13688 20398
rect 13634 20360 13636 20369
rect 13688 20360 13690 20369
rect 13634 20295 13690 20304
rect 14004 19916 14056 19922
rect 14004 19858 14056 19864
rect 14016 19514 14044 19858
rect 14004 19508 14056 19514
rect 14004 19450 14056 19456
rect 13728 18760 13780 18766
rect 13728 18702 13780 18708
rect 13740 18426 13768 18702
rect 13728 18420 13780 18426
rect 13728 18362 13780 18368
rect 13556 18278 13676 18306
rect 13452 18216 13504 18222
rect 13452 18158 13504 18164
rect 13544 18148 13596 18154
rect 13544 18090 13596 18096
rect 13556 17882 13584 18090
rect 13544 17876 13596 17882
rect 13544 17818 13596 17824
rect 13268 17740 13320 17746
rect 13372 17734 13584 17762
rect 13268 17682 13320 17688
rect 13280 16794 13308 17682
rect 13268 16788 13320 16794
rect 13268 16730 13320 16736
rect 13084 16040 13136 16046
rect 13084 15982 13136 15988
rect 12900 15564 12952 15570
rect 12900 15506 12952 15512
rect 12992 15360 13044 15366
rect 12992 15302 13044 15308
rect 13004 13977 13032 15302
rect 13280 15026 13308 16730
rect 13452 16584 13504 16590
rect 13452 16526 13504 16532
rect 13464 15978 13492 16526
rect 13452 15972 13504 15978
rect 13452 15914 13504 15920
rect 13360 15632 13412 15638
rect 13358 15600 13360 15609
rect 13412 15600 13414 15609
rect 13358 15535 13414 15544
rect 13372 15162 13400 15535
rect 13360 15156 13412 15162
rect 13360 15098 13412 15104
rect 13268 15020 13320 15026
rect 13268 14962 13320 14968
rect 13268 14884 13320 14890
rect 13268 14826 13320 14832
rect 13084 14476 13136 14482
rect 13084 14418 13136 14424
rect 13096 14074 13124 14418
rect 13084 14068 13136 14074
rect 13084 14010 13136 14016
rect 12990 13968 13046 13977
rect 12990 13903 13046 13912
rect 12808 13864 12860 13870
rect 12808 13806 12860 13812
rect 12820 13530 12848 13806
rect 12808 13524 12860 13530
rect 12808 13466 12860 13472
rect 13004 12374 13032 13903
rect 12992 12368 13044 12374
rect 12992 12310 13044 12316
rect 13004 11898 13032 12310
rect 13280 12306 13308 14826
rect 13268 12300 13320 12306
rect 13268 12242 13320 12248
rect 12992 11892 13044 11898
rect 12992 11834 13044 11840
rect 13280 11354 13308 12242
rect 13268 11348 13320 11354
rect 13268 11290 13320 11296
rect 13360 11280 13412 11286
rect 12728 11206 12848 11234
rect 13360 11222 13412 11228
rect 12820 11150 12848 11206
rect 12808 11144 12860 11150
rect 12808 11086 12860 11092
rect 12820 10470 12848 11086
rect 13372 10742 13400 11222
rect 13464 10810 13492 15914
rect 13556 13954 13584 17734
rect 13648 15162 13676 18278
rect 13726 18184 13782 18193
rect 13726 18119 13782 18128
rect 13740 17814 13768 18119
rect 13728 17808 13780 17814
rect 13728 17750 13780 17756
rect 13820 17332 13872 17338
rect 13820 17274 13872 17280
rect 13832 16658 13860 17274
rect 14108 16658 14136 28018
rect 14200 23118 14228 29582
rect 14280 29504 14332 29510
rect 14280 29446 14332 29452
rect 14292 29073 14320 29446
rect 14278 29064 14334 29073
rect 14278 28999 14334 29008
rect 14384 28744 14412 31282
rect 14476 30802 14504 36740
rect 14556 36722 14608 36728
rect 14556 36576 14608 36582
rect 14556 36518 14608 36524
rect 14568 36242 14596 36518
rect 14556 36236 14608 36242
rect 14556 36178 14608 36184
rect 14556 35692 14608 35698
rect 14556 35634 14608 35640
rect 14568 35193 14596 35634
rect 14554 35184 14610 35193
rect 14554 35119 14556 35128
rect 14608 35119 14610 35128
rect 14556 35090 14608 35096
rect 14568 34921 14596 35090
rect 14554 34912 14610 34921
rect 14554 34847 14610 34856
rect 14556 34740 14608 34746
rect 14556 34682 14608 34688
rect 14568 34474 14596 34682
rect 14556 34468 14608 34474
rect 14556 34410 14608 34416
rect 14554 33960 14610 33969
rect 14554 33895 14610 33904
rect 14568 33425 14596 33895
rect 14554 33416 14610 33425
rect 14554 33351 14610 33360
rect 14568 33114 14596 33351
rect 14556 33108 14608 33114
rect 14556 33050 14608 33056
rect 14556 32904 14608 32910
rect 14556 32846 14608 32852
rect 14464 30796 14516 30802
rect 14464 30738 14516 30744
rect 14464 30660 14516 30666
rect 14464 30602 14516 30608
rect 14292 28716 14412 28744
rect 14292 26790 14320 28716
rect 14370 28656 14426 28665
rect 14370 28591 14426 28600
rect 14384 28490 14412 28591
rect 14372 28484 14424 28490
rect 14372 28426 14424 28432
rect 14372 28212 14424 28218
rect 14372 28154 14424 28160
rect 14384 28014 14412 28154
rect 14372 28008 14424 28014
rect 14372 27950 14424 27956
rect 14384 27878 14412 27950
rect 14372 27872 14424 27878
rect 14372 27814 14424 27820
rect 14280 26784 14332 26790
rect 14280 26726 14332 26732
rect 14384 24410 14412 27814
rect 14476 27674 14504 30602
rect 14568 28626 14596 32846
rect 14660 31890 14688 37295
rect 14740 37120 14792 37126
rect 14738 37088 14740 37097
rect 14792 37088 14794 37097
rect 14738 37023 14794 37032
rect 14752 36650 14780 37023
rect 15016 36848 15068 36854
rect 15016 36790 15068 36796
rect 14740 36644 14792 36650
rect 14740 36586 14792 36592
rect 14752 36310 14780 36586
rect 15028 36553 15056 36790
rect 15014 36544 15070 36553
rect 15014 36479 15070 36488
rect 15028 36378 15056 36479
rect 15016 36372 15068 36378
rect 15016 36314 15068 36320
rect 14740 36304 14792 36310
rect 14740 36246 14792 36252
rect 15016 36100 15068 36106
rect 15016 36042 15068 36048
rect 14832 36032 14884 36038
rect 14832 35974 14884 35980
rect 14740 35556 14792 35562
rect 14740 35498 14792 35504
rect 14752 35222 14780 35498
rect 14740 35216 14792 35222
rect 14740 35158 14792 35164
rect 14740 34604 14792 34610
rect 14740 34546 14792 34552
rect 14752 34513 14780 34546
rect 14738 34504 14794 34513
rect 14738 34439 14794 34448
rect 14752 34218 14780 34439
rect 14844 34406 14872 35974
rect 14924 35488 14976 35494
rect 14924 35430 14976 35436
rect 14936 35290 14964 35430
rect 14924 35284 14976 35290
rect 14924 35226 14976 35232
rect 14832 34400 14884 34406
rect 14832 34342 14884 34348
rect 14752 34190 14872 34218
rect 14740 34128 14792 34134
rect 14844 34105 14872 34190
rect 14740 34070 14792 34076
rect 14830 34096 14886 34105
rect 14752 33046 14780 34070
rect 14830 34031 14886 34040
rect 14844 33402 14872 34031
rect 14936 33522 14964 35226
rect 15028 34746 15056 36042
rect 15120 35834 15148 38218
rect 15108 35828 15160 35834
rect 15108 35770 15160 35776
rect 15120 35698 15148 35770
rect 15108 35692 15160 35698
rect 15108 35634 15160 35640
rect 15106 35592 15162 35601
rect 15106 35527 15162 35536
rect 15120 35222 15148 35527
rect 15108 35216 15160 35222
rect 15108 35158 15160 35164
rect 15120 34746 15148 35158
rect 15016 34740 15068 34746
rect 15016 34682 15068 34688
rect 15108 34740 15160 34746
rect 15108 34682 15160 34688
rect 15108 34536 15160 34542
rect 15108 34478 15160 34484
rect 15016 34468 15068 34474
rect 15016 34410 15068 34416
rect 15028 34241 15056 34410
rect 15014 34232 15070 34241
rect 15014 34167 15070 34176
rect 15120 34134 15148 34478
rect 15108 34128 15160 34134
rect 15108 34070 15160 34076
rect 15016 33584 15068 33590
rect 15016 33526 15068 33532
rect 15106 33552 15162 33561
rect 14924 33516 14976 33522
rect 14924 33458 14976 33464
rect 14844 33374 14964 33402
rect 14832 33312 14884 33318
rect 14832 33254 14884 33260
rect 14844 33114 14872 33254
rect 14832 33108 14884 33114
rect 14832 33050 14884 33056
rect 14740 33040 14792 33046
rect 14936 32994 14964 33374
rect 14740 32982 14792 32988
rect 14844 32966 14964 32994
rect 14844 32910 14872 32966
rect 14832 32904 14884 32910
rect 14738 32872 14794 32881
rect 14832 32846 14884 32852
rect 14924 32904 14976 32910
rect 14924 32846 14976 32852
rect 14738 32807 14794 32816
rect 14752 32756 14780 32807
rect 14752 32728 14872 32756
rect 14740 32292 14792 32298
rect 14740 32234 14792 32240
rect 14752 32201 14780 32234
rect 14738 32192 14794 32201
rect 14738 32127 14794 32136
rect 14648 31884 14700 31890
rect 14648 31826 14700 31832
rect 14844 31770 14872 32728
rect 14660 31742 14872 31770
rect 14936 31754 14964 32846
rect 15028 32026 15056 33526
rect 15106 33487 15162 33496
rect 15120 33454 15148 33487
rect 15108 33448 15160 33454
rect 15108 33390 15160 33396
rect 15120 33114 15148 33390
rect 15108 33108 15160 33114
rect 15108 33050 15160 33056
rect 15108 32224 15160 32230
rect 15108 32166 15160 32172
rect 15016 32020 15068 32026
rect 15016 31962 15068 31968
rect 15120 31906 15148 32166
rect 15028 31878 15148 31906
rect 14924 31748 14976 31754
rect 14660 29782 14688 31742
rect 14924 31690 14976 31696
rect 14832 31340 14884 31346
rect 14832 31282 14884 31288
rect 14740 30592 14792 30598
rect 14740 30534 14792 30540
rect 14752 30190 14780 30534
rect 14740 30184 14792 30190
rect 14740 30126 14792 30132
rect 14648 29776 14700 29782
rect 14648 29718 14700 29724
rect 14648 29096 14700 29102
rect 14648 29038 14700 29044
rect 14556 28620 14608 28626
rect 14556 28562 14608 28568
rect 14464 27668 14516 27674
rect 14464 27610 14516 27616
rect 14556 27600 14608 27606
rect 14556 27542 14608 27548
rect 14464 27532 14516 27538
rect 14464 27474 14516 27480
rect 14476 26194 14504 27474
rect 14568 27418 14596 27542
rect 14660 27538 14688 29038
rect 14752 28937 14780 30126
rect 14844 29288 14872 31282
rect 15028 30870 15056 31878
rect 15108 31204 15160 31210
rect 15108 31146 15160 31152
rect 15120 30977 15148 31146
rect 15106 30968 15162 30977
rect 15106 30903 15162 30912
rect 15016 30864 15068 30870
rect 15016 30806 15068 30812
rect 14924 30728 14976 30734
rect 14924 30670 14976 30676
rect 14936 30297 14964 30670
rect 15028 30569 15056 30806
rect 15014 30560 15070 30569
rect 15014 30495 15070 30504
rect 14922 30288 14978 30297
rect 14978 30246 15056 30274
rect 14922 30223 14978 30232
rect 14924 30184 14976 30190
rect 14924 30126 14976 30132
rect 14936 29646 14964 30126
rect 15028 30054 15056 30246
rect 15108 30184 15160 30190
rect 15108 30126 15160 30132
rect 15016 30048 15068 30054
rect 15016 29990 15068 29996
rect 15016 29844 15068 29850
rect 15016 29786 15068 29792
rect 14924 29640 14976 29646
rect 14924 29582 14976 29588
rect 14844 29260 14964 29288
rect 14832 29164 14884 29170
rect 14832 29106 14884 29112
rect 14738 28928 14794 28937
rect 14738 28863 14794 28872
rect 14738 28792 14794 28801
rect 14738 28727 14794 28736
rect 14648 27532 14700 27538
rect 14648 27474 14700 27480
rect 14568 27390 14688 27418
rect 14476 26166 14596 26194
rect 14464 26036 14516 26042
rect 14464 25978 14516 25984
rect 14476 24954 14504 25978
rect 14568 25770 14596 26166
rect 14556 25764 14608 25770
rect 14556 25706 14608 25712
rect 14464 24948 14516 24954
rect 14464 24890 14516 24896
rect 14464 24744 14516 24750
rect 14464 24686 14516 24692
rect 14372 24404 14424 24410
rect 14372 24346 14424 24352
rect 14280 24132 14332 24138
rect 14280 24074 14332 24080
rect 14292 23662 14320 24074
rect 14372 24064 14424 24070
rect 14372 24006 14424 24012
rect 14384 23662 14412 24006
rect 14280 23656 14332 23662
rect 14280 23598 14332 23604
rect 14372 23656 14424 23662
rect 14372 23598 14424 23604
rect 14372 23316 14424 23322
rect 14372 23258 14424 23264
rect 14188 23112 14240 23118
rect 14188 23054 14240 23060
rect 14200 21978 14228 23054
rect 14280 22976 14332 22982
rect 14280 22918 14332 22924
rect 14292 22574 14320 22918
rect 14280 22568 14332 22574
rect 14280 22510 14332 22516
rect 14292 22234 14320 22510
rect 14280 22228 14332 22234
rect 14280 22170 14332 22176
rect 14200 21950 14320 21978
rect 14188 21888 14240 21894
rect 14188 21830 14240 21836
rect 14200 21026 14228 21830
rect 14292 21418 14320 21950
rect 14280 21412 14332 21418
rect 14280 21354 14332 21360
rect 14292 21146 14320 21354
rect 14280 21140 14332 21146
rect 14280 21082 14332 21088
rect 14200 21010 14320 21026
rect 14188 21004 14320 21010
rect 14240 20998 14320 21004
rect 14188 20946 14240 20952
rect 14186 20904 14242 20913
rect 14186 20839 14242 20848
rect 14200 20398 14228 20839
rect 14188 20392 14240 20398
rect 14188 20334 14240 20340
rect 14292 20058 14320 20998
rect 14280 20052 14332 20058
rect 14280 19994 14332 20000
rect 14384 19718 14412 23258
rect 14372 19712 14424 19718
rect 14372 19654 14424 19660
rect 14372 19304 14424 19310
rect 14372 19246 14424 19252
rect 14188 18964 14240 18970
rect 14188 18906 14240 18912
rect 14200 17202 14228 18906
rect 14384 18426 14412 19246
rect 14372 18420 14424 18426
rect 14372 18362 14424 18368
rect 14476 17338 14504 24686
rect 14568 24342 14596 25706
rect 14556 24336 14608 24342
rect 14556 24278 14608 24284
rect 14660 23526 14688 27390
rect 14752 25974 14780 28727
rect 14844 26586 14872 29106
rect 14936 29102 14964 29260
rect 14924 29096 14976 29102
rect 14924 29038 14976 29044
rect 14924 28960 14976 28966
rect 14924 28902 14976 28908
rect 14936 28626 14964 28902
rect 14924 28620 14976 28626
rect 14924 28562 14976 28568
rect 14924 28484 14976 28490
rect 14924 28426 14976 28432
rect 14936 28150 14964 28426
rect 14924 28144 14976 28150
rect 14924 28086 14976 28092
rect 14936 28014 14964 28086
rect 14924 28008 14976 28014
rect 14924 27950 14976 27956
rect 14936 27334 14964 27950
rect 14924 27328 14976 27334
rect 14924 27270 14976 27276
rect 15028 27112 15056 29786
rect 15120 29782 15148 30126
rect 15108 29776 15160 29782
rect 15106 29744 15108 29753
rect 15160 29744 15162 29753
rect 15106 29679 15162 29688
rect 15108 29300 15160 29306
rect 15108 29242 15160 29248
rect 15120 29170 15148 29242
rect 15108 29164 15160 29170
rect 15108 29106 15160 29112
rect 15120 28121 15148 29106
rect 15106 28112 15162 28121
rect 15106 28047 15162 28056
rect 15108 28008 15160 28014
rect 15108 27950 15160 27956
rect 15120 27674 15148 27950
rect 15108 27668 15160 27674
rect 15108 27610 15160 27616
rect 15108 27328 15160 27334
rect 15108 27270 15160 27276
rect 14936 27084 15056 27112
rect 14832 26580 14884 26586
rect 14832 26522 14884 26528
rect 14740 25968 14792 25974
rect 14792 25928 14872 25956
rect 14740 25910 14792 25916
rect 14738 25800 14794 25809
rect 14738 25735 14740 25744
rect 14792 25735 14794 25744
rect 14740 25706 14792 25712
rect 14752 24886 14780 25706
rect 14844 25702 14872 25928
rect 14832 25696 14884 25702
rect 14832 25638 14884 25644
rect 14740 24880 14792 24886
rect 14740 24822 14792 24828
rect 14844 23746 14872 25638
rect 14936 25498 14964 27084
rect 15120 27062 15148 27270
rect 15108 27056 15160 27062
rect 15108 26998 15160 27004
rect 15016 26920 15068 26926
rect 15016 26862 15068 26868
rect 15028 26246 15056 26862
rect 15108 26852 15160 26858
rect 15108 26794 15160 26800
rect 15016 26240 15068 26246
rect 15016 26182 15068 26188
rect 14924 25492 14976 25498
rect 14924 25434 14976 25440
rect 14922 24984 14978 24993
rect 14922 24919 14978 24928
rect 14936 24410 14964 24919
rect 14924 24404 14976 24410
rect 14924 24346 14976 24352
rect 14924 24064 14976 24070
rect 14924 24006 14976 24012
rect 14752 23718 14872 23746
rect 14648 23520 14700 23526
rect 14648 23462 14700 23468
rect 14556 23248 14608 23254
rect 14556 23190 14608 23196
rect 14568 19553 14596 23190
rect 14648 23044 14700 23050
rect 14648 22986 14700 22992
rect 14660 22574 14688 22986
rect 14648 22568 14700 22574
rect 14648 22510 14700 22516
rect 14752 22250 14780 23718
rect 14936 23662 14964 24006
rect 14832 23656 14884 23662
rect 14832 23598 14884 23604
rect 14924 23656 14976 23662
rect 14924 23598 14976 23604
rect 14844 23322 14872 23598
rect 14832 23316 14884 23322
rect 14832 23258 14884 23264
rect 14936 23202 14964 23598
rect 14844 23174 14964 23202
rect 14844 22642 14872 23174
rect 14922 22808 14978 22817
rect 14922 22743 14978 22752
rect 14832 22636 14884 22642
rect 14832 22578 14884 22584
rect 14936 22506 14964 22743
rect 14924 22500 14976 22506
rect 14924 22442 14976 22448
rect 14752 22222 14872 22250
rect 14936 22234 14964 22442
rect 14740 22160 14792 22166
rect 14740 22102 14792 22108
rect 14646 21312 14702 21321
rect 14646 21247 14702 21256
rect 14660 21078 14688 21247
rect 14752 21146 14780 22102
rect 14740 21140 14792 21146
rect 14740 21082 14792 21088
rect 14648 21072 14700 21078
rect 14648 21014 14700 21020
rect 14844 20448 14872 22222
rect 14924 22228 14976 22234
rect 14924 22170 14976 22176
rect 15028 22114 15056 26182
rect 15120 25906 15148 26794
rect 15108 25900 15160 25906
rect 15108 25842 15160 25848
rect 15108 24336 15160 24342
rect 15108 24278 15160 24284
rect 15120 23322 15148 24278
rect 15108 23316 15160 23322
rect 15108 23258 15160 23264
rect 15120 22778 15148 23258
rect 15108 22772 15160 22778
rect 15108 22714 15160 22720
rect 15106 22264 15162 22273
rect 15106 22199 15162 22208
rect 14752 20420 14872 20448
rect 14936 22086 15056 22114
rect 14648 20256 14700 20262
rect 14648 20198 14700 20204
rect 14554 19544 14610 19553
rect 14554 19479 14610 19488
rect 14660 19174 14688 20198
rect 14752 20058 14780 20420
rect 14832 20324 14884 20330
rect 14832 20266 14884 20272
rect 14740 20052 14792 20058
rect 14740 19994 14792 20000
rect 14740 19712 14792 19718
rect 14740 19654 14792 19660
rect 14648 19168 14700 19174
rect 14648 19110 14700 19116
rect 14648 18216 14700 18222
rect 14648 18158 14700 18164
rect 14660 17882 14688 18158
rect 14752 18086 14780 19654
rect 14740 18080 14792 18086
rect 14740 18022 14792 18028
rect 14648 17876 14700 17882
rect 14648 17818 14700 17824
rect 14464 17332 14516 17338
rect 14464 17274 14516 17280
rect 14188 17196 14240 17202
rect 14188 17138 14240 17144
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 14096 16652 14148 16658
rect 14096 16594 14148 16600
rect 13832 16250 13860 16594
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 13820 15972 13872 15978
rect 13820 15914 13872 15920
rect 13832 15858 13860 15914
rect 13740 15830 13860 15858
rect 13636 15156 13688 15162
rect 13636 15098 13688 15104
rect 13648 14346 13676 15098
rect 13740 14550 13768 15830
rect 13820 15564 13872 15570
rect 13820 15506 13872 15512
rect 13832 14550 13860 15506
rect 14200 15337 14228 17138
rect 14476 17134 14504 17274
rect 14280 17128 14332 17134
rect 14280 17070 14332 17076
rect 14464 17128 14516 17134
rect 14464 17070 14516 17076
rect 14292 16998 14320 17070
rect 14280 16992 14332 16998
rect 14280 16934 14332 16940
rect 14186 15328 14242 15337
rect 14186 15263 14242 15272
rect 13728 14544 13780 14550
rect 13728 14486 13780 14492
rect 13820 14544 13872 14550
rect 13820 14486 13872 14492
rect 13636 14340 13688 14346
rect 13636 14282 13688 14288
rect 13648 14074 13676 14282
rect 14292 14074 14320 16934
rect 14648 16584 14700 16590
rect 14648 16526 14700 16532
rect 14660 15994 14688 16526
rect 14740 16040 14792 16046
rect 14660 15988 14740 15994
rect 14660 15982 14792 15988
rect 14660 15966 14780 15982
rect 14660 15638 14688 15966
rect 14648 15632 14700 15638
rect 14648 15574 14700 15580
rect 14464 14952 14516 14958
rect 14464 14894 14516 14900
rect 14476 14618 14504 14894
rect 14646 14648 14702 14657
rect 14464 14612 14516 14618
rect 14646 14583 14702 14592
rect 14464 14554 14516 14560
rect 14660 14482 14688 14583
rect 14648 14476 14700 14482
rect 14648 14418 14700 14424
rect 13636 14068 13688 14074
rect 13636 14010 13688 14016
rect 14280 14068 14332 14074
rect 14280 14010 14332 14016
rect 13556 13926 13676 13954
rect 13542 13560 13598 13569
rect 13542 13495 13598 13504
rect 13556 13394 13584 13495
rect 13544 13388 13596 13394
rect 13544 13330 13596 13336
rect 13556 12918 13584 13330
rect 13544 12912 13596 12918
rect 13544 12854 13596 12860
rect 13648 12356 13676 13926
rect 14660 13870 14688 14418
rect 14844 14226 14872 20266
rect 14936 15094 14964 22086
rect 15120 22030 15148 22199
rect 15016 22024 15068 22030
rect 15016 21966 15068 21972
rect 15108 22024 15160 22030
rect 15108 21966 15160 21972
rect 15028 21350 15056 21966
rect 15016 21344 15068 21350
rect 15016 21286 15068 21292
rect 15016 20800 15068 20806
rect 15014 20768 15016 20777
rect 15068 20768 15070 20777
rect 15014 20703 15070 20712
rect 15014 20224 15070 20233
rect 15014 20159 15070 20168
rect 15028 18970 15056 20159
rect 15108 19304 15160 19310
rect 15108 19246 15160 19252
rect 15016 18964 15068 18970
rect 15016 18906 15068 18912
rect 15120 18698 15148 19246
rect 15108 18692 15160 18698
rect 15108 18634 15160 18640
rect 15106 18320 15162 18329
rect 15016 18284 15068 18290
rect 15106 18255 15162 18264
rect 15016 18226 15068 18232
rect 15028 17762 15056 18226
rect 15120 18222 15148 18255
rect 15108 18216 15160 18222
rect 15108 18158 15160 18164
rect 15028 17734 15148 17762
rect 15016 17672 15068 17678
rect 15016 17614 15068 17620
rect 15028 17134 15056 17614
rect 15016 17128 15068 17134
rect 15016 17070 15068 17076
rect 15028 16726 15056 17070
rect 15120 16726 15148 17734
rect 15016 16720 15068 16726
rect 15016 16662 15068 16668
rect 15108 16720 15160 16726
rect 15108 16662 15160 16668
rect 15014 15736 15070 15745
rect 15014 15671 15070 15680
rect 14924 15088 14976 15094
rect 14924 15030 14976 15036
rect 15028 14958 15056 15671
rect 15016 14952 15068 14958
rect 15016 14894 15068 14900
rect 14924 14884 14976 14890
rect 14924 14826 14976 14832
rect 14936 14414 14964 14826
rect 15028 14550 15056 14894
rect 15016 14544 15068 14550
rect 15016 14486 15068 14492
rect 14924 14408 14976 14414
rect 14922 14376 14924 14385
rect 14976 14376 14978 14385
rect 14922 14311 14978 14320
rect 14844 14198 15148 14226
rect 14648 13864 14700 13870
rect 14648 13806 14700 13812
rect 15014 13696 15070 13705
rect 15014 13631 15070 13640
rect 13912 13320 13964 13326
rect 13912 13262 13964 13268
rect 13924 12986 13952 13262
rect 13912 12980 13964 12986
rect 13912 12922 13964 12928
rect 13556 12328 13676 12356
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 13360 10736 13412 10742
rect 13360 10678 13412 10684
rect 12808 10464 12860 10470
rect 12808 10406 12860 10412
rect 12624 9716 12676 9722
rect 12624 9658 12676 9664
rect 12440 9512 12492 9518
rect 12440 9454 12492 9460
rect 12164 8968 12216 8974
rect 12164 8910 12216 8916
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 12176 3505 12204 8910
rect 12452 8090 12480 9454
rect 12636 9042 12664 9658
rect 12624 9036 12676 9042
rect 12624 8978 12676 8984
rect 12636 8634 12664 8978
rect 12624 8628 12676 8634
rect 12624 8570 12676 8576
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12162 3496 12218 3505
rect 12162 3431 12218 3440
rect 12820 2689 12848 10406
rect 13268 9376 13320 9382
rect 13268 9318 13320 9324
rect 12990 9072 13046 9081
rect 12990 9007 12992 9016
rect 13044 9007 13046 9016
rect 12992 8978 13044 8984
rect 13004 8566 13032 8978
rect 13280 8566 13308 9318
rect 12992 8560 13044 8566
rect 12992 8502 13044 8508
rect 13268 8560 13320 8566
rect 13268 8502 13320 8508
rect 13280 8430 13308 8502
rect 13268 8424 13320 8430
rect 13268 8366 13320 8372
rect 13452 8016 13504 8022
rect 13450 7984 13452 7993
rect 13504 7984 13506 7993
rect 13450 7919 13506 7928
rect 13084 7336 13136 7342
rect 13084 7278 13136 7284
rect 13096 6662 13124 7278
rect 13084 6656 13136 6662
rect 13084 6598 13136 6604
rect 13096 5574 13124 6598
rect 13360 5840 13412 5846
rect 13360 5782 13412 5788
rect 13084 5568 13136 5574
rect 13084 5510 13136 5516
rect 13096 5166 13124 5510
rect 13372 5370 13400 5782
rect 13452 5568 13504 5574
rect 13452 5510 13504 5516
rect 13360 5364 13412 5370
rect 13360 5306 13412 5312
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 12898 3496 12954 3505
rect 12898 3431 12954 3440
rect 12806 2680 12862 2689
rect 12806 2615 12862 2624
rect 12440 2508 12492 2514
rect 12440 2450 12492 2456
rect 12452 2310 12480 2450
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 12452 800 12480 2246
rect 12912 800 12940 3431
rect 13096 2446 13124 5102
rect 13464 4049 13492 5510
rect 13556 4758 13584 12328
rect 14188 12096 14240 12102
rect 14188 12038 14240 12044
rect 14922 12064 14978 12073
rect 13728 11620 13780 11626
rect 13728 11562 13780 11568
rect 13636 11212 13688 11218
rect 13636 11154 13688 11160
rect 13648 10810 13676 11154
rect 13636 10804 13688 10810
rect 13636 10746 13688 10752
rect 13740 8616 13768 11562
rect 14002 11384 14058 11393
rect 14002 11319 14058 11328
rect 14016 10169 14044 11319
rect 14002 10160 14058 10169
rect 14002 10095 14058 10104
rect 14096 8832 14148 8838
rect 14096 8774 14148 8780
rect 14004 8628 14056 8634
rect 13740 8588 13860 8616
rect 13728 8492 13780 8498
rect 13728 8434 13780 8440
rect 13740 7449 13768 8434
rect 13832 8362 13860 8588
rect 14004 8570 14056 8576
rect 14016 8498 14044 8570
rect 14004 8492 14056 8498
rect 14004 8434 14056 8440
rect 13820 8356 13872 8362
rect 13820 8298 13872 8304
rect 13832 8090 13860 8298
rect 13820 8084 13872 8090
rect 13820 8026 13872 8032
rect 13726 7440 13782 7449
rect 13832 7410 13860 8026
rect 14016 8022 14044 8434
rect 14108 8430 14136 8774
rect 14096 8424 14148 8430
rect 14096 8366 14148 8372
rect 14004 8016 14056 8022
rect 14004 7958 14056 7964
rect 13726 7375 13782 7384
rect 13820 7404 13872 7410
rect 13820 7346 13872 7352
rect 13820 5772 13872 5778
rect 13820 5714 13872 5720
rect 13728 5704 13780 5710
rect 13728 5646 13780 5652
rect 13636 5024 13688 5030
rect 13636 4966 13688 4972
rect 13648 4826 13676 4966
rect 13636 4820 13688 4826
rect 13636 4762 13688 4768
rect 13544 4752 13596 4758
rect 13544 4694 13596 4700
rect 13740 4690 13768 5646
rect 13832 5030 13860 5714
rect 14016 5710 14044 7958
rect 14108 7546 14136 8366
rect 14096 7540 14148 7546
rect 14096 7482 14148 7488
rect 14200 6458 14228 12038
rect 14922 11999 14978 12008
rect 14936 11898 14964 11999
rect 14924 11892 14976 11898
rect 14924 11834 14976 11840
rect 14922 9616 14978 9625
rect 14922 9551 14924 9560
rect 14976 9551 14978 9560
rect 14924 9522 14976 9528
rect 14464 9512 14516 9518
rect 14462 9480 14464 9489
rect 14516 9480 14518 9489
rect 14462 9415 14518 9424
rect 14554 8120 14610 8129
rect 14554 8055 14610 8064
rect 14568 6662 14596 8055
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 14568 6254 14596 6598
rect 14556 6248 14608 6254
rect 14556 6190 14608 6196
rect 14188 5772 14240 5778
rect 14188 5714 14240 5720
rect 14004 5704 14056 5710
rect 14004 5646 14056 5652
rect 14200 5166 14228 5714
rect 14188 5160 14240 5166
rect 14188 5102 14240 5108
rect 13820 5024 13872 5030
rect 13820 4966 13872 4972
rect 14200 4826 14228 5102
rect 14188 4820 14240 4826
rect 14188 4762 14240 4768
rect 13728 4684 13780 4690
rect 13728 4626 13780 4632
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 13450 4040 13506 4049
rect 13450 3975 13506 3984
rect 13084 2440 13136 2446
rect 13084 2382 13136 2388
rect 13832 800 13860 4082
rect 14002 2680 14058 2689
rect 14002 2615 14004 2624
rect 14056 2615 14058 2624
rect 14004 2586 14056 2592
rect 15028 1034 15056 13631
rect 15120 4146 15148 14198
rect 15212 8265 15240 42248
rect 15488 41290 15516 44152
rect 15752 43716 15804 43722
rect 15752 43658 15804 43664
rect 15764 43450 15792 43658
rect 15752 43444 15804 43450
rect 15752 43386 15804 43392
rect 15660 41472 15712 41478
rect 15660 41414 15712 41420
rect 15488 41262 15608 41290
rect 15292 39500 15344 39506
rect 15292 39442 15344 39448
rect 15304 38962 15332 39442
rect 15292 38956 15344 38962
rect 15292 38898 15344 38904
rect 15292 38820 15344 38826
rect 15292 38762 15344 38768
rect 15304 37806 15332 38762
rect 15476 38752 15528 38758
rect 15476 38694 15528 38700
rect 15384 38208 15436 38214
rect 15384 38150 15436 38156
rect 15396 37874 15424 38150
rect 15488 37913 15516 38694
rect 15474 37904 15530 37913
rect 15384 37868 15436 37874
rect 15474 37839 15530 37848
rect 15384 37810 15436 37816
rect 15292 37800 15344 37806
rect 15292 37742 15344 37748
rect 15292 37664 15344 37670
rect 15292 37606 15344 37612
rect 15304 36854 15332 37606
rect 15384 37460 15436 37466
rect 15384 37402 15436 37408
rect 15292 36848 15344 36854
rect 15292 36790 15344 36796
rect 15292 36576 15344 36582
rect 15292 36518 15344 36524
rect 15304 34950 15332 36518
rect 15292 34944 15344 34950
rect 15292 34886 15344 34892
rect 15292 34060 15344 34066
rect 15292 34002 15344 34008
rect 15304 33289 15332 34002
rect 15396 33590 15424 37402
rect 15488 35601 15516 37839
rect 15580 36530 15608 41262
rect 15672 41138 15700 41414
rect 15750 41304 15806 41313
rect 15750 41239 15806 41248
rect 15660 41132 15712 41138
rect 15660 41074 15712 41080
rect 15672 40390 15700 41074
rect 15764 41002 15792 41239
rect 15752 40996 15804 41002
rect 15752 40938 15804 40944
rect 15660 40384 15712 40390
rect 15660 40326 15712 40332
rect 15672 40089 15700 40326
rect 15658 40080 15714 40089
rect 15658 40015 15714 40024
rect 15752 39296 15804 39302
rect 15752 39238 15804 39244
rect 15660 38956 15712 38962
rect 15660 38898 15712 38904
rect 15672 38758 15700 38898
rect 15660 38752 15712 38758
rect 15660 38694 15712 38700
rect 15672 37942 15700 38694
rect 15764 38282 15792 39238
rect 15752 38276 15804 38282
rect 15752 38218 15804 38224
rect 15752 38004 15804 38010
rect 15752 37946 15804 37952
rect 15660 37936 15712 37942
rect 15660 37878 15712 37884
rect 15660 37800 15712 37806
rect 15660 37742 15712 37748
rect 15672 37398 15700 37742
rect 15764 37738 15792 37946
rect 15752 37732 15804 37738
rect 15752 37674 15804 37680
rect 15660 37392 15712 37398
rect 15764 37369 15792 37674
rect 15660 37334 15712 37340
rect 15750 37360 15806 37369
rect 15672 37262 15700 37334
rect 15750 37295 15806 37304
rect 15660 37256 15712 37262
rect 15660 37198 15712 37204
rect 15660 37120 15712 37126
rect 15752 37120 15804 37126
rect 15660 37062 15712 37068
rect 15750 37088 15752 37097
rect 15804 37088 15806 37097
rect 15672 36922 15700 37062
rect 15750 37023 15806 37032
rect 15660 36916 15712 36922
rect 15660 36858 15712 36864
rect 15580 36502 15792 36530
rect 15658 36408 15714 36417
rect 15658 36343 15714 36352
rect 15566 36136 15622 36145
rect 15566 36071 15622 36080
rect 15474 35592 15530 35601
rect 15474 35527 15530 35536
rect 15476 35488 15528 35494
rect 15476 35430 15528 35436
rect 15384 33584 15436 33590
rect 15384 33526 15436 33532
rect 15384 33448 15436 33454
rect 15488 33425 15516 35430
rect 15580 34474 15608 36071
rect 15672 35086 15700 36343
rect 15660 35080 15712 35086
rect 15660 35022 15712 35028
rect 15568 34468 15620 34474
rect 15568 34410 15620 34416
rect 15568 33856 15620 33862
rect 15568 33798 15620 33804
rect 15660 33856 15712 33862
rect 15660 33798 15712 33804
rect 15580 33658 15608 33798
rect 15568 33652 15620 33658
rect 15568 33594 15620 33600
rect 15384 33390 15436 33396
rect 15474 33416 15530 33425
rect 15290 33280 15346 33289
rect 15290 33215 15346 33224
rect 15396 33130 15424 33390
rect 15474 33351 15530 33360
rect 15304 33102 15424 33130
rect 15476 33108 15528 33114
rect 15304 31890 15332 33102
rect 15476 33050 15528 33056
rect 15384 33040 15436 33046
rect 15384 32982 15436 32988
rect 15292 31884 15344 31890
rect 15292 31826 15344 31832
rect 15304 31482 15332 31826
rect 15396 31793 15424 32982
rect 15488 31822 15516 33050
rect 15566 33008 15622 33017
rect 15566 32943 15568 32952
rect 15620 32943 15622 32952
rect 15568 32914 15620 32920
rect 15580 32570 15608 32914
rect 15568 32564 15620 32570
rect 15568 32506 15620 32512
rect 15566 32464 15622 32473
rect 15566 32399 15568 32408
rect 15620 32399 15622 32408
rect 15568 32370 15620 32376
rect 15568 32224 15620 32230
rect 15568 32166 15620 32172
rect 15580 31929 15608 32166
rect 15566 31920 15622 31929
rect 15566 31855 15622 31864
rect 15476 31816 15528 31822
rect 15382 31784 15438 31793
rect 15476 31758 15528 31764
rect 15382 31719 15438 31728
rect 15568 31680 15620 31686
rect 15568 31622 15620 31628
rect 15474 31512 15530 31521
rect 15292 31476 15344 31482
rect 15474 31447 15530 31456
rect 15292 31418 15344 31424
rect 15304 31113 15332 31418
rect 15290 31104 15346 31113
rect 15290 31039 15346 31048
rect 15292 30796 15344 30802
rect 15292 30738 15344 30744
rect 15384 30796 15436 30802
rect 15384 30738 15436 30744
rect 15304 30326 15332 30738
rect 15396 30394 15424 30738
rect 15384 30388 15436 30394
rect 15384 30330 15436 30336
rect 15292 30320 15344 30326
rect 15292 30262 15344 30268
rect 15304 29306 15332 30262
rect 15384 30048 15436 30054
rect 15384 29990 15436 29996
rect 15396 29782 15424 29990
rect 15384 29776 15436 29782
rect 15384 29718 15436 29724
rect 15384 29504 15436 29510
rect 15384 29446 15436 29452
rect 15292 29300 15344 29306
rect 15292 29242 15344 29248
rect 15396 28762 15424 29446
rect 15384 28756 15436 28762
rect 15384 28698 15436 28704
rect 15292 28688 15344 28694
rect 15292 28630 15344 28636
rect 15304 27674 15332 28630
rect 15384 28552 15436 28558
rect 15384 28494 15436 28500
rect 15396 27878 15424 28494
rect 15384 27872 15436 27878
rect 15384 27814 15436 27820
rect 15488 27690 15516 31447
rect 15580 31142 15608 31622
rect 15672 31464 15700 33798
rect 15764 31657 15792 36502
rect 15856 32434 15884 51224
rect 15956 51164 16252 51184
rect 16012 51162 16036 51164
rect 16092 51162 16116 51164
rect 16172 51162 16196 51164
rect 16034 51110 16036 51162
rect 16098 51110 16110 51162
rect 16172 51110 16174 51162
rect 16012 51108 16036 51110
rect 16092 51108 16116 51110
rect 16172 51108 16196 51110
rect 15956 51088 16252 51108
rect 16316 50998 16344 51342
rect 16304 50992 16356 50998
rect 16304 50934 16356 50940
rect 16316 50522 16344 50934
rect 16304 50516 16356 50522
rect 16304 50458 16356 50464
rect 15956 50076 16252 50096
rect 16012 50074 16036 50076
rect 16092 50074 16116 50076
rect 16172 50074 16196 50076
rect 16034 50022 16036 50074
rect 16098 50022 16110 50074
rect 16172 50022 16174 50074
rect 16012 50020 16036 50022
rect 16092 50020 16116 50022
rect 16172 50020 16196 50022
rect 15956 50000 16252 50020
rect 16028 49768 16080 49774
rect 16028 49710 16080 49716
rect 16040 49609 16068 49710
rect 16026 49600 16082 49609
rect 16026 49535 16082 49544
rect 16304 49360 16356 49366
rect 16304 49302 16356 49308
rect 15956 48988 16252 49008
rect 16012 48986 16036 48988
rect 16092 48986 16116 48988
rect 16172 48986 16196 48988
rect 16034 48934 16036 48986
rect 16098 48934 16110 48986
rect 16172 48934 16174 48986
rect 16012 48932 16036 48934
rect 16092 48932 16116 48934
rect 16172 48932 16196 48934
rect 15956 48912 16252 48932
rect 16316 48754 16344 49302
rect 16304 48748 16356 48754
rect 16304 48690 16356 48696
rect 15956 47900 16252 47920
rect 16012 47898 16036 47900
rect 16092 47898 16116 47900
rect 16172 47898 16196 47900
rect 16034 47846 16036 47898
rect 16098 47846 16110 47898
rect 16172 47846 16174 47898
rect 16012 47844 16036 47846
rect 16092 47844 16116 47846
rect 16172 47844 16196 47846
rect 15956 47824 16252 47844
rect 16302 47696 16358 47705
rect 16302 47631 16358 47640
rect 16316 47598 16344 47631
rect 16304 47592 16356 47598
rect 16304 47534 16356 47540
rect 16212 47524 16264 47530
rect 16212 47466 16264 47472
rect 16118 47016 16174 47025
rect 16224 47002 16252 47466
rect 16316 47122 16344 47534
rect 16304 47116 16356 47122
rect 16304 47058 16356 47064
rect 16224 46974 16344 47002
rect 16118 46951 16120 46960
rect 16172 46951 16174 46960
rect 16120 46922 16172 46928
rect 15956 46812 16252 46832
rect 16012 46810 16036 46812
rect 16092 46810 16116 46812
rect 16172 46810 16196 46812
rect 16034 46758 16036 46810
rect 16098 46758 16110 46810
rect 16172 46758 16174 46810
rect 16012 46756 16036 46758
rect 16092 46756 16116 46758
rect 16172 46756 16196 46758
rect 15956 46736 16252 46756
rect 16120 46572 16172 46578
rect 16120 46514 16172 46520
rect 16132 46170 16160 46514
rect 16212 46504 16264 46510
rect 16316 46492 16344 46974
rect 16264 46464 16344 46492
rect 16212 46446 16264 46452
rect 16224 46170 16252 46446
rect 16120 46164 16172 46170
rect 16120 46106 16172 46112
rect 16212 46164 16264 46170
rect 16212 46106 16264 46112
rect 16118 45928 16174 45937
rect 16118 45863 16120 45872
rect 16172 45863 16174 45872
rect 16120 45834 16172 45840
rect 15956 45724 16252 45744
rect 16012 45722 16036 45724
rect 16092 45722 16116 45724
rect 16172 45722 16196 45724
rect 16034 45670 16036 45722
rect 16098 45670 16110 45722
rect 16172 45670 16174 45722
rect 16012 45668 16036 45670
rect 16092 45668 16116 45670
rect 16172 45668 16196 45670
rect 15956 45648 16252 45668
rect 15956 44636 16252 44656
rect 16012 44634 16036 44636
rect 16092 44634 16116 44636
rect 16172 44634 16196 44636
rect 16034 44582 16036 44634
rect 16098 44582 16110 44634
rect 16172 44582 16174 44634
rect 16012 44580 16036 44582
rect 16092 44580 16116 44582
rect 16172 44580 16196 44582
rect 15956 44560 16252 44580
rect 16118 44296 16174 44305
rect 16118 44231 16174 44240
rect 16132 44198 16160 44231
rect 16120 44192 16172 44198
rect 16120 44134 16172 44140
rect 16132 43722 16160 44134
rect 16304 43852 16356 43858
rect 16304 43794 16356 43800
rect 16120 43716 16172 43722
rect 16120 43658 16172 43664
rect 15956 43548 16252 43568
rect 16012 43546 16036 43548
rect 16092 43546 16116 43548
rect 16172 43546 16196 43548
rect 16034 43494 16036 43546
rect 16098 43494 16110 43546
rect 16172 43494 16174 43546
rect 16012 43492 16036 43494
rect 16092 43492 16116 43494
rect 16172 43492 16196 43494
rect 15956 43472 16252 43492
rect 16316 43450 16344 43794
rect 16304 43444 16356 43450
rect 16304 43386 16356 43392
rect 15956 42460 16252 42480
rect 16012 42458 16036 42460
rect 16092 42458 16116 42460
rect 16172 42458 16196 42460
rect 16034 42406 16036 42458
rect 16098 42406 16110 42458
rect 16172 42406 16174 42458
rect 16012 42404 16036 42406
rect 16092 42404 16116 42406
rect 16172 42404 16196 42406
rect 15956 42384 16252 42404
rect 16408 41698 16436 67594
rect 16500 58546 16528 74734
rect 17038 73400 17094 73409
rect 17038 73335 17094 73344
rect 16578 69048 16634 69057
rect 16578 68983 16634 68992
rect 16592 67658 16620 68983
rect 16580 67652 16632 67658
rect 16580 67594 16632 67600
rect 16948 66632 17000 66638
rect 16948 66574 17000 66580
rect 16960 66026 16988 66574
rect 16948 66020 17000 66026
rect 16948 65962 17000 65968
rect 17052 63986 17080 73335
rect 17406 73264 17462 73273
rect 17406 73199 17462 73208
rect 17224 66700 17276 66706
rect 17224 66642 17276 66648
rect 17236 65958 17264 66642
rect 17224 65952 17276 65958
rect 17224 65894 17276 65900
rect 17236 65074 17264 65894
rect 17224 65068 17276 65074
rect 17224 65010 17276 65016
rect 17040 63980 17092 63986
rect 17040 63922 17092 63928
rect 16762 63472 16818 63481
rect 16762 63407 16818 63416
rect 16672 62280 16724 62286
rect 16672 62222 16724 62228
rect 16580 62212 16632 62218
rect 16580 62154 16632 62160
rect 16592 61674 16620 62154
rect 16580 61668 16632 61674
rect 16580 61610 16632 61616
rect 16684 61606 16712 62222
rect 16672 61600 16724 61606
rect 16672 61542 16724 61548
rect 16580 61056 16632 61062
rect 16580 60998 16632 61004
rect 16592 60654 16620 60998
rect 16580 60648 16632 60654
rect 16580 60590 16632 60596
rect 16592 59265 16620 60590
rect 16684 59537 16712 61542
rect 16670 59528 16726 59537
rect 16670 59463 16726 59472
rect 16578 59256 16634 59265
rect 16578 59191 16634 59200
rect 16672 58948 16724 58954
rect 16672 58890 16724 58896
rect 16488 58540 16540 58546
rect 16488 58482 16540 58488
rect 16488 58404 16540 58410
rect 16488 58346 16540 58352
rect 16500 56914 16528 58346
rect 16578 58304 16634 58313
rect 16578 58239 16634 58248
rect 16592 57050 16620 58239
rect 16580 57044 16632 57050
rect 16580 56986 16632 56992
rect 16684 56953 16712 58890
rect 16670 56944 16726 56953
rect 16488 56908 16540 56914
rect 16488 56850 16540 56856
rect 16580 56908 16632 56914
rect 16670 56879 16726 56888
rect 16580 56850 16632 56856
rect 16592 56522 16620 56850
rect 16672 56772 16724 56778
rect 16672 56714 16724 56720
rect 16500 56494 16620 56522
rect 16500 56234 16528 56494
rect 16580 56432 16632 56438
rect 16578 56400 16580 56409
rect 16632 56400 16634 56409
rect 16684 56370 16712 56714
rect 16578 56335 16634 56344
rect 16672 56364 16724 56370
rect 16672 56306 16724 56312
rect 16488 56228 16540 56234
rect 16488 56170 16540 56176
rect 16500 55706 16528 56170
rect 16670 56128 16726 56137
rect 16670 56063 16726 56072
rect 16500 55678 16620 55706
rect 16488 55616 16540 55622
rect 16486 55584 16488 55593
rect 16540 55584 16542 55593
rect 16486 55519 16542 55528
rect 16500 55418 16528 55519
rect 16488 55412 16540 55418
rect 16488 55354 16540 55360
rect 16592 55214 16620 55678
rect 16684 55418 16712 56063
rect 16672 55412 16724 55418
rect 16672 55354 16724 55360
rect 16580 55208 16632 55214
rect 16580 55150 16632 55156
rect 16488 54664 16540 54670
rect 16488 54606 16540 54612
rect 16500 53242 16528 54606
rect 16592 54330 16620 55150
rect 16670 54904 16726 54913
rect 16670 54839 16726 54848
rect 16684 54806 16712 54839
rect 16672 54800 16724 54806
rect 16672 54742 16724 54748
rect 16672 54596 16724 54602
rect 16672 54538 16724 54544
rect 16580 54324 16632 54330
rect 16580 54266 16632 54272
rect 16684 53666 16712 54538
rect 16592 53638 16712 53666
rect 16592 53446 16620 53638
rect 16672 53508 16724 53514
rect 16672 53450 16724 53456
rect 16580 53440 16632 53446
rect 16580 53382 16632 53388
rect 16578 53272 16634 53281
rect 16488 53236 16540 53242
rect 16578 53207 16634 53216
rect 16488 53178 16540 53184
rect 16500 52601 16528 53178
rect 16486 52592 16542 52601
rect 16486 52527 16542 52536
rect 16488 52488 16540 52494
rect 16592 52476 16620 53207
rect 16540 52448 16620 52476
rect 16488 52430 16540 52436
rect 16500 51882 16528 52430
rect 16580 52352 16632 52358
rect 16580 52294 16632 52300
rect 16488 51876 16540 51882
rect 16488 51818 16540 51824
rect 16592 51626 16620 52294
rect 16684 51950 16712 53450
rect 16672 51944 16724 51950
rect 16672 51886 16724 51892
rect 16500 51598 16620 51626
rect 16672 51604 16724 51610
rect 16500 51270 16528 51598
rect 16672 51546 16724 51552
rect 16684 51513 16712 51546
rect 16670 51504 16726 51513
rect 16670 51439 16726 51448
rect 16672 51400 16724 51406
rect 16672 51342 16724 51348
rect 16580 51332 16632 51338
rect 16580 51274 16632 51280
rect 16488 51264 16540 51270
rect 16488 51206 16540 51212
rect 16500 50318 16528 51206
rect 16592 50862 16620 51274
rect 16580 50856 16632 50862
rect 16580 50798 16632 50804
rect 16684 50522 16712 51342
rect 16672 50516 16724 50522
rect 16672 50458 16724 50464
rect 16488 50312 16540 50318
rect 16488 50254 16540 50260
rect 16672 50312 16724 50318
rect 16672 50254 16724 50260
rect 16488 49768 16540 49774
rect 16488 49710 16540 49716
rect 16500 49434 16528 49710
rect 16488 49428 16540 49434
rect 16488 49370 16540 49376
rect 16500 48686 16528 49370
rect 16580 49292 16632 49298
rect 16580 49234 16632 49240
rect 16592 48822 16620 49234
rect 16580 48816 16632 48822
rect 16580 48758 16632 48764
rect 16488 48680 16540 48686
rect 16488 48622 16540 48628
rect 16488 47660 16540 47666
rect 16488 47602 16540 47608
rect 16500 47025 16528 47602
rect 16486 47016 16542 47025
rect 16486 46951 16542 46960
rect 16592 46034 16620 48758
rect 16684 48142 16712 50254
rect 16672 48136 16724 48142
rect 16672 48078 16724 48084
rect 16684 47054 16712 48078
rect 16672 47048 16724 47054
rect 16672 46990 16724 46996
rect 16580 46028 16632 46034
rect 16500 45966 16528 45997
rect 16580 45970 16632 45976
rect 16488 45960 16540 45966
rect 16486 45928 16488 45937
rect 16540 45928 16542 45937
rect 16684 45898 16712 46990
rect 16486 45863 16542 45872
rect 16672 45892 16724 45898
rect 16500 45422 16528 45863
rect 16672 45834 16724 45840
rect 16488 45416 16540 45422
rect 16488 45358 16540 45364
rect 16672 44940 16724 44946
rect 16672 44882 16724 44888
rect 16684 44402 16712 44882
rect 16672 44396 16724 44402
rect 16672 44338 16724 44344
rect 16488 44328 16540 44334
rect 16488 44270 16540 44276
rect 16580 44328 16632 44334
rect 16580 44270 16632 44276
rect 16500 43994 16528 44270
rect 16488 43988 16540 43994
rect 16488 43930 16540 43936
rect 16488 43852 16540 43858
rect 16592 43840 16620 44270
rect 16672 44192 16724 44198
rect 16672 44134 16724 44140
rect 16540 43812 16620 43840
rect 16488 43794 16540 43800
rect 16500 43382 16528 43794
rect 16488 43376 16540 43382
rect 16488 43318 16540 43324
rect 16408 41670 16528 41698
rect 15956 41372 16252 41392
rect 16012 41370 16036 41372
rect 16092 41370 16116 41372
rect 16172 41370 16196 41372
rect 16034 41318 16036 41370
rect 16098 41318 16110 41370
rect 16172 41318 16174 41370
rect 16012 41316 16036 41318
rect 16092 41316 16116 41318
rect 16172 41316 16196 41318
rect 15956 41296 16252 41316
rect 16500 41206 16528 41670
rect 16488 41200 16540 41206
rect 16488 41142 16540 41148
rect 16580 41064 16632 41070
rect 16580 41006 16632 41012
rect 16592 40458 16620 41006
rect 16580 40452 16632 40458
rect 16580 40394 16632 40400
rect 15956 40284 16252 40304
rect 16012 40282 16036 40284
rect 16092 40282 16116 40284
rect 16172 40282 16196 40284
rect 16034 40230 16036 40282
rect 16098 40230 16110 40282
rect 16172 40230 16174 40282
rect 16012 40228 16036 40230
rect 16092 40228 16116 40230
rect 16172 40228 16196 40230
rect 15956 40208 16252 40228
rect 15934 40080 15990 40089
rect 15934 40015 15936 40024
rect 15988 40015 15990 40024
rect 15936 39986 15988 39992
rect 16592 39302 16620 40394
rect 16684 39438 16712 44134
rect 16776 40662 16804 63407
rect 17040 60716 17092 60722
rect 17092 60676 17172 60704
rect 17040 60658 17092 60664
rect 16856 60240 16908 60246
rect 16856 60182 16908 60188
rect 16868 59090 16896 60182
rect 17040 60172 17092 60178
rect 17040 60114 17092 60120
rect 17052 59430 17080 60114
rect 17040 59424 17092 59430
rect 17038 59392 17040 59401
rect 17092 59392 17094 59401
rect 17038 59327 17094 59336
rect 16856 59084 16908 59090
rect 16856 59026 16908 59032
rect 17144 58410 17172 60676
rect 17236 60178 17264 65010
rect 17224 60172 17276 60178
rect 17224 60114 17276 60120
rect 17316 59968 17368 59974
rect 17316 59910 17368 59916
rect 17328 59566 17356 59910
rect 17316 59560 17368 59566
rect 17316 59502 17368 59508
rect 17328 58954 17356 59502
rect 17316 58948 17368 58954
rect 17316 58890 17368 58896
rect 17132 58404 17184 58410
rect 17132 58346 17184 58352
rect 17224 58336 17276 58342
rect 17224 58278 17276 58284
rect 17040 58064 17092 58070
rect 17040 58006 17092 58012
rect 16856 57996 16908 58002
rect 16856 57938 16908 57944
rect 16868 57254 16896 57938
rect 17052 57798 17080 58006
rect 17040 57792 17092 57798
rect 17040 57734 17092 57740
rect 17132 57792 17184 57798
rect 17132 57734 17184 57740
rect 17052 57458 17080 57734
rect 17040 57452 17092 57458
rect 17040 57394 17092 57400
rect 16948 57384 17000 57390
rect 16948 57326 17000 57332
rect 16856 57248 16908 57254
rect 16856 57190 16908 57196
rect 16868 55826 16896 57190
rect 16960 56778 16988 57326
rect 17052 57322 17080 57394
rect 17040 57316 17092 57322
rect 17040 57258 17092 57264
rect 17144 57254 17172 57734
rect 17132 57248 17184 57254
rect 17132 57190 17184 57196
rect 16948 56772 17000 56778
rect 16948 56714 17000 56720
rect 16948 56160 17000 56166
rect 16948 56102 17000 56108
rect 16960 55865 16988 56102
rect 16946 55856 17002 55865
rect 16856 55820 16908 55826
rect 16946 55791 17002 55800
rect 16856 55762 16908 55768
rect 16868 55214 16896 55762
rect 16960 55758 16988 55791
rect 16948 55752 17000 55758
rect 16948 55694 17000 55700
rect 17038 55720 17094 55729
rect 16960 55418 16988 55694
rect 17144 55706 17172 57190
rect 17236 56982 17264 58278
rect 17314 57216 17370 57225
rect 17314 57151 17370 57160
rect 17224 56976 17276 56982
rect 17224 56918 17276 56924
rect 17224 56704 17276 56710
rect 17224 56646 17276 56652
rect 17094 55678 17172 55706
rect 17038 55655 17040 55664
rect 17092 55655 17094 55664
rect 17040 55626 17092 55632
rect 16948 55412 17000 55418
rect 16948 55354 17000 55360
rect 17052 55350 17080 55626
rect 17132 55616 17184 55622
rect 17236 55593 17264 56646
rect 17132 55558 17184 55564
rect 17222 55584 17278 55593
rect 17040 55344 17092 55350
rect 17040 55286 17092 55292
rect 16856 55208 16908 55214
rect 16856 55150 16908 55156
rect 16868 54806 16896 55150
rect 17052 55146 17080 55286
rect 17040 55140 17092 55146
rect 17040 55082 17092 55088
rect 17144 54874 17172 55558
rect 17222 55519 17278 55528
rect 17132 54868 17184 54874
rect 17132 54810 17184 54816
rect 16856 54800 16908 54806
rect 17328 54754 17356 57151
rect 16856 54742 16908 54748
rect 17144 54726 17356 54754
rect 16856 53984 16908 53990
rect 16856 53926 16908 53932
rect 16868 50946 16896 53926
rect 16948 53576 17000 53582
rect 16948 53518 17000 53524
rect 16960 53281 16988 53518
rect 17040 53440 17092 53446
rect 17040 53382 17092 53388
rect 16946 53272 17002 53281
rect 17052 53242 17080 53382
rect 16946 53207 17002 53216
rect 17040 53236 17092 53242
rect 17040 53178 17092 53184
rect 16948 53168 17000 53174
rect 16948 53110 17000 53116
rect 16960 53009 16988 53110
rect 16946 53000 17002 53009
rect 16946 52935 17002 52944
rect 17144 52884 17172 54726
rect 17316 53576 17368 53582
rect 17316 53518 17368 53524
rect 16960 52856 17172 52884
rect 17224 52896 17276 52902
rect 17222 52864 17224 52873
rect 17276 52864 17278 52873
rect 16960 51785 16988 52856
rect 17222 52799 17278 52808
rect 17040 52556 17092 52562
rect 17040 52498 17092 52504
rect 17052 51950 17080 52498
rect 17224 52488 17276 52494
rect 17224 52430 17276 52436
rect 17040 51944 17092 51950
rect 17040 51886 17092 51892
rect 16946 51776 17002 51785
rect 16946 51711 17002 51720
rect 17052 51542 17080 51886
rect 17040 51536 17092 51542
rect 17092 51484 17172 51490
rect 17040 51478 17172 51484
rect 17052 51462 17172 51478
rect 17052 51413 17080 51462
rect 17040 51332 17092 51338
rect 17040 51274 17092 51280
rect 16868 50918 16988 50946
rect 16960 50862 16988 50918
rect 16948 50856 17000 50862
rect 16948 50798 17000 50804
rect 16856 49904 16908 49910
rect 16854 49872 16856 49881
rect 16908 49872 16910 49881
rect 16854 49807 16910 49816
rect 16856 49292 16908 49298
rect 16856 49234 16908 49240
rect 16868 48890 16896 49234
rect 16856 48884 16908 48890
rect 16856 48826 16908 48832
rect 16960 48686 16988 50798
rect 16948 48680 17000 48686
rect 16948 48622 17000 48628
rect 16946 48512 17002 48521
rect 16946 48447 17002 48456
rect 16856 48000 16908 48006
rect 16856 47942 16908 47948
rect 16868 47802 16896 47942
rect 16856 47796 16908 47802
rect 16856 47738 16908 47744
rect 16854 45656 16910 45665
rect 16854 45591 16910 45600
rect 16868 45082 16896 45591
rect 16856 45076 16908 45082
rect 16856 45018 16908 45024
rect 16960 44198 16988 48447
rect 17052 47802 17080 51274
rect 17144 50930 17172 51462
rect 17132 50924 17184 50930
rect 17132 50866 17184 50872
rect 17236 49298 17264 52430
rect 17328 50561 17356 53518
rect 17314 50552 17370 50561
rect 17314 50487 17370 50496
rect 17328 50386 17356 50487
rect 17316 50380 17368 50386
rect 17316 50322 17368 50328
rect 17328 49910 17356 50322
rect 17316 49904 17368 49910
rect 17316 49846 17368 49852
rect 17316 49700 17368 49706
rect 17316 49642 17368 49648
rect 17224 49292 17276 49298
rect 17224 49234 17276 49240
rect 17130 48920 17186 48929
rect 17130 48855 17186 48864
rect 17144 48754 17172 48855
rect 17132 48748 17184 48754
rect 17132 48690 17184 48696
rect 17040 47796 17092 47802
rect 17040 47738 17092 47744
rect 17144 47190 17172 48690
rect 17236 48278 17264 49234
rect 17328 48550 17356 49642
rect 17316 48544 17368 48550
rect 17316 48486 17368 48492
rect 17224 48272 17276 48278
rect 17224 48214 17276 48220
rect 17132 47184 17184 47190
rect 17132 47126 17184 47132
rect 17132 46436 17184 46442
rect 17132 46378 17184 46384
rect 17040 46028 17092 46034
rect 17040 45970 17092 45976
rect 17052 45082 17080 45970
rect 17040 45076 17092 45082
rect 17040 45018 17092 45024
rect 16948 44192 17000 44198
rect 16948 44134 17000 44140
rect 17040 43240 17092 43246
rect 17040 43182 17092 43188
rect 17052 42906 17080 43182
rect 17040 42900 17092 42906
rect 17040 42842 17092 42848
rect 16948 41064 17000 41070
rect 16948 41006 17000 41012
rect 16764 40656 16816 40662
rect 16764 40598 16816 40604
rect 16776 40186 16804 40598
rect 16764 40180 16816 40186
rect 16764 40122 16816 40128
rect 16764 39840 16816 39846
rect 16764 39782 16816 39788
rect 16776 39506 16804 39782
rect 16856 39636 16908 39642
rect 16856 39578 16908 39584
rect 16764 39500 16816 39506
rect 16764 39442 16816 39448
rect 16672 39432 16724 39438
rect 16672 39374 16724 39380
rect 16396 39296 16448 39302
rect 16396 39238 16448 39244
rect 16580 39296 16632 39302
rect 16580 39238 16632 39244
rect 15956 39196 16252 39216
rect 16012 39194 16036 39196
rect 16092 39194 16116 39196
rect 16172 39194 16196 39196
rect 16034 39142 16036 39194
rect 16098 39142 16110 39194
rect 16172 39142 16174 39194
rect 16012 39140 16036 39142
rect 16092 39140 16116 39142
rect 16172 39140 16196 39142
rect 15956 39120 16252 39140
rect 16408 38894 16436 39238
rect 16776 39098 16804 39442
rect 16764 39092 16816 39098
rect 16764 39034 16816 39040
rect 16396 38888 16448 38894
rect 16396 38830 16448 38836
rect 16486 38856 16542 38865
rect 16408 38486 16436 38830
rect 16486 38791 16542 38800
rect 16500 38554 16528 38791
rect 16488 38548 16540 38554
rect 16488 38490 16540 38496
rect 16396 38480 16448 38486
rect 16396 38422 16448 38428
rect 16580 38412 16632 38418
rect 16580 38354 16632 38360
rect 16488 38344 16540 38350
rect 16488 38286 16540 38292
rect 16304 38276 16356 38282
rect 16304 38218 16356 38224
rect 15956 38108 16252 38128
rect 16012 38106 16036 38108
rect 16092 38106 16116 38108
rect 16172 38106 16196 38108
rect 16034 38054 16036 38106
rect 16098 38054 16110 38106
rect 16172 38054 16174 38106
rect 16012 38052 16036 38054
rect 16092 38052 16116 38054
rect 16172 38052 16196 38054
rect 15956 38032 16252 38052
rect 16120 37936 16172 37942
rect 16120 37878 16172 37884
rect 15936 37732 15988 37738
rect 15936 37674 15988 37680
rect 15948 37233 15976 37674
rect 16132 37233 16160 37878
rect 16316 37670 16344 38218
rect 16396 38208 16448 38214
rect 16396 38150 16448 38156
rect 16408 37942 16436 38150
rect 16396 37936 16448 37942
rect 16396 37878 16448 37884
rect 16396 37800 16448 37806
rect 16396 37742 16448 37748
rect 16304 37664 16356 37670
rect 16304 37606 16356 37612
rect 15934 37224 15990 37233
rect 15934 37159 15990 37168
rect 16118 37224 16174 37233
rect 16118 37159 16174 37168
rect 15956 37020 16252 37040
rect 16012 37018 16036 37020
rect 16092 37018 16116 37020
rect 16172 37018 16196 37020
rect 16034 36966 16036 37018
rect 16098 36966 16110 37018
rect 16172 36966 16174 37018
rect 16012 36964 16036 36966
rect 16092 36964 16116 36966
rect 16172 36964 16196 36966
rect 15956 36944 16252 36964
rect 16316 36802 16344 37606
rect 16408 37097 16436 37742
rect 16394 37088 16450 37097
rect 16394 37023 16450 37032
rect 16396 36916 16448 36922
rect 16396 36858 16448 36864
rect 16224 36774 16344 36802
rect 16120 36644 16172 36650
rect 16120 36586 16172 36592
rect 15936 36576 15988 36582
rect 15936 36518 15988 36524
rect 15948 36242 15976 36518
rect 16132 36417 16160 36586
rect 16118 36408 16174 36417
rect 16118 36343 16174 36352
rect 15936 36236 15988 36242
rect 15936 36178 15988 36184
rect 16132 36106 16160 36343
rect 16224 36281 16252 36774
rect 16304 36712 16356 36718
rect 16304 36654 16356 36660
rect 16316 36310 16344 36654
rect 16304 36304 16356 36310
rect 16210 36272 16266 36281
rect 16304 36246 16356 36252
rect 16210 36207 16266 36216
rect 16224 36106 16252 36207
rect 16120 36100 16172 36106
rect 16120 36042 16172 36048
rect 16212 36100 16264 36106
rect 16212 36042 16264 36048
rect 16408 36038 16436 36858
rect 16500 36582 16528 38286
rect 16592 38010 16620 38354
rect 16868 38350 16896 39578
rect 16856 38344 16908 38350
rect 16856 38286 16908 38292
rect 16764 38208 16816 38214
rect 16764 38150 16816 38156
rect 16580 38004 16632 38010
rect 16580 37946 16632 37952
rect 16580 37868 16632 37874
rect 16580 37810 16632 37816
rect 16592 37777 16620 37810
rect 16578 37768 16634 37777
rect 16776 37738 16804 38150
rect 16868 38049 16896 38286
rect 16854 38040 16910 38049
rect 16854 37975 16910 37984
rect 16578 37703 16634 37712
rect 16764 37732 16816 37738
rect 16764 37674 16816 37680
rect 16764 37324 16816 37330
rect 16764 37266 16816 37272
rect 16856 37324 16908 37330
rect 16856 37266 16908 37272
rect 16672 37120 16724 37126
rect 16672 37062 16724 37068
rect 16580 36848 16632 36854
rect 16580 36790 16632 36796
rect 16488 36576 16540 36582
rect 16488 36518 16540 36524
rect 16488 36168 16540 36174
rect 16488 36110 16540 36116
rect 16396 36032 16448 36038
rect 16396 35974 16448 35980
rect 15956 35932 16252 35952
rect 16012 35930 16036 35932
rect 16092 35930 16116 35932
rect 16172 35930 16196 35932
rect 16034 35878 16036 35930
rect 16098 35878 16110 35930
rect 16172 35878 16174 35930
rect 16012 35876 16036 35878
rect 16092 35876 16116 35878
rect 16172 35876 16196 35878
rect 15956 35856 16252 35876
rect 16408 35873 16436 35974
rect 16394 35864 16450 35873
rect 16394 35799 16450 35808
rect 16304 35760 16356 35766
rect 15934 35728 15990 35737
rect 16304 35702 16356 35708
rect 15934 35663 15936 35672
rect 15988 35663 15990 35672
rect 15936 35634 15988 35640
rect 15948 35290 15976 35634
rect 16028 35624 16080 35630
rect 16026 35592 16028 35601
rect 16080 35592 16082 35601
rect 16026 35527 16082 35536
rect 15936 35284 15988 35290
rect 15936 35226 15988 35232
rect 15956 34844 16252 34864
rect 16012 34842 16036 34844
rect 16092 34842 16116 34844
rect 16172 34842 16196 34844
rect 16034 34790 16036 34842
rect 16098 34790 16110 34842
rect 16172 34790 16174 34842
rect 16012 34788 16036 34790
rect 16092 34788 16116 34790
rect 16172 34788 16196 34790
rect 15956 34768 16252 34788
rect 15936 34536 15988 34542
rect 15936 34478 15988 34484
rect 15948 33930 15976 34478
rect 15936 33924 15988 33930
rect 15936 33866 15988 33872
rect 15956 33756 16252 33776
rect 16012 33754 16036 33756
rect 16092 33754 16116 33756
rect 16172 33754 16196 33756
rect 16034 33702 16036 33754
rect 16098 33702 16110 33754
rect 16172 33702 16174 33754
rect 16012 33700 16036 33702
rect 16092 33700 16116 33702
rect 16172 33700 16196 33702
rect 15956 33680 16252 33700
rect 16212 33516 16264 33522
rect 16212 33458 16264 33464
rect 15936 33448 15988 33454
rect 16224 33425 16252 33458
rect 15936 33390 15988 33396
rect 16210 33416 16266 33425
rect 15948 33318 15976 33390
rect 16210 33351 16266 33360
rect 15936 33312 15988 33318
rect 15936 33254 15988 33260
rect 16026 33280 16082 33289
rect 16026 33215 16082 33224
rect 16040 33046 16068 33215
rect 16224 33114 16252 33351
rect 16212 33108 16264 33114
rect 16212 33050 16264 33056
rect 16028 33040 16080 33046
rect 15934 33008 15990 33017
rect 16028 32982 16080 32988
rect 15934 32943 15936 32952
rect 15988 32943 15990 32952
rect 16316 32960 16344 35702
rect 16500 35562 16528 36110
rect 16488 35556 16540 35562
rect 16488 35498 16540 35504
rect 16500 35290 16528 35498
rect 16488 35284 16540 35290
rect 16488 35226 16540 35232
rect 16592 35170 16620 36790
rect 16684 36650 16712 37062
rect 16776 36786 16804 37266
rect 16868 36786 16896 37266
rect 16764 36780 16816 36786
rect 16764 36722 16816 36728
rect 16856 36780 16908 36786
rect 16856 36722 16908 36728
rect 16672 36644 16724 36650
rect 16672 36586 16724 36592
rect 16856 36168 16908 36174
rect 16856 36110 16908 36116
rect 16672 36032 16724 36038
rect 16672 35974 16724 35980
rect 16762 36000 16818 36009
rect 16684 35222 16712 35974
rect 16762 35935 16818 35944
rect 16776 35562 16804 35935
rect 16868 35698 16896 36110
rect 16856 35692 16908 35698
rect 16856 35634 16908 35640
rect 16764 35556 16816 35562
rect 16764 35498 16816 35504
rect 16396 35148 16448 35154
rect 16396 35090 16448 35096
rect 16500 35142 16620 35170
rect 16672 35216 16724 35222
rect 16672 35158 16724 35164
rect 16854 35184 16910 35193
rect 16408 33674 16436 35090
rect 16500 34610 16528 35142
rect 16854 35119 16910 35128
rect 16868 35086 16896 35119
rect 16856 35080 16908 35086
rect 16856 35022 16908 35028
rect 16580 35012 16632 35018
rect 16580 34954 16632 34960
rect 16764 35012 16816 35018
rect 16764 34954 16816 34960
rect 16592 34746 16620 34954
rect 16672 34944 16724 34950
rect 16672 34886 16724 34892
rect 16580 34740 16632 34746
rect 16580 34682 16632 34688
rect 16488 34604 16540 34610
rect 16488 34546 16540 34552
rect 16488 34468 16540 34474
rect 16488 34410 16540 34416
rect 16500 34184 16528 34410
rect 16684 34406 16712 34886
rect 16672 34400 16724 34406
rect 16672 34342 16724 34348
rect 16776 34202 16804 34954
rect 16868 34202 16896 35022
rect 16960 34406 16988 41006
rect 17040 39432 17092 39438
rect 17040 39374 17092 39380
rect 17052 38758 17080 39374
rect 17040 38752 17092 38758
rect 17040 38694 17092 38700
rect 16948 34400 17000 34406
rect 16948 34342 17000 34348
rect 16764 34196 16816 34202
rect 16500 34156 16620 34184
rect 16500 33998 16528 34156
rect 16488 33992 16540 33998
rect 16488 33934 16540 33940
rect 16488 33856 16540 33862
rect 16486 33824 16488 33833
rect 16540 33824 16542 33833
rect 16486 33759 16542 33768
rect 16408 33646 16528 33674
rect 16500 32994 16528 33646
rect 16592 33114 16620 34156
rect 16764 34138 16816 34144
rect 16856 34196 16908 34202
rect 16856 34138 16908 34144
rect 16672 34060 16724 34066
rect 16672 34002 16724 34008
rect 16580 33108 16632 33114
rect 16580 33050 16632 33056
rect 16500 32966 16620 32994
rect 16316 32932 16436 32960
rect 15936 32914 15988 32920
rect 16304 32836 16356 32842
rect 16304 32778 16356 32784
rect 15956 32668 16252 32688
rect 16012 32666 16036 32668
rect 16092 32666 16116 32668
rect 16172 32666 16196 32668
rect 16034 32614 16036 32666
rect 16098 32614 16110 32666
rect 16172 32614 16174 32666
rect 16012 32612 16036 32614
rect 16092 32612 16116 32614
rect 16172 32612 16196 32614
rect 15956 32592 16252 32612
rect 15844 32428 15896 32434
rect 15844 32370 15896 32376
rect 15844 31884 15896 31890
rect 15844 31826 15896 31832
rect 15856 31754 15884 31826
rect 15844 31748 15896 31754
rect 15844 31690 15896 31696
rect 15750 31648 15806 31657
rect 15750 31583 15806 31592
rect 15956 31580 16252 31600
rect 16012 31578 16036 31580
rect 16092 31578 16116 31580
rect 16172 31578 16196 31580
rect 16034 31526 16036 31578
rect 16098 31526 16110 31578
rect 16172 31526 16174 31578
rect 16012 31524 16036 31526
rect 16092 31524 16116 31526
rect 16172 31524 16196 31526
rect 15956 31504 16252 31524
rect 15672 31436 15792 31464
rect 15658 31376 15714 31385
rect 15658 31311 15714 31320
rect 15568 31136 15620 31142
rect 15568 31078 15620 31084
rect 15580 28082 15608 31078
rect 15672 28642 15700 31311
rect 15764 29850 15792 31436
rect 16316 31346 16344 32778
rect 16408 31521 16436 32932
rect 16488 32904 16540 32910
rect 16488 32846 16540 32852
rect 16394 31512 16450 31521
rect 16394 31447 16396 31456
rect 16448 31447 16450 31456
rect 16396 31418 16448 31424
rect 16408 31387 16436 31418
rect 15844 31340 15896 31346
rect 15844 31282 15896 31288
rect 16304 31340 16356 31346
rect 16304 31282 16356 31288
rect 15752 29844 15804 29850
rect 15752 29786 15804 29792
rect 15752 29504 15804 29510
rect 15750 29472 15752 29481
rect 15804 29472 15806 29481
rect 15750 29407 15806 29416
rect 15750 29336 15806 29345
rect 15750 29271 15806 29280
rect 15764 29102 15792 29271
rect 15752 29096 15804 29102
rect 15752 29038 15804 29044
rect 15752 28960 15804 28966
rect 15752 28902 15804 28908
rect 15764 28762 15792 28902
rect 15752 28756 15804 28762
rect 15752 28698 15804 28704
rect 15672 28614 15792 28642
rect 15660 28552 15712 28558
rect 15660 28494 15712 28500
rect 15568 28076 15620 28082
rect 15568 28018 15620 28024
rect 15568 27940 15620 27946
rect 15568 27882 15620 27888
rect 15292 27668 15344 27674
rect 15292 27610 15344 27616
rect 15396 27662 15516 27690
rect 15292 27328 15344 27334
rect 15292 27270 15344 27276
rect 15304 24750 15332 27270
rect 15292 24744 15344 24750
rect 15292 24686 15344 24692
rect 15292 24336 15344 24342
rect 15292 24278 15344 24284
rect 15304 23730 15332 24278
rect 15292 23724 15344 23730
rect 15292 23666 15344 23672
rect 15292 23588 15344 23594
rect 15292 23530 15344 23536
rect 15304 23322 15332 23530
rect 15292 23316 15344 23322
rect 15292 23258 15344 23264
rect 15290 23216 15346 23225
rect 15290 23151 15346 23160
rect 15304 23118 15332 23151
rect 15292 23112 15344 23118
rect 15292 23054 15344 23060
rect 15304 22574 15332 23054
rect 15396 22681 15424 27662
rect 15476 27600 15528 27606
rect 15476 27542 15528 27548
rect 15488 26926 15516 27542
rect 15580 27305 15608 27882
rect 15566 27296 15622 27305
rect 15566 27231 15622 27240
rect 15568 27124 15620 27130
rect 15568 27066 15620 27072
rect 15476 26920 15528 26926
rect 15476 26862 15528 26868
rect 15488 26518 15516 26862
rect 15476 26512 15528 26518
rect 15476 26454 15528 26460
rect 15580 26450 15608 27066
rect 15568 26444 15620 26450
rect 15568 26386 15620 26392
rect 15476 26376 15528 26382
rect 15476 26318 15528 26324
rect 15488 25702 15516 26318
rect 15476 25696 15528 25702
rect 15476 25638 15528 25644
rect 15488 24070 15516 25638
rect 15580 25498 15608 26386
rect 15568 25492 15620 25498
rect 15568 25434 15620 25440
rect 15566 25120 15622 25129
rect 15566 25055 15622 25064
rect 15580 24614 15608 25055
rect 15672 24993 15700 28494
rect 15764 27130 15792 28614
rect 15752 27124 15804 27130
rect 15752 27066 15804 27072
rect 15856 26908 15884 31282
rect 16500 31278 16528 32846
rect 16592 32774 16620 32966
rect 16580 32768 16632 32774
rect 16580 32710 16632 32716
rect 16592 31414 16620 32710
rect 16684 32570 16712 34002
rect 16776 33969 16804 34138
rect 16856 34060 16908 34066
rect 16856 34002 16908 34008
rect 16948 34060 17000 34066
rect 16948 34002 17000 34008
rect 16762 33960 16818 33969
rect 16762 33895 16818 33904
rect 16868 32910 16896 34002
rect 16960 33386 16988 34002
rect 16948 33380 17000 33386
rect 16948 33322 17000 33328
rect 16856 32904 16908 32910
rect 16856 32846 16908 32852
rect 16672 32564 16724 32570
rect 16672 32506 16724 32512
rect 16856 32360 16908 32366
rect 16856 32302 16908 32308
rect 16670 32192 16726 32201
rect 16670 32127 16726 32136
rect 16580 31408 16632 31414
rect 16580 31350 16632 31356
rect 16488 31272 16540 31278
rect 16580 31272 16632 31278
rect 16488 31214 16540 31220
rect 16578 31240 16580 31249
rect 16632 31240 16634 31249
rect 16578 31175 16634 31184
rect 16394 30968 16450 30977
rect 16684 30938 16712 32127
rect 16762 32056 16818 32065
rect 16762 31991 16818 32000
rect 16776 31482 16804 31991
rect 16868 31890 16896 32302
rect 16948 32224 17000 32230
rect 16948 32166 17000 32172
rect 16856 31884 16908 31890
rect 16856 31826 16908 31832
rect 16764 31476 16816 31482
rect 16764 31418 16816 31424
rect 16856 31204 16908 31210
rect 16856 31146 16908 31152
rect 16394 30903 16450 30912
rect 16672 30932 16724 30938
rect 16304 30660 16356 30666
rect 16304 30602 16356 30608
rect 15956 30492 16252 30512
rect 16012 30490 16036 30492
rect 16092 30490 16116 30492
rect 16172 30490 16196 30492
rect 16034 30438 16036 30490
rect 16098 30438 16110 30490
rect 16172 30438 16174 30490
rect 16012 30436 16036 30438
rect 16092 30436 16116 30438
rect 16172 30436 16196 30438
rect 15956 30416 16252 30436
rect 16316 30326 16344 30602
rect 16304 30320 16356 30326
rect 16304 30262 16356 30268
rect 15936 30184 15988 30190
rect 15934 30152 15936 30161
rect 15988 30152 15990 30161
rect 15934 30087 15990 30096
rect 16212 29776 16264 29782
rect 16212 29718 16264 29724
rect 16224 29617 16252 29718
rect 16304 29640 16356 29646
rect 16210 29608 16266 29617
rect 16304 29582 16356 29588
rect 16210 29543 16266 29552
rect 15956 29404 16252 29424
rect 16012 29402 16036 29404
rect 16092 29402 16116 29404
rect 16172 29402 16196 29404
rect 16034 29350 16036 29402
rect 16098 29350 16110 29402
rect 16172 29350 16174 29402
rect 16012 29348 16036 29350
rect 16092 29348 16116 29350
rect 16172 29348 16196 29350
rect 15956 29328 16252 29348
rect 16120 28960 16172 28966
rect 16120 28902 16172 28908
rect 16026 28792 16082 28801
rect 16026 28727 16082 28736
rect 16040 28694 16068 28727
rect 16028 28688 16080 28694
rect 15934 28656 15990 28665
rect 16028 28630 16080 28636
rect 15934 28591 15990 28600
rect 15948 28490 15976 28591
rect 16132 28490 16160 28902
rect 16316 28762 16344 29582
rect 16408 29306 16436 30903
rect 16672 30874 16724 30880
rect 16762 30832 16818 30841
rect 16762 30767 16818 30776
rect 16580 30728 16632 30734
rect 16672 30728 16724 30734
rect 16580 30670 16632 30676
rect 16670 30696 16672 30705
rect 16724 30696 16726 30705
rect 16486 30288 16542 30297
rect 16486 30223 16542 30232
rect 16500 30190 16528 30223
rect 16488 30184 16540 30190
rect 16488 30126 16540 30132
rect 16592 29714 16620 30670
rect 16670 30631 16726 30640
rect 16670 30560 16726 30569
rect 16670 30495 16726 30504
rect 16684 30122 16712 30495
rect 16672 30116 16724 30122
rect 16672 30058 16724 30064
rect 16488 29708 16540 29714
rect 16488 29650 16540 29656
rect 16580 29708 16632 29714
rect 16580 29650 16632 29656
rect 16396 29300 16448 29306
rect 16396 29242 16448 29248
rect 16408 28801 16436 29242
rect 16394 28792 16450 28801
rect 16304 28756 16356 28762
rect 16394 28727 16450 28736
rect 16500 28778 16528 29650
rect 16672 29640 16724 29646
rect 16672 29582 16724 29588
rect 16578 29336 16634 29345
rect 16578 29271 16634 29280
rect 16592 29102 16620 29271
rect 16580 29096 16632 29102
rect 16580 29038 16632 29044
rect 16500 28762 16620 28778
rect 16500 28756 16632 28762
rect 16500 28750 16580 28756
rect 16304 28698 16356 28704
rect 15936 28484 15988 28490
rect 15936 28426 15988 28432
rect 16120 28484 16172 28490
rect 16120 28426 16172 28432
rect 15956 28316 16252 28336
rect 16012 28314 16036 28316
rect 16092 28314 16116 28316
rect 16172 28314 16196 28316
rect 16034 28262 16036 28314
rect 16098 28262 16110 28314
rect 16172 28262 16174 28314
rect 16012 28260 16036 28262
rect 16092 28260 16116 28262
rect 16172 28260 16196 28262
rect 15956 28240 16252 28260
rect 15934 28112 15990 28121
rect 15934 28047 15990 28056
rect 15948 28014 15976 28047
rect 15936 28008 15988 28014
rect 15936 27950 15988 27956
rect 16212 28008 16264 28014
rect 16212 27950 16264 27956
rect 16224 27674 16252 27950
rect 16212 27668 16264 27674
rect 16212 27610 16264 27616
rect 16224 27441 16252 27610
rect 16316 27606 16344 28698
rect 16396 28620 16448 28626
rect 16396 28562 16448 28568
rect 16408 28218 16436 28562
rect 16396 28212 16448 28218
rect 16396 28154 16448 28160
rect 16408 27713 16436 28154
rect 16394 27704 16450 27713
rect 16394 27639 16450 27648
rect 16304 27600 16356 27606
rect 16304 27542 16356 27548
rect 16396 27600 16448 27606
rect 16396 27542 16448 27548
rect 16210 27432 16266 27441
rect 16210 27367 16266 27376
rect 16304 27328 16356 27334
rect 16304 27270 16356 27276
rect 15956 27228 16252 27248
rect 16012 27226 16036 27228
rect 16092 27226 16116 27228
rect 16172 27226 16196 27228
rect 16034 27174 16036 27226
rect 16098 27174 16110 27226
rect 16172 27174 16174 27226
rect 16012 27172 16036 27174
rect 16092 27172 16116 27174
rect 16172 27172 16196 27174
rect 15956 27152 16252 27172
rect 15764 26880 15884 26908
rect 15658 24984 15714 24993
rect 15658 24919 15714 24928
rect 15568 24608 15620 24614
rect 15568 24550 15620 24556
rect 15476 24064 15528 24070
rect 15476 24006 15528 24012
rect 15488 22982 15516 24006
rect 15476 22976 15528 22982
rect 15476 22918 15528 22924
rect 15382 22672 15438 22681
rect 15382 22607 15438 22616
rect 15292 22568 15344 22574
rect 15292 22510 15344 22516
rect 15476 22500 15528 22506
rect 15476 22442 15528 22448
rect 15384 22432 15436 22438
rect 15384 22374 15436 22380
rect 15290 21992 15346 22001
rect 15290 21927 15346 21936
rect 15304 16182 15332 21927
rect 15396 20482 15424 22374
rect 15488 21010 15516 22442
rect 15580 21185 15608 24550
rect 15660 23248 15712 23254
rect 15660 23190 15712 23196
rect 15672 22574 15700 23190
rect 15660 22568 15712 22574
rect 15660 22510 15712 22516
rect 15672 21593 15700 22510
rect 15658 21584 15714 21593
rect 15658 21519 15714 21528
rect 15660 21412 15712 21418
rect 15660 21354 15712 21360
rect 15566 21176 15622 21185
rect 15566 21111 15622 21120
rect 15476 21004 15528 21010
rect 15476 20946 15528 20952
rect 15568 21004 15620 21010
rect 15568 20946 15620 20952
rect 15488 20602 15516 20946
rect 15476 20596 15528 20602
rect 15476 20538 15528 20544
rect 15396 20454 15516 20482
rect 15382 19544 15438 19553
rect 15382 19479 15438 19488
rect 15396 17338 15424 19479
rect 15384 17332 15436 17338
rect 15384 17274 15436 17280
rect 15488 16658 15516 20454
rect 15580 19174 15608 20946
rect 15672 20806 15700 21354
rect 15660 20800 15712 20806
rect 15660 20742 15712 20748
rect 15568 19168 15620 19174
rect 15568 19110 15620 19116
rect 15580 18222 15608 19110
rect 15568 18216 15620 18222
rect 15568 18158 15620 18164
rect 15566 17912 15622 17921
rect 15566 17847 15568 17856
rect 15620 17847 15622 17856
rect 15568 17818 15620 17824
rect 15672 17762 15700 20742
rect 15764 19922 15792 26880
rect 16316 26382 16344 27270
rect 16408 27169 16436 27542
rect 16394 27160 16450 27169
rect 16394 27095 16396 27104
rect 16448 27095 16450 27104
rect 16396 27066 16448 27072
rect 16500 26586 16528 28750
rect 16580 28698 16632 28704
rect 16684 28642 16712 29582
rect 16776 29578 16804 30767
rect 16868 29889 16896 31146
rect 16854 29880 16910 29889
rect 16854 29815 16910 29824
rect 16856 29708 16908 29714
rect 16856 29650 16908 29656
rect 16764 29572 16816 29578
rect 16764 29514 16816 29520
rect 16776 29306 16804 29514
rect 16868 29306 16896 29650
rect 16764 29300 16816 29306
rect 16764 29242 16816 29248
rect 16856 29300 16908 29306
rect 16856 29242 16908 29248
rect 16854 29064 16910 29073
rect 16854 28999 16910 29008
rect 16762 28928 16818 28937
rect 16762 28863 16818 28872
rect 16592 28614 16712 28642
rect 16592 28422 16620 28614
rect 16580 28416 16632 28422
rect 16580 28358 16632 28364
rect 16592 26994 16620 28358
rect 16670 28248 16726 28257
rect 16776 28218 16804 28863
rect 16868 28558 16896 28999
rect 16856 28552 16908 28558
rect 16856 28494 16908 28500
rect 16670 28183 16726 28192
rect 16764 28212 16816 28218
rect 16684 27946 16712 28183
rect 16764 28154 16816 28160
rect 16762 27976 16818 27985
rect 16672 27940 16724 27946
rect 16762 27911 16818 27920
rect 16672 27882 16724 27888
rect 16670 27568 16726 27577
rect 16670 27503 16672 27512
rect 16724 27503 16726 27512
rect 16672 27474 16724 27480
rect 16670 27432 16726 27441
rect 16670 27367 16726 27376
rect 16580 26988 16632 26994
rect 16580 26930 16632 26936
rect 16488 26580 16540 26586
rect 16488 26522 16540 26528
rect 16684 26450 16712 27367
rect 16672 26444 16724 26450
rect 16672 26386 16724 26392
rect 15844 26376 15896 26382
rect 15844 26318 15896 26324
rect 16304 26376 16356 26382
rect 16304 26318 16356 26324
rect 15856 24721 15884 26318
rect 16672 26240 16724 26246
rect 16672 26182 16724 26188
rect 15956 26140 16252 26160
rect 16012 26138 16036 26140
rect 16092 26138 16116 26140
rect 16172 26138 16196 26140
rect 16034 26086 16036 26138
rect 16098 26086 16110 26138
rect 16172 26086 16174 26138
rect 16012 26084 16036 26086
rect 16092 26084 16116 26086
rect 16172 26084 16196 26086
rect 15956 26064 16252 26084
rect 16684 25838 16712 26182
rect 16672 25832 16724 25838
rect 16672 25774 16724 25780
rect 16028 25764 16080 25770
rect 16028 25706 16080 25712
rect 16040 25498 16068 25706
rect 16212 25696 16264 25702
rect 16210 25664 16212 25673
rect 16304 25696 16356 25702
rect 16264 25664 16266 25673
rect 16304 25638 16356 25644
rect 16210 25599 16266 25608
rect 16028 25492 16080 25498
rect 16028 25434 16080 25440
rect 15956 25052 16252 25072
rect 16012 25050 16036 25052
rect 16092 25050 16116 25052
rect 16172 25050 16196 25052
rect 16034 24998 16036 25050
rect 16098 24998 16110 25050
rect 16172 24998 16174 25050
rect 16012 24996 16036 24998
rect 16092 24996 16116 24998
rect 16172 24996 16196 24998
rect 15956 24976 16252 24996
rect 15842 24712 15898 24721
rect 15842 24647 15898 24656
rect 16316 24274 16344 25638
rect 16396 25288 16448 25294
rect 16396 25230 16448 25236
rect 16408 24750 16436 25230
rect 16580 25152 16632 25158
rect 16580 25094 16632 25100
rect 16592 24954 16620 25094
rect 16580 24948 16632 24954
rect 16580 24890 16632 24896
rect 16684 24834 16712 25774
rect 16776 25702 16804 27911
rect 16868 26586 16896 28494
rect 16960 26976 16988 32166
rect 17052 29170 17080 38694
rect 17040 29164 17092 29170
rect 17040 29106 17092 29112
rect 17040 29028 17092 29034
rect 17040 28970 17092 28976
rect 17052 28937 17080 28970
rect 17038 28928 17094 28937
rect 17038 28863 17094 28872
rect 17052 28694 17080 28863
rect 17040 28688 17092 28694
rect 17040 28630 17092 28636
rect 17040 28416 17092 28422
rect 17040 28358 17092 28364
rect 17052 27334 17080 28358
rect 17040 27328 17092 27334
rect 17040 27270 17092 27276
rect 16960 26948 17080 26976
rect 16948 26852 17000 26858
rect 16948 26794 17000 26800
rect 16960 26586 16988 26794
rect 16856 26580 16908 26586
rect 16856 26522 16908 26528
rect 16948 26580 17000 26586
rect 16948 26522 17000 26528
rect 16948 26308 17000 26314
rect 16948 26250 17000 26256
rect 16856 25832 16908 25838
rect 16856 25774 16908 25780
rect 16764 25696 16816 25702
rect 16764 25638 16816 25644
rect 16764 25356 16816 25362
rect 16764 25298 16816 25304
rect 16776 24954 16804 25298
rect 16868 25158 16896 25774
rect 16856 25152 16908 25158
rect 16856 25094 16908 25100
rect 16764 24948 16816 24954
rect 16764 24890 16816 24896
rect 16500 24806 16712 24834
rect 16396 24744 16448 24750
rect 16396 24686 16448 24692
rect 16304 24268 16356 24274
rect 16304 24210 16356 24216
rect 15956 23964 16252 23984
rect 16012 23962 16036 23964
rect 16092 23962 16116 23964
rect 16172 23962 16196 23964
rect 16034 23910 16036 23962
rect 16098 23910 16110 23962
rect 16172 23910 16174 23962
rect 16012 23908 16036 23910
rect 16092 23908 16116 23910
rect 16172 23908 16196 23910
rect 15956 23888 16252 23908
rect 16316 23866 16344 24210
rect 16304 23860 16356 23866
rect 16304 23802 16356 23808
rect 16396 23860 16448 23866
rect 16396 23802 16448 23808
rect 16304 23656 16356 23662
rect 16304 23598 16356 23604
rect 16316 22982 16344 23598
rect 16304 22976 16356 22982
rect 16304 22918 16356 22924
rect 15956 22876 16252 22896
rect 16012 22874 16036 22876
rect 16092 22874 16116 22876
rect 16172 22874 16196 22876
rect 16034 22822 16036 22874
rect 16098 22822 16110 22874
rect 16172 22822 16174 22874
rect 16012 22820 16036 22822
rect 16092 22820 16116 22822
rect 16172 22820 16196 22822
rect 15956 22800 16252 22820
rect 16304 22704 16356 22710
rect 16304 22646 16356 22652
rect 15844 22432 15896 22438
rect 15844 22374 15896 22380
rect 15752 19916 15804 19922
rect 15752 19858 15804 19864
rect 15764 19514 15792 19858
rect 15752 19508 15804 19514
rect 15752 19450 15804 19456
rect 15764 18970 15792 19450
rect 15752 18964 15804 18970
rect 15752 18906 15804 18912
rect 15764 18358 15792 18906
rect 15752 18352 15804 18358
rect 15752 18294 15804 18300
rect 15580 17734 15700 17762
rect 15580 17377 15608 17734
rect 15752 17672 15804 17678
rect 15752 17614 15804 17620
rect 15566 17368 15622 17377
rect 15566 17303 15568 17312
rect 15620 17303 15622 17312
rect 15568 17274 15620 17280
rect 15764 17134 15792 17614
rect 15752 17128 15804 17134
rect 15752 17070 15804 17076
rect 15568 16788 15620 16794
rect 15568 16730 15620 16736
rect 15476 16652 15528 16658
rect 15476 16594 15528 16600
rect 15292 16176 15344 16182
rect 15292 16118 15344 16124
rect 15382 16008 15438 16017
rect 15382 15943 15438 15952
rect 15396 14074 15424 15943
rect 15488 15638 15516 16594
rect 15580 16046 15608 16730
rect 15856 16658 15884 22374
rect 15956 21788 16252 21808
rect 16012 21786 16036 21788
rect 16092 21786 16116 21788
rect 16172 21786 16196 21788
rect 16034 21734 16036 21786
rect 16098 21734 16110 21786
rect 16172 21734 16174 21786
rect 16012 21732 16036 21734
rect 16092 21732 16116 21734
rect 16172 21732 16196 21734
rect 15956 21712 16252 21732
rect 16316 21690 16344 22646
rect 16408 22438 16436 23802
rect 16500 23798 16528 24806
rect 16856 24608 16908 24614
rect 16856 24550 16908 24556
rect 16868 24138 16896 24550
rect 16856 24132 16908 24138
rect 16856 24074 16908 24080
rect 16488 23792 16540 23798
rect 16486 23760 16488 23769
rect 16540 23760 16542 23769
rect 16486 23695 16542 23704
rect 16670 23760 16726 23769
rect 16670 23695 16726 23704
rect 16486 23624 16542 23633
rect 16486 23559 16542 23568
rect 16500 23186 16528 23559
rect 16488 23180 16540 23186
rect 16488 23122 16540 23128
rect 16500 22710 16528 23122
rect 16488 22704 16540 22710
rect 16488 22646 16540 22652
rect 16684 22506 16712 23695
rect 16856 23520 16908 23526
rect 16856 23462 16908 23468
rect 16764 22976 16816 22982
rect 16764 22918 16816 22924
rect 16672 22500 16724 22506
rect 16592 22438 16620 22469
rect 16672 22442 16724 22448
rect 16396 22432 16448 22438
rect 16580 22432 16632 22438
rect 16396 22374 16448 22380
rect 16578 22400 16580 22409
rect 16632 22400 16634 22409
rect 16578 22335 16634 22344
rect 16592 22234 16620 22335
rect 16580 22228 16632 22234
rect 16580 22170 16632 22176
rect 16776 22098 16804 22918
rect 16580 22092 16632 22098
rect 16580 22034 16632 22040
rect 16764 22092 16816 22098
rect 16764 22034 16816 22040
rect 16488 22024 16540 22030
rect 16488 21966 16540 21972
rect 16304 21684 16356 21690
rect 16304 21626 16356 21632
rect 16396 21684 16448 21690
rect 16396 21626 16448 21632
rect 16210 21448 16266 21457
rect 16210 21383 16266 21392
rect 16224 21350 16252 21383
rect 15936 21344 15988 21350
rect 15936 21286 15988 21292
rect 16212 21344 16264 21350
rect 16212 21286 16264 21292
rect 15948 21010 15976 21286
rect 15936 21004 15988 21010
rect 15936 20946 15988 20952
rect 16304 20936 16356 20942
rect 16304 20878 16356 20884
rect 15956 20700 16252 20720
rect 16012 20698 16036 20700
rect 16092 20698 16116 20700
rect 16172 20698 16196 20700
rect 16034 20646 16036 20698
rect 16098 20646 16110 20698
rect 16172 20646 16174 20698
rect 16012 20644 16036 20646
rect 16092 20644 16116 20646
rect 16172 20644 16196 20646
rect 15956 20624 16252 20644
rect 16212 20460 16264 20466
rect 16212 20402 16264 20408
rect 16224 19700 16252 20402
rect 16316 19922 16344 20878
rect 16304 19916 16356 19922
rect 16304 19858 16356 19864
rect 16224 19672 16344 19700
rect 15956 19612 16252 19632
rect 16012 19610 16036 19612
rect 16092 19610 16116 19612
rect 16172 19610 16196 19612
rect 16034 19558 16036 19610
rect 16098 19558 16110 19610
rect 16172 19558 16174 19610
rect 16012 19556 16036 19558
rect 16092 19556 16116 19558
rect 16172 19556 16196 19558
rect 15956 19536 16252 19556
rect 16316 19496 16344 19672
rect 16224 19468 16344 19496
rect 16224 19310 16252 19468
rect 16212 19304 16264 19310
rect 16212 19246 16264 19252
rect 16224 18970 16252 19246
rect 16212 18964 16264 18970
rect 16212 18906 16264 18912
rect 16304 18828 16356 18834
rect 16304 18770 16356 18776
rect 15956 18524 16252 18544
rect 16012 18522 16036 18524
rect 16092 18522 16116 18524
rect 16172 18522 16196 18524
rect 16034 18470 16036 18522
rect 16098 18470 16110 18522
rect 16172 18470 16174 18522
rect 16012 18468 16036 18470
rect 16092 18468 16116 18470
rect 16172 18468 16196 18470
rect 15956 18448 16252 18468
rect 16316 18426 16344 18770
rect 16304 18420 16356 18426
rect 16304 18362 16356 18368
rect 16316 17882 16344 18362
rect 16304 17876 16356 17882
rect 16304 17818 16356 17824
rect 15956 17436 16252 17456
rect 16012 17434 16036 17436
rect 16092 17434 16116 17436
rect 16172 17434 16196 17436
rect 16034 17382 16036 17434
rect 16098 17382 16110 17434
rect 16172 17382 16174 17434
rect 16012 17380 16036 17382
rect 16092 17380 16116 17382
rect 16172 17380 16196 17382
rect 15956 17360 16252 17380
rect 16316 17338 16344 17818
rect 16304 17332 16356 17338
rect 16304 17274 16356 17280
rect 15844 16652 15896 16658
rect 15844 16594 15896 16600
rect 15856 16250 15884 16594
rect 15956 16348 16252 16368
rect 16012 16346 16036 16348
rect 16092 16346 16116 16348
rect 16172 16346 16196 16348
rect 16034 16294 16036 16346
rect 16098 16294 16110 16346
rect 16172 16294 16174 16346
rect 16012 16292 16036 16294
rect 16092 16292 16116 16294
rect 16172 16292 16196 16294
rect 15956 16272 16252 16292
rect 15844 16244 15896 16250
rect 15844 16186 15896 16192
rect 16210 16144 16266 16153
rect 16210 16079 16266 16088
rect 15568 16040 15620 16046
rect 15568 15982 15620 15988
rect 15844 16040 15896 16046
rect 15844 15982 15896 15988
rect 15856 15706 15884 15982
rect 15844 15700 15896 15706
rect 15844 15642 15896 15648
rect 15476 15632 15528 15638
rect 15474 15600 15476 15609
rect 15528 15600 15530 15609
rect 16224 15570 16252 16079
rect 15474 15535 15530 15544
rect 16212 15564 16264 15570
rect 16264 15524 16344 15552
rect 16212 15506 16264 15512
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 15764 14278 15792 15438
rect 15956 15260 16252 15280
rect 16012 15258 16036 15260
rect 16092 15258 16116 15260
rect 16172 15258 16196 15260
rect 16034 15206 16036 15258
rect 16098 15206 16110 15258
rect 16172 15206 16174 15258
rect 16012 15204 16036 15206
rect 16092 15204 16116 15206
rect 16172 15204 16196 15206
rect 15956 15184 16252 15204
rect 16316 15162 16344 15524
rect 16304 15156 16356 15162
rect 16304 15098 16356 15104
rect 16316 14550 16344 15098
rect 16304 14544 16356 14550
rect 16304 14486 16356 14492
rect 15752 14272 15804 14278
rect 15752 14214 15804 14220
rect 15384 14068 15436 14074
rect 15384 14010 15436 14016
rect 15396 13870 15424 14010
rect 15566 13968 15622 13977
rect 15566 13903 15568 13912
rect 15620 13903 15622 13912
rect 15568 13874 15620 13880
rect 15384 13864 15436 13870
rect 15384 13806 15436 13812
rect 15382 12200 15438 12209
rect 15292 12164 15344 12170
rect 15764 12170 15792 14214
rect 15956 14172 16252 14192
rect 16012 14170 16036 14172
rect 16092 14170 16116 14172
rect 16172 14170 16196 14172
rect 16034 14118 16036 14170
rect 16098 14118 16110 14170
rect 16172 14118 16174 14170
rect 16012 14116 16036 14118
rect 16092 14116 16116 14118
rect 16172 14116 16196 14118
rect 15956 14096 16252 14116
rect 15956 13084 16252 13104
rect 16012 13082 16036 13084
rect 16092 13082 16116 13084
rect 16172 13082 16196 13084
rect 16034 13030 16036 13082
rect 16098 13030 16110 13082
rect 16172 13030 16174 13082
rect 16012 13028 16036 13030
rect 16092 13028 16116 13030
rect 16172 13028 16196 13030
rect 15956 13008 16252 13028
rect 15382 12135 15438 12144
rect 15752 12164 15804 12170
rect 15292 12106 15344 12112
rect 15304 11150 15332 12106
rect 15396 11898 15424 12135
rect 15752 12106 15804 12112
rect 15568 12096 15620 12102
rect 15568 12038 15620 12044
rect 15844 12096 15896 12102
rect 15844 12038 15896 12044
rect 15384 11892 15436 11898
rect 15384 11834 15436 11840
rect 15580 11762 15608 12038
rect 15752 11824 15804 11830
rect 15752 11766 15804 11772
rect 15856 11778 15884 12038
rect 15956 11996 16252 12016
rect 16012 11994 16036 11996
rect 16092 11994 16116 11996
rect 16172 11994 16196 11996
rect 16034 11942 16036 11994
rect 16098 11942 16110 11994
rect 16172 11942 16174 11994
rect 16012 11940 16036 11942
rect 16092 11940 16116 11942
rect 16172 11940 16196 11942
rect 15956 11920 16252 11940
rect 15568 11756 15620 11762
rect 15568 11698 15620 11704
rect 15292 11144 15344 11150
rect 15292 11086 15344 11092
rect 15304 10470 15332 11086
rect 15292 10464 15344 10470
rect 15292 10406 15344 10412
rect 15304 9518 15332 10406
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15304 8956 15332 9454
rect 15488 9110 15516 9522
rect 15476 9104 15528 9110
rect 15476 9046 15528 9052
rect 15304 8928 15516 8956
rect 15488 8838 15516 8928
rect 15476 8832 15528 8838
rect 15476 8774 15528 8780
rect 15198 8256 15254 8265
rect 15198 8191 15254 8200
rect 15488 8129 15516 8774
rect 15580 8634 15608 11698
rect 15660 11620 15712 11626
rect 15660 11562 15712 11568
rect 15672 11218 15700 11562
rect 15660 11212 15712 11218
rect 15660 11154 15712 11160
rect 15672 10810 15700 11154
rect 15660 10804 15712 10810
rect 15660 10746 15712 10752
rect 15764 10062 15792 11766
rect 15856 11750 15976 11778
rect 15948 11694 15976 11750
rect 15936 11688 15988 11694
rect 15936 11630 15988 11636
rect 15948 11354 15976 11630
rect 15936 11348 15988 11354
rect 15936 11290 15988 11296
rect 15956 10908 16252 10928
rect 16012 10906 16036 10908
rect 16092 10906 16116 10908
rect 16172 10906 16196 10908
rect 16034 10854 16036 10906
rect 16098 10854 16110 10906
rect 16172 10854 16174 10906
rect 16012 10852 16036 10854
rect 16092 10852 16116 10854
rect 16172 10852 16196 10854
rect 15956 10832 16252 10852
rect 16408 10282 16436 21626
rect 16500 21486 16528 21966
rect 16488 21480 16540 21486
rect 16488 21422 16540 21428
rect 16488 21344 16540 21350
rect 16488 21286 16540 21292
rect 16500 21146 16528 21286
rect 16488 21140 16540 21146
rect 16488 21082 16540 21088
rect 16500 20534 16528 21082
rect 16488 20528 16540 20534
rect 16488 20470 16540 20476
rect 16592 20398 16620 22034
rect 16672 21888 16724 21894
rect 16672 21830 16724 21836
rect 16684 21486 16712 21830
rect 16776 21690 16804 22034
rect 16764 21684 16816 21690
rect 16764 21626 16816 21632
rect 16672 21480 16724 21486
rect 16672 21422 16724 21428
rect 16684 21146 16712 21422
rect 16764 21412 16816 21418
rect 16764 21354 16816 21360
rect 16672 21140 16724 21146
rect 16672 21082 16724 21088
rect 16672 20936 16724 20942
rect 16670 20904 16672 20913
rect 16776 20924 16804 21354
rect 16724 20904 16804 20924
rect 16726 20896 16804 20904
rect 16868 20856 16896 23462
rect 16960 21298 16988 26250
rect 17052 22030 17080 26948
rect 17040 22024 17092 22030
rect 17040 21966 17092 21972
rect 17144 21876 17172 46378
rect 17236 46170 17264 48214
rect 17328 47977 17356 48486
rect 17314 47968 17370 47977
rect 17314 47903 17370 47912
rect 17316 47728 17368 47734
rect 17316 47670 17368 47676
rect 17328 47122 17356 47670
rect 17316 47116 17368 47122
rect 17316 47058 17368 47064
rect 17328 46714 17356 47058
rect 17316 46708 17368 46714
rect 17316 46650 17368 46656
rect 17420 46186 17448 73199
rect 17590 71088 17646 71097
rect 17590 71023 17646 71032
rect 17604 66570 17632 71023
rect 17682 67824 17738 67833
rect 17682 67759 17738 67768
rect 17592 66564 17644 66570
rect 17592 66506 17644 66512
rect 17592 66020 17644 66026
rect 17592 65962 17644 65968
rect 17604 65550 17632 65962
rect 17592 65544 17644 65550
rect 17592 65486 17644 65492
rect 17604 64938 17632 65486
rect 17592 64932 17644 64938
rect 17592 64874 17644 64880
rect 17500 61192 17552 61198
rect 17500 61134 17552 61140
rect 17512 60722 17540 61134
rect 17500 60716 17552 60722
rect 17500 60658 17552 60664
rect 17512 59770 17540 60658
rect 17500 59764 17552 59770
rect 17500 59706 17552 59712
rect 17604 59242 17632 64874
rect 17696 61826 17724 67759
rect 18616 67674 18644 75239
rect 18786 71496 18842 71505
rect 18786 71431 18842 71440
rect 18616 67646 18736 67674
rect 18602 67552 18658 67561
rect 18602 67487 18658 67496
rect 17868 66700 17920 66706
rect 17868 66642 17920 66648
rect 17880 66178 17908 66642
rect 18052 66496 18104 66502
rect 18052 66438 18104 66444
rect 17880 66150 18000 66178
rect 18064 66162 18092 66438
rect 17774 66056 17830 66065
rect 17774 65991 17776 66000
rect 17828 65991 17830 66000
rect 17776 65962 17828 65968
rect 17972 65618 18000 66150
rect 18052 66156 18104 66162
rect 18052 66098 18104 66104
rect 18616 65686 18644 67487
rect 18604 65680 18656 65686
rect 18604 65622 18656 65628
rect 17868 65612 17920 65618
rect 17868 65554 17920 65560
rect 17960 65612 18012 65618
rect 17960 65554 18012 65560
rect 18236 65612 18288 65618
rect 18236 65554 18288 65560
rect 17880 65210 17908 65554
rect 17868 65204 17920 65210
rect 17868 65146 17920 65152
rect 18248 64977 18276 65554
rect 18708 65521 18736 67646
rect 18694 65512 18750 65521
rect 18694 65447 18750 65456
rect 18234 64968 18290 64977
rect 18234 64903 18236 64912
rect 18288 64903 18290 64912
rect 18236 64874 18288 64880
rect 18602 64016 18658 64025
rect 18602 63951 18604 63960
rect 18656 63951 18658 63960
rect 18604 63922 18656 63928
rect 18800 63481 18828 71431
rect 18892 70417 18920 79200
rect 19812 79098 19840 79200
rect 19812 79070 20116 79098
rect 19340 76968 19392 76974
rect 19340 76910 19392 76916
rect 19352 76820 19380 76910
rect 19260 76792 19380 76820
rect 19260 76430 19288 76792
rect 19248 76424 19300 76430
rect 19248 76366 19300 76372
rect 19156 74792 19208 74798
rect 19260 74746 19288 76366
rect 19208 74740 19288 74746
rect 19156 74734 19288 74740
rect 19168 74718 19288 74734
rect 19260 74458 19288 74718
rect 19248 74452 19300 74458
rect 19248 74394 19300 74400
rect 19706 72720 19762 72729
rect 19706 72655 19762 72664
rect 18878 70408 18934 70417
rect 18878 70343 18934 70352
rect 19062 68912 19118 68921
rect 19062 68847 19118 68856
rect 18880 66496 18932 66502
rect 18880 66438 18932 66444
rect 18892 64025 18920 66438
rect 18878 64016 18934 64025
rect 18878 63951 18934 63960
rect 18892 63918 18920 63951
rect 18880 63912 18932 63918
rect 18880 63854 18932 63860
rect 18892 63578 18920 63854
rect 18880 63572 18932 63578
rect 18880 63514 18932 63520
rect 18786 63472 18842 63481
rect 18786 63407 18842 63416
rect 17958 62792 18014 62801
rect 17958 62727 18014 62736
rect 17868 62212 17920 62218
rect 17868 62154 17920 62160
rect 17696 61798 17816 61826
rect 17684 61600 17736 61606
rect 17684 61542 17736 61548
rect 17696 60314 17724 61542
rect 17788 61146 17816 61798
rect 17880 61334 17908 62154
rect 17868 61328 17920 61334
rect 17868 61270 17920 61276
rect 17788 61118 17908 61146
rect 17972 61130 18000 62727
rect 18052 61600 18104 61606
rect 18052 61542 18104 61548
rect 18788 61600 18840 61606
rect 18788 61542 18840 61548
rect 18064 61266 18092 61542
rect 18052 61260 18104 61266
rect 18052 61202 18104 61208
rect 17684 60308 17736 60314
rect 17684 60250 17736 60256
rect 17684 60036 17736 60042
rect 17684 59978 17736 59984
rect 17696 59702 17724 59978
rect 17684 59696 17736 59702
rect 17684 59638 17736 59644
rect 17512 59214 17632 59242
rect 17512 57769 17540 59214
rect 17592 59152 17644 59158
rect 17590 59120 17592 59129
rect 17644 59120 17646 59129
rect 17696 59090 17724 59638
rect 17590 59055 17646 59064
rect 17684 59084 17736 59090
rect 17684 59026 17736 59032
rect 17774 58984 17830 58993
rect 17774 58919 17830 58928
rect 17684 58404 17736 58410
rect 17684 58346 17736 58352
rect 17592 58064 17644 58070
rect 17592 58006 17644 58012
rect 17604 57934 17632 58006
rect 17592 57928 17644 57934
rect 17592 57870 17644 57876
rect 17592 57792 17644 57798
rect 17498 57760 17554 57769
rect 17592 57734 17644 57740
rect 17498 57695 17554 57704
rect 17604 57254 17632 57734
rect 17696 57594 17724 58346
rect 17788 57934 17816 58919
rect 17776 57928 17828 57934
rect 17776 57870 17828 57876
rect 17684 57588 17736 57594
rect 17684 57530 17736 57536
rect 17592 57248 17644 57254
rect 17592 57190 17644 57196
rect 17604 56710 17632 57190
rect 17776 56840 17828 56846
rect 17776 56782 17828 56788
rect 17500 56704 17552 56710
rect 17500 56646 17552 56652
rect 17592 56704 17644 56710
rect 17592 56646 17644 56652
rect 17512 56438 17540 56646
rect 17500 56432 17552 56438
rect 17500 56374 17552 56380
rect 17512 55962 17540 56374
rect 17500 55956 17552 55962
rect 17500 55898 17552 55904
rect 17500 55140 17552 55146
rect 17500 55082 17552 55088
rect 17512 54670 17540 55082
rect 17604 54874 17632 56646
rect 17788 56370 17816 56782
rect 17776 56364 17828 56370
rect 17776 56306 17828 56312
rect 17776 55888 17828 55894
rect 17774 55856 17776 55865
rect 17828 55856 17830 55865
rect 17774 55791 17830 55800
rect 17774 55448 17830 55457
rect 17774 55383 17830 55392
rect 17592 54868 17644 54874
rect 17592 54810 17644 54816
rect 17500 54664 17552 54670
rect 17500 54606 17552 54612
rect 17604 53582 17632 54810
rect 17684 54800 17736 54806
rect 17684 54742 17736 54748
rect 17696 53990 17724 54742
rect 17684 53984 17736 53990
rect 17684 53926 17736 53932
rect 17592 53576 17644 53582
rect 17592 53518 17644 53524
rect 17592 52964 17644 52970
rect 17592 52906 17644 52912
rect 17604 52340 17632 52906
rect 17512 52312 17632 52340
rect 17512 50454 17540 52312
rect 17590 52184 17646 52193
rect 17590 52119 17646 52128
rect 17604 51338 17632 52119
rect 17592 51332 17644 51338
rect 17592 51274 17644 51280
rect 17592 51060 17644 51066
rect 17592 51002 17644 51008
rect 17500 50448 17552 50454
rect 17500 50390 17552 50396
rect 17512 49978 17540 50390
rect 17500 49972 17552 49978
rect 17500 49914 17552 49920
rect 17512 48385 17540 49914
rect 17604 49366 17632 51002
rect 17696 50833 17724 53926
rect 17788 53718 17816 55383
rect 17776 53712 17828 53718
rect 17776 53654 17828 53660
rect 17776 53440 17828 53446
rect 17776 53382 17828 53388
rect 17788 53242 17816 53382
rect 17776 53236 17828 53242
rect 17776 53178 17828 53184
rect 17788 52562 17816 53178
rect 17776 52556 17828 52562
rect 17776 52498 17828 52504
rect 17776 51468 17828 51474
rect 17776 51410 17828 51416
rect 17682 50824 17738 50833
rect 17682 50759 17738 50768
rect 17592 49360 17644 49366
rect 17592 49302 17644 49308
rect 17696 48618 17724 50759
rect 17788 50454 17816 51410
rect 17776 50448 17828 50454
rect 17776 50390 17828 50396
rect 17776 49768 17828 49774
rect 17776 49710 17828 49716
rect 17788 49434 17816 49710
rect 17776 49428 17828 49434
rect 17776 49370 17828 49376
rect 17684 48612 17736 48618
rect 17684 48554 17736 48560
rect 17498 48376 17554 48385
rect 17696 48328 17724 48554
rect 17776 48544 17828 48550
rect 17776 48486 17828 48492
rect 17498 48311 17554 48320
rect 17512 47410 17540 48311
rect 17604 48300 17724 48328
rect 17604 47734 17632 48300
rect 17684 48204 17736 48210
rect 17684 48146 17736 48152
rect 17592 47728 17644 47734
rect 17592 47670 17644 47676
rect 17592 47592 17644 47598
rect 17590 47560 17592 47569
rect 17644 47560 17646 47569
rect 17590 47495 17646 47504
rect 17512 47382 17632 47410
rect 17500 47252 17552 47258
rect 17500 47194 17552 47200
rect 17224 46164 17276 46170
rect 17224 46106 17276 46112
rect 17328 46158 17448 46186
rect 17512 46170 17540 47194
rect 17604 46986 17632 47382
rect 17696 47297 17724 48146
rect 17682 47288 17738 47297
rect 17682 47223 17738 47232
rect 17788 47190 17816 48486
rect 17776 47184 17828 47190
rect 17776 47126 17828 47132
rect 17592 46980 17644 46986
rect 17592 46922 17644 46928
rect 17684 46708 17736 46714
rect 17684 46650 17736 46656
rect 17500 46164 17552 46170
rect 17236 45626 17264 46106
rect 17224 45620 17276 45626
rect 17224 45562 17276 45568
rect 17224 45416 17276 45422
rect 17224 45358 17276 45364
rect 17236 44713 17264 45358
rect 17222 44704 17278 44713
rect 17222 44639 17278 44648
rect 17222 43888 17278 43897
rect 17222 43823 17278 43832
rect 17236 43625 17264 43823
rect 17222 43616 17278 43625
rect 17222 43551 17278 43560
rect 17224 40520 17276 40526
rect 17224 40462 17276 40468
rect 17236 39982 17264 40462
rect 17224 39976 17276 39982
rect 17224 39918 17276 39924
rect 17236 39438 17264 39918
rect 17328 39642 17356 46158
rect 17500 46106 17552 46112
rect 17696 45626 17724 46650
rect 17774 45792 17830 45801
rect 17774 45727 17830 45736
rect 17684 45620 17736 45626
rect 17684 45562 17736 45568
rect 17788 45558 17816 45727
rect 17776 45552 17828 45558
rect 17776 45494 17828 45500
rect 17408 45484 17460 45490
rect 17408 45426 17460 45432
rect 17420 43450 17448 45426
rect 17592 45348 17644 45354
rect 17592 45290 17644 45296
rect 17498 44432 17554 44441
rect 17498 44367 17500 44376
rect 17552 44367 17554 44376
rect 17500 44338 17552 44344
rect 17604 44010 17632 45290
rect 17684 44940 17736 44946
rect 17684 44882 17736 44888
rect 17696 44198 17724 44882
rect 17776 44804 17828 44810
rect 17776 44746 17828 44752
rect 17684 44192 17736 44198
rect 17682 44160 17684 44169
rect 17736 44160 17738 44169
rect 17682 44095 17738 44104
rect 17500 43988 17552 43994
rect 17604 43982 17724 44010
rect 17500 43930 17552 43936
rect 17408 43444 17460 43450
rect 17408 43386 17460 43392
rect 17512 42906 17540 43930
rect 17592 43920 17644 43926
rect 17590 43888 17592 43897
rect 17644 43888 17646 43897
rect 17696 43858 17724 43982
rect 17788 43858 17816 44746
rect 17590 43823 17646 43832
rect 17684 43852 17736 43858
rect 17684 43794 17736 43800
rect 17776 43852 17828 43858
rect 17776 43794 17828 43800
rect 17696 43450 17724 43794
rect 17684 43444 17736 43450
rect 17684 43386 17736 43392
rect 17684 43308 17736 43314
rect 17684 43250 17736 43256
rect 17500 42900 17552 42906
rect 17500 42842 17552 42848
rect 17696 42770 17724 43250
rect 17788 43246 17816 43794
rect 17776 43240 17828 43246
rect 17776 43182 17828 43188
rect 17684 42764 17736 42770
rect 17684 42706 17736 42712
rect 17696 42294 17724 42706
rect 17788 42362 17816 43182
rect 17776 42356 17828 42362
rect 17776 42298 17828 42304
rect 17684 42288 17736 42294
rect 17684 42230 17736 42236
rect 17696 41818 17724 42230
rect 17408 41812 17460 41818
rect 17408 41754 17460 41760
rect 17684 41812 17736 41818
rect 17684 41754 17736 41760
rect 17420 40526 17448 41754
rect 17408 40520 17460 40526
rect 17408 40462 17460 40468
rect 17316 39636 17368 39642
rect 17316 39578 17368 39584
rect 17224 39432 17276 39438
rect 17224 39374 17276 39380
rect 17788 38962 17816 42298
rect 17776 38956 17828 38962
rect 17776 38898 17828 38904
rect 17408 38208 17460 38214
rect 17408 38150 17460 38156
rect 17316 37800 17368 37806
rect 17316 37742 17368 37748
rect 17222 37360 17278 37369
rect 17222 37295 17278 37304
rect 17236 37126 17264 37295
rect 17224 37120 17276 37126
rect 17224 37062 17276 37068
rect 17236 36854 17264 37062
rect 17224 36848 17276 36854
rect 17224 36790 17276 36796
rect 17236 36106 17264 36790
rect 17224 36100 17276 36106
rect 17224 36042 17276 36048
rect 17236 35834 17264 36042
rect 17224 35828 17276 35834
rect 17224 35770 17276 35776
rect 17236 35630 17264 35770
rect 17224 35624 17276 35630
rect 17224 35566 17276 35572
rect 17224 35216 17276 35222
rect 17328 35204 17356 37742
rect 17420 37670 17448 38150
rect 17500 37732 17552 37738
rect 17500 37674 17552 37680
rect 17408 37664 17460 37670
rect 17408 37606 17460 37612
rect 17408 37324 17460 37330
rect 17408 37266 17460 37272
rect 17276 35176 17356 35204
rect 17224 35158 17276 35164
rect 17236 34513 17264 35158
rect 17222 34504 17278 34513
rect 17222 34439 17278 34448
rect 17224 34400 17276 34406
rect 17224 34342 17276 34348
rect 17236 31793 17264 34342
rect 17316 33992 17368 33998
rect 17316 33934 17368 33940
rect 17222 31784 17278 31793
rect 17222 31719 17278 31728
rect 17222 30288 17278 30297
rect 17222 30223 17224 30232
rect 17276 30223 17278 30232
rect 17224 30194 17276 30200
rect 17236 29238 17264 30194
rect 17224 29232 17276 29238
rect 17224 29174 17276 29180
rect 17224 29096 17276 29102
rect 17224 29038 17276 29044
rect 17236 28694 17264 29038
rect 17224 28688 17276 28694
rect 17224 28630 17276 28636
rect 17224 28552 17276 28558
rect 17222 28520 17224 28529
rect 17276 28520 17278 28529
rect 17222 28455 17278 28464
rect 17236 28218 17264 28455
rect 17224 28212 17276 28218
rect 17224 28154 17276 28160
rect 17224 26920 17276 26926
rect 17224 26862 17276 26868
rect 17236 23526 17264 26862
rect 17224 23520 17276 23526
rect 17224 23462 17276 23468
rect 17144 21848 17264 21876
rect 16960 21270 17172 21298
rect 16946 21176 17002 21185
rect 16946 21111 17002 21120
rect 16670 20839 16726 20848
rect 16776 20828 16896 20856
rect 16672 20800 16724 20806
rect 16672 20742 16724 20748
rect 16684 20602 16712 20742
rect 16672 20596 16724 20602
rect 16672 20538 16724 20544
rect 16670 20496 16726 20505
rect 16670 20431 16726 20440
rect 16580 20392 16632 20398
rect 16500 20352 16580 20380
rect 16500 20058 16528 20352
rect 16580 20334 16632 20340
rect 16488 20052 16540 20058
rect 16488 19994 16540 20000
rect 16580 19984 16632 19990
rect 16580 19926 16632 19932
rect 16488 19848 16540 19854
rect 16488 19790 16540 19796
rect 16500 19378 16528 19790
rect 16488 19372 16540 19378
rect 16488 19314 16540 19320
rect 16592 18834 16620 19926
rect 16684 18850 16712 20431
rect 16776 20262 16804 20828
rect 16856 20392 16908 20398
rect 16856 20334 16908 20340
rect 16764 20256 16816 20262
rect 16764 20198 16816 20204
rect 16764 19848 16816 19854
rect 16764 19790 16816 19796
rect 16776 19281 16804 19790
rect 16868 19718 16896 20334
rect 16856 19712 16908 19718
rect 16856 19654 16908 19660
rect 16868 19514 16896 19654
rect 16856 19508 16908 19514
rect 16856 19450 16908 19456
rect 16856 19372 16908 19378
rect 16856 19314 16908 19320
rect 16762 19272 16818 19281
rect 16762 19207 16818 19216
rect 16776 19174 16804 19207
rect 16764 19168 16816 19174
rect 16764 19110 16816 19116
rect 16580 18828 16632 18834
rect 16684 18822 16804 18850
rect 16580 18770 16632 18776
rect 16488 18624 16540 18630
rect 16488 18566 16540 18572
rect 16580 18624 16632 18630
rect 16580 18566 16632 18572
rect 16500 18358 16528 18566
rect 16488 18352 16540 18358
rect 16488 18294 16540 18300
rect 16500 17882 16528 18294
rect 16592 18290 16620 18566
rect 16580 18284 16632 18290
rect 16580 18226 16632 18232
rect 16488 17876 16540 17882
rect 16540 17836 16620 17864
rect 16488 17818 16540 17824
rect 16488 17740 16540 17746
rect 16488 17682 16540 17688
rect 16500 17270 16528 17682
rect 16488 17264 16540 17270
rect 16488 17206 16540 17212
rect 16592 17202 16620 17836
rect 16580 17196 16632 17202
rect 16580 17138 16632 17144
rect 16672 17060 16724 17066
rect 16672 17002 16724 17008
rect 16684 16794 16712 17002
rect 16672 16788 16724 16794
rect 16672 16730 16724 16736
rect 16776 16658 16804 18822
rect 16580 16652 16632 16658
rect 16580 16594 16632 16600
rect 16764 16652 16816 16658
rect 16764 16594 16816 16600
rect 16592 16250 16620 16594
rect 16580 16244 16632 16250
rect 16580 16186 16632 16192
rect 16868 15745 16896 19314
rect 16960 17202 16988 21111
rect 17038 19952 17094 19961
rect 17038 19887 17094 19896
rect 17052 19281 17080 19887
rect 17144 19514 17172 21270
rect 17132 19508 17184 19514
rect 17132 19450 17184 19456
rect 17130 19408 17186 19417
rect 17130 19343 17186 19352
rect 17038 19272 17094 19281
rect 17038 19207 17094 19216
rect 17144 18630 17172 19343
rect 17132 18624 17184 18630
rect 17132 18566 17184 18572
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 16854 15736 16910 15745
rect 16854 15671 16910 15680
rect 17132 14884 17184 14890
rect 17132 14826 17184 14832
rect 17144 14482 17172 14826
rect 17132 14476 17184 14482
rect 17132 14418 17184 14424
rect 17144 14074 17172 14418
rect 17132 14068 17184 14074
rect 17132 14010 17184 14016
rect 16948 12300 17000 12306
rect 16948 12242 17000 12248
rect 16960 11898 16988 12242
rect 16948 11892 17000 11898
rect 16948 11834 17000 11840
rect 16960 11354 16988 11834
rect 17236 11801 17264 21848
rect 17328 18426 17356 33934
rect 17420 29288 17448 37266
rect 17512 36038 17540 37674
rect 17776 37256 17828 37262
rect 17776 37198 17828 37204
rect 17592 37188 17644 37194
rect 17592 37130 17644 37136
rect 17684 37188 17736 37194
rect 17684 37130 17736 37136
rect 17604 36310 17632 37130
rect 17696 36922 17724 37130
rect 17684 36916 17736 36922
rect 17684 36858 17736 36864
rect 17682 36816 17738 36825
rect 17682 36751 17738 36760
rect 17592 36304 17644 36310
rect 17592 36246 17644 36252
rect 17592 36168 17644 36174
rect 17592 36110 17644 36116
rect 17500 36032 17552 36038
rect 17500 35974 17552 35980
rect 17604 35612 17632 36110
rect 17512 35584 17632 35612
rect 17512 35068 17540 35584
rect 17590 35320 17646 35329
rect 17590 35255 17646 35264
rect 17604 35222 17632 35255
rect 17592 35216 17644 35222
rect 17592 35158 17644 35164
rect 17512 35040 17632 35068
rect 17500 34944 17552 34950
rect 17500 34886 17552 34892
rect 17512 33114 17540 34886
rect 17500 33108 17552 33114
rect 17500 33050 17552 33056
rect 17500 32904 17552 32910
rect 17500 32846 17552 32852
rect 17512 32230 17540 32846
rect 17500 32224 17552 32230
rect 17500 32166 17552 32172
rect 17500 31816 17552 31822
rect 17500 31758 17552 31764
rect 17512 31657 17540 31758
rect 17498 31648 17554 31657
rect 17498 31583 17554 31592
rect 17500 30320 17552 30326
rect 17498 30288 17500 30297
rect 17552 30288 17554 30297
rect 17498 30223 17554 30232
rect 17500 30048 17552 30054
rect 17500 29990 17552 29996
rect 17512 29850 17540 29990
rect 17500 29844 17552 29850
rect 17500 29786 17552 29792
rect 17420 29260 17540 29288
rect 17408 29164 17460 29170
rect 17408 29106 17460 29112
rect 17420 21554 17448 29106
rect 17512 26314 17540 29260
rect 17604 28665 17632 35040
rect 17696 31906 17724 36751
rect 17788 36242 17816 37198
rect 17776 36236 17828 36242
rect 17776 36178 17828 36184
rect 17776 35760 17828 35766
rect 17776 35702 17828 35708
rect 17788 35193 17816 35702
rect 17774 35184 17830 35193
rect 17774 35119 17830 35128
rect 17776 34672 17828 34678
rect 17776 34614 17828 34620
rect 17788 32745 17816 34614
rect 17774 32736 17830 32745
rect 17774 32671 17830 32680
rect 17776 32360 17828 32366
rect 17776 32302 17828 32308
rect 17788 32026 17816 32302
rect 17776 32020 17828 32026
rect 17776 31962 17828 31968
rect 17696 31878 17816 31906
rect 17682 31784 17738 31793
rect 17682 31719 17738 31728
rect 17590 28656 17646 28665
rect 17590 28591 17646 28600
rect 17592 28552 17644 28558
rect 17592 28494 17644 28500
rect 17604 28082 17632 28494
rect 17592 28076 17644 28082
rect 17592 28018 17644 28024
rect 17590 27704 17646 27713
rect 17590 27639 17592 27648
rect 17644 27639 17646 27648
rect 17592 27610 17644 27616
rect 17592 27532 17644 27538
rect 17592 27474 17644 27480
rect 17604 26761 17632 27474
rect 17590 26752 17646 26761
rect 17590 26687 17646 26696
rect 17592 26376 17644 26382
rect 17592 26318 17644 26324
rect 17500 26308 17552 26314
rect 17500 26250 17552 26256
rect 17604 25702 17632 26318
rect 17592 25696 17644 25702
rect 17592 25638 17644 25644
rect 17500 24404 17552 24410
rect 17500 24346 17552 24352
rect 17512 24070 17540 24346
rect 17696 24154 17724 31719
rect 17788 29782 17816 31878
rect 17776 29776 17828 29782
rect 17776 29718 17828 29724
rect 17776 29640 17828 29646
rect 17776 29582 17828 29588
rect 17788 29102 17816 29582
rect 17776 29096 17828 29102
rect 17776 29038 17828 29044
rect 17788 27538 17816 29038
rect 17776 27532 17828 27538
rect 17776 27474 17828 27480
rect 17776 27328 17828 27334
rect 17776 27270 17828 27276
rect 17788 26450 17816 27270
rect 17776 26444 17828 26450
rect 17776 26386 17828 26392
rect 17788 26042 17816 26386
rect 17776 26036 17828 26042
rect 17776 25978 17828 25984
rect 17776 25764 17828 25770
rect 17776 25706 17828 25712
rect 17604 24126 17724 24154
rect 17500 24064 17552 24070
rect 17500 24006 17552 24012
rect 17500 22024 17552 22030
rect 17500 21966 17552 21972
rect 17408 21548 17460 21554
rect 17408 21490 17460 21496
rect 17408 20596 17460 20602
rect 17408 20538 17460 20544
rect 17420 19922 17448 20538
rect 17408 19916 17460 19922
rect 17408 19858 17460 19864
rect 17408 19304 17460 19310
rect 17408 19246 17460 19252
rect 17420 18630 17448 19246
rect 17408 18624 17460 18630
rect 17408 18566 17460 18572
rect 17316 18420 17368 18426
rect 17316 18362 17368 18368
rect 17328 18222 17356 18362
rect 17316 18216 17368 18222
rect 17316 18158 17368 18164
rect 17420 18034 17448 18566
rect 17328 18006 17448 18034
rect 17328 17542 17356 18006
rect 17408 17740 17460 17746
rect 17408 17682 17460 17688
rect 17316 17536 17368 17542
rect 17316 17478 17368 17484
rect 17328 16998 17356 17478
rect 17420 17134 17448 17682
rect 17408 17128 17460 17134
rect 17406 17096 17408 17105
rect 17460 17096 17462 17105
rect 17406 17031 17462 17040
rect 17316 16992 17368 16998
rect 17316 16934 17368 16940
rect 17316 16652 17368 16658
rect 17316 16594 17368 16600
rect 17328 16250 17356 16594
rect 17408 16448 17460 16454
rect 17408 16390 17460 16396
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 17316 15360 17368 15366
rect 17316 15302 17368 15308
rect 17328 14958 17356 15302
rect 17316 14952 17368 14958
rect 17316 14894 17368 14900
rect 17420 14657 17448 16390
rect 17406 14648 17462 14657
rect 17406 14583 17462 14592
rect 17408 14476 17460 14482
rect 17408 14418 17460 14424
rect 17420 14074 17448 14418
rect 17408 14068 17460 14074
rect 17408 14010 17460 14016
rect 17512 13705 17540 21966
rect 17604 14482 17632 24126
rect 17788 21842 17816 25706
rect 17696 21814 17816 21842
rect 17696 21690 17724 21814
rect 17684 21684 17736 21690
rect 17684 21626 17736 21632
rect 17776 21616 17828 21622
rect 17682 21584 17738 21593
rect 17776 21558 17828 21564
rect 17682 21519 17684 21528
rect 17736 21519 17738 21528
rect 17684 21490 17736 21496
rect 17696 20602 17724 21490
rect 17684 20596 17736 20602
rect 17684 20538 17736 20544
rect 17788 19174 17816 21558
rect 17776 19168 17828 19174
rect 17776 19110 17828 19116
rect 17684 18828 17736 18834
rect 17684 18770 17736 18776
rect 17696 18426 17724 18770
rect 17684 18420 17736 18426
rect 17684 18362 17736 18368
rect 17684 15904 17736 15910
rect 17684 15846 17736 15852
rect 17592 14476 17644 14482
rect 17592 14418 17644 14424
rect 17604 14006 17632 14418
rect 17592 14000 17644 14006
rect 17592 13942 17644 13948
rect 17498 13696 17554 13705
rect 17498 13631 17554 13640
rect 17222 11792 17278 11801
rect 17222 11727 17278 11736
rect 16948 11348 17000 11354
rect 16948 11290 17000 11296
rect 16316 10254 16436 10282
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15474 8120 15530 8129
rect 15474 8055 15530 8064
rect 15764 5846 15792 9998
rect 15956 9820 16252 9840
rect 16012 9818 16036 9820
rect 16092 9818 16116 9820
rect 16172 9818 16196 9820
rect 16034 9766 16036 9818
rect 16098 9766 16110 9818
rect 16172 9766 16174 9818
rect 16012 9764 16036 9766
rect 16092 9764 16116 9766
rect 16172 9764 16196 9766
rect 15956 9744 16252 9764
rect 16316 9489 16344 10254
rect 16396 10124 16448 10130
rect 16396 10066 16448 10072
rect 16408 9722 16436 10066
rect 16488 10056 16540 10062
rect 16488 9998 16540 10004
rect 16396 9716 16448 9722
rect 16396 9658 16448 9664
rect 16500 9518 16528 9998
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16488 9512 16540 9518
rect 16302 9480 16358 9489
rect 16488 9454 16540 9460
rect 16302 9415 16358 9424
rect 16592 9042 16620 9862
rect 17038 9072 17094 9081
rect 16580 9036 16632 9042
rect 16580 8978 16632 8984
rect 16948 9036 17000 9042
rect 17604 9042 17632 13942
rect 17038 9007 17040 9016
rect 16948 8978 17000 8984
rect 17092 9007 17094 9016
rect 17592 9036 17644 9042
rect 17040 8978 17092 8984
rect 17592 8978 17644 8984
rect 16488 8900 16540 8906
rect 16488 8842 16540 8848
rect 15956 8732 16252 8752
rect 16012 8730 16036 8732
rect 16092 8730 16116 8732
rect 16172 8730 16196 8732
rect 16034 8678 16036 8730
rect 16098 8678 16110 8730
rect 16172 8678 16174 8730
rect 16012 8676 16036 8678
rect 16092 8676 16116 8678
rect 16172 8676 16196 8678
rect 15956 8656 16252 8676
rect 16500 8537 16528 8842
rect 16592 8634 16620 8978
rect 16854 8936 16910 8945
rect 16854 8871 16910 8880
rect 16580 8628 16632 8634
rect 16580 8570 16632 8576
rect 16486 8528 16542 8537
rect 16486 8463 16542 8472
rect 16868 7954 16896 8871
rect 16960 8634 16988 8978
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 17052 8566 17080 8978
rect 17040 8560 17092 8566
rect 17040 8502 17092 8508
rect 17038 8392 17094 8401
rect 17038 8327 17094 8336
rect 16856 7948 16908 7954
rect 16856 7890 16908 7896
rect 15956 7644 16252 7664
rect 16012 7642 16036 7644
rect 16092 7642 16116 7644
rect 16172 7642 16196 7644
rect 16034 7590 16036 7642
rect 16098 7590 16110 7642
rect 16172 7590 16174 7642
rect 16012 7588 16036 7590
rect 16092 7588 16116 7590
rect 16172 7588 16196 7590
rect 15956 7568 16252 7588
rect 16868 7546 16896 7890
rect 16948 7880 17000 7886
rect 16948 7822 17000 7828
rect 16960 7546 16988 7822
rect 16856 7540 16908 7546
rect 16856 7482 16908 7488
rect 16948 7540 17000 7546
rect 16948 7482 17000 7488
rect 15956 6556 16252 6576
rect 16012 6554 16036 6556
rect 16092 6554 16116 6556
rect 16172 6554 16196 6556
rect 16034 6502 16036 6554
rect 16098 6502 16110 6554
rect 16172 6502 16174 6554
rect 16012 6500 16036 6502
rect 16092 6500 16116 6502
rect 16172 6500 16196 6502
rect 15956 6480 16252 6500
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 15936 6112 15988 6118
rect 15936 6054 15988 6060
rect 15292 5840 15344 5846
rect 15292 5782 15344 5788
rect 15752 5840 15804 5846
rect 15752 5782 15804 5788
rect 15304 5370 15332 5782
rect 15948 5778 15976 6054
rect 16316 5778 16344 6258
rect 15936 5772 15988 5778
rect 15936 5714 15988 5720
rect 16304 5772 16356 5778
rect 16304 5714 16356 5720
rect 15948 5658 15976 5714
rect 15660 5636 15712 5642
rect 15660 5578 15712 5584
rect 15856 5630 15976 5658
rect 15568 5568 15620 5574
rect 15568 5510 15620 5516
rect 15292 5364 15344 5370
rect 15292 5306 15344 5312
rect 15108 4140 15160 4146
rect 15108 4082 15160 4088
rect 15198 4040 15254 4049
rect 15198 3975 15254 3984
rect 14844 1006 15056 1034
rect 14844 898 14872 1006
rect 14752 870 14872 898
rect 14752 800 14780 870
rect 15212 800 15240 3975
rect 15580 3505 15608 5510
rect 15672 5370 15700 5578
rect 15856 5370 15884 5630
rect 15956 5468 16252 5488
rect 16012 5466 16036 5468
rect 16092 5466 16116 5468
rect 16172 5466 16196 5468
rect 16034 5414 16036 5466
rect 16098 5414 16110 5466
rect 16172 5414 16174 5466
rect 16012 5412 16036 5414
rect 16092 5412 16116 5414
rect 16172 5412 16196 5414
rect 15956 5392 16252 5412
rect 15660 5364 15712 5370
rect 15660 5306 15712 5312
rect 15844 5364 15896 5370
rect 15844 5306 15896 5312
rect 16316 4826 16344 5714
rect 16304 4820 16356 4826
rect 16304 4762 16356 4768
rect 15956 4380 16252 4400
rect 16012 4378 16036 4380
rect 16092 4378 16116 4380
rect 16172 4378 16196 4380
rect 16034 4326 16036 4378
rect 16098 4326 16110 4378
rect 16172 4326 16174 4378
rect 16012 4324 16036 4326
rect 16092 4324 16116 4326
rect 16172 4324 16196 4326
rect 15956 4304 16252 4324
rect 16302 4040 16358 4049
rect 16302 3975 16358 3984
rect 15566 3496 15622 3505
rect 15566 3431 15622 3440
rect 15956 3292 16252 3312
rect 16012 3290 16036 3292
rect 16092 3290 16116 3292
rect 16172 3290 16196 3292
rect 16034 3238 16036 3290
rect 16098 3238 16110 3290
rect 16172 3238 16174 3290
rect 16012 3236 16036 3238
rect 16092 3236 16116 3238
rect 16172 3236 16196 3238
rect 15956 3216 16252 3236
rect 15956 2204 16252 2224
rect 16012 2202 16036 2204
rect 16092 2202 16116 2204
rect 16172 2202 16196 2204
rect 16034 2150 16036 2202
rect 16098 2150 16110 2202
rect 16172 2150 16174 2202
rect 16012 2148 16036 2150
rect 16092 2148 16116 2150
rect 16172 2148 16196 2150
rect 15956 2128 16252 2148
rect 16316 1986 16344 3975
rect 16132 1958 16344 1986
rect 16132 800 16160 1958
rect 17052 800 17080 8327
rect 17696 2009 17724 15846
rect 17788 14822 17816 19110
rect 17776 14816 17828 14822
rect 17776 14758 17828 14764
rect 17776 14340 17828 14346
rect 17776 14282 17828 14288
rect 17788 7313 17816 14282
rect 17880 12209 17908 61118
rect 17960 61124 18012 61130
rect 17960 61066 18012 61072
rect 18604 61056 18656 61062
rect 18604 60998 18656 61004
rect 18616 60654 18644 60998
rect 18236 60648 18288 60654
rect 18236 60590 18288 60596
rect 18604 60648 18656 60654
rect 18800 60602 18828 61542
rect 19076 60858 19104 68847
rect 19248 62144 19300 62150
rect 19248 62086 19300 62092
rect 19260 61826 19288 62086
rect 19260 61798 19472 61826
rect 19444 61742 19472 61798
rect 19248 61736 19300 61742
rect 19248 61678 19300 61684
rect 19432 61736 19484 61742
rect 19432 61678 19484 61684
rect 19156 61260 19208 61266
rect 19156 61202 19208 61208
rect 19064 60852 19116 60858
rect 19064 60794 19116 60800
rect 19168 60790 19196 61202
rect 19260 61130 19288 61678
rect 19248 61124 19300 61130
rect 19248 61066 19300 61072
rect 19616 61056 19668 61062
rect 19616 60998 19668 61004
rect 19248 60852 19300 60858
rect 19248 60794 19300 60800
rect 18880 60784 18932 60790
rect 18878 60752 18880 60761
rect 19156 60784 19208 60790
rect 18932 60752 18934 60761
rect 19156 60726 19208 60732
rect 18878 60687 18934 60696
rect 18604 60590 18656 60596
rect 18248 60110 18276 60590
rect 18708 60574 18828 60602
rect 18880 60648 18932 60654
rect 18880 60590 18932 60596
rect 18236 60104 18288 60110
rect 18236 60046 18288 60052
rect 18234 59528 18290 59537
rect 18234 59463 18290 59472
rect 17960 59016 18012 59022
rect 17960 58958 18012 58964
rect 18144 59016 18196 59022
rect 18144 58958 18196 58964
rect 17972 58585 18000 58958
rect 17958 58576 18014 58585
rect 17958 58511 18014 58520
rect 18156 58002 18184 58958
rect 18144 57996 18196 58002
rect 18144 57938 18196 57944
rect 18052 57316 18104 57322
rect 18052 57258 18104 57264
rect 18064 56778 18092 57258
rect 17960 56772 18012 56778
rect 17960 56714 18012 56720
rect 18052 56772 18104 56778
rect 18052 56714 18104 56720
rect 17972 56506 18000 56714
rect 17960 56500 18012 56506
rect 17960 56442 18012 56448
rect 18064 56234 18092 56714
rect 18052 56228 18104 56234
rect 18052 56170 18104 56176
rect 17958 55584 18014 55593
rect 17958 55519 18014 55528
rect 17972 55418 18000 55519
rect 17960 55412 18012 55418
rect 17960 55354 18012 55360
rect 18064 55214 18092 56170
rect 18052 55208 18104 55214
rect 18052 55150 18104 55156
rect 18052 55072 18104 55078
rect 18052 55014 18104 55020
rect 17960 54664 18012 54670
rect 17960 54606 18012 54612
rect 17972 54194 18000 54606
rect 17960 54188 18012 54194
rect 17960 54130 18012 54136
rect 18064 54074 18092 55014
rect 17972 54046 18092 54074
rect 17972 51610 18000 54046
rect 18156 53786 18184 57938
rect 18248 56250 18276 59463
rect 18708 58290 18736 60574
rect 18892 60314 18920 60590
rect 18880 60308 18932 60314
rect 18880 60250 18932 60256
rect 18788 60104 18840 60110
rect 18788 60046 18840 60052
rect 18800 59566 18828 60046
rect 18892 59634 18920 60250
rect 19064 59764 19116 59770
rect 19064 59706 19116 59712
rect 18880 59628 18932 59634
rect 18880 59570 18932 59576
rect 18788 59560 18840 59566
rect 18788 59502 18840 59508
rect 18800 58886 18828 59502
rect 18788 58880 18840 58886
rect 18788 58822 18840 58828
rect 18800 58426 18828 58822
rect 18892 58546 18920 59570
rect 19076 59566 19104 59706
rect 19064 59560 19116 59566
rect 19064 59502 19116 59508
rect 18972 59016 19024 59022
rect 18972 58958 19024 58964
rect 18984 58857 19012 58958
rect 18970 58848 19026 58857
rect 18970 58783 19026 58792
rect 19076 58682 19104 59502
rect 19154 59256 19210 59265
rect 19154 59191 19210 59200
rect 19168 58954 19196 59191
rect 19156 58948 19208 58954
rect 19156 58890 19208 58896
rect 19064 58676 19116 58682
rect 19064 58618 19116 58624
rect 18880 58540 18932 58546
rect 18880 58482 18932 58488
rect 18972 58540 19024 58546
rect 18972 58482 19024 58488
rect 18800 58398 18920 58426
rect 18708 58262 18828 58290
rect 18512 57928 18564 57934
rect 18512 57870 18564 57876
rect 18328 57792 18380 57798
rect 18524 57769 18552 57870
rect 18604 57792 18656 57798
rect 18328 57734 18380 57740
rect 18510 57760 18566 57769
rect 18340 57526 18368 57734
rect 18604 57734 18656 57740
rect 18694 57760 18750 57769
rect 18510 57695 18566 57704
rect 18328 57520 18380 57526
rect 18328 57462 18380 57468
rect 18340 56438 18368 57462
rect 18524 56914 18552 57695
rect 18616 57458 18644 57734
rect 18694 57695 18750 57704
rect 18708 57594 18736 57695
rect 18696 57588 18748 57594
rect 18696 57530 18748 57536
rect 18604 57452 18656 57458
rect 18604 57394 18656 57400
rect 18512 56908 18564 56914
rect 18512 56850 18564 56856
rect 18328 56432 18380 56438
rect 18328 56374 18380 56380
rect 18248 56222 18368 56250
rect 18236 54664 18288 54670
rect 18236 54606 18288 54612
rect 18248 54058 18276 54606
rect 18236 54052 18288 54058
rect 18236 53994 18288 54000
rect 18144 53780 18196 53786
rect 18144 53722 18196 53728
rect 18052 53644 18104 53650
rect 18052 53586 18104 53592
rect 18236 53644 18288 53650
rect 18236 53586 18288 53592
rect 18064 52737 18092 53586
rect 18144 53576 18196 53582
rect 18248 53553 18276 53586
rect 18144 53518 18196 53524
rect 18234 53544 18290 53553
rect 18050 52728 18106 52737
rect 18050 52663 18106 52672
rect 18064 52630 18092 52663
rect 18052 52624 18104 52630
rect 18052 52566 18104 52572
rect 18052 51876 18104 51882
rect 18052 51818 18104 51824
rect 17960 51604 18012 51610
rect 17960 51546 18012 51552
rect 18064 51474 18092 51818
rect 18052 51468 18104 51474
rect 18052 51410 18104 51416
rect 18156 51406 18184 53518
rect 18234 53479 18290 53488
rect 18236 52896 18288 52902
rect 18236 52838 18288 52844
rect 18248 52358 18276 52838
rect 18236 52352 18288 52358
rect 18236 52294 18288 52300
rect 18144 51400 18196 51406
rect 18144 51342 18196 51348
rect 17958 50416 18014 50425
rect 17958 50351 17960 50360
rect 18012 50351 18014 50360
rect 17960 50322 18012 50328
rect 17972 49978 18000 50322
rect 18144 50176 18196 50182
rect 18144 50118 18196 50124
rect 17960 49972 18012 49978
rect 17960 49914 18012 49920
rect 18156 49842 18184 50118
rect 18144 49836 18196 49842
rect 18144 49778 18196 49784
rect 18156 49434 18184 49778
rect 18144 49428 18196 49434
rect 18144 49370 18196 49376
rect 17960 49292 18012 49298
rect 17960 49234 18012 49240
rect 17972 47258 18000 49234
rect 18144 49224 18196 49230
rect 18144 49166 18196 49172
rect 18052 48680 18104 48686
rect 18050 48648 18052 48657
rect 18104 48648 18106 48657
rect 18050 48583 18106 48592
rect 18052 48204 18104 48210
rect 18052 48146 18104 48152
rect 18064 48113 18092 48146
rect 18050 48104 18106 48113
rect 18050 48039 18106 48048
rect 18156 47705 18184 49166
rect 18236 48680 18288 48686
rect 18236 48622 18288 48628
rect 18248 48210 18276 48622
rect 18340 48550 18368 56222
rect 18420 56228 18472 56234
rect 18420 56170 18472 56176
rect 18432 53106 18460 56170
rect 18524 54482 18552 56850
rect 18800 56386 18828 58262
rect 18616 56358 18828 56386
rect 18616 54641 18644 56358
rect 18786 56264 18842 56273
rect 18786 56199 18842 56208
rect 18800 55894 18828 56199
rect 18788 55888 18840 55894
rect 18788 55830 18840 55836
rect 18694 55312 18750 55321
rect 18694 55247 18750 55256
rect 18602 54632 18658 54641
rect 18602 54567 18658 54576
rect 18524 54454 18644 54482
rect 18512 54324 18564 54330
rect 18512 54266 18564 54272
rect 18420 53100 18472 53106
rect 18420 53042 18472 53048
rect 18432 52698 18460 53042
rect 18524 53009 18552 54266
rect 18510 53000 18566 53009
rect 18510 52935 18566 52944
rect 18420 52692 18472 52698
rect 18420 52634 18472 52640
rect 18432 52086 18460 52634
rect 18524 52154 18552 52935
rect 18616 52154 18644 54454
rect 18708 53786 18736 55247
rect 18788 55140 18840 55146
rect 18788 55082 18840 55088
rect 18800 54738 18828 55082
rect 18788 54732 18840 54738
rect 18788 54674 18840 54680
rect 18788 54188 18840 54194
rect 18788 54130 18840 54136
rect 18800 53990 18828 54130
rect 18788 53984 18840 53990
rect 18788 53926 18840 53932
rect 18800 53825 18828 53926
rect 18786 53816 18842 53825
rect 18696 53780 18748 53786
rect 18786 53751 18842 53760
rect 18696 53722 18748 53728
rect 18694 53680 18750 53689
rect 18694 53615 18696 53624
rect 18748 53615 18750 53624
rect 18696 53586 18748 53592
rect 18708 52544 18736 53586
rect 18800 53174 18828 53751
rect 18788 53168 18840 53174
rect 18788 53110 18840 53116
rect 18892 52902 18920 58398
rect 18880 52896 18932 52902
rect 18880 52838 18932 52844
rect 18788 52556 18840 52562
rect 18708 52516 18788 52544
rect 18512 52148 18564 52154
rect 18512 52090 18564 52096
rect 18604 52148 18656 52154
rect 18604 52090 18656 52096
rect 18420 52080 18472 52086
rect 18420 52022 18472 52028
rect 18432 50402 18460 52022
rect 18524 51950 18552 52090
rect 18512 51944 18564 51950
rect 18512 51886 18564 51892
rect 18604 51944 18656 51950
rect 18604 51886 18656 51892
rect 18512 51808 18564 51814
rect 18512 51750 18564 51756
rect 18524 50862 18552 51750
rect 18616 51474 18644 51886
rect 18604 51468 18656 51474
rect 18604 51410 18656 51416
rect 18616 51066 18644 51410
rect 18604 51060 18656 51066
rect 18604 51002 18656 51008
rect 18512 50856 18564 50862
rect 18512 50798 18564 50804
rect 18524 50522 18552 50798
rect 18512 50516 18564 50522
rect 18512 50458 18564 50464
rect 18432 50374 18552 50402
rect 18420 50312 18472 50318
rect 18420 50254 18472 50260
rect 18432 49978 18460 50254
rect 18420 49972 18472 49978
rect 18420 49914 18472 49920
rect 18524 49434 18552 50374
rect 18708 50153 18736 52516
rect 18788 52498 18840 52504
rect 18788 52148 18840 52154
rect 18788 52090 18840 52096
rect 18694 50144 18750 50153
rect 18616 50102 18694 50130
rect 18512 49428 18564 49434
rect 18512 49370 18564 49376
rect 18420 49224 18472 49230
rect 18420 49166 18472 49172
rect 18432 48890 18460 49166
rect 18420 48884 18472 48890
rect 18420 48826 18472 48832
rect 18616 48686 18644 50102
rect 18694 50079 18750 50088
rect 18800 49960 18828 52090
rect 18892 51490 18920 52838
rect 18984 52086 19012 58482
rect 19064 57248 19116 57254
rect 19064 57190 19116 57196
rect 19076 56778 19104 57190
rect 19064 56772 19116 56778
rect 19064 56714 19116 56720
rect 19062 56536 19118 56545
rect 19062 56471 19118 56480
rect 19076 56438 19104 56471
rect 19064 56432 19116 56438
rect 19064 56374 19116 56380
rect 19064 55752 19116 55758
rect 19064 55694 19116 55700
rect 19076 53666 19104 55694
rect 19168 55078 19196 58890
rect 19156 55072 19208 55078
rect 19156 55014 19208 55020
rect 19156 54664 19208 54670
rect 19156 54606 19208 54612
rect 19168 53786 19196 54606
rect 19156 53780 19208 53786
rect 19156 53722 19208 53728
rect 19076 53638 19196 53666
rect 19064 53100 19116 53106
rect 19064 53042 19116 53048
rect 18972 52080 19024 52086
rect 18972 52022 19024 52028
rect 18984 51814 19012 52022
rect 18972 51808 19024 51814
rect 18972 51750 19024 51756
rect 19076 51610 19104 53042
rect 19168 52698 19196 53638
rect 19156 52692 19208 52698
rect 19156 52634 19208 52640
rect 19156 52012 19208 52018
rect 19156 51954 19208 51960
rect 19064 51604 19116 51610
rect 19064 51546 19116 51552
rect 18892 51462 19104 51490
rect 18972 51400 19024 51406
rect 18972 51342 19024 51348
rect 18878 50688 18934 50697
rect 18878 50623 18934 50632
rect 18708 49932 18828 49960
rect 18708 49774 18736 49932
rect 18892 49910 18920 50623
rect 18880 49904 18932 49910
rect 18880 49846 18932 49852
rect 18696 49768 18748 49774
rect 18694 49736 18696 49745
rect 18748 49736 18750 49745
rect 18694 49671 18750 49680
rect 18604 48680 18656 48686
rect 18604 48622 18656 48628
rect 18328 48544 18380 48550
rect 18328 48486 18380 48492
rect 18892 48278 18920 49846
rect 18984 49774 19012 51342
rect 19076 51252 19104 51462
rect 19168 51377 19196 51954
rect 19154 51368 19210 51377
rect 19154 51303 19210 51312
rect 19156 51264 19208 51270
rect 19076 51224 19156 51252
rect 19156 51206 19208 51212
rect 19064 50924 19116 50930
rect 19064 50866 19116 50872
rect 19076 50726 19104 50866
rect 19064 50720 19116 50726
rect 19064 50662 19116 50668
rect 18972 49768 19024 49774
rect 18972 49710 19024 49716
rect 18984 49298 19012 49710
rect 18972 49292 19024 49298
rect 18972 49234 19024 49240
rect 19076 49094 19104 50662
rect 19168 50318 19196 51206
rect 19156 50312 19208 50318
rect 19156 50254 19208 50260
rect 19064 49088 19116 49094
rect 19064 49030 19116 49036
rect 19064 48680 19116 48686
rect 19064 48622 19116 48628
rect 18970 48376 19026 48385
rect 19076 48346 19104 48622
rect 19156 48612 19208 48618
rect 19156 48554 19208 48560
rect 18970 48311 19026 48320
rect 19064 48340 19116 48346
rect 18984 48278 19012 48311
rect 19064 48282 19116 48288
rect 18880 48272 18932 48278
rect 18880 48214 18932 48220
rect 18972 48272 19024 48278
rect 19076 48249 19104 48282
rect 18972 48214 19024 48220
rect 19062 48240 19118 48249
rect 18236 48204 18288 48210
rect 18236 48146 18288 48152
rect 18142 47696 18198 47705
rect 18052 47660 18104 47666
rect 18142 47631 18198 47640
rect 18052 47602 18104 47608
rect 17960 47252 18012 47258
rect 17960 47194 18012 47200
rect 17960 47116 18012 47122
rect 17960 47058 18012 47064
rect 17972 46578 18000 47058
rect 18064 46714 18092 47602
rect 18248 47433 18276 48146
rect 18892 48074 18920 48214
rect 19062 48175 19118 48184
rect 18880 48068 18932 48074
rect 18880 48010 18932 48016
rect 18892 47682 18920 48010
rect 18800 47654 18920 47682
rect 18800 47598 18828 47654
rect 18788 47592 18840 47598
rect 18788 47534 18840 47540
rect 18972 47592 19024 47598
rect 18972 47534 19024 47540
rect 18234 47424 18290 47433
rect 18234 47359 18290 47368
rect 18248 46986 18276 47359
rect 18328 47184 18380 47190
rect 18328 47126 18380 47132
rect 18236 46980 18288 46986
rect 18236 46922 18288 46928
rect 18052 46708 18104 46714
rect 18052 46650 18104 46656
rect 17960 46572 18012 46578
rect 17960 46514 18012 46520
rect 18340 46510 18368 47126
rect 18328 46504 18380 46510
rect 18328 46446 18380 46452
rect 18800 46442 18828 47534
rect 18984 47122 19012 47534
rect 18972 47116 19024 47122
rect 18972 47058 19024 47064
rect 18788 46436 18840 46442
rect 18788 46378 18840 46384
rect 18142 46336 18198 46345
rect 18142 46271 18198 46280
rect 18156 45082 18184 46271
rect 18800 46170 18828 46378
rect 18788 46164 18840 46170
rect 18788 46106 18840 46112
rect 18878 45928 18934 45937
rect 18878 45863 18934 45872
rect 18328 45824 18380 45830
rect 18328 45766 18380 45772
rect 18340 45422 18368 45766
rect 18892 45626 18920 45863
rect 18696 45620 18748 45626
rect 18696 45562 18748 45568
rect 18880 45620 18932 45626
rect 18880 45562 18932 45568
rect 18328 45416 18380 45422
rect 18328 45358 18380 45364
rect 18144 45076 18196 45082
rect 18144 45018 18196 45024
rect 18052 44940 18104 44946
rect 18052 44882 18104 44888
rect 17960 44464 18012 44470
rect 17960 44406 18012 44412
rect 17972 43994 18000 44406
rect 17960 43988 18012 43994
rect 17960 43930 18012 43936
rect 18064 43926 18092 44882
rect 18340 44878 18368 45358
rect 18604 44940 18656 44946
rect 18604 44882 18656 44888
rect 18328 44872 18380 44878
rect 18328 44814 18380 44820
rect 18340 44402 18368 44814
rect 18328 44396 18380 44402
rect 18328 44338 18380 44344
rect 18512 44328 18564 44334
rect 18510 44296 18512 44305
rect 18564 44296 18566 44305
rect 18510 44231 18566 44240
rect 18052 43920 18104 43926
rect 18052 43862 18104 43868
rect 18420 43784 18472 43790
rect 18420 43726 18472 43732
rect 18050 43480 18106 43489
rect 18050 43415 18106 43424
rect 18064 43314 18092 43415
rect 18052 43308 18104 43314
rect 18052 43250 18104 43256
rect 18328 42696 18380 42702
rect 18328 42638 18380 42644
rect 18340 42362 18368 42638
rect 18328 42356 18380 42362
rect 18328 42298 18380 42304
rect 18432 42158 18460 43726
rect 18616 43654 18644 44882
rect 18708 43926 18736 45562
rect 18984 45490 19012 47058
rect 19076 46578 19104 48175
rect 19168 48142 19196 48554
rect 19156 48136 19208 48142
rect 19156 48078 19208 48084
rect 19156 48000 19208 48006
rect 19156 47942 19208 47948
rect 19168 47598 19196 47942
rect 19156 47592 19208 47598
rect 19156 47534 19208 47540
rect 19168 47122 19196 47534
rect 19156 47116 19208 47122
rect 19156 47058 19208 47064
rect 19064 46572 19116 46578
rect 19064 46514 19116 46520
rect 19156 46368 19208 46374
rect 19156 46310 19208 46316
rect 19064 46028 19116 46034
rect 19064 45970 19116 45976
rect 18972 45484 19024 45490
rect 18972 45426 19024 45432
rect 19076 45354 19104 45970
rect 19168 45966 19196 46310
rect 19156 45960 19208 45966
rect 19156 45902 19208 45908
rect 19064 45348 19116 45354
rect 19064 45290 19116 45296
rect 19076 45014 19104 45290
rect 19064 45008 19116 45014
rect 19064 44950 19116 44956
rect 19156 44736 19208 44742
rect 19156 44678 19208 44684
rect 18878 44432 18934 44441
rect 18878 44367 18934 44376
rect 18696 43920 18748 43926
rect 18696 43862 18748 43868
rect 18604 43648 18656 43654
rect 18604 43590 18656 43596
rect 18420 42152 18472 42158
rect 18420 42094 18472 42100
rect 18142 40896 18198 40905
rect 18142 40831 18198 40840
rect 18156 40390 18184 40831
rect 18144 40384 18196 40390
rect 18144 40326 18196 40332
rect 18052 39432 18104 39438
rect 18052 39374 18104 39380
rect 18064 38894 18092 39374
rect 18052 38888 18104 38894
rect 18052 38830 18104 38836
rect 18064 38486 18092 38830
rect 18052 38480 18104 38486
rect 18052 38422 18104 38428
rect 18156 37330 18184 40326
rect 18328 39432 18380 39438
rect 18328 39374 18380 39380
rect 18340 39098 18368 39374
rect 18328 39092 18380 39098
rect 18328 39034 18380 39040
rect 18340 38554 18368 39034
rect 18420 38888 18472 38894
rect 18420 38830 18472 38836
rect 18328 38548 18380 38554
rect 18328 38490 18380 38496
rect 18432 38434 18460 38830
rect 18340 38406 18460 38434
rect 18144 37324 18196 37330
rect 18144 37266 18196 37272
rect 18052 36712 18104 36718
rect 18052 36654 18104 36660
rect 17958 36272 18014 36281
rect 17958 36207 18014 36216
rect 17972 36038 18000 36207
rect 17960 36032 18012 36038
rect 17960 35974 18012 35980
rect 17972 35494 18000 35974
rect 17960 35488 18012 35494
rect 17960 35430 18012 35436
rect 18064 35290 18092 36654
rect 18236 36168 18288 36174
rect 18236 36110 18288 36116
rect 18142 35864 18198 35873
rect 18142 35799 18144 35808
rect 18196 35799 18198 35808
rect 18144 35770 18196 35776
rect 18248 35766 18276 36110
rect 18236 35760 18288 35766
rect 18234 35728 18236 35737
rect 18288 35728 18290 35737
rect 18234 35663 18290 35672
rect 18248 35637 18276 35663
rect 18144 35624 18196 35630
rect 18144 35566 18196 35572
rect 18156 35290 18184 35566
rect 18236 35488 18288 35494
rect 18236 35430 18288 35436
rect 18052 35284 18104 35290
rect 18052 35226 18104 35232
rect 18144 35284 18196 35290
rect 18144 35226 18196 35232
rect 17958 34776 18014 34785
rect 17958 34711 18014 34720
rect 17972 34474 18000 34711
rect 18064 34610 18092 35226
rect 18248 35170 18276 35430
rect 18156 35142 18276 35170
rect 18052 34604 18104 34610
rect 18052 34546 18104 34552
rect 17960 34468 18012 34474
rect 17960 34410 18012 34416
rect 17972 34134 18000 34410
rect 18064 34202 18092 34546
rect 18052 34196 18104 34202
rect 18052 34138 18104 34144
rect 17960 34128 18012 34134
rect 17960 34070 18012 34076
rect 18052 33312 18104 33318
rect 18052 33254 18104 33260
rect 17960 32768 18012 32774
rect 17960 32710 18012 32716
rect 17972 32298 18000 32710
rect 17960 32292 18012 32298
rect 17960 32234 18012 32240
rect 17972 31958 18000 32234
rect 17960 31952 18012 31958
rect 17960 31894 18012 31900
rect 17960 31680 18012 31686
rect 17960 31622 18012 31628
rect 17972 31346 18000 31622
rect 17960 31340 18012 31346
rect 17960 31282 18012 31288
rect 17972 30938 18000 31282
rect 17960 30932 18012 30938
rect 17960 30874 18012 30880
rect 17960 30592 18012 30598
rect 17960 30534 18012 30540
rect 17972 30190 18000 30534
rect 17960 30184 18012 30190
rect 17960 30126 18012 30132
rect 17960 30048 18012 30054
rect 17960 29990 18012 29996
rect 17972 28626 18000 29990
rect 18064 29850 18092 33254
rect 18156 32298 18184 35142
rect 18236 33992 18288 33998
rect 18236 33934 18288 33940
rect 18248 32978 18276 33934
rect 18236 32972 18288 32978
rect 18236 32914 18288 32920
rect 18144 32292 18196 32298
rect 18144 32234 18196 32240
rect 18236 32224 18288 32230
rect 18236 32166 18288 32172
rect 18144 30728 18196 30734
rect 18144 30670 18196 30676
rect 18156 30569 18184 30670
rect 18142 30560 18198 30569
rect 18142 30495 18198 30504
rect 18144 30388 18196 30394
rect 18144 30330 18196 30336
rect 18052 29844 18104 29850
rect 18052 29786 18104 29792
rect 18050 29744 18106 29753
rect 18050 29679 18106 29688
rect 18064 29306 18092 29679
rect 18052 29300 18104 29306
rect 18052 29242 18104 29248
rect 17960 28620 18012 28626
rect 17960 28562 18012 28568
rect 18052 28416 18104 28422
rect 18052 28358 18104 28364
rect 17960 28008 18012 28014
rect 18064 27985 18092 28358
rect 17960 27950 18012 27956
rect 18050 27976 18106 27985
rect 17972 26518 18000 27950
rect 18050 27911 18106 27920
rect 18052 27464 18104 27470
rect 18052 27406 18104 27412
rect 18064 26926 18092 27406
rect 18156 27169 18184 30330
rect 18248 28150 18276 32166
rect 18236 28144 18288 28150
rect 18236 28086 18288 28092
rect 18142 27160 18198 27169
rect 18142 27095 18198 27104
rect 18234 27024 18290 27033
rect 18234 26959 18290 26968
rect 18052 26920 18104 26926
rect 18052 26862 18104 26868
rect 18142 26616 18198 26625
rect 18142 26551 18198 26560
rect 18156 26518 18184 26551
rect 18248 26518 18276 26959
rect 17960 26512 18012 26518
rect 17960 26454 18012 26460
rect 18144 26512 18196 26518
rect 18144 26454 18196 26460
rect 18236 26512 18288 26518
rect 18236 26454 18288 26460
rect 18236 25696 18288 25702
rect 18236 25638 18288 25644
rect 18144 24948 18196 24954
rect 18144 24890 18196 24896
rect 18052 24744 18104 24750
rect 18052 24686 18104 24692
rect 18064 24177 18092 24686
rect 18050 24168 18106 24177
rect 17960 24132 18012 24138
rect 18050 24103 18106 24112
rect 17960 24074 18012 24080
rect 17972 17882 18000 24074
rect 18156 23322 18184 24890
rect 18248 24614 18276 25638
rect 18236 24608 18288 24614
rect 18236 24550 18288 24556
rect 18248 23662 18276 24550
rect 18236 23656 18288 23662
rect 18236 23598 18288 23604
rect 18144 23316 18196 23322
rect 18144 23258 18196 23264
rect 18156 22574 18184 23258
rect 18144 22568 18196 22574
rect 18144 22510 18196 22516
rect 18144 21888 18196 21894
rect 18144 21830 18196 21836
rect 18050 21720 18106 21729
rect 18050 21655 18106 21664
rect 18064 21554 18092 21655
rect 18052 21548 18104 21554
rect 18052 21490 18104 21496
rect 18156 21486 18184 21830
rect 18144 21480 18196 21486
rect 18050 21448 18106 21457
rect 18144 21422 18196 21428
rect 18050 21383 18106 21392
rect 17960 17876 18012 17882
rect 17960 17818 18012 17824
rect 18064 17762 18092 21383
rect 18236 20392 18288 20398
rect 18236 20334 18288 20340
rect 18144 19712 18196 19718
rect 18144 19654 18196 19660
rect 18156 19310 18184 19654
rect 18248 19514 18276 20334
rect 18236 19508 18288 19514
rect 18236 19450 18288 19456
rect 18144 19304 18196 19310
rect 18144 19246 18196 19252
rect 18156 18970 18184 19246
rect 18144 18964 18196 18970
rect 18144 18906 18196 18912
rect 17972 17734 18092 17762
rect 17866 12200 17922 12209
rect 17866 12135 17922 12144
rect 17972 11218 18000 17734
rect 18052 16992 18104 16998
rect 18052 16934 18104 16940
rect 18064 16046 18092 16934
rect 18052 16040 18104 16046
rect 18052 15982 18104 15988
rect 18064 15502 18092 15982
rect 18052 15496 18104 15502
rect 18052 15438 18104 15444
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 17960 11212 18012 11218
rect 17960 11154 18012 11160
rect 17972 11098 18000 11154
rect 17880 11070 18000 11098
rect 17880 10810 17908 11070
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 17960 10260 18012 10266
rect 17960 10202 18012 10208
rect 17972 7562 18000 10202
rect 18064 10130 18092 11290
rect 18052 10124 18104 10130
rect 18052 10066 18104 10072
rect 18142 8256 18198 8265
rect 18142 8191 18198 8200
rect 18156 8090 18184 8191
rect 18144 8084 18196 8090
rect 18144 8026 18196 8032
rect 17880 7546 18000 7562
rect 17868 7540 18000 7546
rect 17920 7534 18000 7540
rect 17868 7482 17920 7488
rect 17774 7304 17830 7313
rect 17774 7239 17830 7248
rect 17972 3602 18000 7534
rect 18340 5545 18368 38406
rect 18510 38040 18566 38049
rect 18510 37975 18512 37984
rect 18564 37975 18566 37984
rect 18512 37946 18564 37952
rect 18512 37868 18564 37874
rect 18512 37810 18564 37816
rect 18420 37324 18472 37330
rect 18420 37266 18472 37272
rect 18432 36922 18460 37266
rect 18420 36916 18472 36922
rect 18420 36858 18472 36864
rect 18432 35698 18460 36858
rect 18420 35692 18472 35698
rect 18420 35634 18472 35640
rect 18432 35222 18460 35634
rect 18420 35216 18472 35222
rect 18420 35158 18472 35164
rect 18432 34746 18460 35158
rect 18420 34740 18472 34746
rect 18420 34682 18472 34688
rect 18524 34626 18552 37810
rect 18432 34598 18552 34626
rect 18432 29170 18460 34598
rect 18512 34400 18564 34406
rect 18512 34342 18564 34348
rect 18524 30394 18552 34342
rect 18616 33114 18644 43590
rect 18892 42294 18920 44367
rect 19168 43994 19196 44678
rect 19156 43988 19208 43994
rect 19156 43930 19208 43936
rect 19168 43382 19196 43930
rect 19156 43376 19208 43382
rect 19156 43318 19208 43324
rect 18972 43240 19024 43246
rect 18972 43182 19024 43188
rect 18984 42566 19012 43182
rect 19062 42800 19118 42809
rect 19062 42735 19118 42744
rect 19156 42764 19208 42770
rect 18972 42560 19024 42566
rect 18972 42502 19024 42508
rect 18880 42288 18932 42294
rect 18880 42230 18932 42236
rect 18984 41818 19012 42502
rect 18972 41812 19024 41818
rect 18972 41754 19024 41760
rect 18970 41032 19026 41041
rect 18970 40967 19026 40976
rect 18694 39264 18750 39273
rect 18694 39199 18750 39208
rect 18604 33108 18656 33114
rect 18604 33050 18656 33056
rect 18708 32586 18736 39199
rect 18880 37664 18932 37670
rect 18880 37606 18932 37612
rect 18788 37120 18840 37126
rect 18788 37062 18840 37068
rect 18800 34377 18828 37062
rect 18892 34542 18920 37606
rect 18880 34536 18932 34542
rect 18880 34478 18932 34484
rect 18786 34368 18842 34377
rect 18786 34303 18842 34312
rect 18800 33833 18828 34303
rect 18786 33824 18842 33833
rect 18786 33759 18842 33768
rect 18892 33697 18920 34478
rect 18878 33688 18934 33697
rect 18878 33623 18934 33632
rect 18892 33454 18920 33623
rect 18880 33448 18932 33454
rect 18880 33390 18932 33396
rect 18788 33380 18840 33386
rect 18788 33322 18840 33328
rect 18616 32558 18736 32586
rect 18616 32230 18644 32558
rect 18696 32496 18748 32502
rect 18696 32438 18748 32444
rect 18604 32224 18656 32230
rect 18604 32166 18656 32172
rect 18512 30388 18564 30394
rect 18512 30330 18564 30336
rect 18512 30252 18564 30258
rect 18512 30194 18564 30200
rect 18524 29306 18552 30194
rect 18604 30184 18656 30190
rect 18604 30126 18656 30132
rect 18512 29300 18564 29306
rect 18512 29242 18564 29248
rect 18420 29164 18472 29170
rect 18420 29106 18472 29112
rect 18432 27112 18460 29106
rect 18512 28620 18564 28626
rect 18512 28562 18564 28568
rect 18524 27674 18552 28562
rect 18512 27668 18564 27674
rect 18512 27610 18564 27616
rect 18432 27084 18552 27112
rect 18418 27024 18474 27033
rect 18418 26959 18420 26968
rect 18472 26959 18474 26968
rect 18420 26930 18472 26936
rect 18418 26072 18474 26081
rect 18418 26007 18420 26016
rect 18472 26007 18474 26016
rect 18420 25978 18472 25984
rect 18432 25809 18460 25978
rect 18418 25800 18474 25809
rect 18418 25735 18474 25744
rect 18524 23746 18552 27084
rect 18432 23718 18552 23746
rect 18432 22642 18460 23718
rect 18510 23624 18566 23633
rect 18510 23559 18566 23568
rect 18420 22636 18472 22642
rect 18420 22578 18472 22584
rect 18432 22234 18460 22578
rect 18420 22228 18472 22234
rect 18420 22170 18472 22176
rect 18420 22024 18472 22030
rect 18420 21966 18472 21972
rect 18432 11665 18460 21966
rect 18524 20534 18552 23559
rect 18616 22098 18644 30126
rect 18708 30025 18736 32438
rect 18800 31385 18828 33322
rect 18880 31884 18932 31890
rect 18880 31826 18932 31832
rect 18786 31376 18842 31385
rect 18786 31311 18842 31320
rect 18892 30122 18920 31826
rect 18984 31822 19012 40967
rect 19076 37126 19104 42735
rect 19156 42706 19208 42712
rect 19168 41546 19196 42706
rect 19156 41540 19208 41546
rect 19156 41482 19208 41488
rect 19064 37120 19116 37126
rect 19064 37062 19116 37068
rect 19076 36718 19104 37062
rect 19064 36712 19116 36718
rect 19064 36654 19116 36660
rect 19076 36242 19104 36654
rect 19064 36236 19116 36242
rect 19064 36178 19116 36184
rect 19076 34785 19104 36178
rect 19156 36032 19208 36038
rect 19156 35974 19208 35980
rect 19168 35737 19196 35974
rect 19154 35728 19210 35737
rect 19154 35663 19210 35672
rect 19168 35562 19196 35663
rect 19156 35556 19208 35562
rect 19156 35498 19208 35504
rect 19062 34776 19118 34785
rect 19062 34711 19118 34720
rect 19062 34640 19118 34649
rect 19062 34575 19064 34584
rect 19116 34575 19118 34584
rect 19064 34546 19116 34552
rect 19260 34066 19288 60794
rect 19340 60580 19392 60586
rect 19340 60522 19392 60528
rect 19352 59226 19380 60522
rect 19432 60308 19484 60314
rect 19432 60250 19484 60256
rect 19340 59220 19392 59226
rect 19340 59162 19392 59168
rect 19338 58032 19394 58041
rect 19338 57967 19340 57976
rect 19392 57967 19394 57976
rect 19340 57938 19392 57944
rect 19338 57080 19394 57089
rect 19338 57015 19394 57024
rect 19352 56914 19380 57015
rect 19340 56908 19392 56914
rect 19340 56850 19392 56856
rect 19352 56438 19380 56850
rect 19340 56432 19392 56438
rect 19340 56374 19392 56380
rect 19352 55894 19380 56374
rect 19340 55888 19392 55894
rect 19340 55830 19392 55836
rect 19352 54874 19380 55830
rect 19340 54868 19392 54874
rect 19340 54810 19392 54816
rect 19338 54632 19394 54641
rect 19338 54567 19394 54576
rect 19352 54330 19380 54567
rect 19340 54324 19392 54330
rect 19340 54266 19392 54272
rect 19340 54052 19392 54058
rect 19340 53994 19392 54000
rect 19352 52850 19380 53994
rect 19444 53650 19472 60250
rect 19524 60172 19576 60178
rect 19524 60114 19576 60120
rect 19536 58886 19564 60114
rect 19628 59242 19656 60998
rect 19720 60042 19748 72655
rect 20088 61810 20116 79070
rect 20272 74746 20300 79200
rect 21192 78010 21220 79200
rect 20732 77982 21220 78010
rect 20272 74718 20668 74746
rect 20352 74656 20404 74662
rect 20352 74598 20404 74604
rect 20364 62393 20392 74598
rect 20640 66314 20668 74718
rect 20732 69057 20760 77982
rect 20956 77820 21252 77840
rect 21012 77818 21036 77820
rect 21092 77818 21116 77820
rect 21172 77818 21196 77820
rect 21034 77766 21036 77818
rect 21098 77766 21110 77818
rect 21172 77766 21174 77818
rect 21012 77764 21036 77766
rect 21092 77764 21116 77766
rect 21172 77764 21196 77766
rect 20956 77744 21252 77764
rect 20956 76732 21252 76752
rect 21012 76730 21036 76732
rect 21092 76730 21116 76732
rect 21172 76730 21196 76732
rect 21034 76678 21036 76730
rect 21098 76678 21110 76730
rect 21172 76678 21174 76730
rect 21012 76676 21036 76678
rect 21092 76676 21116 76678
rect 21172 76676 21196 76678
rect 20956 76656 21252 76676
rect 20812 76492 20864 76498
rect 20812 76434 20864 76440
rect 20824 76090 20852 76434
rect 21364 76424 21416 76430
rect 21270 76392 21326 76401
rect 21364 76366 21416 76372
rect 21270 76327 21326 76336
rect 20812 76084 20864 76090
rect 20812 76026 20864 76032
rect 20824 75721 20852 76026
rect 20810 75712 20866 75721
rect 20810 75647 20866 75656
rect 20956 75644 21252 75664
rect 21012 75642 21036 75644
rect 21092 75642 21116 75644
rect 21172 75642 21196 75644
rect 21034 75590 21036 75642
rect 21098 75590 21110 75642
rect 21172 75590 21174 75642
rect 21012 75588 21036 75590
rect 21092 75588 21116 75590
rect 21172 75588 21196 75590
rect 20956 75568 21252 75588
rect 20810 75304 20866 75313
rect 20810 75239 20866 75248
rect 20824 73409 20852 75239
rect 20956 74556 21252 74576
rect 21012 74554 21036 74556
rect 21092 74554 21116 74556
rect 21172 74554 21196 74556
rect 21034 74502 21036 74554
rect 21098 74502 21110 74554
rect 21172 74502 21174 74554
rect 21012 74500 21036 74502
rect 21092 74500 21116 74502
rect 21172 74500 21196 74502
rect 20956 74480 21252 74500
rect 20956 73468 21252 73488
rect 21012 73466 21036 73468
rect 21092 73466 21116 73468
rect 21172 73466 21196 73468
rect 21034 73414 21036 73466
rect 21098 73414 21110 73466
rect 21172 73414 21174 73466
rect 21012 73412 21036 73414
rect 21092 73412 21116 73414
rect 21172 73412 21196 73414
rect 20810 73400 20866 73409
rect 20956 73392 21252 73412
rect 20810 73335 20866 73344
rect 20956 72380 21252 72400
rect 21012 72378 21036 72380
rect 21092 72378 21116 72380
rect 21172 72378 21196 72380
rect 21034 72326 21036 72378
rect 21098 72326 21110 72378
rect 21172 72326 21174 72378
rect 21012 72324 21036 72326
rect 21092 72324 21116 72326
rect 21172 72324 21196 72326
rect 20956 72304 21252 72324
rect 20812 72140 20864 72146
rect 20812 72082 20864 72088
rect 20824 71398 20852 72082
rect 20812 71392 20864 71398
rect 20812 71334 20864 71340
rect 20718 69048 20774 69057
rect 20718 68983 20774 68992
rect 20640 66286 20760 66314
rect 20536 66020 20588 66026
rect 20536 65962 20588 65968
rect 20444 63844 20496 63850
rect 20444 63786 20496 63792
rect 20350 62384 20406 62393
rect 20350 62319 20406 62328
rect 20166 62248 20222 62257
rect 20166 62183 20222 62192
rect 20076 61804 20128 61810
rect 20076 61746 20128 61752
rect 19800 61736 19852 61742
rect 19800 61678 19852 61684
rect 19812 60178 19840 61678
rect 19800 60172 19852 60178
rect 19800 60114 19852 60120
rect 19708 60036 19760 60042
rect 19708 59978 19760 59984
rect 19800 59492 19852 59498
rect 19800 59434 19852 59440
rect 19628 59214 19748 59242
rect 19616 59084 19668 59090
rect 19616 59026 19668 59032
rect 19628 58993 19656 59026
rect 19614 58984 19670 58993
rect 19614 58919 19670 58928
rect 19524 58880 19576 58886
rect 19720 58834 19748 59214
rect 19524 58822 19576 58828
rect 19536 58410 19564 58822
rect 19628 58806 19748 58834
rect 19628 58478 19656 58806
rect 19616 58472 19668 58478
rect 19616 58414 19668 58420
rect 19524 58404 19576 58410
rect 19524 58346 19576 58352
rect 19708 58404 19760 58410
rect 19708 58346 19760 58352
rect 19536 57594 19564 58346
rect 19720 58002 19748 58346
rect 19708 57996 19760 58002
rect 19708 57938 19760 57944
rect 19616 57860 19668 57866
rect 19616 57802 19668 57808
rect 19524 57588 19576 57594
rect 19524 57530 19576 57536
rect 19524 57384 19576 57390
rect 19524 57326 19576 57332
rect 19536 56778 19564 57326
rect 19524 56772 19576 56778
rect 19524 56714 19576 56720
rect 19628 56522 19656 57802
rect 19720 56914 19748 57938
rect 19708 56908 19760 56914
rect 19708 56850 19760 56856
rect 19708 56772 19760 56778
rect 19708 56714 19760 56720
rect 19536 56494 19656 56522
rect 19432 53644 19484 53650
rect 19432 53586 19484 53592
rect 19444 52970 19472 53586
rect 19432 52964 19484 52970
rect 19432 52906 19484 52912
rect 19352 52822 19472 52850
rect 19340 52488 19392 52494
rect 19340 52430 19392 52436
rect 19352 51950 19380 52430
rect 19444 52426 19472 52822
rect 19432 52420 19484 52426
rect 19432 52362 19484 52368
rect 19536 52057 19564 56494
rect 19616 56364 19668 56370
rect 19616 56306 19668 56312
rect 19628 54874 19656 56306
rect 19616 54868 19668 54874
rect 19616 54810 19668 54816
rect 19628 53718 19656 54810
rect 19720 54058 19748 56714
rect 19708 54052 19760 54058
rect 19708 53994 19760 54000
rect 19616 53712 19668 53718
rect 19616 53654 19668 53660
rect 19628 53106 19656 53654
rect 19708 53644 19760 53650
rect 19708 53586 19760 53592
rect 19616 53100 19668 53106
rect 19616 53042 19668 53048
rect 19720 52902 19748 53586
rect 19708 52896 19760 52902
rect 19708 52838 19760 52844
rect 19522 52048 19578 52057
rect 19522 51983 19578 51992
rect 19340 51944 19392 51950
rect 19392 51892 19656 51898
rect 19340 51886 19656 51892
rect 19352 51870 19656 51886
rect 19524 51604 19576 51610
rect 19524 51546 19576 51552
rect 19432 51536 19484 51542
rect 19432 51478 19484 51484
rect 19340 51468 19392 51474
rect 19340 51410 19392 51416
rect 19352 50930 19380 51410
rect 19444 50998 19472 51478
rect 19536 51066 19564 51546
rect 19524 51060 19576 51066
rect 19524 51002 19576 51008
rect 19432 50992 19484 50998
rect 19432 50934 19484 50940
rect 19340 50924 19392 50930
rect 19340 50866 19392 50872
rect 19340 50788 19392 50794
rect 19340 50730 19392 50736
rect 19352 50386 19380 50730
rect 19432 50720 19484 50726
rect 19432 50662 19484 50668
rect 19340 50380 19392 50386
rect 19340 50322 19392 50328
rect 19352 49842 19380 50322
rect 19340 49836 19392 49842
rect 19340 49778 19392 49784
rect 19444 49722 19472 50662
rect 19352 49694 19472 49722
rect 19524 49700 19576 49706
rect 19352 49230 19380 49694
rect 19524 49642 19576 49648
rect 19432 49292 19484 49298
rect 19432 49234 19484 49240
rect 19340 49224 19392 49230
rect 19340 49166 19392 49172
rect 19340 49088 19392 49094
rect 19340 49030 19392 49036
rect 19352 48793 19380 49030
rect 19444 48890 19472 49234
rect 19432 48884 19484 48890
rect 19432 48826 19484 48832
rect 19338 48784 19394 48793
rect 19338 48719 19394 48728
rect 19352 46442 19380 48719
rect 19430 48512 19486 48521
rect 19430 48447 19486 48456
rect 19444 47161 19472 48447
rect 19430 47152 19486 47161
rect 19430 47087 19486 47096
rect 19340 46436 19392 46442
rect 19340 46378 19392 46384
rect 19432 46028 19484 46034
rect 19432 45970 19484 45976
rect 19444 45914 19472 45970
rect 19352 45886 19472 45914
rect 19352 45286 19380 45886
rect 19432 45416 19484 45422
rect 19432 45358 19484 45364
rect 19340 45280 19392 45286
rect 19340 45222 19392 45228
rect 19352 44334 19380 45222
rect 19444 44946 19472 45358
rect 19432 44940 19484 44946
rect 19432 44882 19484 44888
rect 19340 44328 19392 44334
rect 19340 44270 19392 44276
rect 19352 43330 19380 44270
rect 19430 44024 19486 44033
rect 19430 43959 19486 43968
rect 19444 43450 19472 43959
rect 19432 43444 19484 43450
rect 19432 43386 19484 43392
rect 19352 43302 19472 43330
rect 19338 43208 19394 43217
rect 19444 43178 19472 43302
rect 19338 43143 19394 43152
rect 19432 43172 19484 43178
rect 19352 42090 19380 43143
rect 19432 43114 19484 43120
rect 19340 42084 19392 42090
rect 19340 42026 19392 42032
rect 19352 41818 19380 42026
rect 19340 41812 19392 41818
rect 19340 41754 19392 41760
rect 19352 35834 19380 41754
rect 19444 41682 19472 43114
rect 19432 41676 19484 41682
rect 19432 41618 19484 41624
rect 19430 39944 19486 39953
rect 19430 39879 19486 39888
rect 19444 39642 19472 39879
rect 19432 39636 19484 39642
rect 19432 39578 19484 39584
rect 19536 38865 19564 49642
rect 19628 47666 19656 51870
rect 19812 50538 19840 59434
rect 20076 58472 20128 58478
rect 20076 58414 20128 58420
rect 20088 57798 20116 58414
rect 20076 57792 20128 57798
rect 20076 57734 20128 57740
rect 20088 57390 20116 57734
rect 20076 57384 20128 57390
rect 20076 57326 20128 57332
rect 19984 56976 20036 56982
rect 19984 56918 20036 56924
rect 19996 55962 20024 56918
rect 20076 56840 20128 56846
rect 20076 56782 20128 56788
rect 19984 55956 20036 55962
rect 19984 55898 20036 55904
rect 19984 55072 20036 55078
rect 19984 55014 20036 55020
rect 19996 52698 20024 55014
rect 20088 53938 20116 56782
rect 20180 55842 20208 62183
rect 20258 58848 20314 58857
rect 20258 58783 20314 58792
rect 20272 57866 20300 58783
rect 20260 57860 20312 57866
rect 20260 57802 20312 57808
rect 20272 55962 20300 57802
rect 20456 57594 20484 63786
rect 20444 57588 20496 57594
rect 20444 57530 20496 57536
rect 20352 57384 20404 57390
rect 20352 57326 20404 57332
rect 20364 56302 20392 57326
rect 20444 56908 20496 56914
rect 20444 56850 20496 56856
rect 20352 56296 20404 56302
rect 20352 56238 20404 56244
rect 20456 55962 20484 56850
rect 20260 55956 20312 55962
rect 20260 55898 20312 55904
rect 20444 55956 20496 55962
rect 20444 55898 20496 55904
rect 20180 55814 20484 55842
rect 20352 55752 20404 55758
rect 20352 55694 20404 55700
rect 20168 55684 20220 55690
rect 20168 55626 20220 55632
rect 20180 54874 20208 55626
rect 20168 54868 20220 54874
rect 20168 54810 20220 54816
rect 20364 54534 20392 55694
rect 20352 54528 20404 54534
rect 20352 54470 20404 54476
rect 20088 53910 20300 53938
rect 20168 53644 20220 53650
rect 20168 53586 20220 53592
rect 20076 52896 20128 52902
rect 20076 52838 20128 52844
rect 19984 52692 20036 52698
rect 19984 52634 20036 52640
rect 19984 52420 20036 52426
rect 19984 52362 20036 52368
rect 19996 51270 20024 52362
rect 19984 51264 20036 51270
rect 19984 51206 20036 51212
rect 19996 50862 20024 51206
rect 19984 50856 20036 50862
rect 20088 50833 20116 52838
rect 20180 52698 20208 53586
rect 20168 52692 20220 52698
rect 20168 52634 20220 52640
rect 20180 52494 20208 52634
rect 20168 52488 20220 52494
rect 20168 52430 20220 52436
rect 20168 51944 20220 51950
rect 20168 51886 20220 51892
rect 19984 50798 20036 50804
rect 20074 50824 20130 50833
rect 20074 50759 20130 50768
rect 19812 50510 19932 50538
rect 19708 50312 19760 50318
rect 19708 50254 19760 50260
rect 19616 47660 19668 47666
rect 19616 47602 19668 47608
rect 19720 47274 19748 50254
rect 19800 49428 19852 49434
rect 19800 49370 19852 49376
rect 19812 48686 19840 49370
rect 19800 48680 19852 48686
rect 19904 48657 19932 50510
rect 19984 49088 20036 49094
rect 19984 49030 20036 49036
rect 19996 48929 20024 49030
rect 19982 48920 20038 48929
rect 19982 48855 20038 48864
rect 19996 48754 20024 48855
rect 19984 48748 20036 48754
rect 19984 48690 20036 48696
rect 19800 48622 19852 48628
rect 19890 48648 19946 48657
rect 19812 48346 19840 48622
rect 19890 48583 19946 48592
rect 19996 48362 20024 48690
rect 20088 48521 20116 50759
rect 20074 48512 20130 48521
rect 20074 48447 20130 48456
rect 19800 48340 19852 48346
rect 19996 48334 20116 48362
rect 19800 48282 19852 48288
rect 20088 48210 20116 48334
rect 19892 48204 19944 48210
rect 19892 48146 19944 48152
rect 20076 48204 20128 48210
rect 20076 48146 20128 48152
rect 19800 48136 19852 48142
rect 19800 48078 19852 48084
rect 19812 47802 19840 48078
rect 19904 47802 19932 48146
rect 19984 48136 20036 48142
rect 19984 48078 20036 48084
rect 19996 47841 20024 48078
rect 19982 47832 20038 47841
rect 19800 47796 19852 47802
rect 19800 47738 19852 47744
rect 19892 47796 19944 47802
rect 19982 47767 20038 47776
rect 19892 47738 19944 47744
rect 19628 47246 19748 47274
rect 19522 38856 19578 38865
rect 19522 38791 19578 38800
rect 19432 38208 19484 38214
rect 19432 38150 19484 38156
rect 19444 37126 19472 38150
rect 19524 38004 19576 38010
rect 19524 37946 19576 37952
rect 19536 37466 19564 37946
rect 19524 37460 19576 37466
rect 19524 37402 19576 37408
rect 19432 37120 19484 37126
rect 19432 37062 19484 37068
rect 19444 36242 19472 37062
rect 19628 36825 19656 47246
rect 19708 47116 19760 47122
rect 19708 47058 19760 47064
rect 19720 46578 19748 47058
rect 19708 46572 19760 46578
rect 19708 46514 19760 46520
rect 19812 46442 19840 47738
rect 19984 47728 20036 47734
rect 19984 47670 20036 47676
rect 19892 46912 19944 46918
rect 19892 46854 19944 46860
rect 19904 46510 19932 46854
rect 19892 46504 19944 46510
rect 19892 46446 19944 46452
rect 19708 46436 19760 46442
rect 19708 46378 19760 46384
rect 19800 46436 19852 46442
rect 19800 46378 19852 46384
rect 19720 44878 19748 46378
rect 19812 46170 19840 46378
rect 19800 46164 19852 46170
rect 19800 46106 19852 46112
rect 19800 45552 19852 45558
rect 19800 45494 19852 45500
rect 19708 44872 19760 44878
rect 19708 44814 19760 44820
rect 19812 44810 19840 45494
rect 19800 44804 19852 44810
rect 19800 44746 19852 44752
rect 19706 44704 19762 44713
rect 19706 44639 19762 44648
rect 19720 42770 19748 44639
rect 19812 44538 19840 44746
rect 19800 44532 19852 44538
rect 19800 44474 19852 44480
rect 19904 44169 19932 46446
rect 19996 45642 20024 47670
rect 20076 45824 20128 45830
rect 20074 45792 20076 45801
rect 20128 45792 20130 45801
rect 20074 45727 20130 45736
rect 19996 45614 20116 45642
rect 19984 45416 20036 45422
rect 19984 45358 20036 45364
rect 19996 45014 20024 45358
rect 19984 45008 20036 45014
rect 19984 44950 20036 44956
rect 19996 44742 20024 44950
rect 19984 44736 20036 44742
rect 19984 44678 20036 44684
rect 19890 44160 19946 44169
rect 19890 44095 19946 44104
rect 19904 43994 19932 44095
rect 19892 43988 19944 43994
rect 19892 43930 19944 43936
rect 19892 43852 19944 43858
rect 19892 43794 19944 43800
rect 19708 42764 19760 42770
rect 19708 42706 19760 42712
rect 19904 42634 19932 43794
rect 19996 43654 20024 44678
rect 20088 44198 20116 45614
rect 20076 44192 20128 44198
rect 20076 44134 20128 44140
rect 19984 43648 20036 43654
rect 19984 43590 20036 43596
rect 19996 43246 20024 43590
rect 20088 43382 20116 44134
rect 20076 43376 20128 43382
rect 20076 43318 20128 43324
rect 19984 43240 20036 43246
rect 19984 43182 20036 43188
rect 19892 42628 19944 42634
rect 19720 42588 19892 42616
rect 19720 42362 19748 42588
rect 19892 42570 19944 42576
rect 19996 42514 20024 43182
rect 20076 42764 20128 42770
rect 20076 42706 20128 42712
rect 19812 42486 20024 42514
rect 19708 42356 19760 42362
rect 19708 42298 19760 42304
rect 19720 41206 19748 42298
rect 19812 41274 19840 42486
rect 19890 42392 19946 42401
rect 19890 42327 19946 42336
rect 19904 42294 19932 42327
rect 19892 42288 19944 42294
rect 19892 42230 19944 42236
rect 20088 42158 20116 42706
rect 20076 42152 20128 42158
rect 20076 42094 20128 42100
rect 20074 41984 20130 41993
rect 20074 41919 20130 41928
rect 19892 41812 19944 41818
rect 19892 41754 19944 41760
rect 19800 41268 19852 41274
rect 19800 41210 19852 41216
rect 19708 41200 19760 41206
rect 19708 41142 19760 41148
rect 19798 41168 19854 41177
rect 19798 41103 19854 41112
rect 19614 36816 19670 36825
rect 19614 36751 19670 36760
rect 19614 36680 19670 36689
rect 19614 36615 19670 36624
rect 19628 36378 19656 36615
rect 19616 36372 19668 36378
rect 19616 36314 19668 36320
rect 19432 36236 19484 36242
rect 19432 36178 19484 36184
rect 19340 35828 19392 35834
rect 19340 35770 19392 35776
rect 19444 35601 19472 36178
rect 19430 35592 19486 35601
rect 19430 35527 19486 35536
rect 19338 35456 19394 35465
rect 19338 35391 19394 35400
rect 19352 35290 19380 35391
rect 19340 35284 19392 35290
rect 19340 35226 19392 35232
rect 19444 35154 19472 35527
rect 19432 35148 19484 35154
rect 19432 35090 19484 35096
rect 19430 35048 19486 35057
rect 19430 34983 19486 34992
rect 19444 34746 19472 34983
rect 19432 34740 19484 34746
rect 19432 34682 19484 34688
rect 19616 34468 19668 34474
rect 19616 34410 19668 34416
rect 19248 34060 19300 34066
rect 19248 34002 19300 34008
rect 19260 33658 19288 34002
rect 19248 33652 19300 33658
rect 19248 33594 19300 33600
rect 19628 33454 19656 34410
rect 19616 33448 19668 33454
rect 19616 33390 19668 33396
rect 19432 33312 19484 33318
rect 19430 33280 19432 33289
rect 19484 33280 19486 33289
rect 19430 33215 19486 33224
rect 19628 33114 19656 33390
rect 19706 33280 19762 33289
rect 19706 33215 19762 33224
rect 19616 33108 19668 33114
rect 19616 33050 19668 33056
rect 19156 32972 19208 32978
rect 19156 32914 19208 32920
rect 19168 32366 19196 32914
rect 19156 32360 19208 32366
rect 19156 32302 19208 32308
rect 18972 31816 19024 31822
rect 18972 31758 19024 31764
rect 19064 31748 19116 31754
rect 19064 31690 19116 31696
rect 19076 31278 19104 31690
rect 19064 31272 19116 31278
rect 18970 31240 19026 31249
rect 19064 31214 19116 31220
rect 18970 31175 19026 31184
rect 18880 30116 18932 30122
rect 18880 30058 18932 30064
rect 18694 30016 18750 30025
rect 18694 29951 18750 29960
rect 18708 29764 18736 29951
rect 18880 29776 18932 29782
rect 18708 29736 18880 29764
rect 18708 29238 18736 29736
rect 18880 29718 18932 29724
rect 18880 29504 18932 29510
rect 18880 29446 18932 29452
rect 18892 29238 18920 29446
rect 18696 29232 18748 29238
rect 18696 29174 18748 29180
rect 18880 29232 18932 29238
rect 18880 29174 18932 29180
rect 18696 29096 18748 29102
rect 18696 29038 18748 29044
rect 18708 28762 18736 29038
rect 18892 29034 18920 29174
rect 18880 29028 18932 29034
rect 18880 28970 18932 28976
rect 18878 28792 18934 28801
rect 18696 28756 18748 28762
rect 18878 28727 18880 28736
rect 18696 28698 18748 28704
rect 18932 28727 18934 28736
rect 18880 28698 18932 28704
rect 18696 28008 18748 28014
rect 18696 27950 18748 27956
rect 18788 28008 18840 28014
rect 18788 27950 18840 27956
rect 18708 27577 18736 27950
rect 18800 27674 18828 27950
rect 18788 27668 18840 27674
rect 18788 27610 18840 27616
rect 18694 27568 18750 27577
rect 18694 27503 18750 27512
rect 18696 26920 18748 26926
rect 18696 26862 18748 26868
rect 18708 26042 18736 26862
rect 18696 26036 18748 26042
rect 18696 25978 18748 25984
rect 18708 24954 18736 25978
rect 18696 24948 18748 24954
rect 18696 24890 18748 24896
rect 18604 22092 18656 22098
rect 18604 22034 18656 22040
rect 18616 21078 18644 22034
rect 18800 21622 18828 27610
rect 18880 27532 18932 27538
rect 18880 27474 18932 27480
rect 18892 26586 18920 27474
rect 18880 26580 18932 26586
rect 18880 26522 18932 26528
rect 18880 22228 18932 22234
rect 18880 22170 18932 22176
rect 18892 21962 18920 22170
rect 18880 21956 18932 21962
rect 18880 21898 18932 21904
rect 18788 21616 18840 21622
rect 18788 21558 18840 21564
rect 18604 21072 18656 21078
rect 18604 21014 18656 21020
rect 18984 21010 19012 31175
rect 19076 30734 19104 31214
rect 19168 30802 19196 32302
rect 19524 32020 19576 32026
rect 19524 31962 19576 31968
rect 19536 31822 19564 31962
rect 19616 31884 19668 31890
rect 19616 31826 19668 31832
rect 19524 31816 19576 31822
rect 19524 31758 19576 31764
rect 19156 30796 19208 30802
rect 19156 30738 19208 30744
rect 19064 30728 19116 30734
rect 19064 30670 19116 30676
rect 19064 30592 19116 30598
rect 19064 30534 19116 30540
rect 19076 30190 19104 30534
rect 19064 30184 19116 30190
rect 19064 30126 19116 30132
rect 19064 29708 19116 29714
rect 19064 29650 19116 29656
rect 19076 29481 19104 29650
rect 19168 29646 19196 30738
rect 19340 30660 19392 30666
rect 19340 30602 19392 30608
rect 19248 30320 19300 30326
rect 19246 30288 19248 30297
rect 19300 30288 19302 30297
rect 19246 30223 19302 30232
rect 19352 30138 19380 30602
rect 19536 30580 19564 31758
rect 19628 31482 19656 31826
rect 19616 31476 19668 31482
rect 19616 31418 19668 31424
rect 19616 30592 19668 30598
rect 19536 30552 19616 30580
rect 19616 30534 19668 30540
rect 19260 30122 19380 30138
rect 19248 30116 19380 30122
rect 19300 30110 19380 30116
rect 19430 30152 19486 30161
rect 19430 30087 19432 30096
rect 19248 30058 19300 30064
rect 19484 30087 19486 30096
rect 19432 30058 19484 30064
rect 19340 30048 19392 30054
rect 19260 29996 19340 30002
rect 19260 29990 19392 29996
rect 19260 29974 19380 29990
rect 19156 29640 19208 29646
rect 19156 29582 19208 29588
rect 19062 29472 19118 29481
rect 19062 29407 19118 29416
rect 19064 29232 19116 29238
rect 19064 29174 19116 29180
rect 19076 24274 19104 29174
rect 19168 26926 19196 29582
rect 19260 28098 19288 29974
rect 19340 29504 19392 29510
rect 19340 29446 19392 29452
rect 19352 29238 19380 29446
rect 19340 29232 19392 29238
rect 19340 29174 19392 29180
rect 19444 29102 19472 30058
rect 19628 30054 19656 30534
rect 19616 30048 19668 30054
rect 19616 29990 19668 29996
rect 19432 29096 19484 29102
rect 19432 29038 19484 29044
rect 19432 28960 19484 28966
rect 19338 28928 19394 28937
rect 19432 28902 19484 28908
rect 19338 28863 19394 28872
rect 19352 28762 19380 28863
rect 19340 28756 19392 28762
rect 19340 28698 19392 28704
rect 19444 28626 19472 28902
rect 19432 28620 19484 28626
rect 19432 28562 19484 28568
rect 19444 28218 19472 28562
rect 19616 28416 19668 28422
rect 19616 28358 19668 28364
rect 19628 28257 19656 28358
rect 19614 28248 19670 28257
rect 19432 28212 19484 28218
rect 19614 28183 19670 28192
rect 19432 28154 19484 28160
rect 19444 28121 19472 28154
rect 19430 28112 19486 28121
rect 19260 28070 19380 28098
rect 19248 27940 19300 27946
rect 19248 27882 19300 27888
rect 19260 27554 19288 27882
rect 19352 27826 19380 28070
rect 19430 28047 19486 28056
rect 19352 27798 19472 27826
rect 19260 27526 19380 27554
rect 19352 27470 19380 27526
rect 19340 27464 19392 27470
rect 19340 27406 19392 27412
rect 19444 27316 19472 27798
rect 19260 27288 19472 27316
rect 19156 26920 19208 26926
rect 19156 26862 19208 26868
rect 19260 25265 19288 27288
rect 19524 27124 19576 27130
rect 19524 27066 19576 27072
rect 19246 25256 19302 25265
rect 19246 25191 19302 25200
rect 19154 24848 19210 24857
rect 19154 24783 19210 24792
rect 19064 24268 19116 24274
rect 19064 24210 19116 24216
rect 19076 23866 19104 24210
rect 19064 23860 19116 23866
rect 19064 23802 19116 23808
rect 19064 22024 19116 22030
rect 19064 21966 19116 21972
rect 19076 21321 19104 21966
rect 19062 21312 19118 21321
rect 19062 21247 19118 21256
rect 18972 21004 19024 21010
rect 18972 20946 19024 20952
rect 18512 20528 18564 20534
rect 18512 20470 18564 20476
rect 18696 20392 18748 20398
rect 18696 20334 18748 20340
rect 18708 19854 18736 20334
rect 18984 19990 19012 20946
rect 19076 20806 19104 21247
rect 19064 20800 19116 20806
rect 19064 20742 19116 20748
rect 18972 19984 19024 19990
rect 18972 19926 19024 19932
rect 18696 19848 18748 19854
rect 18696 19790 18748 19796
rect 18984 19514 19012 19926
rect 18972 19508 19024 19514
rect 18972 19450 19024 19456
rect 18418 11656 18474 11665
rect 18418 11591 18474 11600
rect 19062 10568 19118 10577
rect 19062 10503 19064 10512
rect 19116 10503 19118 10512
rect 19064 10474 19116 10480
rect 18788 10124 18840 10130
rect 18788 10066 18840 10072
rect 18800 9722 18828 10066
rect 18788 9716 18840 9722
rect 18788 9658 18840 9664
rect 18326 5536 18382 5545
rect 18326 5471 18382 5480
rect 19168 5273 19196 24783
rect 19260 22030 19288 25191
rect 19340 22432 19392 22438
rect 19340 22374 19392 22380
rect 19352 22098 19380 22374
rect 19340 22092 19392 22098
rect 19340 22034 19392 22040
rect 19248 22024 19300 22030
rect 19248 21966 19300 21972
rect 19260 21146 19288 21966
rect 19352 21690 19380 22034
rect 19340 21684 19392 21690
rect 19340 21626 19392 21632
rect 19248 21140 19300 21146
rect 19248 21082 19300 21088
rect 19248 20800 19300 20806
rect 19246 20768 19248 20777
rect 19300 20768 19302 20777
rect 19246 20703 19302 20712
rect 19536 20482 19564 27066
rect 19616 22772 19668 22778
rect 19616 22714 19668 22720
rect 19444 20454 19564 20482
rect 19248 19848 19300 19854
rect 19248 19790 19300 19796
rect 19260 19378 19288 19790
rect 19248 19372 19300 19378
rect 19248 19314 19300 19320
rect 19444 19310 19472 20454
rect 19522 20360 19578 20369
rect 19522 20295 19578 20304
rect 19536 19990 19564 20295
rect 19524 19984 19576 19990
rect 19524 19926 19576 19932
rect 19432 19304 19484 19310
rect 19432 19246 19484 19252
rect 19248 10668 19300 10674
rect 19248 10610 19300 10616
rect 19260 10266 19288 10610
rect 19248 10260 19300 10266
rect 19248 10202 19300 10208
rect 19430 5536 19486 5545
rect 19430 5471 19486 5480
rect 19154 5264 19210 5273
rect 19154 5199 19210 5208
rect 19444 3738 19472 5471
rect 19432 3732 19484 3738
rect 19432 3674 19484 3680
rect 17960 3596 18012 3602
rect 17960 3538 18012 3544
rect 17972 3126 18000 3538
rect 18144 3528 18196 3534
rect 18144 3470 18196 3476
rect 18156 3194 18184 3470
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 18420 3188 18472 3194
rect 18420 3130 18472 3136
rect 17960 3120 18012 3126
rect 17960 3062 18012 3068
rect 17972 2650 18000 3062
rect 17960 2644 18012 2650
rect 17960 2586 18012 2592
rect 17972 2446 18000 2586
rect 17960 2440 18012 2446
rect 17960 2382 18012 2388
rect 18144 2304 18196 2310
rect 18144 2246 18196 2252
rect 17682 2000 17738 2009
rect 17682 1935 17738 1944
rect 18156 1170 18184 2246
rect 17972 1142 18184 1170
rect 17972 800 18000 1142
rect 18432 800 18460 3130
rect 19628 2632 19656 22714
rect 19720 16250 19748 33215
rect 19812 32434 19840 41103
rect 19904 35290 19932 41754
rect 19984 41676 20036 41682
rect 19984 41618 20036 41624
rect 19996 41274 20024 41618
rect 19984 41268 20036 41274
rect 19984 41210 20036 41216
rect 19982 36544 20038 36553
rect 19982 36479 20038 36488
rect 19996 36378 20024 36479
rect 19984 36372 20036 36378
rect 19984 36314 20036 36320
rect 19892 35284 19944 35290
rect 19892 35226 19944 35232
rect 20088 34746 20116 41919
rect 20076 34740 20128 34746
rect 20076 34682 20128 34688
rect 20088 34542 20116 34682
rect 20076 34536 20128 34542
rect 19890 34504 19946 34513
rect 20076 34478 20128 34484
rect 19890 34439 19946 34448
rect 19800 32428 19852 32434
rect 19800 32370 19852 32376
rect 19904 32314 19932 34439
rect 20076 33856 20128 33862
rect 20076 33798 20128 33804
rect 19984 32768 20036 32774
rect 19982 32736 19984 32745
rect 20036 32736 20038 32745
rect 19982 32671 20038 32680
rect 19812 32286 19932 32314
rect 19812 27130 19840 32286
rect 19892 31952 19944 31958
rect 19892 31894 19944 31900
rect 19904 30954 19932 31894
rect 19996 31822 20024 32671
rect 19984 31816 20036 31822
rect 19984 31758 20036 31764
rect 20088 31657 20116 33798
rect 20074 31648 20130 31657
rect 20074 31583 20130 31592
rect 19984 31136 20036 31142
rect 19982 31104 19984 31113
rect 20036 31104 20038 31113
rect 19982 31039 20038 31048
rect 19904 30926 20024 30954
rect 19892 30728 19944 30734
rect 19892 30670 19944 30676
rect 19904 29714 19932 30670
rect 19892 29708 19944 29714
rect 19892 29650 19944 29656
rect 19890 29336 19946 29345
rect 19890 29271 19892 29280
rect 19944 29271 19946 29280
rect 19892 29242 19944 29248
rect 19996 28082 20024 30926
rect 20088 30190 20116 31583
rect 20076 30184 20128 30190
rect 20076 30126 20128 30132
rect 20088 29850 20116 30126
rect 20076 29844 20128 29850
rect 20076 29786 20128 29792
rect 20088 28762 20116 29786
rect 20076 28756 20128 28762
rect 20076 28698 20128 28704
rect 19984 28076 20036 28082
rect 19984 28018 20036 28024
rect 20076 27872 20128 27878
rect 20074 27840 20076 27849
rect 20128 27840 20130 27849
rect 20074 27775 20130 27784
rect 20074 27568 20130 27577
rect 20074 27503 20076 27512
rect 20128 27503 20130 27512
rect 20076 27474 20128 27480
rect 19892 27328 19944 27334
rect 19892 27270 19944 27276
rect 19800 27124 19852 27130
rect 19800 27066 19852 27072
rect 19904 21457 19932 27270
rect 20088 27130 20116 27474
rect 20076 27124 20128 27130
rect 20076 27066 20128 27072
rect 19890 21448 19946 21457
rect 19890 21383 19946 21392
rect 20180 19553 20208 51886
rect 20272 41449 20300 53910
rect 20364 53514 20392 54470
rect 20352 53508 20404 53514
rect 20352 53450 20404 53456
rect 20456 52408 20484 55814
rect 20548 52476 20576 65962
rect 20732 64530 20760 66286
rect 20720 64524 20772 64530
rect 20720 64466 20772 64472
rect 20718 64016 20774 64025
rect 20718 63951 20774 63960
rect 20732 61402 20760 63951
rect 20720 61396 20772 61402
rect 20720 61338 20772 61344
rect 20732 61282 20760 61338
rect 20640 61254 20760 61282
rect 20640 60722 20668 61254
rect 20824 61062 20852 71334
rect 20956 71292 21252 71312
rect 21012 71290 21036 71292
rect 21092 71290 21116 71292
rect 21172 71290 21196 71292
rect 21034 71238 21036 71290
rect 21098 71238 21110 71290
rect 21172 71238 21174 71290
rect 21012 71236 21036 71238
rect 21092 71236 21116 71238
rect 21172 71236 21196 71238
rect 20956 71216 21252 71236
rect 20996 71052 21048 71058
rect 20996 70994 21048 71000
rect 21008 70938 21036 70994
rect 20916 70910 21036 70938
rect 20916 70582 20944 70910
rect 20904 70576 20956 70582
rect 20902 70544 20904 70553
rect 20956 70544 20958 70553
rect 20902 70479 20958 70488
rect 20956 70204 21252 70224
rect 21012 70202 21036 70204
rect 21092 70202 21116 70204
rect 21172 70202 21196 70204
rect 21034 70150 21036 70202
rect 21098 70150 21110 70202
rect 21172 70150 21174 70202
rect 21012 70148 21036 70150
rect 21092 70148 21116 70150
rect 21172 70148 21196 70150
rect 20956 70128 21252 70148
rect 21284 69737 21312 76327
rect 21376 75750 21404 76366
rect 21364 75744 21416 75750
rect 21364 75686 21416 75692
rect 21376 72078 21404 75686
rect 22112 74746 22140 79200
rect 22112 74718 22232 74746
rect 22100 74656 22152 74662
rect 22100 74598 22152 74604
rect 21364 72072 21416 72078
rect 21364 72014 21416 72020
rect 21376 71398 21404 72014
rect 21364 71392 21416 71398
rect 21364 71334 21416 71340
rect 21376 70990 21404 71334
rect 21364 70984 21416 70990
rect 21364 70926 21416 70932
rect 21376 70446 21404 70926
rect 21364 70440 21416 70446
rect 21364 70382 21416 70388
rect 21732 70440 21784 70446
rect 21732 70382 21784 70388
rect 21270 69728 21326 69737
rect 21270 69663 21326 69672
rect 20956 69116 21252 69136
rect 21012 69114 21036 69116
rect 21092 69114 21116 69116
rect 21172 69114 21196 69116
rect 21034 69062 21036 69114
rect 21098 69062 21110 69114
rect 21172 69062 21174 69114
rect 21012 69060 21036 69062
rect 21092 69060 21116 69062
rect 21172 69060 21196 69062
rect 20956 69040 21252 69060
rect 20956 68028 21252 68048
rect 21012 68026 21036 68028
rect 21092 68026 21116 68028
rect 21172 68026 21196 68028
rect 21034 67974 21036 68026
rect 21098 67974 21110 68026
rect 21172 67974 21174 68026
rect 21012 67972 21036 67974
rect 21092 67972 21116 67974
rect 21172 67972 21196 67974
rect 20956 67952 21252 67972
rect 21454 67688 21510 67697
rect 21454 67623 21510 67632
rect 20956 66940 21252 66960
rect 21012 66938 21036 66940
rect 21092 66938 21116 66940
rect 21172 66938 21196 66940
rect 21034 66886 21036 66938
rect 21098 66886 21110 66938
rect 21172 66886 21174 66938
rect 21012 66884 21036 66886
rect 21092 66884 21116 66886
rect 21172 66884 21196 66886
rect 20956 66864 21252 66884
rect 20956 65852 21252 65872
rect 21012 65850 21036 65852
rect 21092 65850 21116 65852
rect 21172 65850 21196 65852
rect 21034 65798 21036 65850
rect 21098 65798 21110 65850
rect 21172 65798 21174 65850
rect 21012 65796 21036 65798
rect 21092 65796 21116 65798
rect 21172 65796 21196 65798
rect 20956 65776 21252 65796
rect 20956 64764 21252 64784
rect 21012 64762 21036 64764
rect 21092 64762 21116 64764
rect 21172 64762 21196 64764
rect 21034 64710 21036 64762
rect 21098 64710 21110 64762
rect 21172 64710 21174 64762
rect 21012 64708 21036 64710
rect 21092 64708 21116 64710
rect 21172 64708 21196 64710
rect 20956 64688 21252 64708
rect 20956 63676 21252 63696
rect 21012 63674 21036 63676
rect 21092 63674 21116 63676
rect 21172 63674 21196 63676
rect 21034 63622 21036 63674
rect 21098 63622 21110 63674
rect 21172 63622 21174 63674
rect 21012 63620 21036 63622
rect 21092 63620 21116 63622
rect 21172 63620 21196 63622
rect 20956 63600 21252 63620
rect 20956 62588 21252 62608
rect 21012 62586 21036 62588
rect 21092 62586 21116 62588
rect 21172 62586 21196 62588
rect 21034 62534 21036 62586
rect 21098 62534 21110 62586
rect 21172 62534 21174 62586
rect 21012 62532 21036 62534
rect 21092 62532 21116 62534
rect 21172 62532 21196 62534
rect 20956 62512 21252 62532
rect 20956 61500 21252 61520
rect 21012 61498 21036 61500
rect 21092 61498 21116 61500
rect 21172 61498 21196 61500
rect 21034 61446 21036 61498
rect 21098 61446 21110 61498
rect 21172 61446 21174 61498
rect 21012 61444 21036 61446
rect 21092 61444 21116 61446
rect 21172 61444 21196 61446
rect 20956 61424 21252 61444
rect 21468 61334 21496 67623
rect 21744 66842 21772 70382
rect 21914 69864 21970 69873
rect 21914 69799 21970 69808
rect 21732 66836 21784 66842
rect 21732 66778 21784 66784
rect 21744 64546 21772 66778
rect 21824 66700 21876 66706
rect 21824 66642 21876 66648
rect 21836 66298 21864 66642
rect 21824 66292 21876 66298
rect 21824 66234 21876 66240
rect 21836 65210 21864 66234
rect 21824 65204 21876 65210
rect 21824 65146 21876 65152
rect 21548 64524 21600 64530
rect 21548 64466 21600 64472
rect 21652 64518 21772 64546
rect 21560 64122 21588 64466
rect 21652 64462 21680 64518
rect 21640 64456 21692 64462
rect 21640 64398 21692 64404
rect 21652 64122 21680 64398
rect 21548 64116 21600 64122
rect 21548 64058 21600 64064
rect 21640 64116 21692 64122
rect 21640 64058 21692 64064
rect 21652 64025 21680 64058
rect 21638 64016 21694 64025
rect 21638 63951 21694 63960
rect 21822 63608 21878 63617
rect 21822 63543 21878 63552
rect 21456 61328 21508 61334
rect 21456 61270 21508 61276
rect 21364 61192 21416 61198
rect 21364 61134 21416 61140
rect 21272 61124 21324 61130
rect 21272 61066 21324 61072
rect 20812 61056 20864 61062
rect 20812 60998 20864 61004
rect 21284 60722 21312 61066
rect 21376 60722 21404 61134
rect 21456 61056 21508 61062
rect 21456 60998 21508 61004
rect 20628 60716 20680 60722
rect 20628 60658 20680 60664
rect 21272 60716 21324 60722
rect 21272 60658 21324 60664
rect 21364 60716 21416 60722
rect 21364 60658 21416 60664
rect 20720 60648 20772 60654
rect 20720 60590 20772 60596
rect 20628 60172 20680 60178
rect 20628 60114 20680 60120
rect 20640 58070 20668 60114
rect 20732 58138 20760 60590
rect 20956 60412 21252 60432
rect 21012 60410 21036 60412
rect 21092 60410 21116 60412
rect 21172 60410 21196 60412
rect 21034 60358 21036 60410
rect 21098 60358 21110 60410
rect 21172 60358 21174 60410
rect 21012 60356 21036 60358
rect 21092 60356 21116 60358
rect 21172 60356 21196 60358
rect 20956 60336 21252 60356
rect 21376 59566 21404 60658
rect 21272 59560 21324 59566
rect 21272 59502 21324 59508
rect 21364 59560 21416 59566
rect 21364 59502 21416 59508
rect 20956 59324 21252 59344
rect 21012 59322 21036 59324
rect 21092 59322 21116 59324
rect 21172 59322 21196 59324
rect 21034 59270 21036 59322
rect 21098 59270 21110 59322
rect 21172 59270 21174 59322
rect 21012 59268 21036 59270
rect 21092 59268 21116 59270
rect 21172 59268 21196 59270
rect 20956 59248 21252 59268
rect 20996 58948 21048 58954
rect 20996 58890 21048 58896
rect 21008 58478 21036 58890
rect 20996 58472 21048 58478
rect 21284 58449 21312 59502
rect 21376 59158 21404 59502
rect 21364 59152 21416 59158
rect 21364 59094 21416 59100
rect 20996 58414 21048 58420
rect 21270 58440 21326 58449
rect 21270 58375 21326 58384
rect 20956 58236 21252 58256
rect 21012 58234 21036 58236
rect 21092 58234 21116 58236
rect 21172 58234 21196 58236
rect 21034 58182 21036 58234
rect 21098 58182 21110 58234
rect 21172 58182 21174 58234
rect 21012 58180 21036 58182
rect 21092 58180 21116 58182
rect 21172 58180 21196 58182
rect 20956 58160 21252 58180
rect 20720 58132 20772 58138
rect 20720 58074 20772 58080
rect 20628 58064 20680 58070
rect 20628 58006 20680 58012
rect 20996 58064 21048 58070
rect 20996 58006 21048 58012
rect 20732 57934 20760 57965
rect 20720 57928 20772 57934
rect 20718 57896 20720 57905
rect 20772 57896 20774 57905
rect 20718 57831 20774 57840
rect 20732 57390 20760 57831
rect 20812 57588 20864 57594
rect 20812 57530 20864 57536
rect 20720 57384 20772 57390
rect 20720 57326 20772 57332
rect 20628 57248 20680 57254
rect 20628 57190 20680 57196
rect 20640 56386 20668 57190
rect 20732 57050 20760 57326
rect 20720 57044 20772 57050
rect 20720 56986 20772 56992
rect 20718 56536 20774 56545
rect 20718 56471 20720 56480
rect 20772 56471 20774 56480
rect 20720 56442 20772 56448
rect 20640 56358 20760 56386
rect 20732 56302 20760 56358
rect 20720 56296 20772 56302
rect 20718 56264 20720 56273
rect 20772 56264 20774 56273
rect 20718 56199 20774 56208
rect 20626 55584 20682 55593
rect 20626 55519 20682 55528
rect 20640 55214 20668 55519
rect 20628 55208 20680 55214
rect 20628 55150 20680 55156
rect 20720 54664 20772 54670
rect 20720 54606 20772 54612
rect 20628 54052 20680 54058
rect 20628 53994 20680 54000
rect 20640 53666 20668 53994
rect 20732 53786 20760 54606
rect 20720 53780 20772 53786
rect 20720 53722 20772 53728
rect 20640 53638 20760 53666
rect 20732 53242 20760 53638
rect 20720 53236 20772 53242
rect 20720 53178 20772 53184
rect 20628 53100 20680 53106
rect 20628 53042 20680 53048
rect 20640 52601 20668 53042
rect 20720 52964 20772 52970
rect 20720 52906 20772 52912
rect 20732 52698 20760 52906
rect 20720 52692 20772 52698
rect 20720 52634 20772 52640
rect 20626 52592 20682 52601
rect 20626 52527 20682 52536
rect 20720 52488 20772 52494
rect 20548 52448 20668 52476
rect 20456 52380 20576 52408
rect 20352 52352 20404 52358
rect 20352 52294 20404 52300
rect 20364 51814 20392 52294
rect 20352 51808 20404 51814
rect 20352 51750 20404 51756
rect 20364 51406 20392 51750
rect 20352 51400 20404 51406
rect 20352 51342 20404 51348
rect 20364 50522 20392 51342
rect 20444 50720 20496 50726
rect 20444 50662 20496 50668
rect 20352 50516 20404 50522
rect 20352 50458 20404 50464
rect 20352 50312 20404 50318
rect 20352 50254 20404 50260
rect 20364 49978 20392 50254
rect 20352 49972 20404 49978
rect 20352 49914 20404 49920
rect 20364 49881 20392 49914
rect 20350 49872 20406 49881
rect 20350 49807 20406 49816
rect 20456 49774 20484 50662
rect 20444 49768 20496 49774
rect 20444 49710 20496 49716
rect 20352 49292 20404 49298
rect 20352 49234 20404 49240
rect 20364 47734 20392 49234
rect 20352 47728 20404 47734
rect 20352 47670 20404 47676
rect 20456 47462 20484 49710
rect 20444 47456 20496 47462
rect 20444 47398 20496 47404
rect 20352 46368 20404 46374
rect 20352 46310 20404 46316
rect 20364 45422 20392 46310
rect 20352 45416 20404 45422
rect 20352 45358 20404 45364
rect 20364 45082 20392 45358
rect 20352 45076 20404 45082
rect 20352 45018 20404 45024
rect 20352 44872 20404 44878
rect 20350 44840 20352 44849
rect 20404 44840 20406 44849
rect 20350 44775 20406 44784
rect 20456 44470 20484 47398
rect 20352 44464 20404 44470
rect 20352 44406 20404 44412
rect 20444 44464 20496 44470
rect 20444 44406 20496 44412
rect 20364 41818 20392 44406
rect 20444 44328 20496 44334
rect 20444 44270 20496 44276
rect 20456 42770 20484 44270
rect 20444 42764 20496 42770
rect 20444 42706 20496 42712
rect 20442 42664 20498 42673
rect 20442 42599 20444 42608
rect 20496 42599 20498 42608
rect 20444 42570 20496 42576
rect 20444 42288 20496 42294
rect 20444 42230 20496 42236
rect 20352 41812 20404 41818
rect 20352 41754 20404 41760
rect 20258 41440 20314 41449
rect 20258 41375 20314 41384
rect 20260 37800 20312 37806
rect 20260 37742 20312 37748
rect 20350 37768 20406 37777
rect 20272 37466 20300 37742
rect 20350 37703 20352 37712
rect 20404 37703 20406 37712
rect 20352 37674 20404 37680
rect 20260 37460 20312 37466
rect 20260 37402 20312 37408
rect 20456 36378 20484 42230
rect 20548 41313 20576 52380
rect 20534 41304 20590 41313
rect 20534 41239 20590 41248
rect 20534 41168 20590 41177
rect 20534 41103 20590 41112
rect 20548 38185 20576 41103
rect 20534 38176 20590 38185
rect 20534 38111 20590 38120
rect 20444 36372 20496 36378
rect 20444 36314 20496 36320
rect 20258 36136 20314 36145
rect 20258 36071 20260 36080
rect 20312 36071 20314 36080
rect 20260 36042 20312 36048
rect 20640 35816 20668 52448
rect 20720 52430 20772 52436
rect 20732 52154 20760 52430
rect 20720 52148 20772 52154
rect 20720 52090 20772 52096
rect 20824 50998 20852 57530
rect 21008 57361 21036 58006
rect 21364 57928 21416 57934
rect 21364 57870 21416 57876
rect 20994 57352 21050 57361
rect 20994 57287 21050 57296
rect 20956 57148 21252 57168
rect 21012 57146 21036 57148
rect 21092 57146 21116 57148
rect 21172 57146 21196 57148
rect 21034 57094 21036 57146
rect 21098 57094 21110 57146
rect 21172 57094 21174 57146
rect 21012 57092 21036 57094
rect 21092 57092 21116 57094
rect 21172 57092 21196 57094
rect 20956 57072 21252 57092
rect 20996 56908 21048 56914
rect 20996 56850 21048 56856
rect 21008 56506 21036 56850
rect 21376 56846 21404 57870
rect 21364 56840 21416 56846
rect 21364 56782 21416 56788
rect 20996 56500 21048 56506
rect 20996 56442 21048 56448
rect 21008 56409 21036 56442
rect 20994 56400 21050 56409
rect 20994 56335 21050 56344
rect 21364 56296 21416 56302
rect 21364 56238 21416 56244
rect 21272 56228 21324 56234
rect 21272 56170 21324 56176
rect 20956 56060 21252 56080
rect 21012 56058 21036 56060
rect 21092 56058 21116 56060
rect 21172 56058 21196 56060
rect 21034 56006 21036 56058
rect 21098 56006 21110 56058
rect 21172 56006 21174 56058
rect 21012 56004 21036 56006
rect 21092 56004 21116 56006
rect 21172 56004 21196 56006
rect 20956 55984 21252 56004
rect 20902 55856 20958 55865
rect 20902 55791 20904 55800
rect 20956 55791 20958 55800
rect 20904 55762 20956 55768
rect 21088 55616 21140 55622
rect 21088 55558 21140 55564
rect 21100 55321 21128 55558
rect 21284 55321 21312 56170
rect 21376 55457 21404 56238
rect 21362 55448 21418 55457
rect 21362 55383 21418 55392
rect 21086 55312 21142 55321
rect 21086 55247 21142 55256
rect 21270 55312 21326 55321
rect 21270 55247 21326 55256
rect 21362 55040 21418 55049
rect 20956 54972 21252 54992
rect 21362 54975 21418 54984
rect 21012 54970 21036 54972
rect 21092 54970 21116 54972
rect 21172 54970 21196 54972
rect 21034 54918 21036 54970
rect 21098 54918 21110 54970
rect 21172 54918 21174 54970
rect 21012 54916 21036 54918
rect 21092 54916 21116 54918
rect 21172 54916 21196 54918
rect 20956 54896 21252 54916
rect 21086 54768 21142 54777
rect 21086 54703 21088 54712
rect 21140 54703 21142 54712
rect 21088 54674 21140 54680
rect 21376 54670 21404 54975
rect 21364 54664 21416 54670
rect 21364 54606 21416 54612
rect 20956 53884 21252 53904
rect 21012 53882 21036 53884
rect 21092 53882 21116 53884
rect 21172 53882 21196 53884
rect 21034 53830 21036 53882
rect 21098 53830 21110 53882
rect 21172 53830 21174 53882
rect 21012 53828 21036 53830
rect 21092 53828 21116 53830
rect 21172 53828 21196 53830
rect 20956 53808 21252 53828
rect 21088 53644 21140 53650
rect 21088 53586 21140 53592
rect 21100 53009 21128 53586
rect 21364 53576 21416 53582
rect 21364 53518 21416 53524
rect 21086 53000 21142 53009
rect 21086 52935 21088 52944
rect 21140 52935 21142 52944
rect 21088 52906 21140 52912
rect 20956 52796 21252 52816
rect 21012 52794 21036 52796
rect 21092 52794 21116 52796
rect 21172 52794 21196 52796
rect 21034 52742 21036 52794
rect 21098 52742 21110 52794
rect 21172 52742 21174 52794
rect 21012 52740 21036 52742
rect 21092 52740 21116 52742
rect 21172 52740 21196 52742
rect 20956 52720 21252 52740
rect 21376 52562 21404 53518
rect 21364 52556 21416 52562
rect 21364 52498 21416 52504
rect 21376 52154 21404 52498
rect 21364 52148 21416 52154
rect 21364 52090 21416 52096
rect 21364 51944 21416 51950
rect 21364 51886 21416 51892
rect 20956 51708 21252 51728
rect 21012 51706 21036 51708
rect 21092 51706 21116 51708
rect 21172 51706 21196 51708
rect 21034 51654 21036 51706
rect 21098 51654 21110 51706
rect 21172 51654 21174 51706
rect 21012 51652 21036 51654
rect 21092 51652 21116 51654
rect 21172 51652 21196 51654
rect 20956 51632 21252 51652
rect 21376 51610 21404 51886
rect 21364 51604 21416 51610
rect 21284 51564 21364 51592
rect 21178 51504 21234 51513
rect 21178 51439 21234 51448
rect 20812 50992 20864 50998
rect 20812 50934 20864 50940
rect 21192 50794 21220 51439
rect 20812 50788 20864 50794
rect 20812 50730 20864 50736
rect 21180 50788 21232 50794
rect 21180 50730 21232 50736
rect 20720 50720 20772 50726
rect 20720 50662 20772 50668
rect 20732 49638 20760 50662
rect 20824 49706 20852 50730
rect 20956 50620 21252 50640
rect 21012 50618 21036 50620
rect 21092 50618 21116 50620
rect 21172 50618 21196 50620
rect 21034 50566 21036 50618
rect 21098 50566 21110 50618
rect 21172 50566 21174 50618
rect 21012 50564 21036 50566
rect 21092 50564 21116 50566
rect 21172 50564 21196 50566
rect 20956 50544 21252 50564
rect 21284 50522 21312 51564
rect 21364 51546 21416 51552
rect 21468 51490 21496 60998
rect 21548 60648 21600 60654
rect 21548 60590 21600 60596
rect 21560 60178 21588 60590
rect 21548 60172 21600 60178
rect 21548 60114 21600 60120
rect 21560 59650 21588 60114
rect 21836 60110 21864 63543
rect 21824 60104 21876 60110
rect 21824 60046 21876 60052
rect 21560 59622 21680 59650
rect 21928 59634 21956 69799
rect 22008 61260 22060 61266
rect 22008 61202 22060 61208
rect 22020 60858 22048 61202
rect 22008 60852 22060 60858
rect 22008 60794 22060 60800
rect 22112 60738 22140 74598
rect 22204 62257 22232 74718
rect 22572 74662 22600 79200
rect 22744 76900 22796 76906
rect 22744 76842 22796 76848
rect 22652 76288 22704 76294
rect 22652 76230 22704 76236
rect 22560 74656 22612 74662
rect 22560 74598 22612 74604
rect 22558 73536 22614 73545
rect 22558 73471 22614 73480
rect 22572 72214 22600 73471
rect 22560 72208 22612 72214
rect 22560 72150 22612 72156
rect 22282 69728 22338 69737
rect 22282 69663 22338 69672
rect 22190 62248 22246 62257
rect 22190 62183 22246 62192
rect 22020 60710 22140 60738
rect 21652 59566 21680 59622
rect 21916 59628 21968 59634
rect 21916 59570 21968 59576
rect 21640 59560 21692 59566
rect 21640 59502 21692 59508
rect 21546 58576 21602 58585
rect 21546 58511 21602 58520
rect 21560 53145 21588 58511
rect 21652 57526 21680 59502
rect 21824 59084 21876 59090
rect 21824 59026 21876 59032
rect 21836 58682 21864 59026
rect 21824 58676 21876 58682
rect 21824 58618 21876 58624
rect 21836 58342 21864 58618
rect 21824 58336 21876 58342
rect 21824 58278 21876 58284
rect 21640 57520 21692 57526
rect 21640 57462 21692 57468
rect 21652 57050 21680 57462
rect 21824 57316 21876 57322
rect 21824 57258 21876 57264
rect 21836 57225 21864 57258
rect 21822 57216 21878 57225
rect 21822 57151 21878 57160
rect 21640 57044 21692 57050
rect 21640 56986 21692 56992
rect 22020 56930 22048 60710
rect 22192 60036 22244 60042
rect 22192 59978 22244 59984
rect 22204 59430 22232 59978
rect 22192 59424 22244 59430
rect 22192 59366 22244 59372
rect 22100 59016 22152 59022
rect 22100 58958 22152 58964
rect 22112 57934 22140 58958
rect 22100 57928 22152 57934
rect 22100 57870 22152 57876
rect 22112 57594 22140 57870
rect 22100 57588 22152 57594
rect 22100 57530 22152 57536
rect 21744 56902 22048 56930
rect 21640 56160 21692 56166
rect 21640 56102 21692 56108
rect 21652 55962 21680 56102
rect 21640 55956 21692 55962
rect 21640 55898 21692 55904
rect 21640 55820 21692 55826
rect 21640 55762 21692 55768
rect 21652 55078 21680 55762
rect 21640 55072 21692 55078
rect 21640 55014 21692 55020
rect 21546 53136 21602 53145
rect 21546 53071 21602 53080
rect 21548 52148 21600 52154
rect 21548 52090 21600 52096
rect 21376 51462 21496 51490
rect 21560 51474 21588 52090
rect 21548 51468 21600 51474
rect 21272 50516 21324 50522
rect 21272 50458 21324 50464
rect 20904 49904 20956 49910
rect 20902 49872 20904 49881
rect 20956 49872 20958 49881
rect 20902 49807 20958 49816
rect 20812 49700 20864 49706
rect 20812 49642 20864 49648
rect 20720 49632 20772 49638
rect 20720 49574 20772 49580
rect 20718 49464 20774 49473
rect 20718 49399 20774 49408
rect 20732 48260 20760 49399
rect 20824 49201 20852 49642
rect 21272 49632 21324 49638
rect 21272 49574 21324 49580
rect 20956 49532 21252 49552
rect 21012 49530 21036 49532
rect 21092 49530 21116 49532
rect 21172 49530 21196 49532
rect 21034 49478 21036 49530
rect 21098 49478 21110 49530
rect 21172 49478 21174 49530
rect 21012 49476 21036 49478
rect 21092 49476 21116 49478
rect 21172 49476 21196 49478
rect 20956 49456 21252 49476
rect 21284 49434 21312 49574
rect 21272 49428 21324 49434
rect 21272 49370 21324 49376
rect 20810 49192 20866 49201
rect 20810 49127 20866 49136
rect 21284 48890 21312 49370
rect 21272 48884 21324 48890
rect 21272 48826 21324 48832
rect 20956 48444 21252 48464
rect 21012 48442 21036 48444
rect 21092 48442 21116 48444
rect 21172 48442 21196 48444
rect 21034 48390 21036 48442
rect 21098 48390 21110 48442
rect 21172 48390 21174 48442
rect 21012 48388 21036 48390
rect 21092 48388 21116 48390
rect 21172 48388 21196 48390
rect 20956 48368 21252 48388
rect 20732 48232 20852 48260
rect 20720 47592 20772 47598
rect 20720 47534 20772 47540
rect 20732 46578 20760 47534
rect 20720 46572 20772 46578
rect 20720 46514 20772 46520
rect 20732 46034 20760 46514
rect 20720 46028 20772 46034
rect 20720 45970 20772 45976
rect 20720 45620 20772 45626
rect 20720 45562 20772 45568
rect 20732 44810 20760 45562
rect 20720 44804 20772 44810
rect 20720 44746 20772 44752
rect 20732 43314 20760 44746
rect 20720 43308 20772 43314
rect 20720 43250 20772 43256
rect 20720 43172 20772 43178
rect 20720 43114 20772 43120
rect 20732 42362 20760 43114
rect 20720 42356 20772 42362
rect 20720 42298 20772 42304
rect 20720 41744 20772 41750
rect 20718 41712 20720 41721
rect 20772 41712 20774 41721
rect 20718 41647 20774 41656
rect 20718 41576 20774 41585
rect 20718 41511 20774 41520
rect 20732 38554 20760 41511
rect 20824 40905 20852 48232
rect 21272 47592 21324 47598
rect 21272 47534 21324 47540
rect 20956 47356 21252 47376
rect 21012 47354 21036 47356
rect 21092 47354 21116 47356
rect 21172 47354 21196 47356
rect 21034 47302 21036 47354
rect 21098 47302 21110 47354
rect 21172 47302 21174 47354
rect 21012 47300 21036 47302
rect 21092 47300 21116 47302
rect 21172 47300 21196 47302
rect 20956 47280 21252 47300
rect 20996 47116 21048 47122
rect 20996 47058 21048 47064
rect 21008 46442 21036 47058
rect 20996 46436 21048 46442
rect 20996 46378 21048 46384
rect 20956 46268 21252 46288
rect 21012 46266 21036 46268
rect 21092 46266 21116 46268
rect 21172 46266 21196 46268
rect 21034 46214 21036 46266
rect 21098 46214 21110 46266
rect 21172 46214 21174 46266
rect 21012 46212 21036 46214
rect 21092 46212 21116 46214
rect 21172 46212 21196 46214
rect 20956 46192 21252 46212
rect 21088 46028 21140 46034
rect 21088 45970 21140 45976
rect 20904 45824 20956 45830
rect 20904 45766 20956 45772
rect 20916 45422 20944 45766
rect 21100 45626 21128 45970
rect 21088 45620 21140 45626
rect 21088 45562 21140 45568
rect 20904 45416 20956 45422
rect 20904 45358 20956 45364
rect 20956 45180 21252 45200
rect 21012 45178 21036 45180
rect 21092 45178 21116 45180
rect 21172 45178 21196 45180
rect 21034 45126 21036 45178
rect 21098 45126 21110 45178
rect 21172 45126 21174 45178
rect 21012 45124 21036 45126
rect 21092 45124 21116 45126
rect 21172 45124 21196 45126
rect 20956 45104 21252 45124
rect 21284 45014 21312 47534
rect 21272 45008 21324 45014
rect 21272 44950 21324 44956
rect 20904 44872 20956 44878
rect 21180 44872 21232 44878
rect 20904 44814 20956 44820
rect 21178 44840 21180 44849
rect 21232 44840 21234 44849
rect 20916 44538 20944 44814
rect 21178 44775 21234 44784
rect 20904 44532 20956 44538
rect 20904 44474 20956 44480
rect 21192 44402 21220 44775
rect 21180 44396 21232 44402
rect 21180 44338 21232 44344
rect 20956 44092 21252 44112
rect 21012 44090 21036 44092
rect 21092 44090 21116 44092
rect 21172 44090 21196 44092
rect 21034 44038 21036 44090
rect 21098 44038 21110 44090
rect 21172 44038 21174 44090
rect 21012 44036 21036 44038
rect 21092 44036 21116 44038
rect 21172 44036 21196 44038
rect 20956 44016 21252 44036
rect 21086 43888 21142 43897
rect 21086 43823 21088 43832
rect 21140 43823 21142 43832
rect 21088 43794 21140 43800
rect 21100 43450 21128 43794
rect 21088 43444 21140 43450
rect 21088 43386 21140 43392
rect 21272 43308 21324 43314
rect 21272 43250 21324 43256
rect 20956 43004 21252 43024
rect 21012 43002 21036 43004
rect 21092 43002 21116 43004
rect 21172 43002 21196 43004
rect 21034 42950 21036 43002
rect 21098 42950 21110 43002
rect 21172 42950 21174 43002
rect 21012 42948 21036 42950
rect 21092 42948 21116 42950
rect 21172 42948 21196 42950
rect 20956 42928 21252 42948
rect 21284 42906 21312 43250
rect 21272 42900 21324 42906
rect 21272 42842 21324 42848
rect 21272 42356 21324 42362
rect 21272 42298 21324 42304
rect 20956 41916 21252 41936
rect 21012 41914 21036 41916
rect 21092 41914 21116 41916
rect 21172 41914 21196 41916
rect 21034 41862 21036 41914
rect 21098 41862 21110 41914
rect 21172 41862 21174 41914
rect 21012 41860 21036 41862
rect 21092 41860 21116 41862
rect 21172 41860 21196 41862
rect 20956 41840 21252 41860
rect 21284 41682 21312 42298
rect 21272 41676 21324 41682
rect 21272 41618 21324 41624
rect 21178 41168 21234 41177
rect 21178 41103 21180 41112
rect 21232 41103 21234 41112
rect 21180 41074 21232 41080
rect 20810 40896 20866 40905
rect 20810 40831 20866 40840
rect 20956 40828 21252 40848
rect 21012 40826 21036 40828
rect 21092 40826 21116 40828
rect 21172 40826 21196 40828
rect 21034 40774 21036 40826
rect 21098 40774 21110 40826
rect 21172 40774 21174 40826
rect 21012 40772 21036 40774
rect 21092 40772 21116 40774
rect 21172 40772 21196 40774
rect 20956 40752 21252 40772
rect 21284 40730 21312 41618
rect 21272 40724 21324 40730
rect 21272 40666 21324 40672
rect 20996 40588 21048 40594
rect 20996 40530 21048 40536
rect 21008 39914 21036 40530
rect 20996 39908 21048 39914
rect 20996 39850 21048 39856
rect 20956 39740 21252 39760
rect 21012 39738 21036 39740
rect 21092 39738 21116 39740
rect 21172 39738 21196 39740
rect 21034 39686 21036 39738
rect 21098 39686 21110 39738
rect 21172 39686 21174 39738
rect 21012 39684 21036 39686
rect 21092 39684 21116 39686
rect 21172 39684 21196 39686
rect 20956 39664 21252 39684
rect 21178 39536 21234 39545
rect 21178 39471 21234 39480
rect 21192 38894 21220 39471
rect 21180 38888 21232 38894
rect 21180 38830 21232 38836
rect 20956 38652 21252 38672
rect 21012 38650 21036 38652
rect 21092 38650 21116 38652
rect 21172 38650 21196 38652
rect 21034 38598 21036 38650
rect 21098 38598 21110 38650
rect 21172 38598 21174 38650
rect 21012 38596 21036 38598
rect 21092 38596 21116 38598
rect 21172 38596 21196 38598
rect 20956 38576 21252 38596
rect 21376 38570 21404 51462
rect 21548 51410 21600 51416
rect 21548 51332 21600 51338
rect 21548 51274 21600 51280
rect 21456 50992 21508 50998
rect 21456 50934 21508 50940
rect 21468 50522 21496 50934
rect 21560 50794 21588 51274
rect 21548 50788 21600 50794
rect 21548 50730 21600 50736
rect 21456 50516 21508 50522
rect 21456 50458 21508 50464
rect 21468 50017 21496 50458
rect 21560 50289 21588 50730
rect 21546 50280 21602 50289
rect 21546 50215 21602 50224
rect 21548 50176 21600 50182
rect 21546 50144 21548 50153
rect 21600 50144 21602 50153
rect 21546 50079 21602 50088
rect 21454 50008 21510 50017
rect 21454 49943 21510 49952
rect 21468 49706 21496 49943
rect 21456 49700 21508 49706
rect 21456 49642 21508 49648
rect 21652 49586 21680 55014
rect 21744 52850 21772 56902
rect 21824 56840 21876 56846
rect 21824 56782 21876 56788
rect 21836 54874 21864 56782
rect 22100 56160 22152 56166
rect 22204 56148 22232 59366
rect 22152 56120 22232 56148
rect 22100 56102 22152 56108
rect 22112 55593 22140 56102
rect 22098 55584 22154 55593
rect 22098 55519 22154 55528
rect 22008 55208 22060 55214
rect 22008 55150 22060 55156
rect 21916 55072 21968 55078
rect 21916 55014 21968 55020
rect 21824 54868 21876 54874
rect 21824 54810 21876 54816
rect 21928 54738 21956 55014
rect 21824 54732 21876 54738
rect 21824 54674 21876 54680
rect 21916 54732 21968 54738
rect 21916 54674 21968 54680
rect 21836 53786 21864 54674
rect 21928 54330 21956 54674
rect 21916 54324 21968 54330
rect 21916 54266 21968 54272
rect 21824 53780 21876 53786
rect 21824 53722 21876 53728
rect 21836 53446 21864 53722
rect 21824 53440 21876 53446
rect 21824 53382 21876 53388
rect 21916 53032 21968 53038
rect 21916 52974 21968 52980
rect 21744 52822 21864 52850
rect 21732 52624 21784 52630
rect 21732 52566 21784 52572
rect 21744 52494 21772 52566
rect 21732 52488 21784 52494
rect 21732 52430 21784 52436
rect 21744 51950 21772 52430
rect 21732 51944 21784 51950
rect 21732 51886 21784 51892
rect 21732 51808 21784 51814
rect 21732 51750 21784 51756
rect 21744 51542 21772 51750
rect 21732 51536 21784 51542
rect 21732 51478 21784 51484
rect 21732 51264 21784 51270
rect 21732 51206 21784 51212
rect 21468 49558 21680 49586
rect 21468 48686 21496 49558
rect 21640 49156 21692 49162
rect 21560 49116 21640 49144
rect 21456 48680 21508 48686
rect 21456 48622 21508 48628
rect 21456 48544 21508 48550
rect 21456 48486 21508 48492
rect 21468 47598 21496 48486
rect 21560 48278 21588 49116
rect 21640 49098 21692 49104
rect 21638 49056 21694 49065
rect 21638 48991 21694 49000
rect 21548 48272 21600 48278
rect 21548 48214 21600 48220
rect 21548 48136 21600 48142
rect 21546 48104 21548 48113
rect 21600 48104 21602 48113
rect 21546 48039 21602 48048
rect 21548 48000 21600 48006
rect 21546 47968 21548 47977
rect 21600 47968 21602 47977
rect 21546 47903 21602 47912
rect 21652 47598 21680 48991
rect 21456 47592 21508 47598
rect 21456 47534 21508 47540
rect 21640 47592 21692 47598
rect 21640 47534 21692 47540
rect 21548 47456 21600 47462
rect 21548 47398 21600 47404
rect 21456 46912 21508 46918
rect 21456 46854 21508 46860
rect 20720 38548 20772 38554
rect 20720 38490 20772 38496
rect 21284 38542 21404 38570
rect 20732 37806 20760 38490
rect 20812 37868 20864 37874
rect 20812 37810 20864 37816
rect 20720 37800 20772 37806
rect 20720 37742 20772 37748
rect 20720 36712 20772 36718
rect 20720 36654 20772 36660
rect 20732 36378 20760 36654
rect 20720 36372 20772 36378
rect 20720 36314 20772 36320
rect 20720 36168 20772 36174
rect 20720 36110 20772 36116
rect 20364 35788 20668 35816
rect 20260 34536 20312 34542
rect 20260 34478 20312 34484
rect 20272 32745 20300 34478
rect 20364 33522 20392 35788
rect 20626 35728 20682 35737
rect 20626 35663 20682 35672
rect 20536 35556 20588 35562
rect 20536 35498 20588 35504
rect 20548 35290 20576 35498
rect 20536 35284 20588 35290
rect 20536 35226 20588 35232
rect 20444 35216 20496 35222
rect 20444 35158 20496 35164
rect 20352 33516 20404 33522
rect 20352 33458 20404 33464
rect 20456 33454 20484 35158
rect 20548 34610 20576 35226
rect 20536 34604 20588 34610
rect 20536 34546 20588 34552
rect 20640 33658 20668 35663
rect 20732 35494 20760 36110
rect 20720 35488 20772 35494
rect 20720 35430 20772 35436
rect 20732 34474 20760 35430
rect 20720 34468 20772 34474
rect 20720 34410 20772 34416
rect 20824 34202 20852 37810
rect 20956 37564 21252 37584
rect 21012 37562 21036 37564
rect 21092 37562 21116 37564
rect 21172 37562 21196 37564
rect 21034 37510 21036 37562
rect 21098 37510 21110 37562
rect 21172 37510 21174 37562
rect 21012 37508 21036 37510
rect 21092 37508 21116 37510
rect 21172 37508 21196 37510
rect 20956 37488 21252 37508
rect 20956 36476 21252 36496
rect 21012 36474 21036 36476
rect 21092 36474 21116 36476
rect 21172 36474 21196 36476
rect 21034 36422 21036 36474
rect 21098 36422 21110 36474
rect 21172 36422 21174 36474
rect 21012 36420 21036 36422
rect 21092 36420 21116 36422
rect 21172 36420 21196 36422
rect 20956 36400 21252 36420
rect 21180 36236 21232 36242
rect 21180 36178 21232 36184
rect 21192 36038 21220 36178
rect 21180 36032 21232 36038
rect 21180 35974 21232 35980
rect 21192 35737 21220 35974
rect 21178 35728 21234 35737
rect 21178 35663 21234 35672
rect 20956 35388 21252 35408
rect 21012 35386 21036 35388
rect 21092 35386 21116 35388
rect 21172 35386 21196 35388
rect 21034 35334 21036 35386
rect 21098 35334 21110 35386
rect 21172 35334 21174 35386
rect 21012 35332 21036 35334
rect 21092 35332 21116 35334
rect 21172 35332 21196 35334
rect 20956 35312 21252 35332
rect 20902 35184 20958 35193
rect 20902 35119 20958 35128
rect 20916 34474 20944 35119
rect 20904 34468 20956 34474
rect 20904 34410 20956 34416
rect 20956 34300 21252 34320
rect 21012 34298 21036 34300
rect 21092 34298 21116 34300
rect 21172 34298 21196 34300
rect 21034 34246 21036 34298
rect 21098 34246 21110 34298
rect 21172 34246 21174 34298
rect 21012 34244 21036 34246
rect 21092 34244 21116 34246
rect 21172 34244 21196 34246
rect 20956 34224 21252 34244
rect 20812 34196 20864 34202
rect 20864 34156 20944 34184
rect 20812 34138 20864 34144
rect 20810 34096 20866 34105
rect 20720 34060 20772 34066
rect 20810 34031 20866 34040
rect 20720 34002 20772 34008
rect 20732 33862 20760 34002
rect 20824 33998 20852 34031
rect 20812 33992 20864 33998
rect 20812 33934 20864 33940
rect 20720 33856 20772 33862
rect 20720 33798 20772 33804
rect 20628 33652 20680 33658
rect 20628 33594 20680 33600
rect 20628 33516 20680 33522
rect 20628 33458 20680 33464
rect 20444 33448 20496 33454
rect 20444 33390 20496 33396
rect 20352 33380 20404 33386
rect 20352 33322 20404 33328
rect 20258 32736 20314 32745
rect 20258 32671 20314 32680
rect 20258 32464 20314 32473
rect 20258 32399 20314 32408
rect 20272 30326 20300 32399
rect 20260 30320 20312 30326
rect 20260 30262 20312 30268
rect 20364 29832 20392 33322
rect 20456 33289 20484 33390
rect 20442 33280 20498 33289
rect 20442 33215 20498 33224
rect 20442 33144 20498 33153
rect 20442 33079 20498 33088
rect 20456 32026 20484 33079
rect 20536 32768 20588 32774
rect 20536 32710 20588 32716
rect 20444 32020 20496 32026
rect 20444 31962 20496 31968
rect 20548 31521 20576 32710
rect 20534 31512 20590 31521
rect 20534 31447 20590 31456
rect 20548 31278 20576 31447
rect 20536 31272 20588 31278
rect 20536 31214 20588 31220
rect 20272 29804 20392 29832
rect 20272 24857 20300 29804
rect 20352 29708 20404 29714
rect 20352 29650 20404 29656
rect 20364 28762 20392 29650
rect 20352 28756 20404 28762
rect 20352 28698 20404 28704
rect 20364 28218 20392 28698
rect 20352 28212 20404 28218
rect 20352 28154 20404 28160
rect 20258 24848 20314 24857
rect 20258 24783 20314 24792
rect 20166 19544 20222 19553
rect 20166 19479 20222 19488
rect 19708 16244 19760 16250
rect 19708 16186 19760 16192
rect 20640 14550 20668 33458
rect 20732 31958 20760 33798
rect 20824 33368 20852 33934
rect 20916 33522 20944 34156
rect 20904 33516 20956 33522
rect 20904 33458 20956 33464
rect 20904 33380 20956 33386
rect 20824 33340 20904 33368
rect 20824 33114 20852 33340
rect 20904 33322 20956 33328
rect 20956 33212 21252 33232
rect 21012 33210 21036 33212
rect 21092 33210 21116 33212
rect 21172 33210 21196 33212
rect 21034 33158 21036 33210
rect 21098 33158 21110 33210
rect 21172 33158 21174 33210
rect 21012 33156 21036 33158
rect 21092 33156 21116 33158
rect 21172 33156 21196 33158
rect 20956 33136 21252 33156
rect 20812 33108 20864 33114
rect 20812 33050 20864 33056
rect 21180 32904 21232 32910
rect 21180 32846 21232 32852
rect 21192 32570 21220 32846
rect 21180 32564 21232 32570
rect 21180 32506 21232 32512
rect 20956 32124 21252 32144
rect 21012 32122 21036 32124
rect 21092 32122 21116 32124
rect 21172 32122 21196 32124
rect 21034 32070 21036 32122
rect 21098 32070 21110 32122
rect 21172 32070 21174 32122
rect 21012 32068 21036 32070
rect 21092 32068 21116 32070
rect 21172 32068 21196 32070
rect 20956 32048 21252 32068
rect 20720 31952 20772 31958
rect 20720 31894 20772 31900
rect 20812 31816 20864 31822
rect 20812 31758 20864 31764
rect 20824 31278 20852 31758
rect 21180 31680 21232 31686
rect 21180 31622 21232 31628
rect 20902 31376 20958 31385
rect 20902 31311 20958 31320
rect 20916 31278 20944 31311
rect 20812 31272 20864 31278
rect 20812 31214 20864 31220
rect 20904 31272 20956 31278
rect 21192 31249 21220 31622
rect 20904 31214 20956 31220
rect 21178 31240 21234 31249
rect 21178 31175 21234 31184
rect 20810 31104 20866 31113
rect 20810 31039 20866 31048
rect 20718 28656 20774 28665
rect 20718 28591 20774 28600
rect 20732 28150 20760 28591
rect 20720 28144 20772 28150
rect 20720 28086 20772 28092
rect 20720 28008 20772 28014
rect 20720 27950 20772 27956
rect 20732 27606 20760 27950
rect 20824 27606 20852 31039
rect 20956 31036 21252 31056
rect 21012 31034 21036 31036
rect 21092 31034 21116 31036
rect 21172 31034 21196 31036
rect 21034 30982 21036 31034
rect 21098 30982 21110 31034
rect 21172 30982 21174 31034
rect 21012 30980 21036 30982
rect 21092 30980 21116 30982
rect 21172 30980 21196 30982
rect 20956 30960 21252 30980
rect 20902 30832 20958 30841
rect 20902 30767 20904 30776
rect 20956 30767 20958 30776
rect 20904 30738 20956 30744
rect 20916 30394 20944 30738
rect 21086 30696 21142 30705
rect 21086 30631 21088 30640
rect 21140 30631 21142 30640
rect 21088 30602 21140 30608
rect 20904 30388 20956 30394
rect 20904 30330 20956 30336
rect 20956 29948 21252 29968
rect 21012 29946 21036 29948
rect 21092 29946 21116 29948
rect 21172 29946 21196 29948
rect 21034 29894 21036 29946
rect 21098 29894 21110 29946
rect 21172 29894 21174 29946
rect 21012 29892 21036 29894
rect 21092 29892 21116 29894
rect 21172 29892 21196 29894
rect 20956 29872 21252 29892
rect 20994 29472 21050 29481
rect 20994 29407 21050 29416
rect 21008 29306 21036 29407
rect 20996 29300 21048 29306
rect 20996 29242 21048 29248
rect 20956 28860 21252 28880
rect 21012 28858 21036 28860
rect 21092 28858 21116 28860
rect 21172 28858 21196 28860
rect 21034 28806 21036 28858
rect 21098 28806 21110 28858
rect 21172 28806 21174 28858
rect 21012 28804 21036 28806
rect 21092 28804 21116 28806
rect 21172 28804 21196 28806
rect 20956 28784 21252 28804
rect 20956 27772 21252 27792
rect 21012 27770 21036 27772
rect 21092 27770 21116 27772
rect 21172 27770 21196 27772
rect 21034 27718 21036 27770
rect 21098 27718 21110 27770
rect 21172 27718 21174 27770
rect 21012 27716 21036 27718
rect 21092 27716 21116 27718
rect 21172 27716 21196 27718
rect 20956 27696 21252 27716
rect 20720 27600 20772 27606
rect 20720 27542 20772 27548
rect 20812 27600 20864 27606
rect 20812 27542 20864 27548
rect 20812 27464 20864 27470
rect 20732 27424 20812 27452
rect 20444 14544 20496 14550
rect 20444 14486 20496 14492
rect 20628 14544 20680 14550
rect 20628 14486 20680 14492
rect 20456 10554 20484 14486
rect 20536 13388 20588 13394
rect 20536 13330 20588 13336
rect 20548 10674 20576 13330
rect 20536 10668 20588 10674
rect 20536 10610 20588 10616
rect 20456 10526 20668 10554
rect 20536 9648 20588 9654
rect 20536 9590 20588 9596
rect 19352 2604 19656 2632
rect 18604 2440 18656 2446
rect 18604 2382 18656 2388
rect 18616 2009 18644 2382
rect 18602 2000 18658 2009
rect 18602 1935 18658 1944
rect 19352 800 19380 2604
rect 20260 2372 20312 2378
rect 20260 2314 20312 2320
rect 20272 800 20300 2314
rect 20548 921 20576 9590
rect 20640 2378 20668 10526
rect 20732 9654 20760 27424
rect 20812 27406 20864 27412
rect 20956 26684 21252 26704
rect 21012 26682 21036 26684
rect 21092 26682 21116 26684
rect 21172 26682 21196 26684
rect 21034 26630 21036 26682
rect 21098 26630 21110 26682
rect 21172 26630 21174 26682
rect 21012 26628 21036 26630
rect 21092 26628 21116 26630
rect 21172 26628 21196 26630
rect 20956 26608 21252 26628
rect 20956 25596 21252 25616
rect 21012 25594 21036 25596
rect 21092 25594 21116 25596
rect 21172 25594 21196 25596
rect 21034 25542 21036 25594
rect 21098 25542 21110 25594
rect 21172 25542 21174 25594
rect 21012 25540 21036 25542
rect 21092 25540 21116 25542
rect 21172 25540 21196 25542
rect 20956 25520 21252 25540
rect 20956 24508 21252 24528
rect 21012 24506 21036 24508
rect 21092 24506 21116 24508
rect 21172 24506 21196 24508
rect 21034 24454 21036 24506
rect 21098 24454 21110 24506
rect 21172 24454 21174 24506
rect 21012 24452 21036 24454
rect 21092 24452 21116 24454
rect 21172 24452 21196 24454
rect 20956 24432 21252 24452
rect 20956 23420 21252 23440
rect 21012 23418 21036 23420
rect 21092 23418 21116 23420
rect 21172 23418 21196 23420
rect 21034 23366 21036 23418
rect 21098 23366 21110 23418
rect 21172 23366 21174 23418
rect 21012 23364 21036 23366
rect 21092 23364 21116 23366
rect 21172 23364 21196 23366
rect 20956 23344 21252 23364
rect 21284 22778 21312 38542
rect 21364 34060 21416 34066
rect 21364 34002 21416 34008
rect 21376 33318 21404 34002
rect 21364 33312 21416 33318
rect 21364 33254 21416 33260
rect 21364 32768 21416 32774
rect 21364 32710 21416 32716
rect 21272 22772 21324 22778
rect 21272 22714 21324 22720
rect 20956 22332 21252 22352
rect 21012 22330 21036 22332
rect 21092 22330 21116 22332
rect 21172 22330 21196 22332
rect 21034 22278 21036 22330
rect 21098 22278 21110 22330
rect 21172 22278 21174 22330
rect 21012 22276 21036 22278
rect 21092 22276 21116 22278
rect 21172 22276 21196 22278
rect 20956 22256 21252 22276
rect 20956 21244 21252 21264
rect 21012 21242 21036 21244
rect 21092 21242 21116 21244
rect 21172 21242 21196 21244
rect 21034 21190 21036 21242
rect 21098 21190 21110 21242
rect 21172 21190 21174 21242
rect 21012 21188 21036 21190
rect 21092 21188 21116 21190
rect 21172 21188 21196 21190
rect 20956 21168 21252 21188
rect 20956 20156 21252 20176
rect 21012 20154 21036 20156
rect 21092 20154 21116 20156
rect 21172 20154 21196 20156
rect 21034 20102 21036 20154
rect 21098 20102 21110 20154
rect 21172 20102 21174 20154
rect 21012 20100 21036 20102
rect 21092 20100 21116 20102
rect 21172 20100 21196 20102
rect 20956 20080 21252 20100
rect 21178 19544 21234 19553
rect 21178 19479 21234 19488
rect 21192 19224 21220 19479
rect 21192 19196 21312 19224
rect 20956 19068 21252 19088
rect 21012 19066 21036 19068
rect 21092 19066 21116 19068
rect 21172 19066 21196 19068
rect 21034 19014 21036 19066
rect 21098 19014 21110 19066
rect 21172 19014 21174 19066
rect 21012 19012 21036 19014
rect 21092 19012 21116 19014
rect 21172 19012 21196 19014
rect 20956 18992 21252 19012
rect 20956 17980 21252 18000
rect 21012 17978 21036 17980
rect 21092 17978 21116 17980
rect 21172 17978 21196 17980
rect 21034 17926 21036 17978
rect 21098 17926 21110 17978
rect 21172 17926 21174 17978
rect 21012 17924 21036 17926
rect 21092 17924 21116 17926
rect 21172 17924 21196 17926
rect 20956 17904 21252 17924
rect 20956 16892 21252 16912
rect 21012 16890 21036 16892
rect 21092 16890 21116 16892
rect 21172 16890 21196 16892
rect 21034 16838 21036 16890
rect 21098 16838 21110 16890
rect 21172 16838 21174 16890
rect 21012 16836 21036 16838
rect 21092 16836 21116 16838
rect 21172 16836 21196 16838
rect 20956 16816 21252 16836
rect 20956 15804 21252 15824
rect 21012 15802 21036 15804
rect 21092 15802 21116 15804
rect 21172 15802 21196 15804
rect 21034 15750 21036 15802
rect 21098 15750 21110 15802
rect 21172 15750 21174 15802
rect 21012 15748 21036 15750
rect 21092 15748 21116 15750
rect 21172 15748 21196 15750
rect 20956 15728 21252 15748
rect 20956 14716 21252 14736
rect 21012 14714 21036 14716
rect 21092 14714 21116 14716
rect 21172 14714 21196 14716
rect 21034 14662 21036 14714
rect 21098 14662 21110 14714
rect 21172 14662 21174 14714
rect 21012 14660 21036 14662
rect 21092 14660 21116 14662
rect 21172 14660 21196 14662
rect 20956 14640 21252 14660
rect 20956 13628 21252 13648
rect 21012 13626 21036 13628
rect 21092 13626 21116 13628
rect 21172 13626 21196 13628
rect 21034 13574 21036 13626
rect 21098 13574 21110 13626
rect 21172 13574 21174 13626
rect 21012 13572 21036 13574
rect 21092 13572 21116 13574
rect 21172 13572 21196 13574
rect 20956 13552 21252 13572
rect 21284 12782 21312 19196
rect 21272 12776 21324 12782
rect 21272 12718 21324 12724
rect 20956 12540 21252 12560
rect 21012 12538 21036 12540
rect 21092 12538 21116 12540
rect 21172 12538 21196 12540
rect 21034 12486 21036 12538
rect 21098 12486 21110 12538
rect 21172 12486 21174 12538
rect 21012 12484 21036 12486
rect 21092 12484 21116 12486
rect 21172 12484 21196 12486
rect 20956 12464 21252 12484
rect 20956 11452 21252 11472
rect 21012 11450 21036 11452
rect 21092 11450 21116 11452
rect 21172 11450 21196 11452
rect 21034 11398 21036 11450
rect 21098 11398 21110 11450
rect 21172 11398 21174 11450
rect 21012 11396 21036 11398
rect 21092 11396 21116 11398
rect 21172 11396 21196 11398
rect 20956 11376 21252 11396
rect 21376 10810 21404 32710
rect 21468 20233 21496 46854
rect 21560 45082 21588 47398
rect 21652 47258 21680 47534
rect 21640 47252 21692 47258
rect 21640 47194 21692 47200
rect 21640 47116 21692 47122
rect 21640 47058 21692 47064
rect 21652 46424 21680 47058
rect 21744 46918 21772 51206
rect 21836 48804 21864 52822
rect 21928 51474 21956 52974
rect 21916 51468 21968 51474
rect 21916 51410 21968 51416
rect 22020 50930 22048 55150
rect 22192 54120 22244 54126
rect 22190 54088 22192 54097
rect 22244 54088 22246 54097
rect 22190 54023 22246 54032
rect 22100 53440 22152 53446
rect 22100 53382 22152 53388
rect 22112 51542 22140 53382
rect 22192 52964 22244 52970
rect 22192 52906 22244 52912
rect 22204 52358 22232 52906
rect 22192 52352 22244 52358
rect 22192 52294 22244 52300
rect 22100 51536 22152 51542
rect 22100 51478 22152 51484
rect 22100 51400 22152 51406
rect 22100 51342 22152 51348
rect 22112 51066 22140 51342
rect 22100 51060 22152 51066
rect 22100 51002 22152 51008
rect 22008 50924 22060 50930
rect 22008 50866 22060 50872
rect 22006 50824 22062 50833
rect 22006 50759 22008 50768
rect 22060 50759 22062 50768
rect 22008 50730 22060 50736
rect 22296 50538 22324 69663
rect 22468 64932 22520 64938
rect 22468 64874 22520 64880
rect 22376 57860 22428 57866
rect 22376 57802 22428 57808
rect 22388 57594 22416 57802
rect 22376 57588 22428 57594
rect 22376 57530 22428 57536
rect 22376 57384 22428 57390
rect 22376 57326 22428 57332
rect 22388 55944 22416 57326
rect 22480 56545 22508 64874
rect 22664 59129 22692 76230
rect 22756 61849 22784 76842
rect 23492 74610 23520 79200
rect 23848 77376 23900 77382
rect 23848 77318 23900 77324
rect 23664 75336 23716 75342
rect 23664 75278 23716 75284
rect 23676 75002 23704 75278
rect 23664 74996 23716 75002
rect 23664 74938 23716 74944
rect 23662 74760 23718 74769
rect 23662 74695 23718 74704
rect 23400 74582 23520 74610
rect 23110 74352 23166 74361
rect 23110 74287 23166 74296
rect 23124 70990 23152 74287
rect 23202 73808 23258 73817
rect 23202 73743 23258 73752
rect 23112 70984 23164 70990
rect 23112 70926 23164 70932
rect 22926 62384 22982 62393
rect 22926 62319 22982 62328
rect 22742 61840 22798 61849
rect 22742 61775 22798 61784
rect 22836 61192 22888 61198
rect 22836 61134 22888 61140
rect 22848 60858 22876 61134
rect 22836 60852 22888 60858
rect 22836 60794 22888 60800
rect 22940 60178 22968 62319
rect 22744 60172 22796 60178
rect 22744 60114 22796 60120
rect 22928 60172 22980 60178
rect 22928 60114 22980 60120
rect 22756 59430 22784 60114
rect 22836 60104 22888 60110
rect 22836 60046 22888 60052
rect 22848 59702 22876 60046
rect 22836 59696 22888 59702
rect 22836 59638 22888 59644
rect 22744 59424 22796 59430
rect 22744 59366 22796 59372
rect 22650 59120 22706 59129
rect 22650 59055 22706 59064
rect 22560 58472 22612 58478
rect 22560 58414 22612 58420
rect 22572 57798 22600 58414
rect 22560 57792 22612 57798
rect 22558 57760 22560 57769
rect 22612 57760 22614 57769
rect 22558 57695 22614 57704
rect 22756 57610 22784 59366
rect 22848 59090 22876 59638
rect 22836 59084 22888 59090
rect 22836 59026 22888 59032
rect 22848 58682 22876 59026
rect 22836 58676 22888 58682
rect 22836 58618 22888 58624
rect 23112 58132 23164 58138
rect 23112 58074 23164 58080
rect 23020 57792 23072 57798
rect 23020 57734 23072 57740
rect 22572 57582 22784 57610
rect 22466 56536 22522 56545
rect 22466 56471 22522 56480
rect 22480 56234 22508 56471
rect 22468 56228 22520 56234
rect 22468 56170 22520 56176
rect 22388 55916 22508 55944
rect 22376 55820 22428 55826
rect 22376 55762 22428 55768
rect 22388 55350 22416 55762
rect 22376 55344 22428 55350
rect 22376 55286 22428 55292
rect 22388 54874 22416 55286
rect 22376 54868 22428 54874
rect 22376 54810 22428 54816
rect 22376 54120 22428 54126
rect 22376 54062 22428 54068
rect 22388 53802 22416 54062
rect 22480 53990 22508 55916
rect 22468 53984 22520 53990
rect 22468 53926 22520 53932
rect 22572 53802 22600 57582
rect 22744 56908 22796 56914
rect 22744 56850 22796 56856
rect 22756 56166 22784 56850
rect 23032 56506 23060 57734
rect 23020 56500 23072 56506
rect 23020 56442 23072 56448
rect 22836 56228 22888 56234
rect 22836 56170 22888 56176
rect 22744 56160 22796 56166
rect 22744 56102 22796 56108
rect 22756 55894 22784 56102
rect 22744 55888 22796 55894
rect 22744 55830 22796 55836
rect 22744 55752 22796 55758
rect 22744 55694 22796 55700
rect 22652 55616 22704 55622
rect 22652 55558 22704 55564
rect 22664 55282 22692 55558
rect 22652 55276 22704 55282
rect 22652 55218 22704 55224
rect 22664 54126 22692 55218
rect 22756 55049 22784 55694
rect 22742 55040 22798 55049
rect 22742 54975 22798 54984
rect 22652 54120 22704 54126
rect 22652 54062 22704 54068
rect 22388 53786 22600 53802
rect 22376 53780 22600 53786
rect 22428 53774 22600 53780
rect 22376 53722 22428 53728
rect 22466 53680 22522 53689
rect 22466 53615 22522 53624
rect 22376 53576 22428 53582
rect 22376 53518 22428 53524
rect 22112 50510 22324 50538
rect 22008 50448 22060 50454
rect 22006 50416 22008 50425
rect 22060 50416 22062 50425
rect 22006 50351 22062 50360
rect 22008 50312 22060 50318
rect 22006 50280 22008 50289
rect 22060 50280 22062 50289
rect 22006 50215 22062 50224
rect 22008 49904 22060 49910
rect 22008 49846 22060 49852
rect 22020 49745 22048 49846
rect 22006 49736 22062 49745
rect 22006 49671 22062 49680
rect 21916 49360 21968 49366
rect 21916 49302 21968 49308
rect 21928 48906 21956 49302
rect 22112 49280 22140 50510
rect 22192 50380 22244 50386
rect 22192 50322 22244 50328
rect 22204 49978 22232 50322
rect 22284 50176 22336 50182
rect 22284 50118 22336 50124
rect 22192 49972 22244 49978
rect 22192 49914 22244 49920
rect 22204 49881 22232 49914
rect 22190 49872 22246 49881
rect 22190 49807 22246 49816
rect 22112 49252 22232 49280
rect 22100 49156 22152 49162
rect 22020 49116 22100 49144
rect 22020 49065 22048 49116
rect 22100 49098 22152 49104
rect 22006 49056 22062 49065
rect 22006 48991 22062 49000
rect 21928 48878 22140 48906
rect 21836 48776 21956 48804
rect 21822 48512 21878 48521
rect 21822 48447 21878 48456
rect 21732 46912 21784 46918
rect 21732 46854 21784 46860
rect 21732 46640 21784 46646
rect 21730 46608 21732 46617
rect 21784 46608 21786 46617
rect 21730 46543 21786 46552
rect 21652 46396 21772 46424
rect 21744 46073 21772 46396
rect 21836 46209 21864 48447
rect 21822 46200 21878 46209
rect 21822 46135 21878 46144
rect 21730 46064 21786 46073
rect 21730 45999 21786 46008
rect 21744 45948 21772 45999
rect 21744 45920 21864 45948
rect 21732 45280 21784 45286
rect 21732 45222 21784 45228
rect 21548 45076 21600 45082
rect 21548 45018 21600 45024
rect 21548 44940 21600 44946
rect 21548 44882 21600 44888
rect 21560 41177 21588 44882
rect 21640 43920 21692 43926
rect 21640 43862 21692 43868
rect 21652 42362 21680 43862
rect 21744 42838 21772 45222
rect 21836 44266 21864 45920
rect 21824 44260 21876 44266
rect 21824 44202 21876 44208
rect 21732 42832 21784 42838
rect 21732 42774 21784 42780
rect 21640 42356 21692 42362
rect 21640 42298 21692 42304
rect 21640 42220 21692 42226
rect 21640 42162 21692 42168
rect 21652 41206 21680 42162
rect 21640 41200 21692 41206
rect 21546 41168 21602 41177
rect 21640 41142 21692 41148
rect 21546 41103 21602 41112
rect 21548 41064 21600 41070
rect 21548 41006 21600 41012
rect 21640 41064 21692 41070
rect 21640 41006 21692 41012
rect 21560 40730 21588 41006
rect 21548 40724 21600 40730
rect 21548 40666 21600 40672
rect 21560 39953 21588 40666
rect 21652 40594 21680 41006
rect 21640 40588 21692 40594
rect 21640 40530 21692 40536
rect 21652 40186 21680 40530
rect 21640 40180 21692 40186
rect 21640 40122 21692 40128
rect 21546 39944 21602 39953
rect 21744 39930 21772 42774
rect 21824 42152 21876 42158
rect 21824 42094 21876 42100
rect 21836 41818 21864 42094
rect 21824 41812 21876 41818
rect 21824 41754 21876 41760
rect 21836 41070 21864 41754
rect 21928 41313 21956 48776
rect 22008 48680 22060 48686
rect 22008 48622 22060 48628
rect 22020 47122 22048 48622
rect 22008 47116 22060 47122
rect 22008 47058 22060 47064
rect 22008 46912 22060 46918
rect 22008 46854 22060 46860
rect 22020 45422 22048 46854
rect 22112 46646 22140 48878
rect 22204 48113 22232 49252
rect 22296 48249 22324 50118
rect 22388 49858 22416 53518
rect 22480 52154 22508 53615
rect 22560 52896 22612 52902
rect 22560 52838 22612 52844
rect 22572 52562 22600 52838
rect 22560 52556 22612 52562
rect 22560 52498 22612 52504
rect 22468 52148 22520 52154
rect 22468 52090 22520 52096
rect 22480 50454 22508 52090
rect 22572 50930 22600 52498
rect 22560 50924 22612 50930
rect 22560 50866 22612 50872
rect 22664 50810 22692 54062
rect 22744 53168 22796 53174
rect 22744 53110 22796 53116
rect 22572 50782 22692 50810
rect 22468 50448 22520 50454
rect 22468 50390 22520 50396
rect 22480 49978 22508 50390
rect 22468 49972 22520 49978
rect 22468 49914 22520 49920
rect 22388 49830 22508 49858
rect 22572 49842 22600 50782
rect 22756 50726 22784 53110
rect 22744 50720 22796 50726
rect 22744 50662 22796 50668
rect 22848 50538 22876 56170
rect 23124 55418 23152 58074
rect 23112 55412 23164 55418
rect 23112 55354 23164 55360
rect 23124 55214 23152 55354
rect 23112 55208 23164 55214
rect 23112 55150 23164 55156
rect 23216 54806 23244 73743
rect 23400 71126 23428 74582
rect 23388 71120 23440 71126
rect 23388 71062 23440 71068
rect 23388 70984 23440 70990
rect 23388 70926 23440 70932
rect 23296 59016 23348 59022
rect 23296 58958 23348 58964
rect 23308 58682 23336 58958
rect 23296 58676 23348 58682
rect 23296 58618 23348 58624
rect 23296 58472 23348 58478
rect 23296 58414 23348 58420
rect 23308 57050 23336 58414
rect 23296 57044 23348 57050
rect 23296 56986 23348 56992
rect 23296 56704 23348 56710
rect 23296 56646 23348 56652
rect 23204 54800 23256 54806
rect 23204 54742 23256 54748
rect 23112 54664 23164 54670
rect 23112 54606 23164 54612
rect 23124 54058 23152 54606
rect 23112 54052 23164 54058
rect 23112 53994 23164 54000
rect 23020 53984 23072 53990
rect 23020 53926 23072 53932
rect 22926 51232 22982 51241
rect 22926 51167 22982 51176
rect 22664 50510 22876 50538
rect 22376 49632 22428 49638
rect 22376 49574 22428 49580
rect 22388 49298 22416 49574
rect 22376 49292 22428 49298
rect 22376 49234 22428 49240
rect 22388 48890 22416 49234
rect 22376 48884 22428 48890
rect 22376 48826 22428 48832
rect 22480 48770 22508 49830
rect 22560 49836 22612 49842
rect 22560 49778 22612 49784
rect 22560 49292 22612 49298
rect 22560 49234 22612 49240
rect 22388 48742 22508 48770
rect 22282 48240 22338 48249
rect 22282 48175 22338 48184
rect 22190 48104 22246 48113
rect 22190 48039 22246 48048
rect 22100 46640 22152 46646
rect 22100 46582 22152 46588
rect 22204 46374 22232 48039
rect 22388 46889 22416 48742
rect 22468 48680 22520 48686
rect 22468 48622 22520 48628
rect 22480 47190 22508 48622
rect 22572 48346 22600 49234
rect 22560 48340 22612 48346
rect 22560 48282 22612 48288
rect 22664 48249 22692 50510
rect 22836 50448 22888 50454
rect 22836 50390 22888 50396
rect 22744 50380 22796 50386
rect 22744 50322 22796 50328
rect 22756 49978 22784 50322
rect 22744 49972 22796 49978
rect 22744 49914 22796 49920
rect 22744 49836 22796 49842
rect 22744 49778 22796 49784
rect 22650 48240 22706 48249
rect 22650 48175 22652 48184
rect 22704 48175 22706 48184
rect 22652 48146 22704 48152
rect 22664 48115 22692 48146
rect 22756 47977 22784 49778
rect 22848 49094 22876 50390
rect 22836 49088 22888 49094
rect 22836 49030 22888 49036
rect 22940 48754 22968 51167
rect 23032 50862 23060 53926
rect 23124 53650 23152 53994
rect 23112 53644 23164 53650
rect 23112 53586 23164 53592
rect 23124 53242 23152 53586
rect 23112 53236 23164 53242
rect 23112 53178 23164 53184
rect 23308 52562 23336 56646
rect 23296 52556 23348 52562
rect 23296 52498 23348 52504
rect 23112 52488 23164 52494
rect 23112 52430 23164 52436
rect 23124 52154 23152 52430
rect 23204 52420 23256 52426
rect 23204 52362 23256 52368
rect 23112 52148 23164 52154
rect 23112 52090 23164 52096
rect 23216 51474 23244 52362
rect 23308 52018 23336 52498
rect 23296 52012 23348 52018
rect 23296 51954 23348 51960
rect 23204 51468 23256 51474
rect 23204 51410 23256 51416
rect 23308 51406 23336 51954
rect 23112 51400 23164 51406
rect 23296 51400 23348 51406
rect 23112 51342 23164 51348
rect 23202 51368 23258 51377
rect 23020 50856 23072 50862
rect 23020 50798 23072 50804
rect 23020 50720 23072 50726
rect 23020 50662 23072 50668
rect 22928 48748 22980 48754
rect 22928 48690 22980 48696
rect 22940 48278 22968 48690
rect 22928 48272 22980 48278
rect 22928 48214 22980 48220
rect 23032 48090 23060 50662
rect 22836 48068 22888 48074
rect 22836 48010 22888 48016
rect 22940 48062 23060 48090
rect 22742 47968 22798 47977
rect 22742 47903 22798 47912
rect 22652 47728 22704 47734
rect 22652 47670 22704 47676
rect 22560 47524 22612 47530
rect 22560 47466 22612 47472
rect 22468 47184 22520 47190
rect 22468 47126 22520 47132
rect 22374 46880 22430 46889
rect 22374 46815 22430 46824
rect 22468 46640 22520 46646
rect 22468 46582 22520 46588
rect 22376 46572 22428 46578
rect 22296 46532 22376 46560
rect 22100 46368 22152 46374
rect 22100 46310 22152 46316
rect 22192 46368 22244 46374
rect 22192 46310 22244 46316
rect 22112 45830 22140 46310
rect 22190 46200 22246 46209
rect 22190 46135 22246 46144
rect 22100 45824 22152 45830
rect 22100 45766 22152 45772
rect 22008 45416 22060 45422
rect 22008 45358 22060 45364
rect 22008 45076 22060 45082
rect 22008 45018 22060 45024
rect 22020 41732 22048 45018
rect 22204 44946 22232 46135
rect 22192 44940 22244 44946
rect 22192 44882 22244 44888
rect 22100 44872 22152 44878
rect 22296 44826 22324 46532
rect 22376 46514 22428 46520
rect 22480 46374 22508 46582
rect 22468 46368 22520 46374
rect 22468 46310 22520 46316
rect 22572 46050 22600 47466
rect 22664 47258 22692 47670
rect 22756 47258 22784 47903
rect 22652 47252 22704 47258
rect 22652 47194 22704 47200
rect 22744 47252 22796 47258
rect 22744 47194 22796 47200
rect 22744 47116 22796 47122
rect 22744 47058 22796 47064
rect 22756 46442 22784 47058
rect 22744 46436 22796 46442
rect 22744 46378 22796 46384
rect 22756 46102 22784 46378
rect 22480 46022 22600 46050
rect 22744 46096 22796 46102
rect 22744 46038 22796 46044
rect 22376 45416 22428 45422
rect 22376 45358 22428 45364
rect 22100 44814 22152 44820
rect 22112 44334 22140 44814
rect 22204 44798 22324 44826
rect 22100 44328 22152 44334
rect 22100 44270 22152 44276
rect 22112 43654 22140 44270
rect 22204 43790 22232 44798
rect 22284 44736 22336 44742
rect 22284 44678 22336 44684
rect 22296 44334 22324 44678
rect 22284 44328 22336 44334
rect 22284 44270 22336 44276
rect 22192 43784 22244 43790
rect 22192 43726 22244 43732
rect 22100 43648 22152 43654
rect 22100 43590 22152 43596
rect 22204 43489 22232 43726
rect 22190 43480 22246 43489
rect 22190 43415 22246 43424
rect 22296 42922 22324 44270
rect 22388 43722 22416 45358
rect 22480 44810 22508 46022
rect 22560 45960 22612 45966
rect 22560 45902 22612 45908
rect 22572 44946 22600 45902
rect 22744 45620 22796 45626
rect 22744 45562 22796 45568
rect 22652 45348 22704 45354
rect 22652 45290 22704 45296
rect 22560 44940 22612 44946
rect 22560 44882 22612 44888
rect 22468 44804 22520 44810
rect 22468 44746 22520 44752
rect 22480 44538 22508 44746
rect 22468 44532 22520 44538
rect 22468 44474 22520 44480
rect 22480 44198 22508 44474
rect 22572 44334 22600 44882
rect 22664 44577 22692 45290
rect 22650 44568 22706 44577
rect 22650 44503 22706 44512
rect 22664 44334 22692 44503
rect 22560 44328 22612 44334
rect 22560 44270 22612 44276
rect 22652 44328 22704 44334
rect 22652 44270 22704 44276
rect 22468 44192 22520 44198
rect 22468 44134 22520 44140
rect 22376 43716 22428 43722
rect 22376 43658 22428 43664
rect 22468 43648 22520 43654
rect 22468 43590 22520 43596
rect 22204 42894 22416 42922
rect 22204 42702 22232 42894
rect 22282 42800 22338 42809
rect 22282 42735 22284 42744
rect 22336 42735 22338 42744
rect 22284 42706 22336 42712
rect 22192 42696 22244 42702
rect 22192 42638 22244 42644
rect 22284 42560 22336 42566
rect 22284 42502 22336 42508
rect 22192 42288 22244 42294
rect 22192 42230 22244 42236
rect 22204 42090 22232 42230
rect 22192 42084 22244 42090
rect 22192 42026 22244 42032
rect 22100 42016 22152 42022
rect 22100 41958 22152 41964
rect 22112 41800 22140 41958
rect 22112 41772 22232 41800
rect 22020 41704 22140 41732
rect 22008 41608 22060 41614
rect 22008 41550 22060 41556
rect 21914 41304 21970 41313
rect 21914 41239 21970 41248
rect 21916 41200 21968 41206
rect 21916 41142 21968 41148
rect 21824 41064 21876 41070
rect 21824 41006 21876 41012
rect 21822 40760 21878 40769
rect 21822 40695 21878 40704
rect 21546 39879 21602 39888
rect 21652 39902 21772 39930
rect 21560 39642 21588 39879
rect 21548 39636 21600 39642
rect 21548 39578 21600 39584
rect 21548 39500 21600 39506
rect 21548 39442 21600 39448
rect 21560 39030 21588 39442
rect 21548 39024 21600 39030
rect 21548 38966 21600 38972
rect 21548 38888 21600 38894
rect 21548 38830 21600 38836
rect 21560 37369 21588 38830
rect 21546 37360 21602 37369
rect 21546 37295 21602 37304
rect 21652 36786 21680 39902
rect 21732 39840 21784 39846
rect 21732 39782 21784 39788
rect 21744 39506 21772 39782
rect 21732 39500 21784 39506
rect 21732 39442 21784 39448
rect 21744 39098 21772 39442
rect 21732 39092 21784 39098
rect 21732 39034 21784 39040
rect 21730 38856 21786 38865
rect 21730 38791 21786 38800
rect 21744 38350 21772 38791
rect 21732 38344 21784 38350
rect 21732 38286 21784 38292
rect 21640 36780 21692 36786
rect 21640 36722 21692 36728
rect 21548 36644 21600 36650
rect 21548 36586 21600 36592
rect 21560 36174 21588 36586
rect 21548 36168 21600 36174
rect 21548 36110 21600 36116
rect 21546 35864 21602 35873
rect 21652 35834 21680 36722
rect 21836 36530 21864 40695
rect 21928 39574 21956 41142
rect 22020 40730 22048 41550
rect 22008 40724 22060 40730
rect 22008 40666 22060 40672
rect 22008 39976 22060 39982
rect 22008 39918 22060 39924
rect 21916 39568 21968 39574
rect 21916 39510 21968 39516
rect 22020 39302 22048 39918
rect 22008 39296 22060 39302
rect 22008 39238 22060 39244
rect 21916 38888 21968 38894
rect 21916 38830 21968 38836
rect 21928 38729 21956 38830
rect 21914 38720 21970 38729
rect 21914 38655 21970 38664
rect 21744 36502 21864 36530
rect 21546 35799 21602 35808
rect 21640 35828 21692 35834
rect 21560 34610 21588 35799
rect 21640 35770 21692 35776
rect 21652 35630 21680 35770
rect 21640 35624 21692 35630
rect 21640 35566 21692 35572
rect 21640 35080 21692 35086
rect 21640 35022 21692 35028
rect 21548 34604 21600 34610
rect 21548 34546 21600 34552
rect 21652 34542 21680 35022
rect 21640 34536 21692 34542
rect 21560 34484 21640 34490
rect 21560 34478 21692 34484
rect 21560 34462 21680 34478
rect 21560 28218 21588 34462
rect 21640 34400 21692 34406
rect 21640 34342 21692 34348
rect 21652 34241 21680 34342
rect 21638 34232 21694 34241
rect 21638 34167 21694 34176
rect 21652 34134 21680 34167
rect 21640 34128 21692 34134
rect 21640 34070 21692 34076
rect 21640 33992 21692 33998
rect 21640 33934 21692 33940
rect 21652 33425 21680 33934
rect 21638 33416 21694 33425
rect 21638 33351 21694 33360
rect 21640 32904 21692 32910
rect 21744 32892 21772 36502
rect 21822 36408 21878 36417
rect 21822 36343 21878 36352
rect 21836 36310 21864 36343
rect 21824 36304 21876 36310
rect 21824 36246 21876 36252
rect 22020 36174 22048 39238
rect 22112 37466 22140 41704
rect 22204 40594 22232 41772
rect 22192 40588 22244 40594
rect 22192 40530 22244 40536
rect 22204 39642 22232 40530
rect 22296 39982 22324 42502
rect 22388 42158 22416 42894
rect 22480 42702 22508 43590
rect 22468 42696 22520 42702
rect 22468 42638 22520 42644
rect 22376 42152 22428 42158
rect 22376 42094 22428 42100
rect 22388 41750 22416 42094
rect 22480 42022 22508 42638
rect 22572 42566 22600 44270
rect 22652 44192 22704 44198
rect 22652 44134 22704 44140
rect 22664 43194 22692 44134
rect 22756 43858 22784 45562
rect 22744 43852 22796 43858
rect 22744 43794 22796 43800
rect 22756 43314 22784 43794
rect 22744 43308 22796 43314
rect 22744 43250 22796 43256
rect 22664 43166 22784 43194
rect 22756 42770 22784 43166
rect 22848 43081 22876 48010
rect 22940 43625 22968 48062
rect 23124 47954 23152 51342
rect 23296 51342 23348 51348
rect 23202 51303 23258 51312
rect 23216 50454 23244 51303
rect 23296 51264 23348 51270
rect 23296 51206 23348 51212
rect 23308 50833 23336 51206
rect 23294 50824 23350 50833
rect 23294 50759 23350 50768
rect 23296 50720 23348 50726
rect 23296 50662 23348 50668
rect 23204 50448 23256 50454
rect 23204 50390 23256 50396
rect 23204 49836 23256 49842
rect 23204 49778 23256 49784
rect 23032 47926 23152 47954
rect 23032 46753 23060 47926
rect 23110 47832 23166 47841
rect 23110 47767 23112 47776
rect 23164 47767 23166 47776
rect 23112 47738 23164 47744
rect 23216 47530 23244 49778
rect 23204 47524 23256 47530
rect 23204 47466 23256 47472
rect 23308 47410 23336 50662
rect 23124 47382 23336 47410
rect 23018 46744 23074 46753
rect 23018 46679 23074 46688
rect 23124 46050 23152 47382
rect 23294 47288 23350 47297
rect 23294 47223 23350 47232
rect 23204 47184 23256 47190
rect 23204 47126 23256 47132
rect 23216 46646 23244 47126
rect 23308 47122 23336 47223
rect 23296 47116 23348 47122
rect 23296 47058 23348 47064
rect 23204 46640 23256 46646
rect 23204 46582 23256 46588
rect 23216 46170 23244 46582
rect 23204 46164 23256 46170
rect 23204 46106 23256 46112
rect 23032 46022 23152 46050
rect 23204 46028 23256 46034
rect 22926 43616 22982 43625
rect 22926 43551 22982 43560
rect 22940 43450 22968 43551
rect 22928 43444 22980 43450
rect 22928 43386 22980 43392
rect 22834 43072 22890 43081
rect 22834 43007 22890 43016
rect 22928 42832 22980 42838
rect 22928 42774 22980 42780
rect 22652 42764 22704 42770
rect 22652 42706 22704 42712
rect 22744 42764 22796 42770
rect 22744 42706 22796 42712
rect 22560 42560 22612 42566
rect 22560 42502 22612 42508
rect 22664 42090 22692 42706
rect 22652 42084 22704 42090
rect 22652 42026 22704 42032
rect 22468 42016 22520 42022
rect 22468 41958 22520 41964
rect 22756 41818 22784 42706
rect 22468 41812 22520 41818
rect 22468 41754 22520 41760
rect 22744 41812 22796 41818
rect 22744 41754 22796 41760
rect 22376 41744 22428 41750
rect 22376 41686 22428 41692
rect 22480 41546 22508 41754
rect 22940 41721 22968 42774
rect 23032 42294 23060 46022
rect 23204 45970 23256 45976
rect 23110 45928 23166 45937
rect 23110 45863 23166 45872
rect 23124 45014 23152 45863
rect 23216 45098 23244 45970
rect 23296 45824 23348 45830
rect 23296 45766 23348 45772
rect 23308 45393 23336 45766
rect 23294 45384 23350 45393
rect 23294 45319 23350 45328
rect 23294 45112 23350 45121
rect 23216 45070 23294 45098
rect 23294 45047 23296 45056
rect 23348 45047 23350 45056
rect 23296 45018 23348 45024
rect 23112 45008 23164 45014
rect 23112 44950 23164 44956
rect 23124 44538 23152 44950
rect 23112 44532 23164 44538
rect 23112 44474 23164 44480
rect 23110 44024 23166 44033
rect 23110 43959 23166 43968
rect 23124 43858 23152 43959
rect 23112 43852 23164 43858
rect 23112 43794 23164 43800
rect 23124 42838 23152 43794
rect 23112 42832 23164 42838
rect 23112 42774 23164 42780
rect 23020 42288 23072 42294
rect 23020 42230 23072 42236
rect 22926 41712 22982 41721
rect 22560 41676 22612 41682
rect 23032 41682 23060 42230
rect 23296 42016 23348 42022
rect 23296 41958 23348 41964
rect 23202 41712 23258 41721
rect 22926 41647 22982 41656
rect 23020 41676 23072 41682
rect 22560 41618 22612 41624
rect 22468 41540 22520 41546
rect 22468 41482 22520 41488
rect 22480 41274 22508 41482
rect 22468 41268 22520 41274
rect 22468 41210 22520 41216
rect 22572 40662 22600 41618
rect 22560 40656 22612 40662
rect 22560 40598 22612 40604
rect 22284 39976 22336 39982
rect 22284 39918 22336 39924
rect 22376 39908 22428 39914
rect 22376 39850 22428 39856
rect 22192 39636 22244 39642
rect 22192 39578 22244 39584
rect 22388 38962 22416 39850
rect 22560 39840 22612 39846
rect 22560 39782 22612 39788
rect 22376 38956 22428 38962
rect 22376 38898 22428 38904
rect 22572 38894 22600 39782
rect 22560 38888 22612 38894
rect 22560 38830 22612 38836
rect 22652 38344 22704 38350
rect 22652 38286 22704 38292
rect 22100 37460 22152 37466
rect 22100 37402 22152 37408
rect 22112 36922 22140 37402
rect 22560 37324 22612 37330
rect 22560 37266 22612 37272
rect 22468 37256 22520 37262
rect 22468 37198 22520 37204
rect 22374 37088 22430 37097
rect 22374 37023 22430 37032
rect 22100 36916 22152 36922
rect 22100 36858 22152 36864
rect 21824 36168 21876 36174
rect 21824 36110 21876 36116
rect 22008 36168 22060 36174
rect 22008 36110 22060 36116
rect 21836 34082 21864 36110
rect 22284 35556 22336 35562
rect 22284 35498 22336 35504
rect 22192 35284 22244 35290
rect 22192 35226 22244 35232
rect 22006 35184 22062 35193
rect 22006 35119 22008 35128
rect 22060 35119 22062 35128
rect 22008 35090 22060 35096
rect 22020 34746 22048 35090
rect 22204 35086 22232 35226
rect 22296 35222 22324 35498
rect 22284 35216 22336 35222
rect 22284 35158 22336 35164
rect 22192 35080 22244 35086
rect 22192 35022 22244 35028
rect 22204 34746 22232 35022
rect 22008 34740 22060 34746
rect 22008 34682 22060 34688
rect 22192 34740 22244 34746
rect 22192 34682 22244 34688
rect 22296 34678 22324 35158
rect 22284 34672 22336 34678
rect 22190 34640 22246 34649
rect 22284 34614 22336 34620
rect 22190 34575 22246 34584
rect 21836 34054 22048 34082
rect 21822 33688 21878 33697
rect 21822 33623 21878 33632
rect 21836 33289 21864 33623
rect 21916 33312 21968 33318
rect 21822 33280 21878 33289
rect 21916 33254 21968 33260
rect 21822 33215 21878 33224
rect 21692 32864 21772 32892
rect 21640 32846 21692 32852
rect 21730 32736 21786 32745
rect 21730 32671 21786 32680
rect 21744 32366 21772 32671
rect 21928 32586 21956 33254
rect 22020 32774 22048 34054
rect 22008 32768 22060 32774
rect 22008 32710 22060 32716
rect 21928 32558 22140 32586
rect 22006 32464 22062 32473
rect 22006 32399 22062 32408
rect 21732 32360 21784 32366
rect 21732 32302 21784 32308
rect 21640 32224 21692 32230
rect 21640 32166 21692 32172
rect 21652 30122 21680 32166
rect 21744 32026 21772 32302
rect 21732 32020 21784 32026
rect 21732 31962 21784 31968
rect 21732 31884 21784 31890
rect 21732 31826 21784 31832
rect 21744 31482 21772 31826
rect 21732 31476 21784 31482
rect 21732 31418 21784 31424
rect 21732 31204 21784 31210
rect 21732 31146 21784 31152
rect 21640 30116 21692 30122
rect 21640 30058 21692 30064
rect 21638 28928 21694 28937
rect 21638 28863 21694 28872
rect 21548 28212 21600 28218
rect 21548 28154 21600 28160
rect 21652 25809 21680 28863
rect 21638 25800 21694 25809
rect 21638 25735 21694 25744
rect 21744 23769 21772 31146
rect 21916 30932 21968 30938
rect 21916 30874 21968 30880
rect 21928 29850 21956 30874
rect 21916 29844 21968 29850
rect 21916 29786 21968 29792
rect 21824 29708 21876 29714
rect 21824 29650 21876 29656
rect 21836 29306 21864 29650
rect 21824 29300 21876 29306
rect 21824 29242 21876 29248
rect 21916 28076 21968 28082
rect 21916 28018 21968 28024
rect 21824 27940 21876 27946
rect 21824 27882 21876 27888
rect 21730 23760 21786 23769
rect 21730 23695 21786 23704
rect 21730 20632 21786 20641
rect 21730 20567 21786 20576
rect 21454 20224 21510 20233
rect 21454 20159 21510 20168
rect 21638 13696 21694 13705
rect 21638 13631 21694 13640
rect 21548 13388 21600 13394
rect 21652 13376 21680 13631
rect 21600 13348 21680 13376
rect 21548 13330 21600 13336
rect 21456 13320 21508 13326
rect 21456 13262 21508 13268
rect 21468 12986 21496 13262
rect 21652 12986 21680 13348
rect 21456 12980 21508 12986
rect 21456 12922 21508 12928
rect 21640 12980 21692 12986
rect 21640 12922 21692 12928
rect 21364 10804 21416 10810
rect 21364 10746 21416 10752
rect 20956 10364 21252 10384
rect 21012 10362 21036 10364
rect 21092 10362 21116 10364
rect 21172 10362 21196 10364
rect 21034 10310 21036 10362
rect 21098 10310 21110 10362
rect 21172 10310 21174 10362
rect 21012 10308 21036 10310
rect 21092 10308 21116 10310
rect 21172 10308 21196 10310
rect 20956 10288 21252 10308
rect 20720 9648 20772 9654
rect 20720 9590 20772 9596
rect 20956 9276 21252 9296
rect 21012 9274 21036 9276
rect 21092 9274 21116 9276
rect 21172 9274 21196 9276
rect 21034 9222 21036 9274
rect 21098 9222 21110 9274
rect 21172 9222 21174 9274
rect 21012 9220 21036 9222
rect 21092 9220 21116 9222
rect 21172 9220 21196 9222
rect 20956 9200 21252 9220
rect 20956 8188 21252 8208
rect 21012 8186 21036 8188
rect 21092 8186 21116 8188
rect 21172 8186 21196 8188
rect 21034 8134 21036 8186
rect 21098 8134 21110 8186
rect 21172 8134 21174 8186
rect 21012 8132 21036 8134
rect 21092 8132 21116 8134
rect 21172 8132 21196 8134
rect 20956 8112 21252 8132
rect 20956 7100 21252 7120
rect 21012 7098 21036 7100
rect 21092 7098 21116 7100
rect 21172 7098 21196 7100
rect 21034 7046 21036 7098
rect 21098 7046 21110 7098
rect 21172 7046 21174 7098
rect 21012 7044 21036 7046
rect 21092 7044 21116 7046
rect 21172 7044 21196 7046
rect 20956 7024 21252 7044
rect 20956 6012 21252 6032
rect 21012 6010 21036 6012
rect 21092 6010 21116 6012
rect 21172 6010 21196 6012
rect 21034 5958 21036 6010
rect 21098 5958 21110 6010
rect 21172 5958 21174 6010
rect 21012 5956 21036 5958
rect 21092 5956 21116 5958
rect 21172 5956 21196 5958
rect 20956 5936 21252 5956
rect 20956 4924 21252 4944
rect 21012 4922 21036 4924
rect 21092 4922 21116 4924
rect 21172 4922 21196 4924
rect 21034 4870 21036 4922
rect 21098 4870 21110 4922
rect 21172 4870 21174 4922
rect 21012 4868 21036 4870
rect 21092 4868 21116 4870
rect 21172 4868 21196 4870
rect 20956 4848 21252 4868
rect 21468 4865 21496 12922
rect 21744 12866 21772 20567
rect 21652 12838 21772 12866
rect 21454 4856 21510 4865
rect 21454 4791 21510 4800
rect 20956 3836 21252 3856
rect 21012 3834 21036 3836
rect 21092 3834 21116 3836
rect 21172 3834 21196 3836
rect 21034 3782 21036 3834
rect 21098 3782 21110 3834
rect 21172 3782 21174 3834
rect 21012 3780 21036 3782
rect 21092 3780 21116 3782
rect 21172 3780 21196 3782
rect 20956 3760 21252 3780
rect 21652 3641 21680 12838
rect 21732 12776 21784 12782
rect 21732 12718 21784 12724
rect 21744 10305 21772 12718
rect 21730 10296 21786 10305
rect 21730 10231 21786 10240
rect 21836 8401 21864 27882
rect 21928 27606 21956 28018
rect 21916 27600 21968 27606
rect 21916 27542 21968 27548
rect 21914 19272 21970 19281
rect 21914 19207 21970 19216
rect 21822 8392 21878 8401
rect 21822 8327 21878 8336
rect 21638 3632 21694 3641
rect 21638 3567 21694 3576
rect 21928 2938 21956 19207
rect 22020 13977 22048 32399
rect 22112 30666 22140 32558
rect 22204 30870 22232 34575
rect 22388 34202 22416 37023
rect 22480 36650 22508 37198
rect 22468 36644 22520 36650
rect 22468 36586 22520 36592
rect 22480 36174 22508 36586
rect 22468 36168 22520 36174
rect 22468 36110 22520 36116
rect 22480 35834 22508 36110
rect 22468 35828 22520 35834
rect 22468 35770 22520 35776
rect 22572 35601 22600 37266
rect 22558 35592 22614 35601
rect 22558 35527 22614 35536
rect 22468 34944 22520 34950
rect 22468 34886 22520 34892
rect 22480 34785 22508 34886
rect 22466 34776 22522 34785
rect 22466 34711 22522 34720
rect 22376 34196 22428 34202
rect 22296 34156 22376 34184
rect 22296 33454 22324 34156
rect 22376 34138 22428 34144
rect 22374 33824 22430 33833
rect 22374 33759 22430 33768
rect 22284 33448 22336 33454
rect 22284 33390 22336 33396
rect 22296 32994 22324 33390
rect 22388 33386 22416 33759
rect 22558 33552 22614 33561
rect 22558 33487 22560 33496
rect 22612 33487 22614 33496
rect 22560 33458 22612 33464
rect 22376 33380 22428 33386
rect 22376 33322 22428 33328
rect 22296 32966 22416 32994
rect 22284 32904 22336 32910
rect 22282 32872 22284 32881
rect 22336 32872 22338 32881
rect 22282 32807 22338 32816
rect 22284 32496 22336 32502
rect 22284 32438 22336 32444
rect 22192 30864 22244 30870
rect 22192 30806 22244 30812
rect 22192 30728 22244 30734
rect 22192 30670 22244 30676
rect 22100 30660 22152 30666
rect 22100 30602 22152 30608
rect 22204 29782 22232 30670
rect 22192 29776 22244 29782
rect 22192 29718 22244 29724
rect 22296 20641 22324 32438
rect 22388 29510 22416 32966
rect 22560 32360 22612 32366
rect 22560 32302 22612 32308
rect 22572 32026 22600 32302
rect 22560 32020 22612 32026
rect 22560 31962 22612 31968
rect 22664 30025 22692 38286
rect 22742 37360 22798 37369
rect 22742 37295 22744 37304
rect 22796 37295 22798 37304
rect 22744 37266 22796 37272
rect 22756 36922 22784 37266
rect 22744 36916 22796 36922
rect 22744 36858 22796 36864
rect 22836 36236 22888 36242
rect 22836 36178 22888 36184
rect 22848 35494 22876 36178
rect 22836 35488 22888 35494
rect 22834 35456 22836 35465
rect 22888 35456 22890 35465
rect 22834 35391 22890 35400
rect 22836 33992 22888 33998
rect 22836 33934 22888 33940
rect 22742 33008 22798 33017
rect 22742 32943 22798 32952
rect 22756 32502 22784 32943
rect 22744 32496 22796 32502
rect 22744 32438 22796 32444
rect 22650 30016 22706 30025
rect 22650 29951 22706 29960
rect 22376 29504 22428 29510
rect 22376 29446 22428 29452
rect 22560 28416 22612 28422
rect 22560 28358 22612 28364
rect 22572 28014 22600 28358
rect 22560 28008 22612 28014
rect 22560 27950 22612 27956
rect 22468 21004 22520 21010
rect 22468 20946 22520 20952
rect 22480 20890 22508 20946
rect 22388 20862 22508 20890
rect 22282 20632 22338 20641
rect 22282 20567 22338 20576
rect 22388 20262 22416 20862
rect 22376 20256 22428 20262
rect 22376 20198 22428 20204
rect 22006 13968 22062 13977
rect 22006 13903 22062 13912
rect 22020 6225 22048 13903
rect 22006 6216 22062 6225
rect 22006 6151 22062 6160
rect 22388 4049 22416 20198
rect 22468 16584 22520 16590
rect 22468 16526 22520 16532
rect 22744 16584 22796 16590
rect 22744 16526 22796 16532
rect 22480 15910 22508 16526
rect 22756 15910 22784 16526
rect 22468 15904 22520 15910
rect 22468 15846 22520 15852
rect 22744 15904 22796 15910
rect 22744 15846 22796 15852
rect 22480 15337 22508 15846
rect 22466 15328 22522 15337
rect 22466 15263 22522 15272
rect 22558 14376 22614 14385
rect 22558 14311 22614 14320
rect 22572 13530 22600 14311
rect 22756 13705 22784 15846
rect 22742 13696 22798 13705
rect 22742 13631 22798 13640
rect 22560 13524 22612 13530
rect 22560 13466 22612 13472
rect 22558 11792 22614 11801
rect 22558 11727 22614 11736
rect 22374 4040 22430 4049
rect 22374 3975 22430 3984
rect 21928 2910 22048 2938
rect 20956 2748 21252 2768
rect 21012 2746 21036 2748
rect 21092 2746 21116 2748
rect 21172 2746 21196 2748
rect 21034 2694 21036 2746
rect 21098 2694 21110 2746
rect 21172 2694 21174 2746
rect 21012 2692 21036 2694
rect 21092 2692 21116 2694
rect 21172 2692 21196 2694
rect 20956 2672 21252 2692
rect 22020 2666 22048 2910
rect 21456 2644 21508 2650
rect 21456 2586 21508 2592
rect 21652 2638 22048 2666
rect 21468 2446 21496 2586
rect 21456 2440 21508 2446
rect 20902 2408 20958 2417
rect 20628 2372 20680 2378
rect 21456 2382 21508 2388
rect 20902 2343 20904 2352
rect 20628 2314 20680 2320
rect 20956 2343 20958 2352
rect 20904 2314 20956 2320
rect 20534 912 20590 921
rect 20534 847 20590 856
rect 20718 912 20774 921
rect 20718 847 20774 856
rect 20732 800 20760 847
rect 21652 800 21680 2638
rect 22572 800 22600 11727
rect 22848 10713 22876 33934
rect 22940 31890 22968 41647
rect 23202 41647 23258 41656
rect 23020 41618 23072 41624
rect 23032 41274 23060 41618
rect 23216 41614 23244 41647
rect 23204 41608 23256 41614
rect 23204 41550 23256 41556
rect 23202 41440 23258 41449
rect 23202 41375 23258 41384
rect 23020 41268 23072 41274
rect 23020 41210 23072 41216
rect 23216 40730 23244 41375
rect 23204 40724 23256 40730
rect 23204 40666 23256 40672
rect 23308 40526 23336 41958
rect 23296 40520 23348 40526
rect 23296 40462 23348 40468
rect 23308 39846 23336 40462
rect 23296 39840 23348 39846
rect 23296 39782 23348 39788
rect 23020 35624 23072 35630
rect 23020 35566 23072 35572
rect 23032 34950 23060 35566
rect 23400 35154 23428 70926
rect 23480 64320 23532 64326
rect 23480 64262 23532 64268
rect 23492 63034 23520 64262
rect 23676 63510 23704 74695
rect 23664 63504 23716 63510
rect 23664 63446 23716 63452
rect 23480 63028 23532 63034
rect 23480 62970 23532 62976
rect 23478 59120 23534 59129
rect 23478 59055 23480 59064
rect 23532 59055 23534 59064
rect 23480 59026 23532 59032
rect 23492 58138 23520 59026
rect 23756 58676 23808 58682
rect 23756 58618 23808 58624
rect 23664 58540 23716 58546
rect 23664 58482 23716 58488
rect 23572 58336 23624 58342
rect 23572 58278 23624 58284
rect 23480 58132 23532 58138
rect 23480 58074 23532 58080
rect 23584 54754 23612 58278
rect 23676 57594 23704 58482
rect 23768 58002 23796 58618
rect 23756 57996 23808 58002
rect 23756 57938 23808 57944
rect 23768 57594 23796 57938
rect 23664 57588 23716 57594
rect 23664 57530 23716 57536
rect 23756 57588 23808 57594
rect 23756 57530 23808 57536
rect 23860 55826 23888 77318
rect 23940 75336 23992 75342
rect 23940 75278 23992 75284
rect 23952 74662 23980 75278
rect 23940 74656 23992 74662
rect 23940 74598 23992 74604
rect 23952 74497 23980 74598
rect 23938 74488 23994 74497
rect 23938 74423 23994 74432
rect 24412 74361 24440 79200
rect 24398 74352 24454 74361
rect 24398 74287 24454 74296
rect 24490 69048 24546 69057
rect 24490 68983 24546 68992
rect 24216 63436 24268 63442
rect 24216 63378 24268 63384
rect 24400 63436 24452 63442
rect 24400 63378 24452 63384
rect 24032 63368 24084 63374
rect 24032 63310 24084 63316
rect 24044 62694 24072 63310
rect 24228 62830 24256 63378
rect 24412 63034 24440 63378
rect 24400 63028 24452 63034
rect 24400 62970 24452 62976
rect 24216 62824 24268 62830
rect 24216 62766 24268 62772
rect 24032 62688 24084 62694
rect 24032 62630 24084 62636
rect 23938 58440 23994 58449
rect 23938 58375 23994 58384
rect 23952 58002 23980 58375
rect 23940 57996 23992 58002
rect 23940 57938 23992 57944
rect 23952 57526 23980 57938
rect 23940 57520 23992 57526
rect 23940 57462 23992 57468
rect 23952 56710 23980 57462
rect 23940 56704 23992 56710
rect 23940 56646 23992 56652
rect 23848 55820 23900 55826
rect 23848 55762 23900 55768
rect 23860 55418 23888 55762
rect 24044 55434 24072 62630
rect 23848 55412 23900 55418
rect 23848 55354 23900 55360
rect 23952 55406 24072 55434
rect 23584 54726 23796 54754
rect 23572 54664 23624 54670
rect 23572 54606 23624 54612
rect 23584 54126 23612 54606
rect 23572 54120 23624 54126
rect 23478 54088 23534 54097
rect 23572 54062 23624 54068
rect 23664 54120 23716 54126
rect 23664 54062 23716 54068
rect 23478 54023 23534 54032
rect 23492 52018 23520 54023
rect 23480 52012 23532 52018
rect 23480 51954 23532 51960
rect 23480 51400 23532 51406
rect 23480 51342 23532 51348
rect 23492 51066 23520 51342
rect 23480 51060 23532 51066
rect 23480 51002 23532 51008
rect 23492 50776 23520 51002
rect 23584 50969 23612 54062
rect 23676 53990 23704 54062
rect 23664 53984 23716 53990
rect 23664 53926 23716 53932
rect 23768 52544 23796 54726
rect 23952 53786 23980 55406
rect 24032 55276 24084 55282
rect 24032 55218 24084 55224
rect 24044 55078 24072 55218
rect 24124 55208 24176 55214
rect 24124 55150 24176 55156
rect 24032 55072 24084 55078
rect 24032 55014 24084 55020
rect 23940 53780 23992 53786
rect 23860 53740 23940 53768
rect 23860 53242 23888 53740
rect 23940 53722 23992 53728
rect 23940 53644 23992 53650
rect 23940 53586 23992 53592
rect 23848 53236 23900 53242
rect 23848 53178 23900 53184
rect 23952 52902 23980 53586
rect 23940 52896 23992 52902
rect 23940 52838 23992 52844
rect 23952 52698 23980 52838
rect 23940 52692 23992 52698
rect 23940 52634 23992 52640
rect 23768 52516 23980 52544
rect 23754 52456 23810 52465
rect 23754 52391 23756 52400
rect 23808 52391 23810 52400
rect 23756 52362 23808 52368
rect 23848 52352 23900 52358
rect 23848 52294 23900 52300
rect 23756 52080 23808 52086
rect 23756 52022 23808 52028
rect 23664 51876 23716 51882
rect 23664 51818 23716 51824
rect 23676 51513 23704 51818
rect 23768 51542 23796 52022
rect 23860 51882 23888 52294
rect 23952 52086 23980 52516
rect 23940 52080 23992 52086
rect 23940 52022 23992 52028
rect 23848 51876 23900 51882
rect 23848 51818 23900 51824
rect 23860 51610 23888 51818
rect 23940 51808 23992 51814
rect 23940 51750 23992 51756
rect 23952 51610 23980 51750
rect 23848 51604 23900 51610
rect 23848 51546 23900 51552
rect 23940 51604 23992 51610
rect 23940 51546 23992 51552
rect 23756 51536 23808 51542
rect 23662 51504 23718 51513
rect 23756 51478 23808 51484
rect 23662 51439 23718 51448
rect 23570 50960 23626 50969
rect 23570 50895 23626 50904
rect 23768 50862 23796 51478
rect 23848 51332 23900 51338
rect 23848 51274 23900 51280
rect 23756 50856 23808 50862
rect 23756 50798 23808 50804
rect 23492 50748 23704 50776
rect 23570 50688 23626 50697
rect 23570 50623 23626 50632
rect 23584 49978 23612 50623
rect 23572 49972 23624 49978
rect 23572 49914 23624 49920
rect 23584 49774 23612 49914
rect 23572 49768 23624 49774
rect 23572 49710 23624 49716
rect 23480 49088 23532 49094
rect 23480 49030 23532 49036
rect 23492 48006 23520 49030
rect 23676 48754 23704 50748
rect 23754 50688 23810 50697
rect 23754 50623 23810 50632
rect 23664 48748 23716 48754
rect 23664 48690 23716 48696
rect 23572 48204 23624 48210
rect 23572 48146 23624 48152
rect 23584 48113 23612 48146
rect 23570 48104 23626 48113
rect 23570 48039 23626 48048
rect 23480 48000 23532 48006
rect 23480 47942 23532 47948
rect 23492 47598 23520 47942
rect 23572 47728 23624 47734
rect 23572 47670 23624 47676
rect 23480 47592 23532 47598
rect 23480 47534 23532 47540
rect 23492 46646 23520 47534
rect 23584 46866 23612 47670
rect 23676 47580 23704 48690
rect 23768 48142 23796 50623
rect 23756 48136 23808 48142
rect 23756 48078 23808 48084
rect 23768 47734 23796 48078
rect 23756 47728 23808 47734
rect 23756 47670 23808 47676
rect 23756 47592 23808 47598
rect 23676 47552 23756 47580
rect 23676 47258 23704 47552
rect 23756 47534 23808 47540
rect 23664 47252 23716 47258
rect 23664 47194 23716 47200
rect 23584 46838 23704 46866
rect 23572 46708 23624 46714
rect 23572 46650 23624 46656
rect 23480 46640 23532 46646
rect 23478 46608 23480 46617
rect 23532 46608 23534 46617
rect 23478 46543 23534 46552
rect 23480 46504 23532 46510
rect 23480 46446 23532 46452
rect 23492 46170 23520 46446
rect 23584 46374 23612 46650
rect 23572 46368 23624 46374
rect 23572 46310 23624 46316
rect 23480 46164 23532 46170
rect 23480 46106 23532 46112
rect 23480 46028 23532 46034
rect 23480 45970 23532 45976
rect 23492 45626 23520 45970
rect 23480 45620 23532 45626
rect 23480 45562 23532 45568
rect 23584 44946 23612 46310
rect 23676 45626 23704 46838
rect 23860 46186 23888 51274
rect 23952 49366 23980 51546
rect 24044 51338 24072 55014
rect 24136 54874 24164 55150
rect 24124 54868 24176 54874
rect 24124 54810 24176 54816
rect 24136 52562 24164 54810
rect 24228 54738 24256 62766
rect 24308 58880 24360 58886
rect 24308 58822 24360 58828
rect 24320 58478 24348 58822
rect 24308 58472 24360 58478
rect 24308 58414 24360 58420
rect 24400 57860 24452 57866
rect 24400 57802 24452 57808
rect 24308 56160 24360 56166
rect 24308 56102 24360 56108
rect 24216 54732 24268 54738
rect 24216 54674 24268 54680
rect 24124 52556 24176 52562
rect 24124 52498 24176 52504
rect 24214 52320 24270 52329
rect 24214 52255 24270 52264
rect 24124 52080 24176 52086
rect 24124 52022 24176 52028
rect 24136 51474 24164 52022
rect 24124 51468 24176 51474
rect 24124 51410 24176 51416
rect 24032 51332 24084 51338
rect 24032 51274 24084 51280
rect 24136 50998 24164 51410
rect 24124 50992 24176 50998
rect 24124 50934 24176 50940
rect 23940 49360 23992 49366
rect 23940 49302 23992 49308
rect 23940 49224 23992 49230
rect 23940 49166 23992 49172
rect 23952 46374 23980 49166
rect 24030 48512 24086 48521
rect 24030 48447 24086 48456
rect 23940 46368 23992 46374
rect 23940 46310 23992 46316
rect 23768 46158 23888 46186
rect 23664 45620 23716 45626
rect 23664 45562 23716 45568
rect 23664 45484 23716 45490
rect 23664 45426 23716 45432
rect 23676 45082 23704 45426
rect 23664 45076 23716 45082
rect 23664 45018 23716 45024
rect 23572 44940 23624 44946
rect 23572 44882 23624 44888
rect 23584 44441 23612 44882
rect 23664 44872 23716 44878
rect 23664 44814 23716 44820
rect 23570 44432 23626 44441
rect 23570 44367 23626 44376
rect 23584 44198 23612 44367
rect 23572 44192 23624 44198
rect 23572 44134 23624 44140
rect 23480 43920 23532 43926
rect 23480 43862 23532 43868
rect 23492 43382 23520 43862
rect 23480 43376 23532 43382
rect 23478 43344 23480 43353
rect 23532 43344 23534 43353
rect 23478 43279 23534 43288
rect 23584 42566 23612 44134
rect 23676 43450 23704 44814
rect 23664 43444 23716 43450
rect 23664 43386 23716 43392
rect 23572 42560 23624 42566
rect 23572 42502 23624 42508
rect 23676 42265 23704 43386
rect 23662 42256 23718 42265
rect 23662 42191 23718 42200
rect 23572 41472 23624 41478
rect 23572 41414 23624 41420
rect 23478 39944 23534 39953
rect 23478 39879 23480 39888
rect 23532 39879 23534 39888
rect 23480 39850 23532 39856
rect 23480 39296 23532 39302
rect 23480 39238 23532 39244
rect 23492 38758 23520 39238
rect 23480 38752 23532 38758
rect 23480 38694 23532 38700
rect 23492 37262 23520 38694
rect 23584 38010 23612 41414
rect 23676 41070 23704 42191
rect 23664 41064 23716 41070
rect 23664 41006 23716 41012
rect 23676 39846 23704 41006
rect 23768 40118 23796 46158
rect 23940 45824 23992 45830
rect 23940 45766 23992 45772
rect 23848 45348 23900 45354
rect 23848 45290 23900 45296
rect 23860 44985 23888 45290
rect 23846 44976 23902 44985
rect 23846 44911 23902 44920
rect 23848 44328 23900 44334
rect 23848 44270 23900 44276
rect 23860 43994 23888 44270
rect 23848 43988 23900 43994
rect 23848 43930 23900 43936
rect 23848 43784 23900 43790
rect 23848 43726 23900 43732
rect 23860 43246 23888 43726
rect 23848 43240 23900 43246
rect 23848 43182 23900 43188
rect 23860 42770 23888 43182
rect 23848 42764 23900 42770
rect 23848 42706 23900 42712
rect 23952 40934 23980 45766
rect 24044 44520 24072 48447
rect 24136 47705 24164 50934
rect 24122 47696 24178 47705
rect 24122 47631 24178 47640
rect 24124 47524 24176 47530
rect 24124 47466 24176 47472
rect 24136 47258 24164 47466
rect 24124 47252 24176 47258
rect 24124 47194 24176 47200
rect 24122 46064 24178 46073
rect 24122 45999 24124 46008
rect 24176 45999 24178 46008
rect 24124 45970 24176 45976
rect 24044 44492 24164 44520
rect 24032 44396 24084 44402
rect 24032 44338 24084 44344
rect 23940 40928 23992 40934
rect 23940 40870 23992 40876
rect 23756 40112 23808 40118
rect 23756 40054 23808 40060
rect 23664 39840 23716 39846
rect 23664 39782 23716 39788
rect 23676 39506 23704 39782
rect 23664 39500 23716 39506
rect 23664 39442 23716 39448
rect 23676 39098 23704 39442
rect 23664 39092 23716 39098
rect 23664 39034 23716 39040
rect 23662 38448 23718 38457
rect 23662 38383 23664 38392
rect 23716 38383 23718 38392
rect 23664 38354 23716 38360
rect 23572 38004 23624 38010
rect 23572 37946 23624 37952
rect 23584 37806 23612 37946
rect 23676 37874 23704 38354
rect 23768 38010 23796 40054
rect 23952 38010 23980 40870
rect 23756 38004 23808 38010
rect 23756 37946 23808 37952
rect 23940 38004 23992 38010
rect 23940 37946 23992 37952
rect 24044 37890 24072 44338
rect 24136 43790 24164 44492
rect 24228 44402 24256 52255
rect 24320 51066 24348 56102
rect 24308 51060 24360 51066
rect 24308 51002 24360 51008
rect 24320 50862 24348 51002
rect 24308 50856 24360 50862
rect 24308 50798 24360 50804
rect 24308 50720 24360 50726
rect 24308 50662 24360 50668
rect 24320 50522 24348 50662
rect 24308 50516 24360 50522
rect 24308 50458 24360 50464
rect 24308 50380 24360 50386
rect 24308 50322 24360 50328
rect 24320 49774 24348 50322
rect 24308 49768 24360 49774
rect 24308 49710 24360 49716
rect 24320 47297 24348 49710
rect 24412 49230 24440 57802
rect 24504 55214 24532 68983
rect 24582 59392 24638 59401
rect 24582 59327 24638 59336
rect 24596 58546 24624 59327
rect 24584 58540 24636 58546
rect 24584 58482 24636 58488
rect 24596 58002 24624 58482
rect 24584 57996 24636 58002
rect 24584 57938 24636 57944
rect 24688 56166 24716 79591
rect 24858 79200 24914 80000
rect 25778 79200 25834 80000
rect 26698 79200 26754 80000
rect 27618 79200 27674 80000
rect 28078 79200 28134 80000
rect 28998 79200 29054 80000
rect 29918 79200 29974 80000
rect 24768 74996 24820 75002
rect 24768 74938 24820 74944
rect 24780 70428 24808 74938
rect 24872 74633 24900 79200
rect 25792 77058 25820 79200
rect 25870 78296 25926 78305
rect 25870 78231 25926 78240
rect 25884 77382 25912 78231
rect 25872 77376 25924 77382
rect 25872 77318 25924 77324
rect 25956 77276 26252 77296
rect 26012 77274 26036 77276
rect 26092 77274 26116 77276
rect 26172 77274 26196 77276
rect 26034 77222 26036 77274
rect 26098 77222 26110 77274
rect 26172 77222 26174 77274
rect 26012 77220 26036 77222
rect 26092 77220 26116 77222
rect 26172 77220 26196 77222
rect 25956 77200 26252 77220
rect 25700 77030 25820 77058
rect 25134 76392 25190 76401
rect 25134 76327 25190 76336
rect 25042 75984 25098 75993
rect 25042 75919 25098 75928
rect 25056 75546 25084 75919
rect 25044 75540 25096 75546
rect 25044 75482 25096 75488
rect 24858 74624 24914 74633
rect 24858 74559 24914 74568
rect 24860 70440 24912 70446
rect 24780 70400 24860 70428
rect 24860 70382 24912 70388
rect 24860 69352 24912 69358
rect 24860 69294 24912 69300
rect 24768 65204 24820 65210
rect 24872 65192 24900 69294
rect 25148 68921 25176 76327
rect 25226 74896 25282 74905
rect 25226 74831 25282 74840
rect 25240 69057 25268 74831
rect 25700 74769 25728 77030
rect 25778 76936 25834 76945
rect 25778 76871 25834 76880
rect 25686 74760 25742 74769
rect 25686 74695 25742 74704
rect 25502 70136 25558 70145
rect 25502 70071 25558 70080
rect 25226 69048 25282 69057
rect 25226 68983 25282 68992
rect 25134 68912 25190 68921
rect 25134 68847 25190 68856
rect 25516 67833 25544 70071
rect 25502 67824 25558 67833
rect 25502 67759 25558 67768
rect 25502 66736 25558 66745
rect 25502 66671 25558 66680
rect 24952 65544 25004 65550
rect 24952 65486 25004 65492
rect 24820 65164 24900 65192
rect 24768 65146 24820 65152
rect 24872 62830 24900 65164
rect 24860 62824 24912 62830
rect 24860 62766 24912 62772
rect 24964 62098 24992 65486
rect 24780 62070 24992 62098
rect 24676 56160 24728 56166
rect 24676 56102 24728 56108
rect 24780 55944 24808 62070
rect 25516 61962 25544 66671
rect 25792 65550 25820 76871
rect 25956 76188 26252 76208
rect 26012 76186 26036 76188
rect 26092 76186 26116 76188
rect 26172 76186 26196 76188
rect 26034 76134 26036 76186
rect 26098 76134 26110 76186
rect 26172 76134 26174 76186
rect 26012 76132 26036 76134
rect 26092 76132 26116 76134
rect 26172 76132 26196 76134
rect 25956 76112 26252 76132
rect 26712 75313 26740 79200
rect 26698 75304 26754 75313
rect 26698 75239 26754 75248
rect 25956 75100 26252 75120
rect 26012 75098 26036 75100
rect 26092 75098 26116 75100
rect 26172 75098 26196 75100
rect 26034 75046 26036 75098
rect 26098 75046 26110 75098
rect 26172 75046 26174 75098
rect 26012 75044 26036 75046
rect 26092 75044 26116 75046
rect 26172 75044 26196 75046
rect 25956 75024 26252 75044
rect 27632 74746 27660 79200
rect 28092 79098 28120 79200
rect 27816 79070 28120 79098
rect 27632 74718 27752 74746
rect 27620 74656 27672 74662
rect 27620 74598 27672 74604
rect 25956 74012 26252 74032
rect 26012 74010 26036 74012
rect 26092 74010 26116 74012
rect 26172 74010 26196 74012
rect 26034 73958 26036 74010
rect 26098 73958 26110 74010
rect 26172 73958 26174 74010
rect 26012 73956 26036 73958
rect 26092 73956 26116 73958
rect 26172 73956 26196 73958
rect 25956 73936 26252 73956
rect 25956 72924 26252 72944
rect 26012 72922 26036 72924
rect 26092 72922 26116 72924
rect 26172 72922 26196 72924
rect 26034 72870 26036 72922
rect 26098 72870 26110 72922
rect 26172 72870 26174 72922
rect 26012 72868 26036 72870
rect 26092 72868 26116 72870
rect 26172 72868 26196 72870
rect 25956 72848 26252 72868
rect 25956 71836 26252 71856
rect 26012 71834 26036 71836
rect 26092 71834 26116 71836
rect 26172 71834 26196 71836
rect 26034 71782 26036 71834
rect 26098 71782 26110 71834
rect 26172 71782 26174 71834
rect 26012 71780 26036 71782
rect 26092 71780 26116 71782
rect 26172 71780 26196 71782
rect 25956 71760 26252 71780
rect 26422 71768 26478 71777
rect 26422 71703 26478 71712
rect 25956 70748 26252 70768
rect 26012 70746 26036 70748
rect 26092 70746 26116 70748
rect 26172 70746 26196 70748
rect 26034 70694 26036 70746
rect 26098 70694 26110 70746
rect 26172 70694 26174 70746
rect 26012 70692 26036 70694
rect 26092 70692 26116 70694
rect 26172 70692 26196 70694
rect 25956 70672 26252 70692
rect 26436 70514 26464 71703
rect 26424 70508 26476 70514
rect 26424 70450 26476 70456
rect 26148 70440 26200 70446
rect 26148 70382 26200 70388
rect 26160 70106 26188 70382
rect 26424 70304 26476 70310
rect 26424 70246 26476 70252
rect 25872 70100 25924 70106
rect 25872 70042 25924 70048
rect 26148 70100 26200 70106
rect 26148 70042 26200 70048
rect 25884 69358 25912 70042
rect 25956 69660 26252 69680
rect 26012 69658 26036 69660
rect 26092 69658 26116 69660
rect 26172 69658 26196 69660
rect 26034 69606 26036 69658
rect 26098 69606 26110 69658
rect 26172 69606 26174 69658
rect 26012 69604 26036 69606
rect 26092 69604 26116 69606
rect 26172 69604 26196 69606
rect 25956 69584 26252 69604
rect 26436 69426 26464 70246
rect 26424 69420 26476 69426
rect 26424 69362 26476 69368
rect 25872 69352 25924 69358
rect 25872 69294 25924 69300
rect 26240 69352 26292 69358
rect 26240 69294 26292 69300
rect 26252 69018 26280 69294
rect 26240 69012 26292 69018
rect 26240 68954 26292 68960
rect 25956 68572 26252 68592
rect 26012 68570 26036 68572
rect 26092 68570 26116 68572
rect 26172 68570 26196 68572
rect 26034 68518 26036 68570
rect 26098 68518 26110 68570
rect 26172 68518 26174 68570
rect 26012 68516 26036 68518
rect 26092 68516 26116 68518
rect 26172 68516 26196 68518
rect 25956 68496 26252 68516
rect 25956 67484 26252 67504
rect 26012 67482 26036 67484
rect 26092 67482 26116 67484
rect 26172 67482 26196 67484
rect 26034 67430 26036 67482
rect 26098 67430 26110 67482
rect 26172 67430 26174 67482
rect 26012 67428 26036 67430
rect 26092 67428 26116 67430
rect 26172 67428 26196 67430
rect 25956 67408 26252 67428
rect 25956 66396 26252 66416
rect 26012 66394 26036 66396
rect 26092 66394 26116 66396
rect 26172 66394 26196 66396
rect 26034 66342 26036 66394
rect 26098 66342 26110 66394
rect 26172 66342 26174 66394
rect 26012 66340 26036 66342
rect 26092 66340 26116 66342
rect 26172 66340 26196 66342
rect 25956 66320 26252 66340
rect 25780 65544 25832 65550
rect 25780 65486 25832 65492
rect 25956 65308 26252 65328
rect 26012 65306 26036 65308
rect 26092 65306 26116 65308
rect 26172 65306 26196 65308
rect 26034 65254 26036 65306
rect 26098 65254 26110 65306
rect 26172 65254 26174 65306
rect 26012 65252 26036 65254
rect 26092 65252 26116 65254
rect 26172 65252 26196 65254
rect 25956 65232 26252 65252
rect 25594 65104 25650 65113
rect 25594 65039 25650 65048
rect 25608 62937 25636 65039
rect 27632 64818 27660 74598
rect 27724 70378 27752 74718
rect 27712 70372 27764 70378
rect 27712 70314 27764 70320
rect 27712 69216 27764 69222
rect 27712 69158 27764 69164
rect 27724 66298 27752 69158
rect 27712 66292 27764 66298
rect 27712 66234 27764 66240
rect 27540 64790 27660 64818
rect 25870 64696 25926 64705
rect 25870 64631 25926 64640
rect 25778 63336 25834 63345
rect 25778 63271 25834 63280
rect 25594 62928 25650 62937
rect 25594 62863 25650 62872
rect 25516 61934 25728 61962
rect 25594 61840 25650 61849
rect 25594 61775 25650 61784
rect 24950 61296 25006 61305
rect 24950 61231 25006 61240
rect 24596 55916 24808 55944
rect 24492 55208 24544 55214
rect 24492 55150 24544 55156
rect 24490 53136 24546 53145
rect 24490 53071 24492 53080
rect 24544 53071 24546 53080
rect 24492 53042 24544 53048
rect 24492 50788 24544 50794
rect 24492 50730 24544 50736
rect 24504 49842 24532 50730
rect 24492 49836 24544 49842
rect 24492 49778 24544 49784
rect 24400 49224 24452 49230
rect 24400 49166 24452 49172
rect 24400 49088 24452 49094
rect 24400 49030 24452 49036
rect 24412 47666 24440 49030
rect 24492 47796 24544 47802
rect 24492 47738 24544 47744
rect 24400 47660 24452 47666
rect 24400 47602 24452 47608
rect 24306 47288 24362 47297
rect 24306 47223 24362 47232
rect 24308 47048 24360 47054
rect 24308 46990 24360 46996
rect 24216 44396 24268 44402
rect 24216 44338 24268 44344
rect 24320 44248 24348 46990
rect 24412 46646 24440 47602
rect 24504 47598 24532 47738
rect 24492 47592 24544 47598
rect 24492 47534 24544 47540
rect 24504 47161 24532 47534
rect 24490 47152 24546 47161
rect 24490 47087 24546 47096
rect 24492 46980 24544 46986
rect 24492 46922 24544 46928
rect 24400 46640 24452 46646
rect 24400 46582 24452 46588
rect 24412 46170 24440 46582
rect 24400 46164 24452 46170
rect 24400 46106 24452 46112
rect 24504 46050 24532 46922
rect 24412 46022 24532 46050
rect 24412 45830 24440 46022
rect 24492 45960 24544 45966
rect 24492 45902 24544 45908
rect 24400 45824 24452 45830
rect 24400 45766 24452 45772
rect 24504 45626 24532 45902
rect 24492 45620 24544 45626
rect 24492 45562 24544 45568
rect 24492 45416 24544 45422
rect 24492 45358 24544 45364
rect 24228 44220 24348 44248
rect 24124 43784 24176 43790
rect 24124 43726 24176 43732
rect 24136 43450 24164 43726
rect 24124 43444 24176 43450
rect 24124 43386 24176 43392
rect 24124 40384 24176 40390
rect 24124 40326 24176 40332
rect 23664 37868 23716 37874
rect 23664 37810 23716 37816
rect 23768 37862 24072 37890
rect 23572 37800 23624 37806
rect 23572 37742 23624 37748
rect 23664 37664 23716 37670
rect 23664 37606 23716 37612
rect 23676 37330 23704 37606
rect 23664 37324 23716 37330
rect 23664 37266 23716 37272
rect 23480 37256 23532 37262
rect 23480 37198 23532 37204
rect 23572 36032 23624 36038
rect 23572 35974 23624 35980
rect 23584 35630 23612 35974
rect 23572 35624 23624 35630
rect 23572 35566 23624 35572
rect 23388 35148 23440 35154
rect 23388 35090 23440 35096
rect 23020 34944 23072 34950
rect 23020 34886 23072 34892
rect 23032 34542 23060 34886
rect 23400 34746 23428 35090
rect 23480 34944 23532 34950
rect 23480 34886 23532 34892
rect 23388 34740 23440 34746
rect 23388 34682 23440 34688
rect 23020 34536 23072 34542
rect 23020 34478 23072 34484
rect 23492 34184 23520 34886
rect 23308 34156 23520 34184
rect 23570 34232 23626 34241
rect 23570 34167 23626 34176
rect 23204 34128 23256 34134
rect 23204 34070 23256 34076
rect 23020 33992 23072 33998
rect 23020 33934 23072 33940
rect 23032 33658 23060 33934
rect 23216 33658 23244 34070
rect 23020 33652 23072 33658
rect 23020 33594 23072 33600
rect 23204 33652 23256 33658
rect 23204 33594 23256 33600
rect 23032 32366 23060 33594
rect 23112 33584 23164 33590
rect 23112 33526 23164 33532
rect 23124 32434 23152 33526
rect 23308 33386 23336 34156
rect 23386 34096 23442 34105
rect 23386 34031 23388 34040
rect 23440 34031 23442 34040
rect 23388 34002 23440 34008
rect 23296 33380 23348 33386
rect 23296 33322 23348 33328
rect 23308 33046 23336 33322
rect 23400 33114 23428 34002
rect 23480 33856 23532 33862
rect 23480 33798 23532 33804
rect 23388 33108 23440 33114
rect 23388 33050 23440 33056
rect 23296 33040 23348 33046
rect 23296 32982 23348 32988
rect 23492 32570 23520 33798
rect 23584 33658 23612 34167
rect 23572 33652 23624 33658
rect 23572 33594 23624 33600
rect 23480 32564 23532 32570
rect 23480 32506 23532 32512
rect 23112 32428 23164 32434
rect 23112 32370 23164 32376
rect 23020 32360 23072 32366
rect 23020 32302 23072 32308
rect 23124 31958 23152 32370
rect 23492 32026 23520 32506
rect 23480 32020 23532 32026
rect 23400 31980 23480 32008
rect 23112 31952 23164 31958
rect 23112 31894 23164 31900
rect 22928 31884 22980 31890
rect 22928 31826 22980 31832
rect 22940 31278 22968 31826
rect 22928 31272 22980 31278
rect 22926 31240 22928 31249
rect 22980 31240 22982 31249
rect 22926 31175 22982 31184
rect 23400 30734 23428 31980
rect 23480 31962 23532 31968
rect 23676 31890 23704 37266
rect 23768 34542 23796 37862
rect 23848 37732 23900 37738
rect 23848 37674 23900 37680
rect 23756 34536 23808 34542
rect 23756 34478 23808 34484
rect 23754 33280 23810 33289
rect 23754 33215 23810 33224
rect 23768 33114 23796 33215
rect 23756 33108 23808 33114
rect 23756 33050 23808 33056
rect 23756 32904 23808 32910
rect 23756 32846 23808 32852
rect 23480 31884 23532 31890
rect 23480 31826 23532 31832
rect 23664 31884 23716 31890
rect 23664 31826 23716 31832
rect 23388 30728 23440 30734
rect 23388 30670 23440 30676
rect 23388 28076 23440 28082
rect 23492 28064 23520 31826
rect 23768 31278 23796 32846
rect 23756 31272 23808 31278
rect 23756 31214 23808 31220
rect 23768 30938 23796 31214
rect 23756 30932 23808 30938
rect 23756 30874 23808 30880
rect 23440 28036 23520 28064
rect 23388 28018 23440 28024
rect 23664 28008 23716 28014
rect 23664 27950 23716 27956
rect 22926 21176 22982 21185
rect 22926 21111 22982 21120
rect 22940 21010 22968 21111
rect 22928 21004 22980 21010
rect 22928 20946 22980 20952
rect 22940 20602 22968 20946
rect 22928 20596 22980 20602
rect 22928 20538 22980 20544
rect 23676 16794 23704 27950
rect 23860 23225 23888 37674
rect 24032 37324 24084 37330
rect 24032 37266 24084 37272
rect 23938 37088 23994 37097
rect 24044 37074 24072 37266
rect 23994 37046 24072 37074
rect 23938 37023 23994 37032
rect 23952 36922 23980 37023
rect 23940 36916 23992 36922
rect 23940 36858 23992 36864
rect 23938 36136 23994 36145
rect 23938 36071 23994 36080
rect 23952 35698 23980 36071
rect 23940 35692 23992 35698
rect 23940 35634 23992 35640
rect 24032 32904 24084 32910
rect 24032 32846 24084 32852
rect 24044 32230 24072 32846
rect 24032 32224 24084 32230
rect 24032 32166 24084 32172
rect 23938 31376 23994 31385
rect 23938 31311 23940 31320
rect 23992 31311 23994 31320
rect 23940 31282 23992 31288
rect 23846 23216 23902 23225
rect 23846 23151 23902 23160
rect 23756 20800 23808 20806
rect 23754 20768 23756 20777
rect 24044 20777 24072 32166
rect 24136 28665 24164 40326
rect 24122 28656 24178 28665
rect 24122 28591 24178 28600
rect 23808 20768 23810 20777
rect 23754 20703 23810 20712
rect 24030 20768 24086 20777
rect 24030 20703 24086 20712
rect 24228 19281 24256 44220
rect 24504 43761 24532 45358
rect 24490 43752 24546 43761
rect 24490 43687 24546 43696
rect 24596 42770 24624 55916
rect 24860 55616 24912 55622
rect 24860 55558 24912 55564
rect 24676 55140 24728 55146
rect 24676 55082 24728 55088
rect 24688 54874 24716 55082
rect 24872 54890 24900 55558
rect 24676 54868 24728 54874
rect 24676 54810 24728 54816
rect 24780 54862 24900 54890
rect 24780 54806 24808 54862
rect 24768 54800 24820 54806
rect 24768 54742 24820 54748
rect 24676 54732 24728 54738
rect 24676 54674 24728 54680
rect 24688 48362 24716 54674
rect 24768 53440 24820 53446
rect 24768 53382 24820 53388
rect 24780 53038 24808 53382
rect 24768 53032 24820 53038
rect 24768 52974 24820 52980
rect 24780 51270 24808 52974
rect 24872 52154 24900 54862
rect 24860 52148 24912 52154
rect 24860 52090 24912 52096
rect 24872 51882 24900 52090
rect 24860 51876 24912 51882
rect 24860 51818 24912 51824
rect 24768 51264 24820 51270
rect 24768 51206 24820 51212
rect 24780 50930 24808 51206
rect 24768 50924 24820 50930
rect 24768 50866 24820 50872
rect 24768 49292 24820 49298
rect 24768 49234 24820 49240
rect 24780 48890 24808 49234
rect 24768 48884 24820 48890
rect 24768 48826 24820 48832
rect 24688 48334 24808 48362
rect 24676 48204 24728 48210
rect 24676 48146 24728 48152
rect 24688 47802 24716 48146
rect 24676 47796 24728 47802
rect 24676 47738 24728 47744
rect 24780 47240 24808 48334
rect 24860 48000 24912 48006
rect 24858 47968 24860 47977
rect 24912 47968 24914 47977
rect 24858 47903 24914 47912
rect 24688 47212 24808 47240
rect 24688 46170 24716 47212
rect 24768 47116 24820 47122
rect 24768 47058 24820 47064
rect 24780 46492 24808 47058
rect 24860 46504 24912 46510
rect 24780 46464 24860 46492
rect 24860 46446 24912 46452
rect 24768 46368 24820 46374
rect 24768 46310 24820 46316
rect 24676 46164 24728 46170
rect 24676 46106 24728 46112
rect 24688 45558 24716 46106
rect 24676 45552 24728 45558
rect 24676 45494 24728 45500
rect 24676 45280 24728 45286
rect 24676 45222 24728 45228
rect 24688 44470 24716 45222
rect 24780 44470 24808 46310
rect 24860 45892 24912 45898
rect 24860 45834 24912 45840
rect 24872 45082 24900 45834
rect 24860 45076 24912 45082
rect 24860 45018 24912 45024
rect 24676 44464 24728 44470
rect 24676 44406 24728 44412
rect 24768 44464 24820 44470
rect 24768 44406 24820 44412
rect 24860 44396 24912 44402
rect 24860 44338 24912 44344
rect 24676 44328 24728 44334
rect 24676 44270 24728 44276
rect 24688 43897 24716 44270
rect 24872 44248 24900 44338
rect 24780 44220 24900 44248
rect 24674 43888 24730 43897
rect 24674 43823 24730 43832
rect 24688 43654 24716 43823
rect 24676 43648 24728 43654
rect 24676 43590 24728 43596
rect 24584 42764 24636 42770
rect 24584 42706 24636 42712
rect 24308 42560 24360 42566
rect 24308 42502 24360 42508
rect 24320 42158 24348 42502
rect 24308 42152 24360 42158
rect 24308 42094 24360 42100
rect 24306 41848 24362 41857
rect 24596 41818 24624 42706
rect 24780 42378 24808 44220
rect 24860 43240 24912 43246
rect 24860 43182 24912 43188
rect 24688 42350 24808 42378
rect 24688 41857 24716 42350
rect 24768 42288 24820 42294
rect 24768 42230 24820 42236
rect 24674 41848 24730 41857
rect 24306 41783 24362 41792
rect 24584 41812 24636 41818
rect 24320 41002 24348 41783
rect 24674 41783 24730 41792
rect 24584 41754 24636 41760
rect 24584 41676 24636 41682
rect 24584 41618 24636 41624
rect 24400 41608 24452 41614
rect 24400 41550 24452 41556
rect 24308 40996 24360 41002
rect 24308 40938 24360 40944
rect 24306 40896 24362 40905
rect 24306 40831 24362 40840
rect 24320 35193 24348 40831
rect 24306 35184 24362 35193
rect 24306 35119 24362 35128
rect 24320 34785 24348 35119
rect 24306 34776 24362 34785
rect 24306 34711 24362 34720
rect 24308 34400 24360 34406
rect 24308 34342 24360 34348
rect 24320 33862 24348 34342
rect 24308 33856 24360 33862
rect 24308 33798 24360 33804
rect 24320 32978 24348 33798
rect 24308 32972 24360 32978
rect 24308 32914 24360 32920
rect 24214 19272 24270 19281
rect 24214 19207 24270 19216
rect 23664 16788 23716 16794
rect 23664 16730 23716 16736
rect 22834 10704 22890 10713
rect 22834 10639 22890 10648
rect 24412 6905 24440 41550
rect 24596 41449 24624 41618
rect 24688 41614 24716 41783
rect 24676 41608 24728 41614
rect 24676 41550 24728 41556
rect 24582 41440 24638 41449
rect 24582 41375 24638 41384
rect 24676 40996 24728 41002
rect 24676 40938 24728 40944
rect 24492 40588 24544 40594
rect 24492 40530 24544 40536
rect 24504 39914 24532 40530
rect 24584 40452 24636 40458
rect 24584 40394 24636 40400
rect 24596 40050 24624 40394
rect 24584 40044 24636 40050
rect 24584 39986 24636 39992
rect 24492 39908 24544 39914
rect 24492 39850 24544 39856
rect 24504 39642 24532 39850
rect 24596 39846 24624 39986
rect 24584 39840 24636 39846
rect 24584 39782 24636 39788
rect 24492 39636 24544 39642
rect 24492 39578 24544 39584
rect 24596 39506 24624 39782
rect 24688 39642 24716 40938
rect 24676 39636 24728 39642
rect 24676 39578 24728 39584
rect 24584 39500 24636 39506
rect 24584 39442 24636 39448
rect 24490 39128 24546 39137
rect 24490 39063 24492 39072
rect 24544 39063 24546 39072
rect 24492 39034 24544 39040
rect 24780 38321 24808 42230
rect 24766 38312 24822 38321
rect 24766 38247 24822 38256
rect 24768 37800 24820 37806
rect 24768 37742 24820 37748
rect 24676 37256 24728 37262
rect 24780 37210 24808 37742
rect 24728 37204 24808 37210
rect 24676 37198 24808 37204
rect 24688 37182 24808 37198
rect 24780 36922 24808 37182
rect 24768 36916 24820 36922
rect 24768 36858 24820 36864
rect 24676 32224 24728 32230
rect 24676 32166 24728 32172
rect 24688 31278 24716 32166
rect 24676 31272 24728 31278
rect 24676 31214 24728 31220
rect 24398 6896 24454 6905
rect 24398 6831 24454 6840
rect 24872 5273 24900 43182
rect 24964 34950 24992 61231
rect 25504 60852 25556 60858
rect 25504 60794 25556 60800
rect 25042 55176 25098 55185
rect 25042 55111 25098 55120
rect 25056 46560 25084 55111
rect 25410 53816 25466 53825
rect 25410 53751 25466 53760
rect 25318 52456 25374 52465
rect 25318 52391 25374 52400
rect 25226 51640 25282 51649
rect 25226 51575 25282 51584
rect 25136 50720 25188 50726
rect 25136 50662 25188 50668
rect 25148 49298 25176 50662
rect 25240 50425 25268 51575
rect 25226 50416 25282 50425
rect 25226 50351 25282 50360
rect 25228 49632 25280 49638
rect 25228 49574 25280 49580
rect 25136 49292 25188 49298
rect 25136 49234 25188 49240
rect 25240 48793 25268 49574
rect 25226 48784 25282 48793
rect 25226 48719 25282 48728
rect 25240 48686 25268 48719
rect 25228 48680 25280 48686
rect 25228 48622 25280 48628
rect 25136 48272 25188 48278
rect 25134 48240 25136 48249
rect 25188 48240 25190 48249
rect 25134 48175 25190 48184
rect 25332 47122 25360 52391
rect 25424 50402 25452 53751
rect 25516 51610 25544 60794
rect 25504 51604 25556 51610
rect 25504 51546 25556 51552
rect 25424 50374 25544 50402
rect 25410 50280 25466 50289
rect 25410 50215 25466 50224
rect 25424 48890 25452 50215
rect 25412 48884 25464 48890
rect 25412 48826 25464 48832
rect 25412 47456 25464 47462
rect 25412 47398 25464 47404
rect 25320 47116 25372 47122
rect 25320 47058 25372 47064
rect 25056 46532 25268 46560
rect 25136 46436 25188 46442
rect 25136 46378 25188 46384
rect 25044 46368 25096 46374
rect 25044 46310 25096 46316
rect 25056 45422 25084 46310
rect 25148 45665 25176 46378
rect 25134 45656 25190 45665
rect 25134 45591 25190 45600
rect 25044 45416 25096 45422
rect 25044 45358 25096 45364
rect 25134 45384 25190 45393
rect 25134 45319 25136 45328
rect 25188 45319 25190 45328
rect 25136 45290 25188 45296
rect 25044 45280 25096 45286
rect 25044 45222 25096 45228
rect 25056 44577 25084 45222
rect 25148 44878 25176 45290
rect 25240 45286 25268 46532
rect 25332 46170 25360 47058
rect 25320 46164 25372 46170
rect 25320 46106 25372 46112
rect 25228 45280 25280 45286
rect 25228 45222 25280 45228
rect 25424 45098 25452 47398
rect 25240 45070 25452 45098
rect 25136 44872 25188 44878
rect 25136 44814 25188 44820
rect 25042 44568 25098 44577
rect 25148 44538 25176 44814
rect 25042 44503 25098 44512
rect 25136 44532 25188 44538
rect 25136 44474 25188 44480
rect 25044 44464 25096 44470
rect 25044 44406 25096 44412
rect 25056 41857 25084 44406
rect 25136 44260 25188 44266
rect 25136 44202 25188 44208
rect 25148 43761 25176 44202
rect 25134 43752 25190 43761
rect 25134 43687 25190 43696
rect 25136 42560 25188 42566
rect 25136 42502 25188 42508
rect 25042 41848 25098 41857
rect 25042 41783 25098 41792
rect 25044 41540 25096 41546
rect 25044 41482 25096 41488
rect 25056 40730 25084 41482
rect 25044 40724 25096 40730
rect 25044 40666 25096 40672
rect 25148 40594 25176 42502
rect 25136 40588 25188 40594
rect 25136 40530 25188 40536
rect 25148 40050 25176 40530
rect 25136 40044 25188 40050
rect 25136 39986 25188 39992
rect 25134 35456 25190 35465
rect 25134 35391 25190 35400
rect 24952 34944 25004 34950
rect 24952 34886 25004 34892
rect 24952 34740 25004 34746
rect 24952 34682 25004 34688
rect 24964 33998 24992 34682
rect 25044 34604 25096 34610
rect 25044 34546 25096 34552
rect 25056 34105 25084 34546
rect 25042 34096 25098 34105
rect 25042 34031 25098 34040
rect 24952 33992 25004 33998
rect 24952 33934 25004 33940
rect 25044 33992 25096 33998
rect 25044 33934 25096 33940
rect 24964 33590 24992 33934
rect 25056 33658 25084 33934
rect 25044 33652 25096 33658
rect 25044 33594 25096 33600
rect 24952 33584 25004 33590
rect 24952 33526 25004 33532
rect 25148 33114 25176 35391
rect 25136 33108 25188 33114
rect 25136 33050 25188 33056
rect 24950 32056 25006 32065
rect 24950 31991 25006 32000
rect 24964 30297 24992 31991
rect 25044 31136 25096 31142
rect 25044 31078 25096 31084
rect 24950 30288 25006 30297
rect 24950 30223 25006 30232
rect 25056 26081 25084 31078
rect 25134 27670 25190 27679
rect 25134 27605 25190 27614
rect 25148 26246 25176 27605
rect 25136 26240 25188 26246
rect 25136 26182 25188 26188
rect 25042 26072 25098 26081
rect 25042 26007 25098 26016
rect 25044 21412 25096 21418
rect 25044 21354 25096 21360
rect 25056 13190 25084 21354
rect 25044 13184 25096 13190
rect 25044 13126 25096 13132
rect 25240 11665 25268 45070
rect 25412 44940 25464 44946
rect 25412 44882 25464 44888
rect 25424 44849 25452 44882
rect 25410 44840 25466 44849
rect 25410 44775 25466 44784
rect 25318 44568 25374 44577
rect 25318 44503 25374 44512
rect 25332 41834 25360 44503
rect 25424 43994 25452 44775
rect 25412 43988 25464 43994
rect 25412 43930 25464 43936
rect 25410 43072 25466 43081
rect 25410 43007 25466 43016
rect 25424 41993 25452 43007
rect 25410 41984 25466 41993
rect 25410 41919 25466 41928
rect 25332 41806 25452 41834
rect 25320 41064 25372 41070
rect 25320 41006 25372 41012
rect 25332 35680 25360 41006
rect 25424 38010 25452 41806
rect 25516 41585 25544 50374
rect 25608 42770 25636 61775
rect 25700 52714 25728 61934
rect 25792 61810 25820 63271
rect 25884 62898 25912 64631
rect 25956 64220 26252 64240
rect 26012 64218 26036 64220
rect 26092 64218 26116 64220
rect 26172 64218 26196 64220
rect 26034 64166 26036 64218
rect 26098 64166 26110 64218
rect 26172 64166 26174 64218
rect 26012 64164 26036 64166
rect 26092 64164 26116 64166
rect 26172 64164 26196 64166
rect 25956 64144 26252 64164
rect 27540 63617 27568 64790
rect 27526 63608 27582 63617
rect 27526 63543 27582 63552
rect 25956 63132 26252 63152
rect 26012 63130 26036 63132
rect 26092 63130 26116 63132
rect 26172 63130 26196 63132
rect 26034 63078 26036 63130
rect 26098 63078 26110 63130
rect 26172 63078 26174 63130
rect 26012 63076 26036 63078
rect 26092 63076 26116 63078
rect 26172 63076 26196 63078
rect 25956 63056 26252 63076
rect 27816 62898 27844 79070
rect 29012 74662 29040 79200
rect 29000 74656 29052 74662
rect 29000 74598 29052 74604
rect 29932 72593 29960 79200
rect 29918 72584 29974 72593
rect 29918 72519 29974 72528
rect 27896 70372 27948 70378
rect 27896 70314 27948 70320
rect 25872 62892 25924 62898
rect 25872 62834 25924 62840
rect 27620 62892 27672 62898
rect 27620 62834 27672 62840
rect 27804 62892 27856 62898
rect 27804 62834 27856 62840
rect 26148 62824 26200 62830
rect 26148 62766 26200 62772
rect 26160 62490 26188 62766
rect 25872 62484 25924 62490
rect 25872 62426 25924 62432
rect 26148 62484 26200 62490
rect 26148 62426 26200 62432
rect 25780 61804 25832 61810
rect 25780 61746 25832 61752
rect 25884 61742 25912 62426
rect 25956 62044 26252 62064
rect 26012 62042 26036 62044
rect 26092 62042 26116 62044
rect 26172 62042 26196 62044
rect 26034 61990 26036 62042
rect 26098 61990 26110 62042
rect 26172 61990 26174 62042
rect 26012 61988 26036 61990
rect 26092 61988 26116 61990
rect 26172 61988 26196 61990
rect 25956 61968 26252 61988
rect 26698 61976 26754 61985
rect 26698 61911 26754 61920
rect 25872 61736 25924 61742
rect 25872 61678 25924 61684
rect 25884 61402 25912 61678
rect 25872 61396 25924 61402
rect 25872 61338 25924 61344
rect 25778 59664 25834 59673
rect 25778 59599 25834 59608
rect 25792 56506 25820 59599
rect 25780 56500 25832 56506
rect 25780 56442 25832 56448
rect 25792 56302 25820 56442
rect 25884 56370 25912 61338
rect 26712 61334 26740 61911
rect 26700 61328 26752 61334
rect 26700 61270 26752 61276
rect 27344 61260 27396 61266
rect 27344 61202 27396 61208
rect 26516 61192 26568 61198
rect 26516 61134 26568 61140
rect 26884 61192 26936 61198
rect 26884 61134 26936 61140
rect 25956 60956 26252 60976
rect 26012 60954 26036 60956
rect 26092 60954 26116 60956
rect 26172 60954 26196 60956
rect 26034 60902 26036 60954
rect 26098 60902 26110 60954
rect 26172 60902 26174 60954
rect 26012 60900 26036 60902
rect 26092 60900 26116 60902
rect 26172 60900 26196 60902
rect 25956 60880 26252 60900
rect 26528 60722 26556 61134
rect 26896 60858 26924 61134
rect 27356 60858 27384 61202
rect 26884 60852 26936 60858
rect 26884 60794 26936 60800
rect 27344 60852 27396 60858
rect 27344 60794 27396 60800
rect 26516 60716 26568 60722
rect 26516 60658 26568 60664
rect 25956 59868 26252 59888
rect 26012 59866 26036 59868
rect 26092 59866 26116 59868
rect 26172 59866 26196 59868
rect 26034 59814 26036 59866
rect 26098 59814 26110 59866
rect 26172 59814 26174 59866
rect 26012 59812 26036 59814
rect 26092 59812 26116 59814
rect 26172 59812 26196 59814
rect 25956 59792 26252 59812
rect 26528 59401 26556 60658
rect 26514 59392 26570 59401
rect 26514 59327 26570 59336
rect 25956 58780 26252 58800
rect 26012 58778 26036 58780
rect 26092 58778 26116 58780
rect 26172 58778 26196 58780
rect 26034 58726 26036 58778
rect 26098 58726 26110 58778
rect 26172 58726 26174 58778
rect 26012 58724 26036 58726
rect 26092 58724 26116 58726
rect 26172 58724 26196 58726
rect 25956 58704 26252 58724
rect 25956 57692 26252 57712
rect 26012 57690 26036 57692
rect 26092 57690 26116 57692
rect 26172 57690 26196 57692
rect 26034 57638 26036 57690
rect 26098 57638 26110 57690
rect 26172 57638 26174 57690
rect 26012 57636 26036 57638
rect 26092 57636 26116 57638
rect 26172 57636 26196 57638
rect 25956 57616 26252 57636
rect 25956 56604 26252 56624
rect 26012 56602 26036 56604
rect 26092 56602 26116 56604
rect 26172 56602 26196 56604
rect 26034 56550 26036 56602
rect 26098 56550 26110 56602
rect 26172 56550 26174 56602
rect 26012 56548 26036 56550
rect 26092 56548 26116 56550
rect 26172 56548 26196 56550
rect 25956 56528 26252 56548
rect 25962 56400 26018 56409
rect 25872 56364 25924 56370
rect 25962 56335 26018 56344
rect 25872 56306 25924 56312
rect 25780 56296 25832 56302
rect 25780 56238 25832 56244
rect 25884 55962 25912 56306
rect 25872 55956 25924 55962
rect 25872 55898 25924 55904
rect 25976 55706 26004 56335
rect 25884 55678 26004 55706
rect 26332 55752 26384 55758
rect 26332 55694 26384 55700
rect 25884 54194 25912 55678
rect 25956 55516 26252 55536
rect 26012 55514 26036 55516
rect 26092 55514 26116 55516
rect 26172 55514 26196 55516
rect 26034 55462 26036 55514
rect 26098 55462 26110 55514
rect 26172 55462 26174 55514
rect 26012 55460 26036 55462
rect 26092 55460 26116 55462
rect 26172 55460 26196 55462
rect 25956 55440 26252 55460
rect 26240 55208 26292 55214
rect 26344 55196 26372 55694
rect 27632 55298 27660 62834
rect 27804 62756 27856 62762
rect 27804 62698 27856 62704
rect 27816 61266 27844 62698
rect 27804 61260 27856 61266
rect 27804 61202 27856 61208
rect 27712 56160 27764 56166
rect 27712 56102 27764 56108
rect 27540 55282 27660 55298
rect 27528 55276 27660 55282
rect 27580 55270 27660 55276
rect 27528 55218 27580 55224
rect 26292 55168 26372 55196
rect 26240 55150 26292 55156
rect 26344 54534 26372 55168
rect 26606 55040 26662 55049
rect 26606 54975 26662 54984
rect 26620 54670 26648 54975
rect 27724 54738 27752 56102
rect 27712 54732 27764 54738
rect 27712 54674 27764 54680
rect 26608 54664 26660 54670
rect 26608 54606 26660 54612
rect 26976 54664 27028 54670
rect 26976 54606 27028 54612
rect 27528 54664 27580 54670
rect 27528 54606 27580 54612
rect 26332 54528 26384 54534
rect 26332 54470 26384 54476
rect 25956 54428 26252 54448
rect 26012 54426 26036 54428
rect 26092 54426 26116 54428
rect 26172 54426 26196 54428
rect 26034 54374 26036 54426
rect 26098 54374 26110 54426
rect 26172 54374 26174 54426
rect 26012 54372 26036 54374
rect 26092 54372 26116 54374
rect 26172 54372 26196 54374
rect 25956 54352 26252 54372
rect 25872 54188 25924 54194
rect 25872 54130 25924 54136
rect 26344 54126 26372 54470
rect 25964 54120 26016 54126
rect 25964 54062 26016 54068
rect 26332 54120 26384 54126
rect 26332 54062 26384 54068
rect 25976 53582 26004 54062
rect 26620 53786 26648 54606
rect 26608 53780 26660 53786
rect 26608 53722 26660 53728
rect 25964 53576 26016 53582
rect 25964 53518 26016 53524
rect 25956 53340 26252 53360
rect 26012 53338 26036 53340
rect 26092 53338 26116 53340
rect 26172 53338 26196 53340
rect 26034 53286 26036 53338
rect 26098 53286 26110 53338
rect 26172 53286 26174 53338
rect 26012 53284 26036 53286
rect 26092 53284 26116 53286
rect 26172 53284 26196 53286
rect 25956 53264 26252 53284
rect 25700 52686 25820 52714
rect 25686 52592 25742 52601
rect 25686 52527 25742 52536
rect 25700 51785 25728 52527
rect 25792 52329 25820 52686
rect 25778 52320 25834 52329
rect 25778 52255 25834 52264
rect 25956 52252 26252 52272
rect 26012 52250 26036 52252
rect 26092 52250 26116 52252
rect 26172 52250 26196 52252
rect 26034 52198 26036 52250
rect 26098 52198 26110 52250
rect 26172 52198 26174 52250
rect 26012 52196 26036 52198
rect 26092 52196 26116 52198
rect 26172 52196 26196 52198
rect 25956 52176 26252 52196
rect 25686 51776 25742 51785
rect 25686 51711 25742 51720
rect 25688 51604 25740 51610
rect 25688 51546 25740 51552
rect 25700 47122 25728 51546
rect 25780 51264 25832 51270
rect 25780 51206 25832 51212
rect 25792 47666 25820 51206
rect 25956 51164 26252 51184
rect 26012 51162 26036 51164
rect 26092 51162 26116 51164
rect 26172 51162 26196 51164
rect 26034 51110 26036 51162
rect 26098 51110 26110 51162
rect 26172 51110 26174 51162
rect 26012 51108 26036 51110
rect 26092 51108 26116 51110
rect 26172 51108 26196 51110
rect 25956 51088 26252 51108
rect 25956 50076 26252 50096
rect 26012 50074 26036 50076
rect 26092 50074 26116 50076
rect 26172 50074 26196 50076
rect 26034 50022 26036 50074
rect 26098 50022 26110 50074
rect 26172 50022 26174 50074
rect 26012 50020 26036 50022
rect 26092 50020 26116 50022
rect 26172 50020 26196 50022
rect 25956 50000 26252 50020
rect 25956 48988 26252 49008
rect 26012 48986 26036 48988
rect 26092 48986 26116 48988
rect 26172 48986 26196 48988
rect 26034 48934 26036 48986
rect 26098 48934 26110 48986
rect 26172 48934 26174 48986
rect 26012 48932 26036 48934
rect 26092 48932 26116 48934
rect 26172 48932 26196 48934
rect 25956 48912 26252 48932
rect 26332 48000 26384 48006
rect 26332 47942 26384 47948
rect 25956 47900 26252 47920
rect 26012 47898 26036 47900
rect 26092 47898 26116 47900
rect 26172 47898 26196 47900
rect 26034 47846 26036 47898
rect 26098 47846 26110 47898
rect 26172 47846 26174 47898
rect 26012 47844 26036 47846
rect 26092 47844 26116 47846
rect 26172 47844 26196 47846
rect 25956 47824 26252 47844
rect 26344 47666 26372 47942
rect 26698 47696 26754 47705
rect 25780 47660 25832 47666
rect 25780 47602 25832 47608
rect 26332 47660 26384 47666
rect 26698 47631 26754 47640
rect 26884 47660 26936 47666
rect 26332 47602 26384 47608
rect 25872 47592 25924 47598
rect 25872 47534 25924 47540
rect 25884 47297 25912 47534
rect 25870 47288 25926 47297
rect 26712 47258 26740 47631
rect 26884 47602 26936 47608
rect 25870 47223 25926 47232
rect 26700 47252 26752 47258
rect 25688 47116 25740 47122
rect 25688 47058 25740 47064
rect 25686 47016 25742 47025
rect 25686 46951 25742 46960
rect 25596 42764 25648 42770
rect 25596 42706 25648 42712
rect 25608 42294 25636 42706
rect 25596 42288 25648 42294
rect 25596 42230 25648 42236
rect 25502 41576 25558 41585
rect 25502 41511 25558 41520
rect 25502 38584 25558 38593
rect 25502 38519 25558 38528
rect 25412 38004 25464 38010
rect 25412 37946 25464 37952
rect 25516 37466 25544 38519
rect 25594 38176 25650 38185
rect 25594 38111 25650 38120
rect 25504 37460 25556 37466
rect 25504 37402 25556 37408
rect 25332 35652 25452 35680
rect 25320 35556 25372 35562
rect 25320 35498 25372 35504
rect 25332 34746 25360 35498
rect 25320 34740 25372 34746
rect 25320 34682 25372 34688
rect 25318 34640 25374 34649
rect 25318 34575 25374 34584
rect 25332 34066 25360 34575
rect 25320 34060 25372 34066
rect 25320 34002 25372 34008
rect 25332 33522 25360 34002
rect 25320 33516 25372 33522
rect 25320 33458 25372 33464
rect 25424 27713 25452 35652
rect 25504 34944 25556 34950
rect 25504 34886 25556 34892
rect 25516 33658 25544 34886
rect 25504 33652 25556 33658
rect 25504 33594 25556 33600
rect 25608 33425 25636 38111
rect 25700 33810 25728 46951
rect 25884 46918 25912 47223
rect 26700 47194 26752 47200
rect 26514 47152 26570 47161
rect 26514 47087 26516 47096
rect 26568 47087 26570 47096
rect 26516 47058 26568 47064
rect 25872 46912 25924 46918
rect 25872 46854 25924 46860
rect 25884 46492 25912 46854
rect 25956 46812 26252 46832
rect 26012 46810 26036 46812
rect 26092 46810 26116 46812
rect 26172 46810 26196 46812
rect 26034 46758 26036 46810
rect 26098 46758 26110 46810
rect 26172 46758 26174 46810
rect 26012 46756 26036 46758
rect 26092 46756 26116 46758
rect 26172 46756 26196 46758
rect 25956 46736 26252 46756
rect 26528 46714 26556 47058
rect 26516 46708 26568 46714
rect 26516 46650 26568 46656
rect 25964 46504 26016 46510
rect 25884 46464 25964 46492
rect 25964 46446 26016 46452
rect 25780 46096 25832 46102
rect 25780 46038 25832 46044
rect 25792 45286 25820 46038
rect 25976 46034 26004 46446
rect 26516 46436 26568 46442
rect 26516 46378 26568 46384
rect 26332 46368 26384 46374
rect 26332 46310 26384 46316
rect 25964 46028 26016 46034
rect 25964 45970 26016 45976
rect 25872 45824 25924 45830
rect 25872 45766 25924 45772
rect 25780 45280 25832 45286
rect 25780 45222 25832 45228
rect 25792 45082 25820 45222
rect 25780 45076 25832 45082
rect 25780 45018 25832 45024
rect 25884 44962 25912 45766
rect 25956 45724 26252 45744
rect 26012 45722 26036 45724
rect 26092 45722 26116 45724
rect 26172 45722 26196 45724
rect 26034 45670 26036 45722
rect 26098 45670 26110 45722
rect 26172 45670 26174 45722
rect 26012 45668 26036 45670
rect 26092 45668 26116 45670
rect 26172 45668 26196 45670
rect 25956 45648 26252 45668
rect 26344 45608 26372 46310
rect 26528 45937 26556 46378
rect 26514 45928 26570 45937
rect 26514 45863 26570 45872
rect 26252 45580 26372 45608
rect 26056 45280 26108 45286
rect 26056 45222 26108 45228
rect 25792 44934 25912 44962
rect 26068 44946 26096 45222
rect 26252 44996 26280 45580
rect 26422 45520 26478 45529
rect 26422 45455 26478 45464
rect 26332 45348 26384 45354
rect 26332 45290 26384 45296
rect 26344 45121 26372 45290
rect 26330 45112 26386 45121
rect 26330 45047 26386 45056
rect 26252 44968 26372 44996
rect 26056 44940 26108 44946
rect 25792 43450 25820 44934
rect 26056 44882 26108 44888
rect 25956 44636 26252 44656
rect 26012 44634 26036 44636
rect 26092 44634 26116 44636
rect 26172 44634 26196 44636
rect 26034 44582 26036 44634
rect 26098 44582 26110 44634
rect 26172 44582 26174 44634
rect 26012 44580 26036 44582
rect 26092 44580 26116 44582
rect 26172 44580 26196 44582
rect 25956 44560 26252 44580
rect 25872 43784 25924 43790
rect 25872 43726 25924 43732
rect 25780 43444 25832 43450
rect 25780 43386 25832 43392
rect 25780 42696 25832 42702
rect 25780 42638 25832 42644
rect 25792 41818 25820 42638
rect 25884 42226 25912 43726
rect 25956 43548 26252 43568
rect 26012 43546 26036 43548
rect 26092 43546 26116 43548
rect 26172 43546 26196 43548
rect 26034 43494 26036 43546
rect 26098 43494 26110 43546
rect 26172 43494 26174 43546
rect 26012 43492 26036 43494
rect 26092 43492 26116 43494
rect 26172 43492 26196 43494
rect 25956 43472 26252 43492
rect 26344 43246 26372 44968
rect 26436 44402 26464 45455
rect 26608 45280 26660 45286
rect 26608 45222 26660 45228
rect 26620 45014 26648 45222
rect 26700 45076 26752 45082
rect 26700 45018 26752 45024
rect 26608 45008 26660 45014
rect 26608 44950 26660 44956
rect 26516 44872 26568 44878
rect 26620 44849 26648 44950
rect 26516 44814 26568 44820
rect 26606 44840 26662 44849
rect 26424 44396 26476 44402
rect 26424 44338 26476 44344
rect 26528 43926 26556 44814
rect 26606 44775 26662 44784
rect 26608 44396 26660 44402
rect 26608 44338 26660 44344
rect 26516 43920 26568 43926
rect 26516 43862 26568 43868
rect 26528 43450 26556 43862
rect 26516 43444 26568 43450
rect 26516 43386 26568 43392
rect 26332 43240 26384 43246
rect 26332 43182 26384 43188
rect 26620 42888 26648 44338
rect 26712 44334 26740 45018
rect 26792 44940 26844 44946
rect 26792 44882 26844 44888
rect 26700 44328 26752 44334
rect 26700 44270 26752 44276
rect 26712 43994 26740 44270
rect 26804 43994 26832 44882
rect 26896 44742 26924 47602
rect 26884 44736 26936 44742
rect 26884 44678 26936 44684
rect 26896 44402 26924 44678
rect 26884 44396 26936 44402
rect 26884 44338 26936 44344
rect 26700 43988 26752 43994
rect 26700 43930 26752 43936
rect 26792 43988 26844 43994
rect 26792 43930 26844 43936
rect 26712 43450 26740 43930
rect 26804 43858 26832 43930
rect 26884 43920 26936 43926
rect 26882 43888 26884 43897
rect 26936 43888 26938 43897
rect 26792 43852 26844 43858
rect 26882 43823 26938 43832
rect 26792 43794 26844 43800
rect 26700 43444 26752 43450
rect 26700 43386 26752 43392
rect 26804 42906 26832 43794
rect 26896 43382 26924 43823
rect 26884 43376 26936 43382
rect 26884 43318 26936 43324
rect 26528 42860 26648 42888
rect 26792 42900 26844 42906
rect 25956 42460 26252 42480
rect 26012 42458 26036 42460
rect 26092 42458 26116 42460
rect 26172 42458 26196 42460
rect 26034 42406 26036 42458
rect 26098 42406 26110 42458
rect 26172 42406 26174 42458
rect 26012 42404 26036 42406
rect 26092 42404 26116 42406
rect 26172 42404 26196 42406
rect 25956 42384 26252 42404
rect 25964 42288 26016 42294
rect 25962 42256 25964 42265
rect 26016 42256 26018 42265
rect 25872 42220 25924 42226
rect 26528 42226 26556 42860
rect 26792 42842 26844 42848
rect 26608 42764 26660 42770
rect 26608 42706 26660 42712
rect 26620 42265 26648 42706
rect 26792 42560 26844 42566
rect 26792 42502 26844 42508
rect 26804 42362 26832 42502
rect 26792 42356 26844 42362
rect 26792 42298 26844 42304
rect 26606 42256 26662 42265
rect 25962 42191 26018 42200
rect 26332 42220 26384 42226
rect 25872 42162 25924 42168
rect 26332 42162 26384 42168
rect 26516 42220 26568 42226
rect 26606 42191 26662 42200
rect 26516 42162 26568 42168
rect 25872 42084 25924 42090
rect 25872 42026 25924 42032
rect 25780 41812 25832 41818
rect 25780 41754 25832 41760
rect 25884 40934 25912 42026
rect 26344 41818 26372 42162
rect 26514 42120 26570 42129
rect 26514 42055 26570 42064
rect 26332 41812 26384 41818
rect 26332 41754 26384 41760
rect 26528 41750 26556 42055
rect 26516 41744 26568 41750
rect 26516 41686 26568 41692
rect 25956 41372 26252 41392
rect 26012 41370 26036 41372
rect 26092 41370 26116 41372
rect 26172 41370 26196 41372
rect 26034 41318 26036 41370
rect 26098 41318 26110 41370
rect 26172 41318 26174 41370
rect 26012 41316 26036 41318
rect 26092 41316 26116 41318
rect 26172 41316 26196 41318
rect 25956 41296 26252 41316
rect 26896 41274 26924 43318
rect 26884 41268 26936 41274
rect 26884 41210 26936 41216
rect 25872 40928 25924 40934
rect 25872 40870 25924 40876
rect 25884 40730 25912 40870
rect 25872 40724 25924 40730
rect 25792 40684 25872 40712
rect 25792 38894 25820 40684
rect 25872 40666 25924 40672
rect 25956 40284 26252 40304
rect 26012 40282 26036 40284
rect 26092 40282 26116 40284
rect 26172 40282 26196 40284
rect 26034 40230 26036 40282
rect 26098 40230 26110 40282
rect 26172 40230 26174 40282
rect 26012 40228 26036 40230
rect 26092 40228 26116 40230
rect 26172 40228 26196 40230
rect 25956 40208 26252 40228
rect 25870 40080 25926 40089
rect 25870 40015 25926 40024
rect 25780 38888 25832 38894
rect 25780 38830 25832 38836
rect 25884 36786 25912 40015
rect 25956 39196 26252 39216
rect 26012 39194 26036 39196
rect 26092 39194 26116 39196
rect 26172 39194 26196 39196
rect 26034 39142 26036 39194
rect 26098 39142 26110 39194
rect 26172 39142 26174 39194
rect 26012 39140 26036 39142
rect 26092 39140 26116 39142
rect 26172 39140 26196 39142
rect 25956 39120 26252 39140
rect 26148 38888 26200 38894
rect 26424 38888 26476 38894
rect 26148 38830 26200 38836
rect 26422 38856 26424 38865
rect 26476 38856 26478 38865
rect 26160 38554 26188 38830
rect 26422 38791 26478 38800
rect 26148 38548 26200 38554
rect 26148 38490 26200 38496
rect 26160 38298 26188 38490
rect 26160 38270 26372 38298
rect 25956 38108 26252 38128
rect 26012 38106 26036 38108
rect 26092 38106 26116 38108
rect 26172 38106 26196 38108
rect 26034 38054 26036 38106
rect 26098 38054 26110 38106
rect 26172 38054 26174 38106
rect 26012 38052 26036 38054
rect 26092 38052 26116 38054
rect 26172 38052 26196 38054
rect 25956 38032 26252 38052
rect 26344 37890 26372 38270
rect 26252 37862 26372 37890
rect 26252 37806 26280 37862
rect 26240 37800 26292 37806
rect 26240 37742 26292 37748
rect 26252 37466 26280 37742
rect 26240 37460 26292 37466
rect 26240 37402 26292 37408
rect 25956 37020 26252 37040
rect 26012 37018 26036 37020
rect 26092 37018 26116 37020
rect 26172 37018 26196 37020
rect 26034 36966 26036 37018
rect 26098 36966 26110 37018
rect 26172 36966 26174 37018
rect 26012 36964 26036 36966
rect 26092 36964 26116 36966
rect 26172 36964 26196 36966
rect 25956 36944 26252 36964
rect 25872 36780 25924 36786
rect 25872 36722 25924 36728
rect 26332 36780 26384 36786
rect 26332 36722 26384 36728
rect 26344 36038 26372 36722
rect 26332 36032 26384 36038
rect 26332 35974 26384 35980
rect 25956 35932 26252 35952
rect 26012 35930 26036 35932
rect 26092 35930 26116 35932
rect 26172 35930 26196 35932
rect 26034 35878 26036 35930
rect 26098 35878 26110 35930
rect 26172 35878 26174 35930
rect 26012 35876 26036 35878
rect 26092 35876 26116 35878
rect 26172 35876 26196 35878
rect 25956 35856 26252 35876
rect 26344 35698 26372 35974
rect 26332 35692 26384 35698
rect 26332 35634 26384 35640
rect 26344 34950 26372 35634
rect 26332 34944 26384 34950
rect 26332 34886 26384 34892
rect 25956 34844 26252 34864
rect 26012 34842 26036 34844
rect 26092 34842 26116 34844
rect 26172 34842 26196 34844
rect 26034 34790 26036 34842
rect 26098 34790 26110 34842
rect 26172 34790 26174 34842
rect 26012 34788 26036 34790
rect 26092 34788 26116 34790
rect 26172 34788 26196 34790
rect 25956 34768 26252 34788
rect 26240 34536 26292 34542
rect 26344 34524 26372 34886
rect 26292 34496 26372 34524
rect 26240 34478 26292 34484
rect 26344 33862 26372 34496
rect 26332 33856 26384 33862
rect 25700 33782 25912 33810
rect 26332 33798 26384 33804
rect 25594 33416 25650 33425
rect 25594 33351 25650 33360
rect 25780 31272 25832 31278
rect 25780 31214 25832 31220
rect 25686 30696 25742 30705
rect 25686 30631 25742 30640
rect 25410 27704 25466 27713
rect 25410 27639 25466 27648
rect 25502 26616 25558 26625
rect 25502 26551 25558 26560
rect 25320 26240 25372 26246
rect 25320 26182 25372 26188
rect 25332 21418 25360 26182
rect 25320 21412 25372 21418
rect 25320 21354 25372 21360
rect 25516 17898 25544 26551
rect 25700 26217 25728 30631
rect 25792 30598 25820 31214
rect 25780 30592 25832 30598
rect 25780 30534 25832 30540
rect 25686 26208 25742 26217
rect 25686 26143 25742 26152
rect 25792 22234 25820 30534
rect 25884 28937 25912 33782
rect 25956 33756 26252 33776
rect 26012 33754 26036 33756
rect 26092 33754 26116 33756
rect 26172 33754 26196 33756
rect 26034 33702 26036 33754
rect 26098 33702 26110 33754
rect 26172 33702 26174 33754
rect 26012 33700 26036 33702
rect 26092 33700 26116 33702
rect 26172 33700 26196 33702
rect 25956 33680 26252 33700
rect 26344 33522 26372 33798
rect 26332 33516 26384 33522
rect 26332 33458 26384 33464
rect 26344 32774 26372 33458
rect 26332 32768 26384 32774
rect 26332 32710 26384 32716
rect 25956 32668 26252 32688
rect 26012 32666 26036 32668
rect 26092 32666 26116 32668
rect 26172 32666 26196 32668
rect 26034 32614 26036 32666
rect 26098 32614 26110 32666
rect 26172 32614 26174 32666
rect 26012 32612 26036 32614
rect 26092 32612 26116 32614
rect 26172 32612 26196 32614
rect 25956 32592 26252 32612
rect 25956 31580 26252 31600
rect 26012 31578 26036 31580
rect 26092 31578 26116 31580
rect 26172 31578 26196 31580
rect 26034 31526 26036 31578
rect 26098 31526 26110 31578
rect 26172 31526 26174 31578
rect 26012 31524 26036 31526
rect 26092 31524 26116 31526
rect 26172 31524 26196 31526
rect 25956 31504 26252 31524
rect 26344 31362 26372 32710
rect 26252 31334 26372 31362
rect 26252 31278 26280 31334
rect 26240 31272 26292 31278
rect 26240 31214 26292 31220
rect 26424 31272 26476 31278
rect 26424 31214 26476 31220
rect 25956 30492 26252 30512
rect 26012 30490 26036 30492
rect 26092 30490 26116 30492
rect 26172 30490 26196 30492
rect 26034 30438 26036 30490
rect 26098 30438 26110 30490
rect 26172 30438 26174 30490
rect 26012 30436 26036 30438
rect 26092 30436 26116 30438
rect 26172 30436 26196 30438
rect 25956 30416 26252 30436
rect 25956 29404 26252 29424
rect 26012 29402 26036 29404
rect 26092 29402 26116 29404
rect 26172 29402 26196 29404
rect 26034 29350 26036 29402
rect 26098 29350 26110 29402
rect 26172 29350 26174 29402
rect 26012 29348 26036 29350
rect 26092 29348 26116 29350
rect 26172 29348 26196 29350
rect 25956 29328 26252 29348
rect 25870 28928 25926 28937
rect 25870 28863 25926 28872
rect 25956 28316 26252 28336
rect 26012 28314 26036 28316
rect 26092 28314 26116 28316
rect 26172 28314 26196 28316
rect 26034 28262 26036 28314
rect 26098 28262 26110 28314
rect 26172 28262 26174 28314
rect 26012 28260 26036 28262
rect 26092 28260 26116 28262
rect 26172 28260 26196 28262
rect 25956 28240 26252 28260
rect 25956 27228 26252 27248
rect 26012 27226 26036 27228
rect 26092 27226 26116 27228
rect 26172 27226 26196 27228
rect 26034 27174 26036 27226
rect 26098 27174 26110 27226
rect 26172 27174 26174 27226
rect 26012 27172 26036 27174
rect 26092 27172 26116 27174
rect 26172 27172 26196 27174
rect 25956 27152 26252 27172
rect 25956 26140 26252 26160
rect 26012 26138 26036 26140
rect 26092 26138 26116 26140
rect 26172 26138 26196 26140
rect 26034 26086 26036 26138
rect 26098 26086 26110 26138
rect 26172 26086 26174 26138
rect 26012 26084 26036 26086
rect 26092 26084 26116 26086
rect 26172 26084 26196 26086
rect 25956 26064 26252 26084
rect 25870 25256 25926 25265
rect 25870 25191 25926 25200
rect 25884 22642 25912 25191
rect 25956 25052 26252 25072
rect 26012 25050 26036 25052
rect 26092 25050 26116 25052
rect 26172 25050 26196 25052
rect 26034 24998 26036 25050
rect 26098 24998 26110 25050
rect 26172 24998 26174 25050
rect 26012 24996 26036 24998
rect 26092 24996 26116 24998
rect 26172 24996 26196 24998
rect 25956 24976 26252 24996
rect 25956 23964 26252 23984
rect 26012 23962 26036 23964
rect 26092 23962 26116 23964
rect 26172 23962 26196 23964
rect 26034 23910 26036 23962
rect 26098 23910 26110 23962
rect 26172 23910 26174 23962
rect 26012 23908 26036 23910
rect 26092 23908 26116 23910
rect 26172 23908 26196 23910
rect 25956 23888 26252 23908
rect 25956 22876 26252 22896
rect 26012 22874 26036 22876
rect 26092 22874 26116 22876
rect 26172 22874 26196 22876
rect 26034 22822 26036 22874
rect 26098 22822 26110 22874
rect 26172 22822 26174 22874
rect 26012 22820 26036 22822
rect 26092 22820 26116 22822
rect 26172 22820 26196 22822
rect 25956 22800 26252 22820
rect 25872 22636 25924 22642
rect 25872 22578 25924 22584
rect 26148 22568 26200 22574
rect 26148 22510 26200 22516
rect 26160 22234 26188 22510
rect 25780 22228 25832 22234
rect 25780 22170 25832 22176
rect 26148 22228 26200 22234
rect 26148 22170 26200 22176
rect 25792 21185 25820 22170
rect 26330 21856 26386 21865
rect 25956 21788 26252 21808
rect 26330 21791 26386 21800
rect 26012 21786 26036 21788
rect 26092 21786 26116 21788
rect 26172 21786 26196 21788
rect 26034 21734 26036 21786
rect 26098 21734 26110 21786
rect 26172 21734 26174 21786
rect 26012 21732 26036 21734
rect 26092 21732 26116 21734
rect 26172 21732 26196 21734
rect 25956 21712 26252 21732
rect 25778 21176 25834 21185
rect 25778 21111 25834 21120
rect 26344 21049 26372 21791
rect 26330 21040 26386 21049
rect 26330 20975 26386 20984
rect 25956 20700 26252 20720
rect 26012 20698 26036 20700
rect 26092 20698 26116 20700
rect 26172 20698 26196 20700
rect 26034 20646 26036 20698
rect 26098 20646 26110 20698
rect 26172 20646 26174 20698
rect 26012 20644 26036 20646
rect 26092 20644 26116 20646
rect 26172 20644 26196 20646
rect 25956 20624 26252 20644
rect 25594 20224 25650 20233
rect 25594 20159 25650 20168
rect 25608 18737 25636 20159
rect 25956 19612 26252 19632
rect 26012 19610 26036 19612
rect 26092 19610 26116 19612
rect 26172 19610 26196 19612
rect 26034 19558 26036 19610
rect 26098 19558 26110 19610
rect 26172 19558 26174 19610
rect 26012 19556 26036 19558
rect 26092 19556 26116 19558
rect 26172 19556 26196 19558
rect 25956 19536 26252 19556
rect 25594 18728 25650 18737
rect 25594 18663 25650 18672
rect 25956 18524 26252 18544
rect 26012 18522 26036 18524
rect 26092 18522 26116 18524
rect 26172 18522 26196 18524
rect 26034 18470 26036 18522
rect 26098 18470 26110 18522
rect 26172 18470 26174 18522
rect 26012 18468 26036 18470
rect 26092 18468 26116 18470
rect 26172 18468 26196 18470
rect 25956 18448 26252 18468
rect 25424 17870 25544 17898
rect 25424 13433 25452 17870
rect 25502 17776 25558 17785
rect 25502 17711 25558 17720
rect 25410 13424 25466 13433
rect 25410 13359 25466 13368
rect 25226 11656 25282 11665
rect 25226 11591 25282 11600
rect 24950 7440 25006 7449
rect 24950 7375 25006 7384
rect 24858 5264 24914 5273
rect 24858 5199 24914 5208
rect 23938 4040 23994 4049
rect 23938 3975 23994 3984
rect 23018 3768 23074 3777
rect 23018 3703 23074 3712
rect 23032 800 23060 3703
rect 23952 800 23980 3975
rect 24860 2304 24912 2310
rect 24860 2246 24912 2252
rect 24872 800 24900 2246
rect 3146 776 3202 785
rect 3146 711 3202 720
rect 3698 0 3754 800
rect 4618 0 4674 800
rect 5078 0 5134 800
rect 5998 0 6054 800
rect 6918 0 6974 800
rect 7378 0 7434 800
rect 8298 0 8354 800
rect 9218 0 9274 800
rect 10138 0 10194 800
rect 10598 0 10654 800
rect 11518 0 11574 800
rect 12438 0 12494 800
rect 12898 0 12954 800
rect 13818 0 13874 800
rect 14738 0 14794 800
rect 15198 0 15254 800
rect 16118 0 16174 800
rect 17038 0 17094 800
rect 17958 0 18014 800
rect 18418 0 18474 800
rect 19338 0 19394 800
rect 20258 0 20314 800
rect 20718 0 20774 800
rect 21638 0 21694 800
rect 22558 0 22614 800
rect 23018 0 23074 800
rect 23938 0 23994 800
rect 24858 0 24914 800
rect 24964 785 24992 7375
rect 25318 6896 25374 6905
rect 25318 6831 25374 6840
rect 25332 4185 25360 6831
rect 25318 4176 25374 4185
rect 25318 4111 25374 4120
rect 25318 2680 25374 2689
rect 25318 2615 25374 2624
rect 25332 800 25360 2615
rect 24950 776 25006 785
rect 24950 711 25006 720
rect 25318 0 25374 800
rect 25516 105 25544 17711
rect 25956 17436 26252 17456
rect 26012 17434 26036 17436
rect 26092 17434 26116 17436
rect 26172 17434 26196 17436
rect 26034 17382 26036 17434
rect 26098 17382 26110 17434
rect 26172 17382 26174 17434
rect 26012 17380 26036 17382
rect 26092 17380 26116 17382
rect 26172 17380 26196 17382
rect 25956 17360 26252 17380
rect 25956 16348 26252 16368
rect 26012 16346 26036 16348
rect 26092 16346 26116 16348
rect 26172 16346 26196 16348
rect 26034 16294 26036 16346
rect 26098 16294 26110 16346
rect 26172 16294 26174 16346
rect 26012 16292 26036 16294
rect 26092 16292 26116 16294
rect 26172 16292 26196 16294
rect 25956 16272 26252 16292
rect 25956 15260 26252 15280
rect 26012 15258 26036 15260
rect 26092 15258 26116 15260
rect 26172 15258 26196 15260
rect 26034 15206 26036 15258
rect 26098 15206 26110 15258
rect 26172 15206 26174 15258
rect 26012 15204 26036 15206
rect 26092 15204 26116 15206
rect 26172 15204 26196 15206
rect 25956 15184 26252 15204
rect 25956 14172 26252 14192
rect 26012 14170 26036 14172
rect 26092 14170 26116 14172
rect 26172 14170 26196 14172
rect 26034 14118 26036 14170
rect 26098 14118 26110 14170
rect 26172 14118 26174 14170
rect 26012 14116 26036 14118
rect 26092 14116 26116 14118
rect 26172 14116 26196 14118
rect 25956 14096 26252 14116
rect 26238 13832 26294 13841
rect 26238 13767 26240 13776
rect 26292 13767 26294 13776
rect 26240 13738 26292 13744
rect 26252 13530 26280 13738
rect 26240 13524 26292 13530
rect 26240 13466 26292 13472
rect 25956 13084 26252 13104
rect 26012 13082 26036 13084
rect 26092 13082 26116 13084
rect 26172 13082 26196 13084
rect 26034 13030 26036 13082
rect 26098 13030 26110 13082
rect 26172 13030 26174 13082
rect 26012 13028 26036 13030
rect 26092 13028 26116 13030
rect 26172 13028 26196 13030
rect 25956 13008 26252 13028
rect 25956 11996 26252 12016
rect 26012 11994 26036 11996
rect 26092 11994 26116 11996
rect 26172 11994 26196 11996
rect 26034 11942 26036 11994
rect 26098 11942 26110 11994
rect 26172 11942 26174 11994
rect 26012 11940 26036 11942
rect 26092 11940 26116 11942
rect 26172 11940 26196 11942
rect 25956 11920 26252 11940
rect 26330 11520 26386 11529
rect 26330 11455 26386 11464
rect 25956 10908 26252 10928
rect 26012 10906 26036 10908
rect 26092 10906 26116 10908
rect 26172 10906 26196 10908
rect 26034 10854 26036 10906
rect 26098 10854 26110 10906
rect 26172 10854 26174 10906
rect 26012 10852 26036 10854
rect 26092 10852 26116 10854
rect 26172 10852 26196 10854
rect 25956 10832 26252 10852
rect 25956 9820 26252 9840
rect 26012 9818 26036 9820
rect 26092 9818 26116 9820
rect 26172 9818 26196 9820
rect 26034 9766 26036 9818
rect 26098 9766 26110 9818
rect 26172 9766 26174 9818
rect 26012 9764 26036 9766
rect 26092 9764 26116 9766
rect 26172 9764 26196 9766
rect 25956 9744 26252 9764
rect 25956 8732 26252 8752
rect 26012 8730 26036 8732
rect 26092 8730 26116 8732
rect 26172 8730 26196 8732
rect 26034 8678 26036 8730
rect 26098 8678 26110 8730
rect 26172 8678 26174 8730
rect 26012 8676 26036 8678
rect 26092 8676 26116 8678
rect 26172 8676 26196 8678
rect 25956 8656 26252 8676
rect 25956 7644 26252 7664
rect 26012 7642 26036 7644
rect 26092 7642 26116 7644
rect 26172 7642 26196 7644
rect 26034 7590 26036 7642
rect 26098 7590 26110 7642
rect 26172 7590 26174 7642
rect 26012 7588 26036 7590
rect 26092 7588 26116 7590
rect 26172 7588 26196 7590
rect 25956 7568 26252 7588
rect 25956 6556 26252 6576
rect 26012 6554 26036 6556
rect 26092 6554 26116 6556
rect 26172 6554 26196 6556
rect 26034 6502 26036 6554
rect 26098 6502 26110 6554
rect 26172 6502 26174 6554
rect 26012 6500 26036 6502
rect 26092 6500 26116 6502
rect 26172 6500 26196 6502
rect 25956 6480 26252 6500
rect 25956 5468 26252 5488
rect 26012 5466 26036 5468
rect 26092 5466 26116 5468
rect 26172 5466 26196 5468
rect 26034 5414 26036 5466
rect 26098 5414 26110 5466
rect 26172 5414 26174 5466
rect 26012 5412 26036 5414
rect 26092 5412 26116 5414
rect 26172 5412 26196 5414
rect 25956 5392 26252 5412
rect 25956 4380 26252 4400
rect 26012 4378 26036 4380
rect 26092 4378 26116 4380
rect 26172 4378 26196 4380
rect 26034 4326 26036 4378
rect 26098 4326 26110 4378
rect 26172 4326 26174 4378
rect 26012 4324 26036 4326
rect 26092 4324 26116 4326
rect 26172 4324 26196 4326
rect 25956 4304 26252 4324
rect 25956 3292 26252 3312
rect 26012 3290 26036 3292
rect 26092 3290 26116 3292
rect 26172 3290 26196 3292
rect 26034 3238 26036 3290
rect 26098 3238 26110 3290
rect 26172 3238 26174 3290
rect 26012 3236 26036 3238
rect 26092 3236 26116 3238
rect 26172 3236 26196 3238
rect 25956 3216 26252 3236
rect 25956 2204 26252 2224
rect 26012 2202 26036 2204
rect 26092 2202 26116 2204
rect 26172 2202 26196 2204
rect 26034 2150 26036 2202
rect 26098 2150 26110 2202
rect 26172 2150 26174 2202
rect 26012 2148 26036 2150
rect 26092 2148 26116 2150
rect 26172 2148 26196 2150
rect 25956 2128 26252 2148
rect 26344 1986 26372 11455
rect 26252 1958 26372 1986
rect 26436 1986 26464 31214
rect 26988 23905 27016 54606
rect 27344 53984 27396 53990
rect 27344 53926 27396 53932
rect 27356 52465 27384 53926
rect 27540 53718 27568 54606
rect 27724 54330 27752 54674
rect 27712 54324 27764 54330
rect 27712 54266 27764 54272
rect 27528 53712 27580 53718
rect 27528 53654 27580 53660
rect 27908 53009 27936 70314
rect 27988 66292 28040 66298
rect 27988 66234 28040 66240
rect 28000 66201 28028 66234
rect 27986 66192 28042 66201
rect 27986 66127 28042 66136
rect 28080 61668 28132 61674
rect 28080 61610 28132 61616
rect 27986 56672 28042 56681
rect 27986 56607 28042 56616
rect 27894 53000 27950 53009
rect 27894 52935 27950 52944
rect 28000 52884 28028 56607
rect 27816 52856 28028 52884
rect 27342 52456 27398 52465
rect 27342 52391 27398 52400
rect 27710 49600 27766 49609
rect 27710 49535 27766 49544
rect 27724 47802 27752 49535
rect 27712 47796 27764 47802
rect 27712 47738 27764 47744
rect 27068 44872 27120 44878
rect 27068 44814 27120 44820
rect 27080 41721 27108 44814
rect 27712 44192 27764 44198
rect 27712 44134 27764 44140
rect 27526 44024 27582 44033
rect 27526 43959 27582 43968
rect 27252 43784 27304 43790
rect 27252 43726 27304 43732
rect 27264 43353 27292 43726
rect 27540 43654 27568 43959
rect 27528 43648 27580 43654
rect 27528 43590 27580 43596
rect 27344 43444 27396 43450
rect 27344 43386 27396 43392
rect 27250 43344 27306 43353
rect 27250 43279 27306 43288
rect 27356 42809 27384 43386
rect 27540 43314 27568 43590
rect 27528 43308 27580 43314
rect 27528 43250 27580 43256
rect 27342 42800 27398 42809
rect 27342 42735 27398 42744
rect 27724 42673 27752 44134
rect 27710 42664 27766 42673
rect 27710 42599 27766 42608
rect 27528 42152 27580 42158
rect 27528 42094 27580 42100
rect 27160 42016 27212 42022
rect 27160 41958 27212 41964
rect 27066 41712 27122 41721
rect 27172 41682 27200 41958
rect 27540 41818 27568 42094
rect 27528 41812 27580 41818
rect 27528 41754 27580 41760
rect 27066 41647 27122 41656
rect 27160 41676 27212 41682
rect 27160 41618 27212 41624
rect 27172 41206 27200 41618
rect 27160 41200 27212 41206
rect 27160 41142 27212 41148
rect 27528 37664 27580 37670
rect 27528 37606 27580 37612
rect 27540 32502 27568 37606
rect 27712 36576 27764 36582
rect 27712 36518 27764 36524
rect 27724 36145 27752 36518
rect 27710 36136 27766 36145
rect 27710 36071 27766 36080
rect 27710 35728 27766 35737
rect 27816 35698 27844 52856
rect 28092 48521 28120 61610
rect 28078 48512 28134 48521
rect 28078 48447 28134 48456
rect 27710 35663 27766 35672
rect 27804 35692 27856 35698
rect 27724 34746 27752 35663
rect 27804 35634 27856 35640
rect 27804 35556 27856 35562
rect 27804 35498 27856 35504
rect 27712 34740 27764 34746
rect 27712 34682 27764 34688
rect 27816 33289 27844 35498
rect 27802 33280 27858 33289
rect 27802 33215 27858 33224
rect 27528 32496 27580 32502
rect 27528 32438 27580 32444
rect 27620 31340 27672 31346
rect 27620 31282 27672 31288
rect 27632 31249 27660 31282
rect 27618 31240 27674 31249
rect 27618 31175 27674 31184
rect 26974 23896 27030 23905
rect 26974 23831 27030 23840
rect 27712 22432 27764 22438
rect 27712 22374 27764 22380
rect 27724 20369 27752 22374
rect 27710 20360 27766 20369
rect 27710 20295 27766 20304
rect 27618 13968 27674 13977
rect 27618 13903 27620 13912
rect 27672 13903 27674 13912
rect 27620 13874 27672 13880
rect 26516 13864 26568 13870
rect 26514 13832 26516 13841
rect 26568 13832 26570 13841
rect 26514 13767 26570 13776
rect 26516 13184 26568 13190
rect 26516 13126 26568 13132
rect 26528 2145 26556 13126
rect 29458 8528 29514 8537
rect 29458 8463 29514 8472
rect 28538 4856 28594 4865
rect 28538 4791 28594 4800
rect 26514 2136 26570 2145
rect 26514 2071 26570 2080
rect 28078 2000 28134 2009
rect 26436 1958 27108 1986
rect 26252 800 26280 1958
rect 27080 898 27108 1958
rect 28078 1935 28134 1944
rect 27080 870 27200 898
rect 27172 800 27200 870
rect 28092 800 28120 1935
rect 28552 800 28580 4791
rect 29472 800 29500 8463
rect 25502 96 25558 105
rect 25502 31 25558 40
rect 26238 0 26294 800
rect 27158 0 27214 800
rect 28078 0 28134 800
rect 28538 0 28594 800
rect 29458 0 29514 800
<< via2 >>
rect 4066 79600 4122 79656
rect 110 72664 166 72720
rect 2318 75792 2374 75848
rect 2962 75520 3018 75576
rect 1398 73616 1454 73672
rect 1766 72120 1822 72176
rect 1674 69300 1676 69320
rect 1676 69300 1728 69320
rect 1728 69300 1730 69320
rect 1674 69264 1730 69300
rect 1674 57160 1730 57216
rect 1674 53760 1730 53816
rect 1582 50904 1638 50960
rect 2778 71440 2834 71496
rect 2042 69420 2098 69456
rect 2042 69400 2044 69420
rect 2044 69400 2096 69420
rect 2096 69400 2098 69420
rect 2778 61920 2834 61976
rect 1950 45600 2006 45656
rect 1766 44920 1822 44976
rect 1766 41520 1822 41576
rect 1674 37440 1730 37496
rect 1582 35400 1638 35456
rect 1582 26560 1638 26616
rect 1306 21528 1362 21584
rect 1950 23840 2006 23896
rect 1858 20440 1914 20496
rect 1490 17040 1546 17096
rect 1674 17196 1730 17232
rect 1674 17176 1676 17196
rect 1676 17176 1728 17196
rect 1728 17176 1730 17196
rect 2870 59880 2926 59936
rect 2686 57452 2742 57488
rect 3330 78240 3386 78296
rect 24674 79600 24730 79656
rect 4066 77424 4122 77480
rect 3238 74840 3294 74896
rect 3422 74704 3478 74760
rect 3238 68720 3294 68776
rect 3054 58520 3110 58576
rect 2686 57432 2688 57452
rect 2688 57432 2740 57452
rect 2740 57432 2742 57452
rect 2226 57160 2282 57216
rect 2962 44532 3018 44568
rect 2962 44512 2964 44532
rect 2964 44512 3016 44532
rect 3016 44512 3018 44532
rect 2134 40160 2190 40216
rect 2042 13640 2098 13696
rect 1582 12280 1638 12336
rect 2042 9036 2098 9072
rect 2042 9016 2044 9036
rect 2044 9016 2096 9036
rect 2096 9016 2098 9036
rect 18 7928 74 7984
rect 1582 7520 1638 7576
rect 2318 41384 2374 41440
rect 2870 35692 2926 35728
rect 2870 35672 2872 35692
rect 2872 35672 2924 35692
rect 2924 35672 2926 35692
rect 2778 34040 2834 34096
rect 2870 33360 2926 33416
rect 2686 25200 2742 25256
rect 3146 43732 3148 43752
rect 3148 43732 3200 43752
rect 3200 43732 3202 43752
rect 3146 43696 3202 43732
rect 3146 43188 3148 43208
rect 3148 43188 3200 43208
rect 3200 43188 3202 43208
rect 3146 43152 3202 43188
rect 5354 75792 5410 75848
rect 5956 77274 6012 77276
rect 6036 77274 6092 77276
rect 6116 77274 6172 77276
rect 6196 77274 6252 77276
rect 5956 77222 5982 77274
rect 5982 77222 6012 77274
rect 6036 77222 6046 77274
rect 6046 77222 6092 77274
rect 6116 77222 6162 77274
rect 6162 77222 6172 77274
rect 6196 77222 6226 77274
rect 6226 77222 6252 77274
rect 5956 77220 6012 77222
rect 6036 77220 6092 77222
rect 6116 77220 6172 77222
rect 6196 77220 6252 77222
rect 5956 76186 6012 76188
rect 6036 76186 6092 76188
rect 6116 76186 6172 76188
rect 6196 76186 6252 76188
rect 5956 76134 5982 76186
rect 5982 76134 6012 76186
rect 6036 76134 6046 76186
rect 6046 76134 6092 76186
rect 6116 76134 6162 76186
rect 6162 76134 6172 76186
rect 6196 76134 6226 76186
rect 6226 76134 6252 76186
rect 5956 76132 6012 76134
rect 6036 76132 6092 76134
rect 6116 76132 6172 76134
rect 6196 76132 6252 76134
rect 5956 75098 6012 75100
rect 6036 75098 6092 75100
rect 6116 75098 6172 75100
rect 6196 75098 6252 75100
rect 5956 75046 5982 75098
rect 5982 75046 6012 75098
rect 6036 75046 6046 75098
rect 6046 75046 6092 75098
rect 6116 75046 6162 75098
rect 6162 75046 6172 75098
rect 6196 75046 6226 75098
rect 6226 75046 6252 75098
rect 5956 75044 6012 75046
rect 6036 75044 6092 75046
rect 6116 75044 6172 75046
rect 6196 75044 6252 75046
rect 5630 74840 5686 74896
rect 5354 73072 5410 73128
rect 4066 66680 4122 66736
rect 4066 66000 4122 66056
rect 4802 65184 4858 65240
rect 4802 64504 4858 64560
rect 3790 63280 3846 63336
rect 3422 62736 3478 62792
rect 3330 57876 3332 57896
rect 3332 57876 3384 57896
rect 3384 57876 3386 57896
rect 3330 57840 3386 57876
rect 3330 57160 3386 57216
rect 3606 57160 3662 57216
rect 3422 55800 3478 55856
rect 3698 49000 3754 49056
rect 3514 48592 3570 48648
rect 3422 43560 3478 43616
rect 3330 43016 3386 43072
rect 3238 41384 3294 41440
rect 3146 39480 3202 39536
rect 3146 38936 3202 38992
rect 3238 30504 3294 30560
rect 3146 29144 3202 29200
rect 2778 21528 2834 21584
rect 3238 24656 3294 24712
rect 3146 21528 3202 21584
rect 2962 19896 3018 19952
rect 2318 10648 2374 10704
rect 478 6160 534 6216
rect 3238 18400 3294 18456
rect 3054 13368 3110 13424
rect 3330 13232 3386 13288
rect 3606 48184 3662 48240
rect 5538 74704 5594 74760
rect 5538 71032 5594 71088
rect 6918 75248 6974 75304
rect 7470 74704 7526 74760
rect 5956 74010 6012 74012
rect 6036 74010 6092 74012
rect 6116 74010 6172 74012
rect 6196 74010 6252 74012
rect 5956 73958 5982 74010
rect 5982 73958 6012 74010
rect 6036 73958 6046 74010
rect 6046 73958 6092 74010
rect 6116 73958 6162 74010
rect 6162 73958 6172 74010
rect 6196 73958 6226 74010
rect 6226 73958 6252 74010
rect 5956 73956 6012 73958
rect 6036 73956 6092 73958
rect 6116 73956 6172 73958
rect 6196 73956 6252 73958
rect 6918 73752 6974 73808
rect 5956 72922 6012 72924
rect 6036 72922 6092 72924
rect 6116 72922 6172 72924
rect 6196 72922 6252 72924
rect 5956 72870 5982 72922
rect 5982 72870 6012 72922
rect 6036 72870 6046 72922
rect 6046 72870 6092 72922
rect 6116 72870 6162 72922
rect 6162 72870 6172 72922
rect 6196 72870 6226 72922
rect 6226 72870 6252 72922
rect 5956 72868 6012 72870
rect 6036 72868 6092 72870
rect 6116 72868 6172 72870
rect 6196 72868 6252 72870
rect 7286 72528 7342 72584
rect 5956 71834 6012 71836
rect 6036 71834 6092 71836
rect 6116 71834 6172 71836
rect 6196 71834 6252 71836
rect 5956 71782 5982 71834
rect 5982 71782 6012 71834
rect 6036 71782 6046 71834
rect 6046 71782 6092 71834
rect 6116 71782 6162 71834
rect 6162 71782 6172 71834
rect 6196 71782 6226 71834
rect 6226 71782 6252 71834
rect 5956 71780 6012 71782
rect 6036 71780 6092 71782
rect 6116 71780 6172 71782
rect 6196 71780 6252 71782
rect 5956 70746 6012 70748
rect 6036 70746 6092 70748
rect 6116 70746 6172 70748
rect 6196 70746 6252 70748
rect 5956 70694 5982 70746
rect 5982 70694 6012 70746
rect 6036 70694 6046 70746
rect 6046 70694 6092 70746
rect 6116 70694 6162 70746
rect 6162 70694 6172 70746
rect 6196 70694 6226 70746
rect 6226 70694 6252 70746
rect 5956 70692 6012 70694
rect 6036 70692 6092 70694
rect 6116 70692 6172 70694
rect 6196 70692 6252 70694
rect 5630 69808 5686 69864
rect 5956 69658 6012 69660
rect 6036 69658 6092 69660
rect 6116 69658 6172 69660
rect 6196 69658 6252 69660
rect 5956 69606 5982 69658
rect 5982 69606 6012 69658
rect 6036 69606 6046 69658
rect 6046 69606 6092 69658
rect 6116 69606 6162 69658
rect 6162 69606 6172 69658
rect 6196 69606 6226 69658
rect 6226 69606 6252 69658
rect 5956 69604 6012 69606
rect 6036 69604 6092 69606
rect 6116 69604 6172 69606
rect 6196 69604 6252 69606
rect 5956 68570 6012 68572
rect 6036 68570 6092 68572
rect 6116 68570 6172 68572
rect 6196 68570 6252 68572
rect 5956 68518 5982 68570
rect 5982 68518 6012 68570
rect 6036 68518 6046 68570
rect 6046 68518 6092 68570
rect 6116 68518 6162 68570
rect 6162 68518 6172 68570
rect 6196 68518 6226 68570
rect 6226 68518 6252 68570
rect 5956 68516 6012 68518
rect 6036 68516 6092 68518
rect 6116 68516 6172 68518
rect 6196 68516 6252 68518
rect 5956 67482 6012 67484
rect 6036 67482 6092 67484
rect 6116 67482 6172 67484
rect 6196 67482 6252 67484
rect 5956 67430 5982 67482
rect 5982 67430 6012 67482
rect 6036 67430 6046 67482
rect 6046 67430 6092 67482
rect 6116 67430 6162 67482
rect 6162 67430 6172 67482
rect 6196 67430 6226 67482
rect 6226 67430 6252 67482
rect 5956 67428 6012 67430
rect 6036 67428 6092 67430
rect 6116 67428 6172 67430
rect 6196 67428 6252 67430
rect 5956 66394 6012 66396
rect 6036 66394 6092 66396
rect 6116 66394 6172 66396
rect 6196 66394 6252 66396
rect 5956 66342 5982 66394
rect 5982 66342 6012 66394
rect 6036 66342 6046 66394
rect 6046 66342 6092 66394
rect 6116 66342 6162 66394
rect 6162 66342 6172 66394
rect 6196 66342 6226 66394
rect 6226 66342 6252 66394
rect 5956 66340 6012 66342
rect 6036 66340 6092 66342
rect 6116 66340 6172 66342
rect 6196 66340 6252 66342
rect 5956 65306 6012 65308
rect 6036 65306 6092 65308
rect 6116 65306 6172 65308
rect 6196 65306 6252 65308
rect 5956 65254 5982 65306
rect 5982 65254 6012 65306
rect 6036 65254 6046 65306
rect 6046 65254 6092 65306
rect 6116 65254 6162 65306
rect 6162 65254 6172 65306
rect 6196 65254 6226 65306
rect 6226 65254 6252 65306
rect 5956 65252 6012 65254
rect 6036 65252 6092 65254
rect 6116 65252 6172 65254
rect 6196 65252 6252 65254
rect 5956 64218 6012 64220
rect 6036 64218 6092 64220
rect 6116 64218 6172 64220
rect 6196 64218 6252 64220
rect 5956 64166 5982 64218
rect 5982 64166 6012 64218
rect 6036 64166 6046 64218
rect 6046 64166 6092 64218
rect 6116 64166 6162 64218
rect 6162 64166 6172 64218
rect 6196 64166 6226 64218
rect 6226 64166 6252 64218
rect 5956 64164 6012 64166
rect 6036 64164 6092 64166
rect 6116 64164 6172 64166
rect 6196 64164 6252 64166
rect 5956 63130 6012 63132
rect 6036 63130 6092 63132
rect 6116 63130 6172 63132
rect 6196 63130 6252 63132
rect 5956 63078 5982 63130
rect 5982 63078 6012 63130
rect 6036 63078 6046 63130
rect 6046 63078 6092 63130
rect 6116 63078 6162 63130
rect 6162 63078 6172 63130
rect 6196 63078 6226 63130
rect 6226 63078 6252 63130
rect 5956 63076 6012 63078
rect 6036 63076 6092 63078
rect 6116 63076 6172 63078
rect 6196 63076 6252 63078
rect 5956 62042 6012 62044
rect 6036 62042 6092 62044
rect 6116 62042 6172 62044
rect 6196 62042 6252 62044
rect 5956 61990 5982 62042
rect 5982 61990 6012 62042
rect 6036 61990 6046 62042
rect 6046 61990 6092 62042
rect 6116 61990 6162 62042
rect 6162 61990 6172 62042
rect 6196 61990 6226 62042
rect 6226 61990 6252 62042
rect 5956 61988 6012 61990
rect 6036 61988 6092 61990
rect 6116 61988 6172 61990
rect 6196 61988 6252 61990
rect 5956 60954 6012 60956
rect 6036 60954 6092 60956
rect 6116 60954 6172 60956
rect 6196 60954 6252 60956
rect 5956 60902 5982 60954
rect 5982 60902 6012 60954
rect 6036 60902 6046 60954
rect 6046 60902 6092 60954
rect 6116 60902 6162 60954
rect 6162 60902 6172 60954
rect 6196 60902 6226 60954
rect 6226 60902 6252 60954
rect 5956 60900 6012 60902
rect 6036 60900 6092 60902
rect 6116 60900 6172 60902
rect 6196 60900 6252 60902
rect 5446 60696 5502 60752
rect 5956 59866 6012 59868
rect 6036 59866 6092 59868
rect 6116 59866 6172 59868
rect 6196 59866 6252 59868
rect 5956 59814 5982 59866
rect 5982 59814 6012 59866
rect 6036 59814 6046 59866
rect 6046 59814 6092 59866
rect 6116 59814 6162 59866
rect 6162 59814 6172 59866
rect 6196 59814 6226 59866
rect 6226 59814 6252 59866
rect 5956 59812 6012 59814
rect 6036 59812 6092 59814
rect 6116 59812 6172 59814
rect 6196 59812 6252 59814
rect 5956 58778 6012 58780
rect 6036 58778 6092 58780
rect 6116 58778 6172 58780
rect 6196 58778 6252 58780
rect 5956 58726 5982 58778
rect 5982 58726 6012 58778
rect 6036 58726 6046 58778
rect 6046 58726 6092 58778
rect 6116 58726 6162 58778
rect 6162 58726 6172 58778
rect 6196 58726 6226 58778
rect 6226 58726 6252 58778
rect 5956 58724 6012 58726
rect 6036 58724 6092 58726
rect 6116 58724 6172 58726
rect 6196 58724 6252 58726
rect 7010 57840 7066 57896
rect 5956 57690 6012 57692
rect 6036 57690 6092 57692
rect 6116 57690 6172 57692
rect 6196 57690 6252 57692
rect 5956 57638 5982 57690
rect 5982 57638 6012 57690
rect 6036 57638 6046 57690
rect 6046 57638 6092 57690
rect 6116 57638 6162 57690
rect 6162 57638 6172 57690
rect 6196 57638 6226 57690
rect 6226 57638 6252 57690
rect 5956 57636 6012 57638
rect 6036 57636 6092 57638
rect 6116 57636 6172 57638
rect 6196 57636 6252 57638
rect 5956 56602 6012 56604
rect 6036 56602 6092 56604
rect 6116 56602 6172 56604
rect 6196 56602 6252 56604
rect 5956 56550 5982 56602
rect 5982 56550 6012 56602
rect 6036 56550 6046 56602
rect 6046 56550 6092 56602
rect 6116 56550 6162 56602
rect 6162 56550 6172 56602
rect 6196 56550 6226 56602
rect 6226 56550 6252 56602
rect 5956 56548 6012 56550
rect 6036 56548 6092 56550
rect 6116 56548 6172 56550
rect 6196 56548 6252 56550
rect 5956 55514 6012 55516
rect 6036 55514 6092 55516
rect 6116 55514 6172 55516
rect 6196 55514 6252 55516
rect 5956 55462 5982 55514
rect 5982 55462 6012 55514
rect 6036 55462 6046 55514
rect 6046 55462 6092 55514
rect 6116 55462 6162 55514
rect 6162 55462 6172 55514
rect 6196 55462 6226 55514
rect 6226 55462 6252 55514
rect 5956 55460 6012 55462
rect 6036 55460 6092 55462
rect 6116 55460 6172 55462
rect 6196 55460 6252 55462
rect 5956 54426 6012 54428
rect 6036 54426 6092 54428
rect 6116 54426 6172 54428
rect 6196 54426 6252 54428
rect 5956 54374 5982 54426
rect 5982 54374 6012 54426
rect 6036 54374 6046 54426
rect 6046 54374 6092 54426
rect 6116 54374 6162 54426
rect 6162 54374 6172 54426
rect 6196 54374 6226 54426
rect 6226 54374 6252 54426
rect 5956 54372 6012 54374
rect 6036 54372 6092 54374
rect 6116 54372 6172 54374
rect 6196 54372 6252 54374
rect 5956 53338 6012 53340
rect 6036 53338 6092 53340
rect 6116 53338 6172 53340
rect 6196 53338 6252 53340
rect 5956 53286 5982 53338
rect 5982 53286 6012 53338
rect 6036 53286 6046 53338
rect 6046 53286 6092 53338
rect 6116 53286 6162 53338
rect 6162 53286 6172 53338
rect 6196 53286 6226 53338
rect 6226 53286 6252 53338
rect 5956 53284 6012 53286
rect 6036 53284 6092 53286
rect 6116 53284 6172 53286
rect 6196 53284 6252 53286
rect 4066 52556 4122 52592
rect 4066 52536 4068 52556
rect 4068 52536 4120 52556
rect 4120 52536 4122 52556
rect 5956 52250 6012 52252
rect 6036 52250 6092 52252
rect 6116 52250 6172 52252
rect 6196 52250 6252 52252
rect 5956 52198 5982 52250
rect 5982 52198 6012 52250
rect 6036 52198 6046 52250
rect 6046 52198 6092 52250
rect 6116 52198 6162 52250
rect 6162 52198 6172 52250
rect 6196 52198 6226 52250
rect 6226 52198 6252 52250
rect 5956 52196 6012 52198
rect 6036 52196 6092 52198
rect 6116 52196 6172 52198
rect 6196 52196 6252 52198
rect 6274 51312 6330 51368
rect 5956 51162 6012 51164
rect 6036 51162 6092 51164
rect 6116 51162 6172 51164
rect 6196 51162 6252 51164
rect 5956 51110 5982 51162
rect 5982 51110 6012 51162
rect 6036 51110 6046 51162
rect 6046 51110 6092 51162
rect 6116 51110 6162 51162
rect 6162 51110 6172 51162
rect 6196 51110 6226 51162
rect 6226 51110 6252 51162
rect 5956 51108 6012 51110
rect 6036 51108 6092 51110
rect 6116 51108 6172 51110
rect 6196 51108 6252 51110
rect 5814 50904 5870 50960
rect 4066 50360 4122 50416
rect 5956 50074 6012 50076
rect 6036 50074 6092 50076
rect 6116 50074 6172 50076
rect 6196 50074 6252 50076
rect 5956 50022 5982 50074
rect 5982 50022 6012 50074
rect 6036 50022 6046 50074
rect 6046 50022 6092 50074
rect 6116 50022 6162 50074
rect 6162 50022 6172 50074
rect 6196 50022 6226 50074
rect 6226 50022 6252 50074
rect 5956 50020 6012 50022
rect 6036 50020 6092 50022
rect 6116 50020 6172 50022
rect 6196 50020 6252 50022
rect 4066 49680 4122 49736
rect 5956 48986 6012 48988
rect 6036 48986 6092 48988
rect 6116 48986 6172 48988
rect 6196 48986 6252 48988
rect 5956 48934 5982 48986
rect 5982 48934 6012 48986
rect 6036 48934 6046 48986
rect 6046 48934 6092 48986
rect 6116 48934 6162 48986
rect 6162 48934 6172 48986
rect 6196 48934 6226 48986
rect 6226 48934 6252 48986
rect 5956 48932 6012 48934
rect 6036 48932 6092 48934
rect 6116 48932 6172 48934
rect 6196 48932 6252 48934
rect 4066 48320 4122 48376
rect 3790 48048 3846 48104
rect 7194 48184 7250 48240
rect 5956 47898 6012 47900
rect 6036 47898 6092 47900
rect 6116 47898 6172 47900
rect 6196 47898 6252 47900
rect 5956 47846 5982 47898
rect 5982 47846 6012 47898
rect 6036 47846 6046 47898
rect 6046 47846 6092 47898
rect 6116 47846 6162 47898
rect 6162 47846 6172 47898
rect 6196 47846 6226 47898
rect 6226 47846 6252 47898
rect 5956 47844 6012 47846
rect 6036 47844 6092 47846
rect 6116 47844 6172 47846
rect 6196 47844 6252 47846
rect 5956 46810 6012 46812
rect 6036 46810 6092 46812
rect 6116 46810 6172 46812
rect 6196 46810 6252 46812
rect 5956 46758 5982 46810
rect 5982 46758 6012 46810
rect 6036 46758 6046 46810
rect 6046 46758 6092 46810
rect 6116 46758 6162 46810
rect 6162 46758 6172 46810
rect 6196 46758 6226 46810
rect 6226 46758 6252 46810
rect 5956 46756 6012 46758
rect 6036 46756 6092 46758
rect 6116 46756 6172 46758
rect 6196 46756 6252 46758
rect 4066 46416 4122 46472
rect 6274 45872 6330 45928
rect 5956 45722 6012 45724
rect 6036 45722 6092 45724
rect 6116 45722 6172 45724
rect 6196 45722 6252 45724
rect 5956 45670 5982 45722
rect 5982 45670 6012 45722
rect 6036 45670 6046 45722
rect 6046 45670 6092 45722
rect 6116 45670 6162 45722
rect 6162 45670 6172 45722
rect 6196 45670 6226 45722
rect 6226 45670 6252 45722
rect 5956 45668 6012 45670
rect 6036 45668 6092 45670
rect 6116 45668 6172 45670
rect 6196 45668 6252 45670
rect 5956 44634 6012 44636
rect 6036 44634 6092 44636
rect 6116 44634 6172 44636
rect 6196 44634 6252 44636
rect 5956 44582 5982 44634
rect 5982 44582 6012 44634
rect 6036 44582 6046 44634
rect 6046 44582 6092 44634
rect 6116 44582 6162 44634
rect 6162 44582 6172 44634
rect 6196 44582 6226 44634
rect 6226 44582 6252 44634
rect 5956 44580 6012 44582
rect 6036 44580 6092 44582
rect 6116 44580 6172 44582
rect 6196 44580 6252 44582
rect 4066 43832 4122 43888
rect 5956 43546 6012 43548
rect 6036 43546 6092 43548
rect 6116 43546 6172 43548
rect 6196 43546 6252 43548
rect 5956 43494 5982 43546
rect 5982 43494 6012 43546
rect 6036 43494 6046 43546
rect 6046 43494 6092 43546
rect 6116 43494 6162 43546
rect 6162 43494 6172 43546
rect 6196 43494 6226 43546
rect 6226 43494 6252 43546
rect 5956 43492 6012 43494
rect 6036 43492 6092 43494
rect 6116 43492 6172 43494
rect 6196 43492 6252 43494
rect 5956 42458 6012 42460
rect 6036 42458 6092 42460
rect 6116 42458 6172 42460
rect 6196 42458 6252 42460
rect 5956 42406 5982 42458
rect 5982 42406 6012 42458
rect 6036 42406 6046 42458
rect 6046 42406 6092 42458
rect 6116 42406 6162 42458
rect 6162 42406 6172 42458
rect 6196 42406 6226 42458
rect 6226 42406 6252 42458
rect 5956 42404 6012 42406
rect 6036 42404 6092 42406
rect 6116 42404 6172 42406
rect 6196 42404 6252 42406
rect 5956 41370 6012 41372
rect 6036 41370 6092 41372
rect 6116 41370 6172 41372
rect 6196 41370 6252 41372
rect 5956 41318 5982 41370
rect 5982 41318 6012 41370
rect 6036 41318 6046 41370
rect 6046 41318 6092 41370
rect 6116 41318 6162 41370
rect 6162 41318 6172 41370
rect 6196 41318 6226 41370
rect 6226 41318 6252 41370
rect 5956 41316 6012 41318
rect 6036 41316 6092 41318
rect 6116 41316 6172 41318
rect 6196 41316 6252 41318
rect 5956 40282 6012 40284
rect 6036 40282 6092 40284
rect 6116 40282 6172 40284
rect 6196 40282 6252 40284
rect 5956 40230 5982 40282
rect 5982 40230 6012 40282
rect 6036 40230 6046 40282
rect 6046 40230 6092 40282
rect 6116 40230 6162 40282
rect 6162 40230 6172 40282
rect 6196 40230 6226 40282
rect 6226 40230 6252 40282
rect 5956 40228 6012 40230
rect 6036 40228 6092 40230
rect 6116 40228 6172 40230
rect 6196 40228 6252 40230
rect 5956 39194 6012 39196
rect 6036 39194 6092 39196
rect 6116 39194 6172 39196
rect 6196 39194 6252 39196
rect 5956 39142 5982 39194
rect 5982 39142 6012 39194
rect 6036 39142 6046 39194
rect 6046 39142 6092 39194
rect 6116 39142 6162 39194
rect 6162 39142 6172 39194
rect 6196 39142 6226 39194
rect 6226 39142 6252 39194
rect 5956 39140 6012 39142
rect 6036 39140 6092 39142
rect 6116 39140 6172 39142
rect 6196 39140 6252 39142
rect 5956 38106 6012 38108
rect 6036 38106 6092 38108
rect 6116 38106 6172 38108
rect 6196 38106 6252 38108
rect 5956 38054 5982 38106
rect 5982 38054 6012 38106
rect 6036 38054 6046 38106
rect 6046 38054 6092 38106
rect 6116 38054 6162 38106
rect 6162 38054 6172 38106
rect 6196 38054 6226 38106
rect 6226 38054 6252 38106
rect 5956 38052 6012 38054
rect 6036 38052 6092 38054
rect 6116 38052 6172 38054
rect 6196 38052 6252 38054
rect 4618 36352 4674 36408
rect 5078 37168 5134 37224
rect 4618 35284 4674 35320
rect 4618 35264 4620 35284
rect 4620 35264 4672 35284
rect 4672 35264 4674 35284
rect 5956 37018 6012 37020
rect 6036 37018 6092 37020
rect 6116 37018 6172 37020
rect 6196 37018 6252 37020
rect 5956 36966 5982 37018
rect 5982 36966 6012 37018
rect 6036 36966 6046 37018
rect 6046 36966 6092 37018
rect 6116 36966 6162 37018
rect 6162 36966 6172 37018
rect 6196 36966 6226 37018
rect 6226 36966 6252 37018
rect 5956 36964 6012 36966
rect 6036 36964 6092 36966
rect 6116 36964 6172 36966
rect 6196 36964 6252 36966
rect 5446 36080 5502 36136
rect 3882 34604 3938 34640
rect 3882 34584 3884 34604
rect 3884 34584 3936 34604
rect 3936 34584 3938 34604
rect 3882 33380 3938 33416
rect 3882 33360 3884 33380
rect 3884 33360 3936 33380
rect 3936 33360 3938 33380
rect 3882 32408 3938 32464
rect 4342 34448 4398 34504
rect 4342 34040 4398 34096
rect 4618 33108 4674 33144
rect 4618 33088 4620 33108
rect 4620 33088 4672 33108
rect 4672 33088 4674 33108
rect 4894 32816 4950 32872
rect 3974 31184 4030 31240
rect 3606 30640 3662 30696
rect 5354 34176 5410 34232
rect 5956 35930 6012 35932
rect 6036 35930 6092 35932
rect 6116 35930 6172 35932
rect 6196 35930 6252 35932
rect 5956 35878 5982 35930
rect 5982 35878 6012 35930
rect 6036 35878 6046 35930
rect 6046 35878 6092 35930
rect 6116 35878 6162 35930
rect 6162 35878 6172 35930
rect 6196 35878 6226 35930
rect 6226 35878 6252 35930
rect 5956 35876 6012 35878
rect 6036 35876 6092 35878
rect 6116 35876 6172 35878
rect 6196 35876 6252 35878
rect 6182 35572 6184 35592
rect 6184 35572 6236 35592
rect 6236 35572 6238 35592
rect 6182 35536 6238 35572
rect 5998 35028 6000 35048
rect 6000 35028 6052 35048
rect 6052 35028 6054 35048
rect 5998 34992 6054 35028
rect 5956 34842 6012 34844
rect 6036 34842 6092 34844
rect 6116 34842 6172 34844
rect 6196 34842 6252 34844
rect 5956 34790 5982 34842
rect 5982 34790 6012 34842
rect 6036 34790 6046 34842
rect 6046 34790 6092 34842
rect 6116 34790 6162 34842
rect 6162 34790 6172 34842
rect 6196 34790 6226 34842
rect 6226 34790 6252 34842
rect 5956 34788 6012 34790
rect 6036 34788 6092 34790
rect 6116 34788 6172 34790
rect 6196 34788 6252 34790
rect 5906 34604 5962 34640
rect 5906 34584 5908 34604
rect 5908 34584 5960 34604
rect 5960 34584 5962 34604
rect 5354 33516 5410 33552
rect 5354 33496 5356 33516
rect 5356 33496 5408 33516
rect 5408 33496 5410 33516
rect 6182 33940 6184 33960
rect 6184 33940 6236 33960
rect 6236 33940 6238 33960
rect 6182 33904 6238 33940
rect 5956 33754 6012 33756
rect 6036 33754 6092 33756
rect 6116 33754 6172 33756
rect 6196 33754 6252 33756
rect 5956 33702 5982 33754
rect 5982 33702 6012 33754
rect 6036 33702 6046 33754
rect 6046 33702 6092 33754
rect 6116 33702 6162 33754
rect 6162 33702 6172 33754
rect 6196 33702 6226 33754
rect 6226 33702 6252 33754
rect 5956 33700 6012 33702
rect 6036 33700 6092 33702
rect 6116 33700 6172 33702
rect 6196 33700 6252 33702
rect 5262 32020 5318 32056
rect 5262 32000 5264 32020
rect 5264 32000 5316 32020
rect 5316 32000 5318 32020
rect 5722 32952 5778 33008
rect 5906 32952 5962 33008
rect 5956 32666 6012 32668
rect 6036 32666 6092 32668
rect 6116 32666 6172 32668
rect 6196 32666 6252 32668
rect 5956 32614 5982 32666
rect 5982 32614 6012 32666
rect 6036 32614 6046 32666
rect 6046 32614 6092 32666
rect 6116 32614 6162 32666
rect 6162 32614 6172 32666
rect 6196 32614 6226 32666
rect 6226 32614 6252 32666
rect 5956 32612 6012 32614
rect 6036 32612 6092 32614
rect 6116 32612 6172 32614
rect 6196 32612 6252 32614
rect 5630 32292 5686 32328
rect 5630 32272 5632 32292
rect 5632 32272 5684 32292
rect 5684 32272 5686 32292
rect 5722 31900 5724 31920
rect 5724 31900 5776 31920
rect 5776 31900 5778 31920
rect 5722 31864 5778 31900
rect 5906 32172 5908 32192
rect 5908 32172 5960 32192
rect 5960 32172 5962 32192
rect 5906 32136 5962 32172
rect 5538 31356 5540 31376
rect 5540 31356 5592 31376
rect 5592 31356 5594 31376
rect 5538 31320 5594 31356
rect 5262 30640 5318 30696
rect 4986 29688 5042 29744
rect 4066 27648 4122 27704
rect 4710 28600 4766 28656
rect 4158 27240 4214 27296
rect 5956 31578 6012 31580
rect 6036 31578 6092 31580
rect 6116 31578 6172 31580
rect 6196 31578 6252 31580
rect 5956 31526 5982 31578
rect 5982 31526 6012 31578
rect 6036 31526 6046 31578
rect 6046 31526 6092 31578
rect 6116 31526 6162 31578
rect 6162 31526 6172 31578
rect 6196 31526 6226 31578
rect 6226 31526 6252 31578
rect 5956 31524 6012 31526
rect 6036 31524 6092 31526
rect 6116 31524 6172 31526
rect 6196 31524 6252 31526
rect 5630 30504 5686 30560
rect 5956 30490 6012 30492
rect 6036 30490 6092 30492
rect 6116 30490 6172 30492
rect 6196 30490 6252 30492
rect 5956 30438 5982 30490
rect 5982 30438 6012 30490
rect 6036 30438 6046 30490
rect 6046 30438 6092 30490
rect 6116 30438 6162 30490
rect 6162 30438 6172 30490
rect 6196 30438 6226 30490
rect 6226 30438 6252 30490
rect 5956 30436 6012 30438
rect 6036 30436 6092 30438
rect 6116 30436 6172 30438
rect 6196 30436 6252 30438
rect 5814 29960 5870 30016
rect 5956 29402 6012 29404
rect 6036 29402 6092 29404
rect 6116 29402 6172 29404
rect 6196 29402 6252 29404
rect 5956 29350 5982 29402
rect 5982 29350 6012 29402
rect 6036 29350 6046 29402
rect 6046 29350 6092 29402
rect 6116 29350 6162 29402
rect 6162 29350 6172 29402
rect 6196 29350 6226 29402
rect 6226 29350 6252 29402
rect 5956 29348 6012 29350
rect 6036 29348 6092 29350
rect 6116 29348 6172 29350
rect 6196 29348 6252 29350
rect 6182 29144 6238 29200
rect 5956 28314 6012 28316
rect 6036 28314 6092 28316
rect 6116 28314 6172 28316
rect 6196 28314 6252 28316
rect 5956 28262 5982 28314
rect 5982 28262 6012 28314
rect 6036 28262 6046 28314
rect 6046 28262 6092 28314
rect 6116 28262 6162 28314
rect 6162 28262 6172 28314
rect 6196 28262 6226 28314
rect 6226 28262 6252 28314
rect 5956 28260 6012 28262
rect 6036 28260 6092 28262
rect 6116 28260 6172 28262
rect 6196 28260 6252 28262
rect 5956 27226 6012 27228
rect 6036 27226 6092 27228
rect 6116 27226 6172 27228
rect 6196 27226 6252 27228
rect 5956 27174 5982 27226
rect 5982 27174 6012 27226
rect 6036 27174 6046 27226
rect 6046 27174 6092 27226
rect 6116 27174 6162 27226
rect 6162 27174 6172 27226
rect 6196 27174 6226 27226
rect 6226 27174 6252 27226
rect 5956 27172 6012 27174
rect 6036 27172 6092 27174
rect 6116 27172 6172 27174
rect 6196 27172 6252 27174
rect 5956 26138 6012 26140
rect 6036 26138 6092 26140
rect 6116 26138 6172 26140
rect 6196 26138 6252 26140
rect 5956 26086 5982 26138
rect 5982 26086 6012 26138
rect 6036 26086 6046 26138
rect 6046 26086 6092 26138
rect 6116 26086 6162 26138
rect 6162 26086 6172 26138
rect 6196 26086 6226 26138
rect 6226 26086 6252 26138
rect 5956 26084 6012 26086
rect 6036 26084 6092 26086
rect 6116 26084 6172 26086
rect 6196 26084 6252 26086
rect 5814 25608 5870 25664
rect 5956 25050 6012 25052
rect 6036 25050 6092 25052
rect 6116 25050 6172 25052
rect 6196 25050 6252 25052
rect 5956 24998 5982 25050
rect 5982 24998 6012 25050
rect 6036 24998 6046 25050
rect 6046 24998 6092 25050
rect 6116 24998 6162 25050
rect 6162 24998 6172 25050
rect 6196 24998 6226 25050
rect 6226 24998 6252 25050
rect 5956 24996 6012 24998
rect 6036 24996 6092 24998
rect 6116 24996 6172 24998
rect 6196 24996 6252 24998
rect 6734 44784 6790 44840
rect 6550 36796 6552 36816
rect 6552 36796 6604 36816
rect 6604 36796 6606 36816
rect 6550 36760 6606 36796
rect 6642 35148 6698 35184
rect 6642 35128 6644 35148
rect 6644 35128 6696 35148
rect 6696 35128 6698 35148
rect 6458 34040 6514 34096
rect 6458 33768 6514 33824
rect 6642 33652 6698 33688
rect 6642 33632 6644 33652
rect 6644 33632 6696 33652
rect 6696 33632 6698 33652
rect 6550 33224 6606 33280
rect 6550 32408 6606 32464
rect 6366 31592 6422 31648
rect 6642 31728 6698 31784
rect 6642 31476 6698 31512
rect 6642 31456 6644 31476
rect 6644 31456 6696 31476
rect 6696 31456 6698 31476
rect 6642 29552 6698 29608
rect 6550 28756 6606 28792
rect 6550 28736 6552 28756
rect 6552 28736 6604 28756
rect 6604 28736 6606 28756
rect 6458 28600 6514 28656
rect 6366 27104 6422 27160
rect 6274 24656 6330 24712
rect 5956 23962 6012 23964
rect 6036 23962 6092 23964
rect 6116 23962 6172 23964
rect 6196 23962 6252 23964
rect 5956 23910 5982 23962
rect 5982 23910 6012 23962
rect 6036 23910 6046 23962
rect 6046 23910 6092 23962
rect 6116 23910 6162 23962
rect 6162 23910 6172 23962
rect 6196 23910 6226 23962
rect 6226 23910 6252 23962
rect 5956 23908 6012 23910
rect 6036 23908 6092 23910
rect 6116 23908 6172 23910
rect 6196 23908 6252 23910
rect 5956 22874 6012 22876
rect 6036 22874 6092 22876
rect 6116 22874 6172 22876
rect 6196 22874 6252 22876
rect 5956 22822 5982 22874
rect 5982 22822 6012 22874
rect 6036 22822 6046 22874
rect 6046 22822 6092 22874
rect 6116 22822 6162 22874
rect 6162 22822 6172 22874
rect 6196 22822 6226 22874
rect 6226 22822 6252 22874
rect 5956 22820 6012 22822
rect 6036 22820 6092 22822
rect 6116 22820 6172 22822
rect 6196 22820 6252 22822
rect 5538 22072 5594 22128
rect 5956 21786 6012 21788
rect 6036 21786 6092 21788
rect 6116 21786 6172 21788
rect 6196 21786 6252 21788
rect 5956 21734 5982 21786
rect 5982 21734 6012 21786
rect 6036 21734 6046 21786
rect 6046 21734 6092 21786
rect 6116 21734 6162 21786
rect 6162 21734 6172 21786
rect 6196 21734 6226 21786
rect 6226 21734 6252 21786
rect 5956 21732 6012 21734
rect 6036 21732 6092 21734
rect 6116 21732 6172 21734
rect 6196 21732 6252 21734
rect 6550 27648 6606 27704
rect 6550 26016 6606 26072
rect 6458 21664 6514 21720
rect 6366 21564 6368 21584
rect 6368 21564 6420 21584
rect 6420 21564 6422 21584
rect 6366 21528 6422 21564
rect 5956 20698 6012 20700
rect 6036 20698 6092 20700
rect 6116 20698 6172 20700
rect 6196 20698 6252 20700
rect 5956 20646 5982 20698
rect 5982 20646 6012 20698
rect 6036 20646 6046 20698
rect 6046 20646 6092 20698
rect 6116 20646 6162 20698
rect 6162 20646 6172 20698
rect 6196 20646 6226 20698
rect 6226 20646 6252 20698
rect 5956 20644 6012 20646
rect 6036 20644 6092 20646
rect 6116 20644 6172 20646
rect 6196 20644 6252 20646
rect 5956 19610 6012 19612
rect 6036 19610 6092 19612
rect 6116 19610 6172 19612
rect 6196 19610 6252 19612
rect 5956 19558 5982 19610
rect 5982 19558 6012 19610
rect 6036 19558 6046 19610
rect 6046 19558 6092 19610
rect 6116 19558 6162 19610
rect 6162 19558 6172 19610
rect 6196 19558 6226 19610
rect 6226 19558 6252 19610
rect 5956 19556 6012 19558
rect 6036 19556 6092 19558
rect 6116 19556 6172 19558
rect 6196 19556 6252 19558
rect 6826 36916 6882 36952
rect 6826 36896 6828 36916
rect 6828 36896 6880 36916
rect 6880 36896 6882 36916
rect 6918 34856 6974 34912
rect 6826 33904 6882 33960
rect 7102 34312 7158 34368
rect 6918 33088 6974 33144
rect 7102 33496 7158 33552
rect 7378 50904 7434 50960
rect 7378 46960 7434 47016
rect 6918 30368 6974 30424
rect 6826 29280 6882 29336
rect 7102 29960 7158 30016
rect 7102 27956 7104 27976
rect 7104 27956 7156 27976
rect 7156 27956 7158 27976
rect 7102 27920 7158 27956
rect 7746 73616 7802 73672
rect 7562 73072 7618 73128
rect 9586 77016 9642 77072
rect 9586 76336 9642 76392
rect 10956 77818 11012 77820
rect 11036 77818 11092 77820
rect 11116 77818 11172 77820
rect 11196 77818 11252 77820
rect 10956 77766 10982 77818
rect 10982 77766 11012 77818
rect 11036 77766 11046 77818
rect 11046 77766 11092 77818
rect 11116 77766 11162 77818
rect 11162 77766 11172 77818
rect 11196 77766 11226 77818
rect 11226 77766 11252 77818
rect 10956 77764 11012 77766
rect 11036 77764 11092 77766
rect 11116 77764 11172 77766
rect 11196 77764 11252 77766
rect 10138 75792 10194 75848
rect 9678 74704 9734 74760
rect 7930 60560 7986 60616
rect 7838 51312 7894 51368
rect 7838 48048 7894 48104
rect 7746 44376 7802 44432
rect 7194 26152 7250 26208
rect 7470 26288 7526 26344
rect 7378 25336 7434 25392
rect 6826 23704 6882 23760
rect 7378 21664 7434 21720
rect 6734 19080 6790 19136
rect 5956 18522 6012 18524
rect 6036 18522 6092 18524
rect 6116 18522 6172 18524
rect 6196 18522 6252 18524
rect 5956 18470 5982 18522
rect 5982 18470 6012 18522
rect 6036 18470 6046 18522
rect 6046 18470 6092 18522
rect 6116 18470 6162 18522
rect 6162 18470 6172 18522
rect 6196 18470 6226 18522
rect 6226 18470 6252 18522
rect 5956 18468 6012 18470
rect 6036 18468 6092 18470
rect 6116 18468 6172 18470
rect 6196 18468 6252 18470
rect 5956 17434 6012 17436
rect 6036 17434 6092 17436
rect 6116 17434 6172 17436
rect 6196 17434 6252 17436
rect 5956 17382 5982 17434
rect 5982 17382 6012 17434
rect 6036 17382 6046 17434
rect 6046 17382 6092 17434
rect 6116 17382 6162 17434
rect 6162 17382 6172 17434
rect 6196 17382 6226 17434
rect 6226 17382 6252 17434
rect 5956 17380 6012 17382
rect 6036 17380 6092 17382
rect 6116 17380 6172 17382
rect 6196 17380 6252 17382
rect 3514 10240 3570 10296
rect 3330 8880 3386 8936
rect 5956 16346 6012 16348
rect 6036 16346 6092 16348
rect 6116 16346 6172 16348
rect 6196 16346 6252 16348
rect 5956 16294 5982 16346
rect 5982 16294 6012 16346
rect 6036 16294 6046 16346
rect 6046 16294 6092 16346
rect 6116 16294 6162 16346
rect 6162 16294 6172 16346
rect 6196 16294 6226 16346
rect 6226 16294 6252 16346
rect 5956 16292 6012 16294
rect 6036 16292 6092 16294
rect 6116 16292 6172 16294
rect 6196 16292 6252 16294
rect 3974 11192 4030 11248
rect 3882 10512 3938 10568
rect 3882 6840 3938 6896
rect 5956 15258 6012 15260
rect 6036 15258 6092 15260
rect 6116 15258 6172 15260
rect 6196 15258 6252 15260
rect 5956 15206 5982 15258
rect 5982 15206 6012 15258
rect 6036 15206 6046 15258
rect 6046 15206 6092 15258
rect 6116 15206 6162 15258
rect 6162 15206 6172 15258
rect 6196 15206 6226 15258
rect 6226 15206 6252 15258
rect 5956 15204 6012 15206
rect 6036 15204 6092 15206
rect 6116 15204 6172 15206
rect 6196 15204 6252 15206
rect 5956 14170 6012 14172
rect 6036 14170 6092 14172
rect 6116 14170 6172 14172
rect 6196 14170 6252 14172
rect 5956 14118 5982 14170
rect 5982 14118 6012 14170
rect 6036 14118 6046 14170
rect 6046 14118 6092 14170
rect 6116 14118 6162 14170
rect 6162 14118 6172 14170
rect 6196 14118 6226 14170
rect 6226 14118 6252 14170
rect 5956 14116 6012 14118
rect 6036 14116 6092 14118
rect 6116 14116 6172 14118
rect 6196 14116 6252 14118
rect 5956 13082 6012 13084
rect 6036 13082 6092 13084
rect 6116 13082 6172 13084
rect 6196 13082 6252 13084
rect 5956 13030 5982 13082
rect 5982 13030 6012 13082
rect 6036 13030 6046 13082
rect 6046 13030 6092 13082
rect 6116 13030 6162 13082
rect 6162 13030 6172 13082
rect 6196 13030 6226 13082
rect 6226 13030 6252 13082
rect 5956 13028 6012 13030
rect 6036 13028 6092 13030
rect 6116 13028 6172 13030
rect 6196 13028 6252 13030
rect 5956 11994 6012 11996
rect 6036 11994 6092 11996
rect 6116 11994 6172 11996
rect 6196 11994 6252 11996
rect 5956 11942 5982 11994
rect 5982 11942 6012 11994
rect 6036 11942 6046 11994
rect 6046 11942 6092 11994
rect 6116 11942 6162 11994
rect 6162 11942 6172 11994
rect 6196 11942 6226 11994
rect 6226 11942 6252 11994
rect 5956 11940 6012 11942
rect 6036 11940 6092 11942
rect 6116 11940 6172 11942
rect 6196 11940 6252 11942
rect 7286 15680 7342 15736
rect 7746 35400 7802 35456
rect 7654 34040 7710 34096
rect 7838 34992 7894 35048
rect 7930 34720 7986 34776
rect 7746 33088 7802 33144
rect 7654 32544 7710 32600
rect 7654 25200 7710 25256
rect 7562 15000 7618 15056
rect 6918 11192 6974 11248
rect 4618 11056 4674 11112
rect 5814 11056 5870 11112
rect 4066 10920 4122 10976
rect 4066 10104 4122 10160
rect 4066 6976 4122 7032
rect 3974 4120 4030 4176
rect 4066 3440 4122 3496
rect 3146 1944 3202 2000
rect 2962 856 3018 912
rect 3698 856 3754 912
rect 5956 10906 6012 10908
rect 6036 10906 6092 10908
rect 6116 10906 6172 10908
rect 6196 10906 6252 10908
rect 5956 10854 5982 10906
rect 5982 10854 6012 10906
rect 6036 10854 6046 10906
rect 6046 10854 6092 10906
rect 6116 10854 6162 10906
rect 6162 10854 6172 10906
rect 6196 10854 6226 10906
rect 6226 10854 6252 10906
rect 5956 10852 6012 10854
rect 6036 10852 6092 10854
rect 6116 10852 6172 10854
rect 6196 10852 6252 10854
rect 5956 9818 6012 9820
rect 6036 9818 6092 9820
rect 6116 9818 6172 9820
rect 6196 9818 6252 9820
rect 5956 9766 5982 9818
rect 5982 9766 6012 9818
rect 6036 9766 6046 9818
rect 6046 9766 6092 9818
rect 6116 9766 6162 9818
rect 6162 9766 6172 9818
rect 6196 9766 6226 9818
rect 6226 9766 6252 9818
rect 5956 9764 6012 9766
rect 6036 9764 6092 9766
rect 6116 9764 6172 9766
rect 6196 9764 6252 9766
rect 5956 8730 6012 8732
rect 6036 8730 6092 8732
rect 6116 8730 6172 8732
rect 6196 8730 6252 8732
rect 5956 8678 5982 8730
rect 5982 8678 6012 8730
rect 6036 8678 6046 8730
rect 6046 8678 6092 8730
rect 6116 8678 6162 8730
rect 6162 8678 6172 8730
rect 6196 8678 6226 8730
rect 6226 8678 6252 8730
rect 5956 8676 6012 8678
rect 6036 8676 6092 8678
rect 6116 8676 6172 8678
rect 6196 8676 6252 8678
rect 5956 7642 6012 7644
rect 6036 7642 6092 7644
rect 6116 7642 6172 7644
rect 6196 7642 6252 7644
rect 5956 7590 5982 7642
rect 5982 7590 6012 7642
rect 6036 7590 6046 7642
rect 6046 7590 6092 7642
rect 6116 7590 6162 7642
rect 6162 7590 6172 7642
rect 6196 7590 6226 7642
rect 6226 7590 6252 7642
rect 5956 7588 6012 7590
rect 6036 7588 6092 7590
rect 6116 7588 6172 7590
rect 6196 7588 6252 7590
rect 7654 7520 7710 7576
rect 7930 28872 7986 28928
rect 7838 28500 7840 28520
rect 7840 28500 7892 28520
rect 7892 28500 7894 28520
rect 7838 28464 7894 28500
rect 7930 28328 7986 28384
rect 7838 22752 7894 22808
rect 9126 69400 9182 69456
rect 8206 66136 8262 66192
rect 8758 57160 8814 57216
rect 8390 52148 8446 52184
rect 8390 52128 8392 52148
rect 8392 52128 8444 52148
rect 8444 52128 8446 52148
rect 8206 48184 8262 48240
rect 8298 46552 8354 46608
rect 8942 50224 8998 50280
rect 10956 76730 11012 76732
rect 11036 76730 11092 76732
rect 11116 76730 11172 76732
rect 11196 76730 11252 76732
rect 10956 76678 10982 76730
rect 10982 76678 11012 76730
rect 11036 76678 11046 76730
rect 11046 76678 11092 76730
rect 11116 76678 11162 76730
rect 11162 76678 11172 76730
rect 11196 76678 11226 76730
rect 11226 76678 11252 76730
rect 10956 76676 11012 76678
rect 11036 76676 11092 76678
rect 11116 76676 11172 76678
rect 11196 76676 11252 76678
rect 10956 75642 11012 75644
rect 11036 75642 11092 75644
rect 11116 75642 11172 75644
rect 11196 75642 11252 75644
rect 10956 75590 10982 75642
rect 10982 75590 11012 75642
rect 11036 75590 11046 75642
rect 11046 75590 11092 75642
rect 11116 75590 11162 75642
rect 11162 75590 11172 75642
rect 11196 75590 11226 75642
rect 11226 75590 11252 75642
rect 10956 75588 11012 75590
rect 11036 75588 11092 75590
rect 11116 75588 11172 75590
rect 11196 75588 11252 75590
rect 10956 74554 11012 74556
rect 11036 74554 11092 74556
rect 11116 74554 11172 74556
rect 11196 74554 11252 74556
rect 10956 74502 10982 74554
rect 10982 74502 11012 74554
rect 11036 74502 11046 74554
rect 11046 74502 11092 74554
rect 11116 74502 11162 74554
rect 11162 74502 11172 74554
rect 11196 74502 11226 74554
rect 11226 74502 11252 74554
rect 10956 74500 11012 74502
rect 11036 74500 11092 74502
rect 11116 74500 11172 74502
rect 11196 74500 11252 74502
rect 10956 73466 11012 73468
rect 11036 73466 11092 73468
rect 11116 73466 11172 73468
rect 11196 73466 11252 73468
rect 10956 73414 10982 73466
rect 10982 73414 11012 73466
rect 11036 73414 11046 73466
rect 11046 73414 11092 73466
rect 11116 73414 11162 73466
rect 11162 73414 11172 73466
rect 11196 73414 11226 73466
rect 11226 73414 11252 73466
rect 10956 73412 11012 73414
rect 11036 73412 11092 73414
rect 11116 73412 11172 73414
rect 11196 73412 11252 73414
rect 11518 73208 11574 73264
rect 10956 72378 11012 72380
rect 11036 72378 11092 72380
rect 11116 72378 11172 72380
rect 11196 72378 11252 72380
rect 10956 72326 10982 72378
rect 10982 72326 11012 72378
rect 11036 72326 11046 72378
rect 11046 72326 11092 72378
rect 11116 72326 11162 72378
rect 11162 72326 11172 72378
rect 11196 72326 11226 72378
rect 11226 72326 11252 72378
rect 10956 72324 11012 72326
rect 11036 72324 11092 72326
rect 11116 72324 11172 72326
rect 11196 72324 11252 72326
rect 10956 71290 11012 71292
rect 11036 71290 11092 71292
rect 11116 71290 11172 71292
rect 11196 71290 11252 71292
rect 10956 71238 10982 71290
rect 10982 71238 11012 71290
rect 11036 71238 11046 71290
rect 11046 71238 11092 71290
rect 11116 71238 11162 71290
rect 11162 71238 11172 71290
rect 11196 71238 11226 71290
rect 11226 71238 11252 71290
rect 10956 71236 11012 71238
rect 11036 71236 11092 71238
rect 11116 71236 11172 71238
rect 11196 71236 11252 71238
rect 10956 70202 11012 70204
rect 11036 70202 11092 70204
rect 11116 70202 11172 70204
rect 11196 70202 11252 70204
rect 10956 70150 10982 70202
rect 10982 70150 11012 70202
rect 11036 70150 11046 70202
rect 11046 70150 11092 70202
rect 11116 70150 11162 70202
rect 11162 70150 11172 70202
rect 11196 70150 11226 70202
rect 11226 70150 11252 70202
rect 10956 70148 11012 70150
rect 11036 70148 11092 70150
rect 11116 70148 11172 70150
rect 11196 70148 11252 70150
rect 10782 69400 10838 69456
rect 10956 69114 11012 69116
rect 11036 69114 11092 69116
rect 11116 69114 11172 69116
rect 11196 69114 11252 69116
rect 10956 69062 10982 69114
rect 10982 69062 11012 69114
rect 11036 69062 11046 69114
rect 11046 69062 11092 69114
rect 11116 69062 11162 69114
rect 11162 69062 11172 69114
rect 11196 69062 11226 69114
rect 11226 69062 11252 69114
rect 10956 69060 11012 69062
rect 11036 69060 11092 69062
rect 11116 69060 11172 69062
rect 11196 69060 11252 69062
rect 11518 68856 11574 68912
rect 10956 68026 11012 68028
rect 11036 68026 11092 68028
rect 11116 68026 11172 68028
rect 11196 68026 11252 68028
rect 10956 67974 10982 68026
rect 10982 67974 11012 68026
rect 11036 67974 11046 68026
rect 11046 67974 11092 68026
rect 11116 67974 11162 68026
rect 11162 67974 11172 68026
rect 11196 67974 11226 68026
rect 11226 67974 11252 68026
rect 10956 67972 11012 67974
rect 11036 67972 11092 67974
rect 11116 67972 11172 67974
rect 11196 67972 11252 67974
rect 12162 75828 12164 75848
rect 12164 75828 12216 75848
rect 12216 75828 12218 75848
rect 12162 75792 12218 75828
rect 11242 67652 11298 67688
rect 11242 67632 11244 67652
rect 11244 67632 11296 67652
rect 11296 67632 11298 67652
rect 11610 67632 11666 67688
rect 11978 67652 12034 67688
rect 11978 67632 11980 67652
rect 11980 67632 12032 67652
rect 12032 67632 12034 67652
rect 13726 76356 13782 76392
rect 13726 76336 13728 76356
rect 13728 76336 13780 76356
rect 13780 76336 13782 76356
rect 13358 75792 13414 75848
rect 13358 75692 13360 75712
rect 13360 75692 13412 75712
rect 13412 75692 13414 75712
rect 13358 75656 13414 75692
rect 15106 75792 15162 75848
rect 12622 70352 12678 70408
rect 12254 67496 12310 67552
rect 11518 67360 11574 67416
rect 10956 66938 11012 66940
rect 11036 66938 11092 66940
rect 11116 66938 11172 66940
rect 11196 66938 11252 66940
rect 10956 66886 10982 66938
rect 10982 66886 11012 66938
rect 11036 66886 11046 66938
rect 11046 66886 11092 66938
rect 11116 66886 11162 66938
rect 11162 66886 11172 66938
rect 11196 66886 11226 66938
rect 11226 66886 11252 66938
rect 10956 66884 11012 66886
rect 11036 66884 11092 66886
rect 11116 66884 11172 66886
rect 11196 66884 11252 66886
rect 10956 65850 11012 65852
rect 11036 65850 11092 65852
rect 11116 65850 11172 65852
rect 11196 65850 11252 65852
rect 10956 65798 10982 65850
rect 10982 65798 11012 65850
rect 11036 65798 11046 65850
rect 11046 65798 11092 65850
rect 11116 65798 11162 65850
rect 11162 65798 11172 65850
rect 11196 65798 11226 65850
rect 11226 65798 11252 65850
rect 10956 65796 11012 65798
rect 11036 65796 11092 65798
rect 11116 65796 11172 65798
rect 11196 65796 11252 65798
rect 10956 64762 11012 64764
rect 11036 64762 11092 64764
rect 11116 64762 11172 64764
rect 11196 64762 11252 64764
rect 10956 64710 10982 64762
rect 10982 64710 11012 64762
rect 11036 64710 11046 64762
rect 11046 64710 11092 64762
rect 11116 64710 11162 64762
rect 11162 64710 11172 64762
rect 11196 64710 11226 64762
rect 11226 64710 11252 64762
rect 10956 64708 11012 64710
rect 11036 64708 11092 64710
rect 11116 64708 11172 64710
rect 11196 64708 11252 64710
rect 10956 63674 11012 63676
rect 11036 63674 11092 63676
rect 11116 63674 11172 63676
rect 11196 63674 11252 63676
rect 10956 63622 10982 63674
rect 10982 63622 11012 63674
rect 11036 63622 11046 63674
rect 11046 63622 11092 63674
rect 11116 63622 11162 63674
rect 11162 63622 11172 63674
rect 11196 63622 11226 63674
rect 11226 63622 11252 63674
rect 10956 63620 11012 63622
rect 11036 63620 11092 63622
rect 11116 63620 11172 63622
rect 11196 63620 11252 63622
rect 10956 62586 11012 62588
rect 11036 62586 11092 62588
rect 11116 62586 11172 62588
rect 11196 62586 11252 62588
rect 10956 62534 10982 62586
rect 10982 62534 11012 62586
rect 11036 62534 11046 62586
rect 11046 62534 11092 62586
rect 11116 62534 11162 62586
rect 11162 62534 11172 62586
rect 11196 62534 11226 62586
rect 11226 62534 11252 62586
rect 10956 62532 11012 62534
rect 11036 62532 11092 62534
rect 11116 62532 11172 62534
rect 11196 62532 11252 62534
rect 10956 61498 11012 61500
rect 11036 61498 11092 61500
rect 11116 61498 11172 61500
rect 11196 61498 11252 61500
rect 10956 61446 10982 61498
rect 10982 61446 11012 61498
rect 11036 61446 11046 61498
rect 11046 61446 11092 61498
rect 11116 61446 11162 61498
rect 11162 61446 11172 61498
rect 11196 61446 11226 61498
rect 11226 61446 11252 61498
rect 10956 61444 11012 61446
rect 11036 61444 11092 61446
rect 11116 61444 11172 61446
rect 11196 61444 11252 61446
rect 10956 60410 11012 60412
rect 11036 60410 11092 60412
rect 11116 60410 11172 60412
rect 11196 60410 11252 60412
rect 10956 60358 10982 60410
rect 10982 60358 11012 60410
rect 11036 60358 11046 60410
rect 11046 60358 11092 60410
rect 11116 60358 11162 60410
rect 11162 60358 11172 60410
rect 11196 60358 11226 60410
rect 11226 60358 11252 60410
rect 10956 60356 11012 60358
rect 11036 60356 11092 60358
rect 11116 60356 11172 60358
rect 11196 60356 11252 60358
rect 10956 59322 11012 59324
rect 11036 59322 11092 59324
rect 11116 59322 11172 59324
rect 11196 59322 11252 59324
rect 10956 59270 10982 59322
rect 10982 59270 11012 59322
rect 11036 59270 11046 59322
rect 11046 59270 11092 59322
rect 11116 59270 11162 59322
rect 11162 59270 11172 59322
rect 11196 59270 11226 59322
rect 11226 59270 11252 59322
rect 10956 59268 11012 59270
rect 11036 59268 11092 59270
rect 11116 59268 11172 59270
rect 11196 59268 11252 59270
rect 10956 58234 11012 58236
rect 11036 58234 11092 58236
rect 11116 58234 11172 58236
rect 11196 58234 11252 58236
rect 10956 58182 10982 58234
rect 10982 58182 11012 58234
rect 11036 58182 11046 58234
rect 11046 58182 11092 58234
rect 11116 58182 11162 58234
rect 11162 58182 11172 58234
rect 11196 58182 11226 58234
rect 11226 58182 11252 58234
rect 10956 58180 11012 58182
rect 11036 58180 11092 58182
rect 11116 58180 11172 58182
rect 11196 58180 11252 58182
rect 11518 57976 11574 58032
rect 10956 57146 11012 57148
rect 11036 57146 11092 57148
rect 11116 57146 11172 57148
rect 11196 57146 11252 57148
rect 10956 57094 10982 57146
rect 10982 57094 11012 57146
rect 11036 57094 11046 57146
rect 11046 57094 11092 57146
rect 11116 57094 11162 57146
rect 11162 57094 11172 57146
rect 11196 57094 11226 57146
rect 11226 57094 11252 57146
rect 10956 57092 11012 57094
rect 11036 57092 11092 57094
rect 11116 57092 11172 57094
rect 11196 57092 11252 57094
rect 10956 56058 11012 56060
rect 11036 56058 11092 56060
rect 11116 56058 11172 56060
rect 11196 56058 11252 56060
rect 10956 56006 10982 56058
rect 10982 56006 11012 56058
rect 11036 56006 11046 56058
rect 11046 56006 11092 56058
rect 11116 56006 11162 56058
rect 11162 56006 11172 56058
rect 11196 56006 11226 56058
rect 11226 56006 11252 56058
rect 10956 56004 11012 56006
rect 11036 56004 11092 56006
rect 11116 56004 11172 56006
rect 11196 56004 11252 56006
rect 10956 54970 11012 54972
rect 11036 54970 11092 54972
rect 11116 54970 11172 54972
rect 11196 54970 11252 54972
rect 10956 54918 10982 54970
rect 10982 54918 11012 54970
rect 11036 54918 11046 54970
rect 11046 54918 11092 54970
rect 11116 54918 11162 54970
rect 11162 54918 11172 54970
rect 11196 54918 11226 54970
rect 11226 54918 11252 54970
rect 10956 54916 11012 54918
rect 11036 54916 11092 54918
rect 11116 54916 11172 54918
rect 11196 54916 11252 54918
rect 11518 54032 11574 54088
rect 10956 53882 11012 53884
rect 11036 53882 11092 53884
rect 11116 53882 11172 53884
rect 11196 53882 11252 53884
rect 10956 53830 10982 53882
rect 10982 53830 11012 53882
rect 11036 53830 11046 53882
rect 11046 53830 11092 53882
rect 11116 53830 11162 53882
rect 11162 53830 11172 53882
rect 11196 53830 11226 53882
rect 11226 53830 11252 53882
rect 10956 53828 11012 53830
rect 11036 53828 11092 53830
rect 11116 53828 11172 53830
rect 11196 53828 11252 53830
rect 11610 53624 11666 53680
rect 11426 53388 11428 53408
rect 11428 53388 11480 53408
rect 11480 53388 11482 53408
rect 11426 53352 11482 53388
rect 10956 52794 11012 52796
rect 11036 52794 11092 52796
rect 11116 52794 11172 52796
rect 11196 52794 11252 52796
rect 10956 52742 10982 52794
rect 10982 52742 11012 52794
rect 11036 52742 11046 52794
rect 11046 52742 11092 52794
rect 11116 52742 11162 52794
rect 11162 52742 11172 52794
rect 11196 52742 11226 52794
rect 11226 52742 11252 52794
rect 10956 52740 11012 52742
rect 11036 52740 11092 52742
rect 11116 52740 11172 52742
rect 11196 52740 11252 52742
rect 11334 52672 11390 52728
rect 10414 51312 10470 51368
rect 10966 52264 11022 52320
rect 10956 51706 11012 51708
rect 11036 51706 11092 51708
rect 11116 51706 11172 51708
rect 11196 51706 11252 51708
rect 10956 51654 10982 51706
rect 10982 51654 11012 51706
rect 11036 51654 11046 51706
rect 11046 51654 11092 51706
rect 11116 51654 11162 51706
rect 11162 51654 11172 51706
rect 11196 51654 11226 51706
rect 11226 51654 11252 51706
rect 10956 51652 11012 51654
rect 11036 51652 11092 51654
rect 11116 51652 11172 51654
rect 11196 51652 11252 51654
rect 11610 52400 11666 52456
rect 12070 56752 12126 56808
rect 12162 55800 12218 55856
rect 11794 55664 11850 55720
rect 12070 55392 12126 55448
rect 11886 54188 11942 54224
rect 11886 54168 11888 54188
rect 11888 54168 11940 54188
rect 11940 54168 11942 54188
rect 11886 53896 11942 53952
rect 11702 52128 11758 52184
rect 11518 50940 11520 50960
rect 11520 50940 11572 50960
rect 11572 50940 11574 50960
rect 11518 50904 11574 50940
rect 10956 50618 11012 50620
rect 11036 50618 11092 50620
rect 11116 50618 11172 50620
rect 11196 50618 11252 50620
rect 10956 50566 10982 50618
rect 10982 50566 11012 50618
rect 11036 50566 11046 50618
rect 11046 50566 11092 50618
rect 11116 50566 11162 50618
rect 11162 50566 11172 50618
rect 11196 50566 11226 50618
rect 11226 50566 11252 50618
rect 10956 50564 11012 50566
rect 11036 50564 11092 50566
rect 11116 50564 11172 50566
rect 11196 50564 11252 50566
rect 10506 49816 10562 49872
rect 10956 49530 11012 49532
rect 11036 49530 11092 49532
rect 11116 49530 11172 49532
rect 11196 49530 11252 49532
rect 10956 49478 10982 49530
rect 10982 49478 11012 49530
rect 11036 49478 11046 49530
rect 11046 49478 11092 49530
rect 11116 49478 11162 49530
rect 11162 49478 11172 49530
rect 11196 49478 11226 49530
rect 11226 49478 11252 49530
rect 10956 49476 11012 49478
rect 11036 49476 11092 49478
rect 11116 49476 11172 49478
rect 11196 49476 11252 49478
rect 10956 48442 11012 48444
rect 11036 48442 11092 48444
rect 11116 48442 11172 48444
rect 11196 48442 11252 48444
rect 10956 48390 10982 48442
rect 10982 48390 11012 48442
rect 11036 48390 11046 48442
rect 11046 48390 11092 48442
rect 11116 48390 11162 48442
rect 11162 48390 11172 48442
rect 11196 48390 11226 48442
rect 11226 48390 11252 48442
rect 10956 48388 11012 48390
rect 11036 48388 11092 48390
rect 11116 48388 11172 48390
rect 11196 48388 11252 48390
rect 11426 48184 11482 48240
rect 9402 48048 9458 48104
rect 8574 43852 8630 43888
rect 8574 43832 8576 43852
rect 8576 43832 8628 43852
rect 8628 43832 8630 43852
rect 8758 43852 8814 43888
rect 8758 43832 8760 43852
rect 8760 43832 8812 43852
rect 8812 43832 8814 43852
rect 9218 42100 9220 42120
rect 9220 42100 9272 42120
rect 9272 42100 9274 42120
rect 8298 38800 8354 38856
rect 8206 37748 8208 37768
rect 8208 37748 8260 37768
rect 8260 37748 8262 37768
rect 8206 37712 8262 37748
rect 8666 38392 8722 38448
rect 8298 37032 8354 37088
rect 8206 36760 8262 36816
rect 8206 33396 8208 33416
rect 8208 33396 8260 33416
rect 8260 33396 8262 33416
rect 8206 33360 8262 33396
rect 8482 37304 8538 37360
rect 8574 36352 8630 36408
rect 8482 34720 8538 34776
rect 8298 32428 8354 32464
rect 8298 32408 8300 32428
rect 8300 32408 8352 32428
rect 8352 32408 8354 32428
rect 8206 31184 8262 31240
rect 8206 29416 8262 29472
rect 8298 29144 8354 29200
rect 8114 29028 8170 29064
rect 8114 29008 8116 29028
rect 8116 29008 8168 29028
rect 8168 29008 8170 29028
rect 8666 34484 8668 34504
rect 8668 34484 8720 34504
rect 8720 34484 8722 34504
rect 8666 34448 8722 34484
rect 9218 42064 9274 42100
rect 9034 41420 9036 41440
rect 9036 41420 9088 41440
rect 9088 41420 9090 41440
rect 9034 41384 9090 41420
rect 9034 38120 9090 38176
rect 10956 47354 11012 47356
rect 11036 47354 11092 47356
rect 11116 47354 11172 47356
rect 11196 47354 11252 47356
rect 10956 47302 10982 47354
rect 10982 47302 11012 47354
rect 11036 47302 11046 47354
rect 11046 47302 11092 47354
rect 11116 47302 11162 47354
rect 11162 47302 11172 47354
rect 11196 47302 11226 47354
rect 11226 47302 11252 47354
rect 10956 47300 11012 47302
rect 11036 47300 11092 47302
rect 11116 47300 11172 47302
rect 11196 47300 11252 47302
rect 9770 46960 9826 47016
rect 9494 46416 9550 46472
rect 10956 46266 11012 46268
rect 11036 46266 11092 46268
rect 11116 46266 11172 46268
rect 11196 46266 11252 46268
rect 10956 46214 10982 46266
rect 10982 46214 11012 46266
rect 11036 46214 11046 46266
rect 11046 46214 11092 46266
rect 11116 46214 11162 46266
rect 11162 46214 11172 46266
rect 11196 46214 11226 46266
rect 11226 46214 11252 46266
rect 10956 46212 11012 46214
rect 11036 46212 11092 46214
rect 11116 46212 11172 46214
rect 11196 46212 11252 46214
rect 10956 45178 11012 45180
rect 11036 45178 11092 45180
rect 11116 45178 11172 45180
rect 11196 45178 11252 45180
rect 10956 45126 10982 45178
rect 10982 45126 11012 45178
rect 11036 45126 11046 45178
rect 11046 45126 11092 45178
rect 11116 45126 11162 45178
rect 11162 45126 11172 45178
rect 11196 45126 11226 45178
rect 11226 45126 11252 45178
rect 10956 45124 11012 45126
rect 11036 45124 11092 45126
rect 11116 45124 11172 45126
rect 11196 45124 11252 45126
rect 10598 43052 10600 43072
rect 10600 43052 10652 43072
rect 10652 43052 10654 43072
rect 10598 43016 10654 43052
rect 9402 37984 9458 38040
rect 8850 36216 8906 36272
rect 8574 31728 8630 31784
rect 9126 35672 9182 35728
rect 8942 34992 8998 35048
rect 8942 34720 8998 34776
rect 8850 32000 8906 32056
rect 9126 34856 9182 34912
rect 9126 32988 9128 33008
rect 9128 32988 9180 33008
rect 9180 32988 9182 33008
rect 9126 32952 9182 32988
rect 9034 32136 9090 32192
rect 8850 31728 8906 31784
rect 8390 28736 8446 28792
rect 8942 31628 8944 31648
rect 8944 31628 8996 31648
rect 8996 31628 8998 31648
rect 8942 31592 8998 31628
rect 8850 31048 8906 31104
rect 8666 30504 8722 30560
rect 8758 29688 8814 29744
rect 8390 27648 8446 27704
rect 8114 27376 8170 27432
rect 8666 27240 8722 27296
rect 9494 35400 9550 35456
rect 10956 44090 11012 44092
rect 11036 44090 11092 44092
rect 11116 44090 11172 44092
rect 11196 44090 11252 44092
rect 10956 44038 10982 44090
rect 10982 44038 11012 44090
rect 11036 44038 11046 44090
rect 11046 44038 11092 44090
rect 11116 44038 11162 44090
rect 11162 44038 11172 44090
rect 11196 44038 11226 44090
rect 11226 44038 11252 44090
rect 10956 44036 11012 44038
rect 11036 44036 11092 44038
rect 11116 44036 11172 44038
rect 11196 44036 11252 44038
rect 10956 43002 11012 43004
rect 11036 43002 11092 43004
rect 11116 43002 11172 43004
rect 11196 43002 11252 43004
rect 10956 42950 10982 43002
rect 10982 42950 11012 43002
rect 11036 42950 11046 43002
rect 11046 42950 11092 43002
rect 11116 42950 11162 43002
rect 11162 42950 11172 43002
rect 11196 42950 11226 43002
rect 11226 42950 11252 43002
rect 10956 42948 11012 42950
rect 11036 42948 11092 42950
rect 11116 42948 11172 42950
rect 11196 42948 11252 42950
rect 10782 42064 10838 42120
rect 10956 41914 11012 41916
rect 11036 41914 11092 41916
rect 11116 41914 11172 41916
rect 11196 41914 11252 41916
rect 10956 41862 10982 41914
rect 10982 41862 11012 41914
rect 11036 41862 11046 41914
rect 11046 41862 11092 41914
rect 11116 41862 11162 41914
rect 11162 41862 11172 41914
rect 11196 41862 11226 41914
rect 11226 41862 11252 41914
rect 10956 41860 11012 41862
rect 11036 41860 11092 41862
rect 11116 41860 11172 41862
rect 11196 41860 11252 41862
rect 10414 41384 10470 41440
rect 9954 40044 10010 40080
rect 9954 40024 9956 40044
rect 9956 40024 10008 40044
rect 10008 40024 10010 40044
rect 9862 37612 9864 37632
rect 9864 37612 9916 37632
rect 9916 37612 9918 37632
rect 9862 37576 9918 37612
rect 9678 35944 9734 36000
rect 9954 35400 10010 35456
rect 10230 37712 10286 37768
rect 9678 34720 9734 34776
rect 9586 34312 9642 34368
rect 9586 32972 9642 33008
rect 9586 32952 9588 32972
rect 9588 32952 9640 32972
rect 9640 32952 9642 32972
rect 9310 32000 9366 32056
rect 9494 31592 9550 31648
rect 9126 28636 9128 28656
rect 9128 28636 9180 28656
rect 9180 28636 9182 28656
rect 9126 28600 9182 28636
rect 8942 28212 8998 28248
rect 8942 28192 8944 28212
rect 8944 28192 8996 28212
rect 8996 28192 8998 28212
rect 8482 25064 8538 25120
rect 8574 24112 8630 24168
rect 8114 21392 8170 21448
rect 8206 20304 8262 20360
rect 8758 26288 8814 26344
rect 9586 31184 9642 31240
rect 9126 25744 9182 25800
rect 10138 34312 10194 34368
rect 10322 35264 10378 35320
rect 10956 40826 11012 40828
rect 11036 40826 11092 40828
rect 11116 40826 11172 40828
rect 11196 40826 11252 40828
rect 10956 40774 10982 40826
rect 10982 40774 11012 40826
rect 11036 40774 11046 40826
rect 11046 40774 11092 40826
rect 11116 40774 11162 40826
rect 11162 40774 11172 40826
rect 11196 40774 11226 40826
rect 11226 40774 11252 40826
rect 10956 40772 11012 40774
rect 11036 40772 11092 40774
rect 11116 40772 11172 40774
rect 11196 40772 11252 40774
rect 10956 39738 11012 39740
rect 11036 39738 11092 39740
rect 11116 39738 11172 39740
rect 11196 39738 11252 39740
rect 10956 39686 10982 39738
rect 10982 39686 11012 39738
rect 11036 39686 11046 39738
rect 11046 39686 11092 39738
rect 11116 39686 11162 39738
rect 11162 39686 11172 39738
rect 11196 39686 11226 39738
rect 11226 39686 11252 39738
rect 10956 39684 11012 39686
rect 11036 39684 11092 39686
rect 11116 39684 11172 39686
rect 11196 39684 11252 39686
rect 11426 39616 11482 39672
rect 10956 38650 11012 38652
rect 11036 38650 11092 38652
rect 11116 38650 11172 38652
rect 11196 38650 11252 38652
rect 10956 38598 10982 38650
rect 10982 38598 11012 38650
rect 11036 38598 11046 38650
rect 11046 38598 11092 38650
rect 11116 38598 11162 38650
rect 11162 38598 11172 38650
rect 11196 38598 11226 38650
rect 11226 38598 11252 38650
rect 10956 38596 11012 38598
rect 11036 38596 11092 38598
rect 11116 38596 11172 38598
rect 11196 38596 11252 38598
rect 10874 38412 10930 38448
rect 10874 38392 10876 38412
rect 10876 38392 10928 38412
rect 10928 38392 10930 38412
rect 11334 37984 11390 38040
rect 10956 37562 11012 37564
rect 11036 37562 11092 37564
rect 11116 37562 11172 37564
rect 11196 37562 11252 37564
rect 10956 37510 10982 37562
rect 10982 37510 11012 37562
rect 11036 37510 11046 37562
rect 11046 37510 11092 37562
rect 11116 37510 11162 37562
rect 11162 37510 11172 37562
rect 11196 37510 11226 37562
rect 11226 37510 11252 37562
rect 10956 37508 11012 37510
rect 11036 37508 11092 37510
rect 11116 37508 11172 37510
rect 11196 37508 11252 37510
rect 10874 37340 10876 37360
rect 10876 37340 10928 37360
rect 10928 37340 10930 37360
rect 10874 37304 10930 37340
rect 11242 37168 11298 37224
rect 11058 36916 11114 36952
rect 11058 36896 11060 36916
rect 11060 36896 11112 36916
rect 11112 36896 11114 36916
rect 11150 36780 11206 36816
rect 11150 36760 11152 36780
rect 11152 36760 11204 36780
rect 11204 36760 11206 36780
rect 10956 36474 11012 36476
rect 11036 36474 11092 36476
rect 11116 36474 11172 36476
rect 11196 36474 11252 36476
rect 10956 36422 10982 36474
rect 10982 36422 11012 36474
rect 11036 36422 11046 36474
rect 11046 36422 11092 36474
rect 11116 36422 11162 36474
rect 11162 36422 11172 36474
rect 11196 36422 11226 36474
rect 11226 36422 11252 36474
rect 10956 36420 11012 36422
rect 11036 36420 11092 36422
rect 11116 36420 11172 36422
rect 11196 36420 11252 36422
rect 10598 35028 10600 35048
rect 10600 35028 10652 35048
rect 10652 35028 10654 35048
rect 10598 34992 10654 35028
rect 10690 34856 10746 34912
rect 10506 34584 10562 34640
rect 10506 34196 10562 34232
rect 10506 34176 10508 34196
rect 10508 34176 10560 34196
rect 10560 34176 10562 34196
rect 10322 32972 10378 33008
rect 10322 32952 10324 32972
rect 10324 32952 10376 32972
rect 10376 32952 10378 32972
rect 10046 32020 10102 32056
rect 10046 32000 10048 32020
rect 10048 32000 10100 32020
rect 10100 32000 10102 32020
rect 9954 31048 10010 31104
rect 9954 30776 10010 30832
rect 11426 35808 11482 35864
rect 10956 35386 11012 35388
rect 11036 35386 11092 35388
rect 11116 35386 11172 35388
rect 11196 35386 11252 35388
rect 10956 35334 10982 35386
rect 10982 35334 11012 35386
rect 11036 35334 11046 35386
rect 11046 35334 11092 35386
rect 11116 35334 11162 35386
rect 11162 35334 11172 35386
rect 11196 35334 11226 35386
rect 11226 35334 11252 35386
rect 10956 35332 11012 35334
rect 11036 35332 11092 35334
rect 11116 35332 11172 35334
rect 11196 35332 11252 35334
rect 10956 34298 11012 34300
rect 11036 34298 11092 34300
rect 11116 34298 11172 34300
rect 11196 34298 11252 34300
rect 10956 34246 10982 34298
rect 10982 34246 11012 34298
rect 11036 34246 11046 34298
rect 11046 34246 11092 34298
rect 11116 34246 11162 34298
rect 11162 34246 11172 34298
rect 11196 34246 11226 34298
rect 11226 34246 11252 34298
rect 10956 34244 11012 34246
rect 11036 34244 11092 34246
rect 11116 34244 11172 34246
rect 11196 34244 11252 34246
rect 10782 33224 10838 33280
rect 10782 32544 10838 32600
rect 10506 31884 10562 31920
rect 10506 31864 10508 31884
rect 10508 31864 10560 31884
rect 10560 31864 10562 31884
rect 10230 31456 10286 31512
rect 10506 31220 10508 31240
rect 10508 31220 10560 31240
rect 10560 31220 10562 31240
rect 10506 31184 10562 31220
rect 10322 30776 10378 30832
rect 9678 28464 9734 28520
rect 8942 21528 8998 21584
rect 8114 15544 8170 15600
rect 8666 15952 8722 16008
rect 8390 13232 8446 13288
rect 7930 9016 7986 9072
rect 8942 19508 8998 19544
rect 8942 19488 8944 19508
rect 8944 19488 8996 19508
rect 8996 19488 8998 19508
rect 9034 19216 9090 19272
rect 9218 23160 9274 23216
rect 9310 20304 9366 20360
rect 9494 20596 9550 20632
rect 9494 20576 9496 20596
rect 9496 20576 9548 20596
rect 9548 20576 9550 20596
rect 9770 27784 9826 27840
rect 10138 29996 10140 30016
rect 10140 29996 10192 30016
rect 10192 29996 10194 30016
rect 10138 29960 10194 29996
rect 10138 29688 10194 29744
rect 10138 29008 10194 29064
rect 10046 28328 10102 28384
rect 9770 22888 9826 22944
rect 10046 25200 10102 25256
rect 9954 21972 9956 21992
rect 9956 21972 10008 21992
rect 10008 21972 10010 21992
rect 9954 21936 10010 21972
rect 9862 21392 9918 21448
rect 9678 20440 9734 20496
rect 9678 20168 9734 20224
rect 9770 19216 9826 19272
rect 9586 17720 9642 17776
rect 9494 17040 9550 17096
rect 10414 27376 10470 27432
rect 10690 28736 10746 28792
rect 10690 28464 10746 28520
rect 10322 26152 10378 26208
rect 10322 25880 10378 25936
rect 10322 21664 10378 21720
rect 10230 19488 10286 19544
rect 10046 15544 10102 15600
rect 9770 13232 9826 13288
rect 10690 25644 10692 25664
rect 10692 25644 10744 25664
rect 10744 25644 10746 25664
rect 10690 25608 10746 25644
rect 10598 22480 10654 22536
rect 10956 33210 11012 33212
rect 11036 33210 11092 33212
rect 11116 33210 11172 33212
rect 11196 33210 11252 33212
rect 10956 33158 10982 33210
rect 10982 33158 11012 33210
rect 11036 33158 11046 33210
rect 11046 33158 11092 33210
rect 11116 33158 11162 33210
rect 11162 33158 11172 33210
rect 11196 33158 11226 33210
rect 11226 33158 11252 33210
rect 10956 33156 11012 33158
rect 11036 33156 11092 33158
rect 11116 33156 11172 33158
rect 11196 33156 11252 33158
rect 11242 32408 11298 32464
rect 10956 32122 11012 32124
rect 11036 32122 11092 32124
rect 11116 32122 11172 32124
rect 11196 32122 11252 32124
rect 10956 32070 10982 32122
rect 10982 32070 11012 32122
rect 11036 32070 11046 32122
rect 11046 32070 11092 32122
rect 11116 32070 11162 32122
rect 11162 32070 11172 32122
rect 11196 32070 11226 32122
rect 11226 32070 11252 32122
rect 10956 32068 11012 32070
rect 11036 32068 11092 32070
rect 11116 32068 11172 32070
rect 11196 32068 11252 32070
rect 11150 31864 11206 31920
rect 11242 31184 11298 31240
rect 10956 31034 11012 31036
rect 11036 31034 11092 31036
rect 11116 31034 11172 31036
rect 11196 31034 11252 31036
rect 10956 30982 10982 31034
rect 10982 30982 11012 31034
rect 11036 30982 11046 31034
rect 11046 30982 11092 31034
rect 11116 30982 11162 31034
rect 11162 30982 11172 31034
rect 11196 30982 11226 31034
rect 11226 30982 11252 31034
rect 10956 30980 11012 30982
rect 11036 30980 11092 30982
rect 11116 30980 11172 30982
rect 11196 30980 11252 30982
rect 10966 30812 10968 30832
rect 10968 30812 11020 30832
rect 11020 30812 11022 30832
rect 10966 30776 11022 30812
rect 10956 29946 11012 29948
rect 11036 29946 11092 29948
rect 11116 29946 11172 29948
rect 11196 29946 11252 29948
rect 10956 29894 10982 29946
rect 10982 29894 11012 29946
rect 11036 29894 11046 29946
rect 11046 29894 11092 29946
rect 11116 29894 11162 29946
rect 11162 29894 11172 29946
rect 11196 29894 11226 29946
rect 11226 29894 11252 29946
rect 10956 29892 11012 29894
rect 11036 29892 11092 29894
rect 11116 29892 11172 29894
rect 11196 29892 11252 29894
rect 10874 29144 10930 29200
rect 10956 28858 11012 28860
rect 11036 28858 11092 28860
rect 11116 28858 11172 28860
rect 11196 28858 11252 28860
rect 10956 28806 10982 28858
rect 10982 28806 11012 28858
rect 11036 28806 11046 28858
rect 11046 28806 11092 28858
rect 11116 28806 11162 28858
rect 11162 28806 11172 28858
rect 11196 28806 11226 28858
rect 11226 28806 11252 28858
rect 10956 28804 11012 28806
rect 11036 28804 11092 28806
rect 11116 28804 11172 28806
rect 11196 28804 11252 28806
rect 10874 28056 10930 28112
rect 10874 27920 10930 27976
rect 10956 27770 11012 27772
rect 11036 27770 11092 27772
rect 11116 27770 11172 27772
rect 11196 27770 11252 27772
rect 10956 27718 10982 27770
rect 10982 27718 11012 27770
rect 11036 27718 11046 27770
rect 11046 27718 11092 27770
rect 11116 27718 11162 27770
rect 11162 27718 11172 27770
rect 11196 27718 11226 27770
rect 11226 27718 11252 27770
rect 10956 27716 11012 27718
rect 11036 27716 11092 27718
rect 11116 27716 11172 27718
rect 11196 27716 11252 27718
rect 10956 26682 11012 26684
rect 11036 26682 11092 26684
rect 11116 26682 11172 26684
rect 11196 26682 11252 26684
rect 10956 26630 10982 26682
rect 10982 26630 11012 26682
rect 11036 26630 11046 26682
rect 11046 26630 11092 26682
rect 11116 26630 11162 26682
rect 11162 26630 11172 26682
rect 11196 26630 11226 26682
rect 11226 26630 11252 26682
rect 10956 26628 11012 26630
rect 11036 26628 11092 26630
rect 11116 26628 11172 26630
rect 11196 26628 11252 26630
rect 11242 26324 11244 26344
rect 11244 26324 11296 26344
rect 11296 26324 11298 26344
rect 11242 26288 11298 26324
rect 11150 25880 11206 25936
rect 11242 25744 11298 25800
rect 10956 25594 11012 25596
rect 11036 25594 11092 25596
rect 11116 25594 11172 25596
rect 11196 25594 11252 25596
rect 10956 25542 10982 25594
rect 10982 25542 11012 25594
rect 11036 25542 11046 25594
rect 11046 25542 11092 25594
rect 11116 25542 11162 25594
rect 11162 25542 11172 25594
rect 11196 25542 11226 25594
rect 11226 25542 11252 25594
rect 10956 25540 11012 25542
rect 11036 25540 11092 25542
rect 11116 25540 11172 25542
rect 11196 25540 11252 25542
rect 11978 49544 12034 49600
rect 12254 52556 12310 52592
rect 12254 52536 12256 52556
rect 12256 52536 12308 52556
rect 12308 52536 12310 52556
rect 12254 50632 12310 50688
rect 12622 52264 12678 52320
rect 12438 51448 12494 51504
rect 12070 48592 12126 48648
rect 11978 47504 12034 47560
rect 11702 41248 11758 41304
rect 11886 41112 11942 41168
rect 11518 31592 11574 31648
rect 11426 31456 11482 31512
rect 11702 34176 11758 34232
rect 11978 38528 12034 38584
rect 12714 51468 12770 51504
rect 12714 51448 12716 51468
rect 12716 51448 12768 51468
rect 12768 51448 12770 51468
rect 12622 49680 12678 49736
rect 13266 56108 13268 56128
rect 13268 56108 13320 56128
rect 13320 56108 13322 56128
rect 13266 56072 13322 56108
rect 13174 54576 13230 54632
rect 13174 54032 13230 54088
rect 13082 50632 13138 50688
rect 13082 50360 13138 50416
rect 12806 48492 12808 48512
rect 12808 48492 12860 48512
rect 12860 48492 12862 48512
rect 12806 48456 12862 48492
rect 13174 48592 13230 48648
rect 12898 48048 12954 48104
rect 13082 48048 13138 48104
rect 14370 73244 14372 73264
rect 14372 73244 14424 73264
rect 14424 73244 14426 73264
rect 14370 73208 14426 73244
rect 15198 68856 15254 68912
rect 15106 66136 15162 66192
rect 13726 56380 13728 56400
rect 13728 56380 13780 56400
rect 13780 56380 13782 56400
rect 13726 56344 13782 56380
rect 13542 56208 13598 56264
rect 13450 54068 13452 54088
rect 13452 54068 13504 54088
rect 13504 54068 13506 54088
rect 13450 54032 13506 54068
rect 14002 53896 14058 53952
rect 14002 52672 14058 52728
rect 13542 51992 13598 52048
rect 13818 50904 13874 50960
rect 14002 50768 14058 50824
rect 13542 49136 13598 49192
rect 13634 48864 13690 48920
rect 14002 47252 14058 47288
rect 14462 59336 14518 59392
rect 14370 59064 14426 59120
rect 14646 58520 14702 58576
rect 14830 58284 14832 58304
rect 14832 58284 14884 58304
rect 14884 58284 14886 58304
rect 14830 58248 14886 58284
rect 14646 57024 14702 57080
rect 14186 56344 14242 56400
rect 14186 56208 14242 56264
rect 14278 55800 14334 55856
rect 14278 52808 14334 52864
rect 14554 55392 14610 55448
rect 14462 53488 14518 53544
rect 14186 50380 14242 50416
rect 14186 50360 14188 50380
rect 14188 50360 14240 50380
rect 14240 50360 14242 50380
rect 14278 49136 14334 49192
rect 14002 47232 14004 47252
rect 14004 47232 14056 47252
rect 14056 47232 14058 47252
rect 12162 35808 12218 35864
rect 12070 34856 12126 34912
rect 11978 34312 12034 34368
rect 11702 33904 11758 33960
rect 11794 33768 11850 33824
rect 11702 31592 11758 31648
rect 11610 31048 11666 31104
rect 11518 30640 11574 30696
rect 11518 29688 11574 29744
rect 11518 29416 11574 29472
rect 12070 33632 12126 33688
rect 11978 32408 12034 32464
rect 11978 31864 12034 31920
rect 11518 28192 11574 28248
rect 11702 28056 11758 28112
rect 10956 24506 11012 24508
rect 11036 24506 11092 24508
rect 11116 24506 11172 24508
rect 11196 24506 11252 24508
rect 10956 24454 10982 24506
rect 10982 24454 11012 24506
rect 11036 24454 11046 24506
rect 11046 24454 11092 24506
rect 11116 24454 11162 24506
rect 11162 24454 11172 24506
rect 11196 24454 11226 24506
rect 11226 24454 11252 24506
rect 10956 24452 11012 24454
rect 11036 24452 11092 24454
rect 11116 24452 11172 24454
rect 11196 24452 11252 24454
rect 10874 24012 10876 24032
rect 10876 24012 10928 24032
rect 10928 24012 10930 24032
rect 10874 23976 10930 24012
rect 10782 21684 10838 21720
rect 10782 21664 10784 21684
rect 10784 21664 10836 21684
rect 10836 21664 10838 21684
rect 10956 23418 11012 23420
rect 11036 23418 11092 23420
rect 11116 23418 11172 23420
rect 11196 23418 11252 23420
rect 10956 23366 10982 23418
rect 10982 23366 11012 23418
rect 11036 23366 11046 23418
rect 11046 23366 11092 23418
rect 11116 23366 11162 23418
rect 11162 23366 11172 23418
rect 11196 23366 11226 23418
rect 11226 23366 11252 23418
rect 10956 23364 11012 23366
rect 11036 23364 11092 23366
rect 11116 23364 11172 23366
rect 11196 23364 11252 23366
rect 11426 23568 11482 23624
rect 11334 22616 11390 22672
rect 10956 22330 11012 22332
rect 11036 22330 11092 22332
rect 11116 22330 11172 22332
rect 11196 22330 11252 22332
rect 10956 22278 10982 22330
rect 10982 22278 11012 22330
rect 11036 22278 11046 22330
rect 11046 22278 11092 22330
rect 11116 22278 11162 22330
rect 11162 22278 11172 22330
rect 11196 22278 11226 22330
rect 11226 22278 11252 22330
rect 10956 22276 11012 22278
rect 11036 22276 11092 22278
rect 11116 22276 11172 22278
rect 11196 22276 11252 22278
rect 10956 21242 11012 21244
rect 11036 21242 11092 21244
rect 11116 21242 11172 21244
rect 11196 21242 11252 21244
rect 10956 21190 10982 21242
rect 10982 21190 11012 21242
rect 11036 21190 11046 21242
rect 11046 21190 11092 21242
rect 11116 21190 11162 21242
rect 11162 21190 11172 21242
rect 11196 21190 11226 21242
rect 11226 21190 11252 21242
rect 10956 21188 11012 21190
rect 11036 21188 11092 21190
rect 11116 21188 11172 21190
rect 11196 21188 11252 21190
rect 10782 20712 10838 20768
rect 10506 18808 10562 18864
rect 10506 17720 10562 17776
rect 11058 20576 11114 20632
rect 10956 20154 11012 20156
rect 11036 20154 11092 20156
rect 11116 20154 11172 20156
rect 11196 20154 11252 20156
rect 10956 20102 10982 20154
rect 10982 20102 11012 20154
rect 11036 20102 11046 20154
rect 11046 20102 11092 20154
rect 11116 20102 11162 20154
rect 11162 20102 11172 20154
rect 11196 20102 11226 20154
rect 11226 20102 11252 20154
rect 10956 20100 11012 20102
rect 11036 20100 11092 20102
rect 11116 20100 11172 20102
rect 11196 20100 11252 20102
rect 11150 19760 11206 19816
rect 10956 19066 11012 19068
rect 11036 19066 11092 19068
rect 11116 19066 11172 19068
rect 11196 19066 11252 19068
rect 10956 19014 10982 19066
rect 10982 19014 11012 19066
rect 11036 19014 11046 19066
rect 11046 19014 11092 19066
rect 11116 19014 11162 19066
rect 11162 19014 11172 19066
rect 11196 19014 11226 19066
rect 11226 19014 11252 19066
rect 10956 19012 11012 19014
rect 11036 19012 11092 19014
rect 11116 19012 11172 19014
rect 11196 19012 11252 19014
rect 10782 18128 10838 18184
rect 13082 40876 13084 40896
rect 13084 40876 13136 40896
rect 13136 40876 13138 40896
rect 13082 40840 13138 40876
rect 12530 38120 12586 38176
rect 12990 38528 13046 38584
rect 12438 35556 12494 35592
rect 12438 35536 12440 35556
rect 12440 35536 12492 35556
rect 12492 35536 12494 35556
rect 12530 35164 12532 35184
rect 12532 35164 12584 35184
rect 12584 35164 12586 35184
rect 12530 35128 12586 35164
rect 12346 33224 12402 33280
rect 12162 32000 12218 32056
rect 12530 33224 12586 33280
rect 12254 31864 12310 31920
rect 12254 31084 12256 31104
rect 12256 31084 12308 31104
rect 12308 31084 12310 31104
rect 12254 31048 12310 31084
rect 13266 42880 13322 42936
rect 13174 37868 13230 37904
rect 13174 37848 13176 37868
rect 13176 37848 13228 37868
rect 13228 37848 13230 37868
rect 12714 35944 12770 36000
rect 12806 34992 12862 35048
rect 13082 37712 13138 37768
rect 12990 36760 13046 36816
rect 12990 35128 13046 35184
rect 12898 34448 12954 34504
rect 12898 33924 12954 33960
rect 12898 33904 12900 33924
rect 12900 33904 12952 33924
rect 12952 33904 12954 33924
rect 13082 34312 13138 34368
rect 13082 34040 13138 34096
rect 12714 33088 12770 33144
rect 13082 33224 13138 33280
rect 13082 32272 13138 32328
rect 12806 31764 12808 31784
rect 12808 31764 12860 31784
rect 12860 31764 12862 31784
rect 12806 31728 12862 31764
rect 12530 31184 12586 31240
rect 12346 29960 12402 30016
rect 12806 31320 12862 31376
rect 12254 27784 12310 27840
rect 12622 28464 12678 28520
rect 12162 26016 12218 26072
rect 11794 24520 11850 24576
rect 11702 20984 11758 21040
rect 11334 18264 11390 18320
rect 10956 17978 11012 17980
rect 11036 17978 11092 17980
rect 11116 17978 11172 17980
rect 11196 17978 11252 17980
rect 10956 17926 10982 17978
rect 10982 17926 11012 17978
rect 11036 17926 11046 17978
rect 11046 17926 11092 17978
rect 11116 17926 11162 17978
rect 11162 17926 11172 17978
rect 11196 17926 11226 17978
rect 11226 17926 11252 17978
rect 10956 17924 11012 17926
rect 11036 17924 11092 17926
rect 11116 17924 11172 17926
rect 11196 17924 11252 17926
rect 11242 17040 11298 17096
rect 10956 16890 11012 16892
rect 11036 16890 11092 16892
rect 11116 16890 11172 16892
rect 11196 16890 11252 16892
rect 10956 16838 10982 16890
rect 10982 16838 11012 16890
rect 11036 16838 11046 16890
rect 11046 16838 11092 16890
rect 11116 16838 11162 16890
rect 11162 16838 11172 16890
rect 11196 16838 11226 16890
rect 11226 16838 11252 16890
rect 10956 16836 11012 16838
rect 11036 16836 11092 16838
rect 11116 16836 11172 16838
rect 11196 16836 11252 16838
rect 11426 17176 11482 17232
rect 10322 15272 10378 15328
rect 9954 14320 10010 14376
rect 9678 9036 9734 9072
rect 9678 9016 9680 9036
rect 9680 9016 9732 9036
rect 9732 9016 9734 9036
rect 10598 16088 10654 16144
rect 10956 15802 11012 15804
rect 11036 15802 11092 15804
rect 11116 15802 11172 15804
rect 11196 15802 11252 15804
rect 10956 15750 10982 15802
rect 10982 15750 11012 15802
rect 11036 15750 11046 15802
rect 11046 15750 11092 15802
rect 11116 15750 11162 15802
rect 11162 15750 11172 15802
rect 11196 15750 11226 15802
rect 11226 15750 11252 15802
rect 10956 15748 11012 15750
rect 11036 15748 11092 15750
rect 11116 15748 11172 15750
rect 11196 15748 11252 15750
rect 10956 14714 11012 14716
rect 11036 14714 11092 14716
rect 11116 14714 11172 14716
rect 11196 14714 11252 14716
rect 10956 14662 10982 14714
rect 10982 14662 11012 14714
rect 11036 14662 11046 14714
rect 11046 14662 11092 14714
rect 11116 14662 11162 14714
rect 11162 14662 11172 14714
rect 11196 14662 11226 14714
rect 11226 14662 11252 14714
rect 10956 14660 11012 14662
rect 11036 14660 11092 14662
rect 11116 14660 11172 14662
rect 11196 14660 11252 14662
rect 10956 13626 11012 13628
rect 11036 13626 11092 13628
rect 11116 13626 11172 13628
rect 11196 13626 11252 13628
rect 10956 13574 10982 13626
rect 10982 13574 11012 13626
rect 11036 13574 11046 13626
rect 11046 13574 11092 13626
rect 11116 13574 11162 13626
rect 11162 13574 11172 13626
rect 11196 13574 11226 13626
rect 11226 13574 11252 13626
rect 10956 13572 11012 13574
rect 11036 13572 11092 13574
rect 11116 13572 11172 13574
rect 11196 13572 11252 13574
rect 10506 9696 10562 9752
rect 8298 7520 8354 7576
rect 6274 7384 6330 7440
rect 7746 7384 7802 7440
rect 5956 6554 6012 6556
rect 6036 6554 6092 6556
rect 6116 6554 6172 6556
rect 6196 6554 6252 6556
rect 5956 6502 5982 6554
rect 5982 6502 6012 6554
rect 6036 6502 6046 6554
rect 6046 6502 6092 6554
rect 6116 6502 6162 6554
rect 6162 6502 6172 6554
rect 6196 6502 6226 6554
rect 6226 6502 6252 6554
rect 5956 6500 6012 6502
rect 6036 6500 6092 6502
rect 6116 6500 6172 6502
rect 6196 6500 6252 6502
rect 5956 5466 6012 5468
rect 6036 5466 6092 5468
rect 6116 5466 6172 5468
rect 6196 5466 6252 5468
rect 5956 5414 5982 5466
rect 5982 5414 6012 5466
rect 6036 5414 6046 5466
rect 6046 5414 6092 5466
rect 6116 5414 6162 5466
rect 6162 5414 6172 5466
rect 6196 5414 6226 5466
rect 6226 5414 6252 5466
rect 5956 5412 6012 5414
rect 6036 5412 6092 5414
rect 6116 5412 6172 5414
rect 6196 5412 6252 5414
rect 5956 4378 6012 4380
rect 6036 4378 6092 4380
rect 6116 4378 6172 4380
rect 6196 4378 6252 4380
rect 5956 4326 5982 4378
rect 5982 4326 6012 4378
rect 6036 4326 6046 4378
rect 6046 4326 6092 4378
rect 6116 4326 6162 4378
rect 6162 4326 6172 4378
rect 6196 4326 6226 4378
rect 6226 4326 6252 4378
rect 5956 4324 6012 4326
rect 6036 4324 6092 4326
rect 6116 4324 6172 4326
rect 6196 4324 6252 4326
rect 5078 3576 5134 3632
rect 5956 3290 6012 3292
rect 6036 3290 6092 3292
rect 6116 3290 6172 3292
rect 6196 3290 6252 3292
rect 5956 3238 5982 3290
rect 5982 3238 6012 3290
rect 6036 3238 6046 3290
rect 6046 3238 6092 3290
rect 6116 3238 6162 3290
rect 6162 3238 6172 3290
rect 6196 3238 6226 3290
rect 6226 3238 6252 3290
rect 5956 3236 6012 3238
rect 6036 3236 6092 3238
rect 6116 3236 6172 3238
rect 6196 3236 6252 3238
rect 5956 2202 6012 2204
rect 6036 2202 6092 2204
rect 6116 2202 6172 2204
rect 6196 2202 6252 2204
rect 5956 2150 5982 2202
rect 5982 2150 6012 2202
rect 6036 2150 6046 2202
rect 6046 2150 6092 2202
rect 6116 2150 6162 2202
rect 6162 2150 6172 2202
rect 6196 2150 6226 2202
rect 6226 2150 6252 2202
rect 5956 2148 6012 2150
rect 6036 2148 6092 2150
rect 6116 2148 6172 2150
rect 6196 2148 6252 2150
rect 6918 3304 6974 3360
rect 7378 3168 7434 3224
rect 11426 15408 11482 15464
rect 10956 12538 11012 12540
rect 11036 12538 11092 12540
rect 11116 12538 11172 12540
rect 11196 12538 11252 12540
rect 10956 12486 10982 12538
rect 10982 12486 11012 12538
rect 11036 12486 11046 12538
rect 11046 12486 11092 12538
rect 11116 12486 11162 12538
rect 11162 12486 11172 12538
rect 11196 12486 11226 12538
rect 11226 12486 11252 12538
rect 10956 12484 11012 12486
rect 11036 12484 11092 12486
rect 11116 12484 11172 12486
rect 11196 12484 11252 12486
rect 12070 23976 12126 24032
rect 11978 23160 12034 23216
rect 12070 22888 12126 22944
rect 12714 27784 12770 27840
rect 12622 27240 12678 27296
rect 12898 30504 12954 30560
rect 12898 30232 12954 30288
rect 12898 29552 12954 29608
rect 12806 26968 12862 27024
rect 12530 26016 12586 26072
rect 12438 24676 12494 24712
rect 12438 24656 12440 24676
rect 12440 24656 12492 24676
rect 12492 24656 12494 24676
rect 12254 22480 12310 22536
rect 12438 22636 12494 22672
rect 12438 22616 12440 22636
rect 12440 22616 12492 22636
rect 12492 22616 12494 22636
rect 12346 22208 12402 22264
rect 12254 20868 12310 20904
rect 12254 20848 12256 20868
rect 12256 20848 12308 20868
rect 12308 20848 12310 20868
rect 12438 17040 12494 17096
rect 12714 18128 12770 18184
rect 12530 15952 12586 16008
rect 12254 15544 12310 15600
rect 12438 15544 12494 15600
rect 10956 11450 11012 11452
rect 11036 11450 11092 11452
rect 11116 11450 11172 11452
rect 11196 11450 11252 11452
rect 10956 11398 10982 11450
rect 10982 11398 11012 11450
rect 11036 11398 11046 11450
rect 11046 11398 11092 11450
rect 11116 11398 11162 11450
rect 11162 11398 11172 11450
rect 11196 11398 11226 11450
rect 11226 11398 11252 11450
rect 10956 11396 11012 11398
rect 11036 11396 11092 11398
rect 11116 11396 11172 11398
rect 11196 11396 11252 11398
rect 10956 10362 11012 10364
rect 11036 10362 11092 10364
rect 11116 10362 11172 10364
rect 11196 10362 11252 10364
rect 10956 10310 10982 10362
rect 10982 10310 11012 10362
rect 11036 10310 11046 10362
rect 11046 10310 11092 10362
rect 11116 10310 11162 10362
rect 11162 10310 11172 10362
rect 11196 10310 11226 10362
rect 11226 10310 11252 10362
rect 10956 10308 11012 10310
rect 11036 10308 11092 10310
rect 11116 10308 11172 10310
rect 11196 10308 11252 10310
rect 10956 9274 11012 9276
rect 11036 9274 11092 9276
rect 11116 9274 11172 9276
rect 11196 9274 11252 9276
rect 10956 9222 10982 9274
rect 10982 9222 11012 9274
rect 11036 9222 11046 9274
rect 11046 9222 11092 9274
rect 11116 9222 11162 9274
rect 11162 9222 11172 9274
rect 11196 9222 11226 9274
rect 11226 9222 11252 9274
rect 10956 9220 11012 9222
rect 11036 9220 11092 9222
rect 11116 9220 11172 9222
rect 11196 9220 11252 9222
rect 10956 8186 11012 8188
rect 11036 8186 11092 8188
rect 11116 8186 11172 8188
rect 11196 8186 11252 8188
rect 10956 8134 10982 8186
rect 10982 8134 11012 8186
rect 11036 8134 11046 8186
rect 11046 8134 11092 8186
rect 11116 8134 11162 8186
rect 11162 8134 11172 8186
rect 11196 8134 11226 8186
rect 11226 8134 11252 8186
rect 10956 8132 11012 8134
rect 11036 8132 11092 8134
rect 11116 8132 11172 8134
rect 11196 8132 11252 8134
rect 9862 7928 9918 7984
rect 9034 6976 9090 7032
rect 9218 5480 9274 5536
rect 10956 7098 11012 7100
rect 11036 7098 11092 7100
rect 11116 7098 11172 7100
rect 11196 7098 11252 7100
rect 10956 7046 10982 7098
rect 10982 7046 11012 7098
rect 11036 7046 11046 7098
rect 11046 7046 11092 7098
rect 11116 7046 11162 7098
rect 11162 7046 11172 7098
rect 11196 7046 11226 7098
rect 11226 7046 11252 7098
rect 10956 7044 11012 7046
rect 11036 7044 11092 7046
rect 11116 7044 11172 7046
rect 11196 7044 11252 7046
rect 10956 6010 11012 6012
rect 11036 6010 11092 6012
rect 11116 6010 11172 6012
rect 11196 6010 11252 6012
rect 10956 5958 10982 6010
rect 10982 5958 11012 6010
rect 11036 5958 11046 6010
rect 11046 5958 11092 6010
rect 11116 5958 11162 6010
rect 11162 5958 11172 6010
rect 11196 5958 11226 6010
rect 11226 5958 11252 6010
rect 10956 5956 11012 5958
rect 11036 5956 11092 5958
rect 11116 5956 11172 5958
rect 11196 5956 11252 5958
rect 10956 4922 11012 4924
rect 11036 4922 11092 4924
rect 11116 4922 11172 4924
rect 11196 4922 11252 4924
rect 10956 4870 10982 4922
rect 10982 4870 11012 4922
rect 11036 4870 11046 4922
rect 11046 4870 11092 4922
rect 11116 4870 11162 4922
rect 11162 4870 11172 4922
rect 11196 4870 11226 4922
rect 11226 4870 11252 4922
rect 10956 4868 11012 4870
rect 11036 4868 11092 4870
rect 11116 4868 11172 4870
rect 11196 4868 11252 4870
rect 10956 3834 11012 3836
rect 11036 3834 11092 3836
rect 11116 3834 11172 3836
rect 11196 3834 11252 3836
rect 10956 3782 10982 3834
rect 10982 3782 11012 3834
rect 11036 3782 11046 3834
rect 11046 3782 11092 3834
rect 11116 3782 11162 3834
rect 11162 3782 11172 3834
rect 11196 3782 11226 3834
rect 11226 3782 11252 3834
rect 10956 3780 11012 3782
rect 11036 3780 11092 3782
rect 11116 3780 11172 3782
rect 11196 3780 11252 3782
rect 11610 10784 11666 10840
rect 10956 2746 11012 2748
rect 11036 2746 11092 2748
rect 11116 2746 11172 2748
rect 11196 2746 11252 2748
rect 10956 2694 10982 2746
rect 10982 2694 11012 2746
rect 11036 2694 11046 2746
rect 11046 2694 11092 2746
rect 11116 2694 11162 2746
rect 11162 2694 11172 2746
rect 11196 2694 11226 2746
rect 11226 2694 11252 2746
rect 10956 2692 11012 2694
rect 11036 2692 11092 2694
rect 11116 2692 11172 2694
rect 11196 2692 11252 2694
rect 11978 13232 12034 13288
rect 12622 15000 12678 15056
rect 14462 50904 14518 50960
rect 15106 55256 15162 55312
rect 14922 54848 14978 54904
rect 15956 77274 16012 77276
rect 16036 77274 16092 77276
rect 16116 77274 16172 77276
rect 16196 77274 16252 77276
rect 15956 77222 15982 77274
rect 15982 77222 16012 77274
rect 16036 77222 16046 77274
rect 16046 77222 16092 77274
rect 16116 77222 16162 77274
rect 16162 77222 16172 77274
rect 16196 77222 16226 77274
rect 16226 77222 16252 77274
rect 15956 77220 16012 77222
rect 16036 77220 16092 77222
rect 16116 77220 16172 77222
rect 16196 77220 16252 77222
rect 15956 76186 16012 76188
rect 16036 76186 16092 76188
rect 16116 76186 16172 76188
rect 16196 76186 16252 76188
rect 15956 76134 15982 76186
rect 15982 76134 16012 76186
rect 16036 76134 16046 76186
rect 16046 76134 16092 76186
rect 16116 76134 16162 76186
rect 16162 76134 16172 76186
rect 16196 76134 16226 76186
rect 16226 76134 16252 76186
rect 15956 76132 16012 76134
rect 16036 76132 16092 76134
rect 16116 76132 16172 76134
rect 16196 76132 16252 76134
rect 16578 75792 16634 75848
rect 15956 75098 16012 75100
rect 16036 75098 16092 75100
rect 16116 75098 16172 75100
rect 16196 75098 16252 75100
rect 15956 75046 15982 75098
rect 15982 75046 16012 75098
rect 16036 75046 16046 75098
rect 16046 75046 16092 75098
rect 16116 75046 16162 75098
rect 16162 75046 16172 75098
rect 16196 75046 16226 75098
rect 16226 75046 16252 75098
rect 15956 75044 16012 75046
rect 16036 75044 16092 75046
rect 16116 75044 16172 75046
rect 16196 75044 16252 75046
rect 18602 75248 18658 75304
rect 15956 74010 16012 74012
rect 16036 74010 16092 74012
rect 16116 74010 16172 74012
rect 16196 74010 16252 74012
rect 15956 73958 15982 74010
rect 15982 73958 16012 74010
rect 16036 73958 16046 74010
rect 16046 73958 16092 74010
rect 16116 73958 16162 74010
rect 16162 73958 16172 74010
rect 16196 73958 16226 74010
rect 16226 73958 16252 74010
rect 15956 73956 16012 73958
rect 16036 73956 16092 73958
rect 16116 73956 16172 73958
rect 16196 73956 16252 73958
rect 15956 72922 16012 72924
rect 16036 72922 16092 72924
rect 16116 72922 16172 72924
rect 16196 72922 16252 72924
rect 15956 72870 15982 72922
rect 15982 72870 16012 72922
rect 16036 72870 16046 72922
rect 16046 72870 16092 72922
rect 16116 72870 16162 72922
rect 16162 72870 16172 72922
rect 16196 72870 16226 72922
rect 16226 72870 16252 72922
rect 15956 72868 16012 72870
rect 16036 72868 16092 72870
rect 16116 72868 16172 72870
rect 16196 72868 16252 72870
rect 15956 71834 16012 71836
rect 16036 71834 16092 71836
rect 16116 71834 16172 71836
rect 16196 71834 16252 71836
rect 15956 71782 15982 71834
rect 15982 71782 16012 71834
rect 16036 71782 16046 71834
rect 16046 71782 16092 71834
rect 16116 71782 16162 71834
rect 16162 71782 16172 71834
rect 16196 71782 16226 71834
rect 16226 71782 16252 71834
rect 15956 71780 16012 71782
rect 16036 71780 16092 71782
rect 16116 71780 16172 71782
rect 16196 71780 16252 71782
rect 15956 70746 16012 70748
rect 16036 70746 16092 70748
rect 16116 70746 16172 70748
rect 16196 70746 16252 70748
rect 15956 70694 15982 70746
rect 15982 70694 16012 70746
rect 16036 70694 16046 70746
rect 16046 70694 16092 70746
rect 16116 70694 16162 70746
rect 16162 70694 16172 70746
rect 16196 70694 16226 70746
rect 16226 70694 16252 70746
rect 15956 70692 16012 70694
rect 16036 70692 16092 70694
rect 16116 70692 16172 70694
rect 16196 70692 16252 70694
rect 15956 69658 16012 69660
rect 16036 69658 16092 69660
rect 16116 69658 16172 69660
rect 16196 69658 16252 69660
rect 15956 69606 15982 69658
rect 15982 69606 16012 69658
rect 16036 69606 16046 69658
rect 16046 69606 16092 69658
rect 16116 69606 16162 69658
rect 16162 69606 16172 69658
rect 16196 69606 16226 69658
rect 16226 69606 16252 69658
rect 15956 69604 16012 69606
rect 16036 69604 16092 69606
rect 16116 69604 16172 69606
rect 16196 69604 16252 69606
rect 15956 68570 16012 68572
rect 16036 68570 16092 68572
rect 16116 68570 16172 68572
rect 16196 68570 16252 68572
rect 15956 68518 15982 68570
rect 15982 68518 16012 68570
rect 16036 68518 16046 68570
rect 16046 68518 16092 68570
rect 16116 68518 16162 68570
rect 16162 68518 16172 68570
rect 16196 68518 16226 68570
rect 16226 68518 16252 68570
rect 15956 68516 16012 68518
rect 16036 68516 16092 68518
rect 16116 68516 16172 68518
rect 16196 68516 16252 68518
rect 15382 67496 15438 67552
rect 15956 67482 16012 67484
rect 16036 67482 16092 67484
rect 16116 67482 16172 67484
rect 16196 67482 16252 67484
rect 15956 67430 15982 67482
rect 15982 67430 16012 67482
rect 16036 67430 16046 67482
rect 16046 67430 16092 67482
rect 16116 67430 16162 67482
rect 16162 67430 16172 67482
rect 16196 67430 16226 67482
rect 16226 67430 16252 67482
rect 15956 67428 16012 67430
rect 16036 67428 16092 67430
rect 16116 67428 16172 67430
rect 16196 67428 16252 67430
rect 15956 66394 16012 66396
rect 16036 66394 16092 66396
rect 16116 66394 16172 66396
rect 16196 66394 16252 66396
rect 15956 66342 15982 66394
rect 15982 66342 16012 66394
rect 16036 66342 16046 66394
rect 16046 66342 16092 66394
rect 16116 66342 16162 66394
rect 16162 66342 16172 66394
rect 16196 66342 16226 66394
rect 16226 66342 16252 66394
rect 15956 66340 16012 66342
rect 16036 66340 16092 66342
rect 16116 66340 16172 66342
rect 16196 66340 16252 66342
rect 15474 64912 15530 64968
rect 15956 65306 16012 65308
rect 16036 65306 16092 65308
rect 16116 65306 16172 65308
rect 16196 65306 16252 65308
rect 15956 65254 15982 65306
rect 15982 65254 16012 65306
rect 16036 65254 16046 65306
rect 16046 65254 16092 65306
rect 16116 65254 16162 65306
rect 16162 65254 16172 65306
rect 16196 65254 16226 65306
rect 16226 65254 16252 65306
rect 15956 65252 16012 65254
rect 16036 65252 16092 65254
rect 16116 65252 16172 65254
rect 16196 65252 16252 65254
rect 15382 57876 15384 57896
rect 15384 57876 15436 57896
rect 15436 57876 15438 57896
rect 15382 57840 15438 57876
rect 14738 53624 14794 53680
rect 14646 53352 14702 53408
rect 14830 52944 14886 53000
rect 15198 54052 15254 54088
rect 15198 54032 15200 54052
rect 15200 54032 15252 54052
rect 15252 54032 15254 54052
rect 15106 53388 15108 53408
rect 15108 53388 15160 53408
rect 15160 53388 15162 53408
rect 15106 53352 15162 53388
rect 15014 52672 15070 52728
rect 15198 52536 15254 52592
rect 15290 52012 15346 52048
rect 15290 51992 15292 52012
rect 15292 51992 15344 52012
rect 15344 51992 15346 52012
rect 15014 51040 15070 51096
rect 15198 51040 15254 51096
rect 14738 47368 14794 47424
rect 14002 43968 14058 44024
rect 14646 42744 14702 42800
rect 15290 49716 15292 49736
rect 15292 49716 15344 49736
rect 15344 49716 15346 49736
rect 15290 49680 15346 49716
rect 15290 49136 15346 49192
rect 15014 47096 15070 47152
rect 15956 64218 16012 64220
rect 16036 64218 16092 64220
rect 16116 64218 16172 64220
rect 16196 64218 16252 64220
rect 15956 64166 15982 64218
rect 15982 64166 16012 64218
rect 16036 64166 16046 64218
rect 16046 64166 16092 64218
rect 16116 64166 16162 64218
rect 16162 64166 16172 64218
rect 16196 64166 16226 64218
rect 16226 64166 16252 64218
rect 15956 64164 16012 64166
rect 16036 64164 16092 64166
rect 16116 64164 16172 64166
rect 16196 64164 16252 64166
rect 15956 63130 16012 63132
rect 16036 63130 16092 63132
rect 16116 63130 16172 63132
rect 16196 63130 16252 63132
rect 15956 63078 15982 63130
rect 15982 63078 16012 63130
rect 16036 63078 16046 63130
rect 16046 63078 16092 63130
rect 16116 63078 16162 63130
rect 16162 63078 16172 63130
rect 16196 63078 16226 63130
rect 16226 63078 16252 63130
rect 15956 63076 16012 63078
rect 16036 63076 16092 63078
rect 16116 63076 16172 63078
rect 16196 63076 16252 63078
rect 15956 62042 16012 62044
rect 16036 62042 16092 62044
rect 16116 62042 16172 62044
rect 16196 62042 16252 62044
rect 15956 61990 15982 62042
rect 15982 61990 16012 62042
rect 16036 61990 16046 62042
rect 16046 61990 16092 62042
rect 16116 61990 16162 62042
rect 16162 61990 16172 62042
rect 16196 61990 16226 62042
rect 16226 61990 16252 62042
rect 15956 61988 16012 61990
rect 16036 61988 16092 61990
rect 16116 61988 16172 61990
rect 16196 61988 16252 61990
rect 15474 56480 15530 56536
rect 15566 50632 15622 50688
rect 15474 48864 15530 48920
rect 15474 48320 15530 48376
rect 15750 56616 15806 56672
rect 15750 56480 15806 56536
rect 15956 60954 16012 60956
rect 16036 60954 16092 60956
rect 16116 60954 16172 60956
rect 16196 60954 16252 60956
rect 15956 60902 15982 60954
rect 15982 60902 16012 60954
rect 16036 60902 16046 60954
rect 16046 60902 16092 60954
rect 16116 60902 16162 60954
rect 16162 60902 16172 60954
rect 16196 60902 16226 60954
rect 16226 60902 16252 60954
rect 15956 60900 16012 60902
rect 16036 60900 16092 60902
rect 16116 60900 16172 60902
rect 16196 60900 16252 60902
rect 15956 59866 16012 59868
rect 16036 59866 16092 59868
rect 16116 59866 16172 59868
rect 16196 59866 16252 59868
rect 15956 59814 15982 59866
rect 15982 59814 16012 59866
rect 16036 59814 16046 59866
rect 16046 59814 16092 59866
rect 16116 59814 16162 59866
rect 16162 59814 16172 59866
rect 16196 59814 16226 59866
rect 16226 59814 16252 59866
rect 15956 59812 16012 59814
rect 16036 59812 16092 59814
rect 16116 59812 16172 59814
rect 16196 59812 16252 59814
rect 16210 59508 16212 59528
rect 16212 59508 16264 59528
rect 16264 59508 16266 59528
rect 16210 59472 16266 59508
rect 15956 58778 16012 58780
rect 16036 58778 16092 58780
rect 16116 58778 16172 58780
rect 16196 58778 16252 58780
rect 15956 58726 15982 58778
rect 15982 58726 16012 58778
rect 16036 58726 16046 58778
rect 16046 58726 16092 58778
rect 16116 58726 16162 58778
rect 16162 58726 16172 58778
rect 16196 58726 16226 58778
rect 16226 58726 16252 58778
rect 15956 58724 16012 58726
rect 16036 58724 16092 58726
rect 16116 58724 16172 58726
rect 16196 58724 16252 58726
rect 16210 58520 16266 58576
rect 15956 57690 16012 57692
rect 16036 57690 16092 57692
rect 16116 57690 16172 57692
rect 16196 57690 16252 57692
rect 15956 57638 15982 57690
rect 15982 57638 16012 57690
rect 16036 57638 16046 57690
rect 16046 57638 16092 57690
rect 16116 57638 16162 57690
rect 16162 57638 16172 57690
rect 16196 57638 16226 57690
rect 16226 57638 16252 57690
rect 15956 57636 16012 57638
rect 16036 57636 16092 57638
rect 16116 57636 16172 57638
rect 16196 57636 16252 57638
rect 15956 56602 16012 56604
rect 16036 56602 16092 56604
rect 16116 56602 16172 56604
rect 16196 56602 16252 56604
rect 15956 56550 15982 56602
rect 15982 56550 16012 56602
rect 16036 56550 16046 56602
rect 16046 56550 16092 56602
rect 16116 56550 16162 56602
rect 16162 56550 16172 56602
rect 16196 56550 16226 56602
rect 16226 56550 16252 56602
rect 15956 56548 16012 56550
rect 16036 56548 16092 56550
rect 16116 56548 16172 56550
rect 16196 56548 16252 56550
rect 15956 55514 16012 55516
rect 16036 55514 16092 55516
rect 16116 55514 16172 55516
rect 16196 55514 16252 55516
rect 15956 55462 15982 55514
rect 15982 55462 16012 55514
rect 16036 55462 16046 55514
rect 16046 55462 16092 55514
rect 16116 55462 16162 55514
rect 16162 55462 16172 55514
rect 16196 55462 16226 55514
rect 16226 55462 16252 55514
rect 15956 55460 16012 55462
rect 16036 55460 16092 55462
rect 16116 55460 16172 55462
rect 16196 55460 16252 55462
rect 15956 54426 16012 54428
rect 16036 54426 16092 54428
rect 16116 54426 16172 54428
rect 16196 54426 16252 54428
rect 15956 54374 15982 54426
rect 15982 54374 16012 54426
rect 16036 54374 16046 54426
rect 16046 54374 16092 54426
rect 16116 54374 16162 54426
rect 16162 54374 16172 54426
rect 16196 54374 16226 54426
rect 16226 54374 16252 54426
rect 15956 54372 16012 54374
rect 16036 54372 16092 54374
rect 16116 54372 16172 54374
rect 16196 54372 16252 54374
rect 16026 54204 16028 54224
rect 16028 54204 16080 54224
rect 16080 54204 16082 54224
rect 16026 54168 16082 54204
rect 15956 53338 16012 53340
rect 16036 53338 16092 53340
rect 16116 53338 16172 53340
rect 16196 53338 16252 53340
rect 15956 53286 15982 53338
rect 15982 53286 16012 53338
rect 16036 53286 16046 53338
rect 16046 53286 16092 53338
rect 16116 53286 16162 53338
rect 16162 53286 16172 53338
rect 16196 53286 16226 53338
rect 16226 53286 16252 53338
rect 15956 53284 16012 53286
rect 16036 53284 16092 53286
rect 16116 53284 16172 53286
rect 16196 53284 16252 53286
rect 15956 52250 16012 52252
rect 16036 52250 16092 52252
rect 16116 52250 16172 52252
rect 16196 52250 16252 52252
rect 15956 52198 15982 52250
rect 15982 52198 16012 52250
rect 16036 52198 16046 52250
rect 16046 52198 16092 52250
rect 16116 52198 16162 52250
rect 16162 52198 16172 52250
rect 16196 52198 16226 52250
rect 16226 52198 16252 52250
rect 15956 52196 16012 52198
rect 16036 52196 16092 52198
rect 16116 52196 16172 52198
rect 16196 52196 16252 52198
rect 15842 51312 15898 51368
rect 15750 49544 15806 49600
rect 15566 46316 15568 46336
rect 15568 46316 15620 46336
rect 15620 46316 15622 46336
rect 15566 46280 15622 46316
rect 15658 44784 15714 44840
rect 14830 42200 14886 42256
rect 15106 42084 15162 42120
rect 15106 42064 15108 42084
rect 15108 42064 15160 42084
rect 15160 42064 15162 42084
rect 14002 41792 14058 41848
rect 15106 41112 15162 41168
rect 13450 39888 13506 39944
rect 13634 39788 13636 39808
rect 13636 39788 13688 39808
rect 13688 39788 13690 39808
rect 13634 39752 13690 39788
rect 13542 38836 13544 38856
rect 13544 38836 13596 38856
rect 13596 38836 13598 38856
rect 13542 38800 13598 38836
rect 13726 38392 13782 38448
rect 13266 36896 13322 36952
rect 13542 37712 13598 37768
rect 13450 37168 13506 37224
rect 13358 36352 13414 36408
rect 13266 34604 13322 34640
rect 13266 34584 13268 34604
rect 13268 34584 13320 34604
rect 13320 34584 13322 34604
rect 13266 32000 13322 32056
rect 13082 31592 13138 31648
rect 13174 30796 13230 30832
rect 13174 30776 13176 30796
rect 13176 30776 13228 30796
rect 13228 30776 13230 30796
rect 13082 30504 13138 30560
rect 13358 30640 13414 30696
rect 13818 36216 13874 36272
rect 13818 35400 13874 35456
rect 13726 35264 13782 35320
rect 13634 35128 13690 35184
rect 13634 34448 13690 34504
rect 13542 32816 13598 32872
rect 13634 31864 13690 31920
rect 13818 34720 13874 34776
rect 14278 37576 14334 37632
rect 14002 34040 14058 34096
rect 13542 31728 13598 31784
rect 13174 29044 13176 29064
rect 13176 29044 13228 29064
rect 13228 29044 13230 29064
rect 13174 29008 13230 29044
rect 13266 28500 13268 28520
rect 13268 28500 13320 28520
rect 13320 28500 13322 28520
rect 13266 28464 13322 28500
rect 13358 28056 13414 28112
rect 13174 26696 13230 26752
rect 13910 32816 13966 32872
rect 13910 32680 13966 32736
rect 14462 37576 14518 37632
rect 14922 37460 14978 37496
rect 14922 37440 14924 37460
rect 14924 37440 14976 37460
rect 14976 37440 14978 37460
rect 14646 37304 14702 37360
rect 14186 33224 14242 33280
rect 13910 30912 13966 30968
rect 13818 30640 13874 30696
rect 14370 32952 14426 33008
rect 14278 31048 14334 31104
rect 13726 29280 13782 29336
rect 13726 29008 13782 29064
rect 13910 28736 13966 28792
rect 13634 28600 13690 28656
rect 13910 28364 13912 28384
rect 13912 28364 13964 28384
rect 13964 28364 13966 28384
rect 13910 28328 13966 28364
rect 14094 29688 14150 29744
rect 14002 27648 14058 27704
rect 13542 26560 13598 26616
rect 13910 27104 13966 27160
rect 13910 26832 13966 26888
rect 13542 24928 13598 24984
rect 13726 25100 13728 25120
rect 13728 25100 13780 25120
rect 13780 25100 13782 25120
rect 13726 25064 13782 25100
rect 13082 20440 13138 20496
rect 12990 17332 13046 17368
rect 12990 17312 12992 17332
rect 12992 17312 13044 17332
rect 13044 17312 13046 17332
rect 13726 23160 13782 23216
rect 13358 22208 13414 22264
rect 13266 17856 13322 17912
rect 13450 19352 13506 19408
rect 13634 20340 13636 20360
rect 13636 20340 13688 20360
rect 13688 20340 13690 20360
rect 13634 20304 13690 20340
rect 13358 15580 13360 15600
rect 13360 15580 13412 15600
rect 13412 15580 13414 15600
rect 13358 15544 13414 15580
rect 12990 13912 13046 13968
rect 13726 18128 13782 18184
rect 14278 29008 14334 29064
rect 14554 35148 14610 35184
rect 14554 35128 14556 35148
rect 14556 35128 14608 35148
rect 14608 35128 14610 35148
rect 14554 34856 14610 34912
rect 14554 33904 14610 33960
rect 14554 33360 14610 33416
rect 14370 28600 14426 28656
rect 14738 37068 14740 37088
rect 14740 37068 14792 37088
rect 14792 37068 14794 37088
rect 14738 37032 14794 37068
rect 15014 36488 15070 36544
rect 14738 34448 14794 34504
rect 14830 34040 14886 34096
rect 15106 35536 15162 35592
rect 15014 34176 15070 34232
rect 14738 32816 14794 32872
rect 14738 32136 14794 32192
rect 15106 33496 15162 33552
rect 15106 30912 15162 30968
rect 15014 30504 15070 30560
rect 14922 30232 14978 30288
rect 14738 28872 14794 28928
rect 14738 28736 14794 28792
rect 14186 20848 14242 20904
rect 15106 29724 15108 29744
rect 15108 29724 15160 29744
rect 15160 29724 15162 29744
rect 15106 29688 15162 29724
rect 15106 28056 15162 28112
rect 14738 25764 14794 25800
rect 14738 25744 14740 25764
rect 14740 25744 14792 25764
rect 14792 25744 14794 25764
rect 14922 24928 14978 24984
rect 14922 22752 14978 22808
rect 14646 21256 14702 21312
rect 15106 22208 15162 22264
rect 14554 19488 14610 19544
rect 14186 15272 14242 15328
rect 14646 14592 14702 14648
rect 13542 13504 13598 13560
rect 15014 20748 15016 20768
rect 15016 20748 15068 20768
rect 15068 20748 15070 20768
rect 15014 20712 15070 20748
rect 15014 20168 15070 20224
rect 15106 18264 15162 18320
rect 15014 15680 15070 15736
rect 14922 14356 14924 14376
rect 14924 14356 14976 14376
rect 14976 14356 14978 14376
rect 14922 14320 14978 14356
rect 15014 13640 15070 13696
rect 12162 3440 12218 3496
rect 12990 9036 13046 9072
rect 12990 9016 12992 9036
rect 12992 9016 13044 9036
rect 13044 9016 13046 9036
rect 13450 7964 13452 7984
rect 13452 7964 13504 7984
rect 13504 7964 13506 7984
rect 13450 7928 13506 7964
rect 12898 3440 12954 3496
rect 12806 2624 12862 2680
rect 14002 11328 14058 11384
rect 14002 10104 14058 10160
rect 13726 7384 13782 7440
rect 14922 12008 14978 12064
rect 14922 9580 14978 9616
rect 14922 9560 14924 9580
rect 14924 9560 14976 9580
rect 14976 9560 14978 9580
rect 14462 9460 14464 9480
rect 14464 9460 14516 9480
rect 14516 9460 14518 9480
rect 14462 9424 14518 9460
rect 14554 8064 14610 8120
rect 13450 3984 13506 4040
rect 14002 2644 14058 2680
rect 14002 2624 14004 2644
rect 14004 2624 14056 2644
rect 14056 2624 14058 2644
rect 15474 37848 15530 37904
rect 15750 41248 15806 41304
rect 15658 40024 15714 40080
rect 15750 37304 15806 37360
rect 15750 37068 15752 37088
rect 15752 37068 15804 37088
rect 15804 37068 15806 37088
rect 15750 37032 15806 37068
rect 15658 36352 15714 36408
rect 15566 36080 15622 36136
rect 15474 35536 15530 35592
rect 15290 33224 15346 33280
rect 15474 33360 15530 33416
rect 15566 32972 15622 33008
rect 15566 32952 15568 32972
rect 15568 32952 15620 32972
rect 15620 32952 15622 32972
rect 15566 32428 15622 32464
rect 15566 32408 15568 32428
rect 15568 32408 15620 32428
rect 15620 32408 15622 32428
rect 15566 31864 15622 31920
rect 15382 31728 15438 31784
rect 15474 31456 15530 31512
rect 15290 31048 15346 31104
rect 15956 51162 16012 51164
rect 16036 51162 16092 51164
rect 16116 51162 16172 51164
rect 16196 51162 16252 51164
rect 15956 51110 15982 51162
rect 15982 51110 16012 51162
rect 16036 51110 16046 51162
rect 16046 51110 16092 51162
rect 16116 51110 16162 51162
rect 16162 51110 16172 51162
rect 16196 51110 16226 51162
rect 16226 51110 16252 51162
rect 15956 51108 16012 51110
rect 16036 51108 16092 51110
rect 16116 51108 16172 51110
rect 16196 51108 16252 51110
rect 15956 50074 16012 50076
rect 16036 50074 16092 50076
rect 16116 50074 16172 50076
rect 16196 50074 16252 50076
rect 15956 50022 15982 50074
rect 15982 50022 16012 50074
rect 16036 50022 16046 50074
rect 16046 50022 16092 50074
rect 16116 50022 16162 50074
rect 16162 50022 16172 50074
rect 16196 50022 16226 50074
rect 16226 50022 16252 50074
rect 15956 50020 16012 50022
rect 16036 50020 16092 50022
rect 16116 50020 16172 50022
rect 16196 50020 16252 50022
rect 16026 49544 16082 49600
rect 15956 48986 16012 48988
rect 16036 48986 16092 48988
rect 16116 48986 16172 48988
rect 16196 48986 16252 48988
rect 15956 48934 15982 48986
rect 15982 48934 16012 48986
rect 16036 48934 16046 48986
rect 16046 48934 16092 48986
rect 16116 48934 16162 48986
rect 16162 48934 16172 48986
rect 16196 48934 16226 48986
rect 16226 48934 16252 48986
rect 15956 48932 16012 48934
rect 16036 48932 16092 48934
rect 16116 48932 16172 48934
rect 16196 48932 16252 48934
rect 15956 47898 16012 47900
rect 16036 47898 16092 47900
rect 16116 47898 16172 47900
rect 16196 47898 16252 47900
rect 15956 47846 15982 47898
rect 15982 47846 16012 47898
rect 16036 47846 16046 47898
rect 16046 47846 16092 47898
rect 16116 47846 16162 47898
rect 16162 47846 16172 47898
rect 16196 47846 16226 47898
rect 16226 47846 16252 47898
rect 15956 47844 16012 47846
rect 16036 47844 16092 47846
rect 16116 47844 16172 47846
rect 16196 47844 16252 47846
rect 16302 47640 16358 47696
rect 16118 46980 16174 47016
rect 16118 46960 16120 46980
rect 16120 46960 16172 46980
rect 16172 46960 16174 46980
rect 15956 46810 16012 46812
rect 16036 46810 16092 46812
rect 16116 46810 16172 46812
rect 16196 46810 16252 46812
rect 15956 46758 15982 46810
rect 15982 46758 16012 46810
rect 16036 46758 16046 46810
rect 16046 46758 16092 46810
rect 16116 46758 16162 46810
rect 16162 46758 16172 46810
rect 16196 46758 16226 46810
rect 16226 46758 16252 46810
rect 15956 46756 16012 46758
rect 16036 46756 16092 46758
rect 16116 46756 16172 46758
rect 16196 46756 16252 46758
rect 16118 45892 16174 45928
rect 16118 45872 16120 45892
rect 16120 45872 16172 45892
rect 16172 45872 16174 45892
rect 15956 45722 16012 45724
rect 16036 45722 16092 45724
rect 16116 45722 16172 45724
rect 16196 45722 16252 45724
rect 15956 45670 15982 45722
rect 15982 45670 16012 45722
rect 16036 45670 16046 45722
rect 16046 45670 16092 45722
rect 16116 45670 16162 45722
rect 16162 45670 16172 45722
rect 16196 45670 16226 45722
rect 16226 45670 16252 45722
rect 15956 45668 16012 45670
rect 16036 45668 16092 45670
rect 16116 45668 16172 45670
rect 16196 45668 16252 45670
rect 15956 44634 16012 44636
rect 16036 44634 16092 44636
rect 16116 44634 16172 44636
rect 16196 44634 16252 44636
rect 15956 44582 15982 44634
rect 15982 44582 16012 44634
rect 16036 44582 16046 44634
rect 16046 44582 16092 44634
rect 16116 44582 16162 44634
rect 16162 44582 16172 44634
rect 16196 44582 16226 44634
rect 16226 44582 16252 44634
rect 15956 44580 16012 44582
rect 16036 44580 16092 44582
rect 16116 44580 16172 44582
rect 16196 44580 16252 44582
rect 16118 44240 16174 44296
rect 15956 43546 16012 43548
rect 16036 43546 16092 43548
rect 16116 43546 16172 43548
rect 16196 43546 16252 43548
rect 15956 43494 15982 43546
rect 15982 43494 16012 43546
rect 16036 43494 16046 43546
rect 16046 43494 16092 43546
rect 16116 43494 16162 43546
rect 16162 43494 16172 43546
rect 16196 43494 16226 43546
rect 16226 43494 16252 43546
rect 15956 43492 16012 43494
rect 16036 43492 16092 43494
rect 16116 43492 16172 43494
rect 16196 43492 16252 43494
rect 15956 42458 16012 42460
rect 16036 42458 16092 42460
rect 16116 42458 16172 42460
rect 16196 42458 16252 42460
rect 15956 42406 15982 42458
rect 15982 42406 16012 42458
rect 16036 42406 16046 42458
rect 16046 42406 16092 42458
rect 16116 42406 16162 42458
rect 16162 42406 16172 42458
rect 16196 42406 16226 42458
rect 16226 42406 16252 42458
rect 15956 42404 16012 42406
rect 16036 42404 16092 42406
rect 16116 42404 16172 42406
rect 16196 42404 16252 42406
rect 17038 73344 17094 73400
rect 16578 68992 16634 69048
rect 17406 73208 17462 73264
rect 16762 63416 16818 63472
rect 16670 59472 16726 59528
rect 16578 59200 16634 59256
rect 16578 58248 16634 58304
rect 16670 56888 16726 56944
rect 16578 56380 16580 56400
rect 16580 56380 16632 56400
rect 16632 56380 16634 56400
rect 16578 56344 16634 56380
rect 16670 56072 16726 56128
rect 16486 55564 16488 55584
rect 16488 55564 16540 55584
rect 16540 55564 16542 55584
rect 16486 55528 16542 55564
rect 16670 54848 16726 54904
rect 16578 53216 16634 53272
rect 16486 52536 16542 52592
rect 16670 51448 16726 51504
rect 16486 46960 16542 47016
rect 16486 45908 16488 45928
rect 16488 45908 16540 45928
rect 16540 45908 16542 45928
rect 16486 45872 16542 45908
rect 15956 41370 16012 41372
rect 16036 41370 16092 41372
rect 16116 41370 16172 41372
rect 16196 41370 16252 41372
rect 15956 41318 15982 41370
rect 15982 41318 16012 41370
rect 16036 41318 16046 41370
rect 16046 41318 16092 41370
rect 16116 41318 16162 41370
rect 16162 41318 16172 41370
rect 16196 41318 16226 41370
rect 16226 41318 16252 41370
rect 15956 41316 16012 41318
rect 16036 41316 16092 41318
rect 16116 41316 16172 41318
rect 16196 41316 16252 41318
rect 15956 40282 16012 40284
rect 16036 40282 16092 40284
rect 16116 40282 16172 40284
rect 16196 40282 16252 40284
rect 15956 40230 15982 40282
rect 15982 40230 16012 40282
rect 16036 40230 16046 40282
rect 16046 40230 16092 40282
rect 16116 40230 16162 40282
rect 16162 40230 16172 40282
rect 16196 40230 16226 40282
rect 16226 40230 16252 40282
rect 15956 40228 16012 40230
rect 16036 40228 16092 40230
rect 16116 40228 16172 40230
rect 16196 40228 16252 40230
rect 15934 40044 15990 40080
rect 15934 40024 15936 40044
rect 15936 40024 15988 40044
rect 15988 40024 15990 40044
rect 17038 59372 17040 59392
rect 17040 59372 17092 59392
rect 17092 59372 17094 59392
rect 17038 59336 17094 59372
rect 16946 55800 17002 55856
rect 17038 55684 17094 55720
rect 17314 57160 17370 57216
rect 17038 55664 17040 55684
rect 17040 55664 17092 55684
rect 17092 55664 17094 55684
rect 17222 55528 17278 55584
rect 16946 53216 17002 53272
rect 16946 52944 17002 53000
rect 17222 52844 17224 52864
rect 17224 52844 17276 52864
rect 17276 52844 17278 52864
rect 17222 52808 17278 52844
rect 16946 51720 17002 51776
rect 16854 49852 16856 49872
rect 16856 49852 16908 49872
rect 16908 49852 16910 49872
rect 16854 49816 16910 49852
rect 16946 48456 17002 48512
rect 16854 45600 16910 45656
rect 17314 50496 17370 50552
rect 17130 48864 17186 48920
rect 15956 39194 16012 39196
rect 16036 39194 16092 39196
rect 16116 39194 16172 39196
rect 16196 39194 16252 39196
rect 15956 39142 15982 39194
rect 15982 39142 16012 39194
rect 16036 39142 16046 39194
rect 16046 39142 16092 39194
rect 16116 39142 16162 39194
rect 16162 39142 16172 39194
rect 16196 39142 16226 39194
rect 16226 39142 16252 39194
rect 15956 39140 16012 39142
rect 16036 39140 16092 39142
rect 16116 39140 16172 39142
rect 16196 39140 16252 39142
rect 16486 38800 16542 38856
rect 15956 38106 16012 38108
rect 16036 38106 16092 38108
rect 16116 38106 16172 38108
rect 16196 38106 16252 38108
rect 15956 38054 15982 38106
rect 15982 38054 16012 38106
rect 16036 38054 16046 38106
rect 16046 38054 16092 38106
rect 16116 38054 16162 38106
rect 16162 38054 16172 38106
rect 16196 38054 16226 38106
rect 16226 38054 16252 38106
rect 15956 38052 16012 38054
rect 16036 38052 16092 38054
rect 16116 38052 16172 38054
rect 16196 38052 16252 38054
rect 15934 37168 15990 37224
rect 16118 37168 16174 37224
rect 15956 37018 16012 37020
rect 16036 37018 16092 37020
rect 16116 37018 16172 37020
rect 16196 37018 16252 37020
rect 15956 36966 15982 37018
rect 15982 36966 16012 37018
rect 16036 36966 16046 37018
rect 16046 36966 16092 37018
rect 16116 36966 16162 37018
rect 16162 36966 16172 37018
rect 16196 36966 16226 37018
rect 16226 36966 16252 37018
rect 15956 36964 16012 36966
rect 16036 36964 16092 36966
rect 16116 36964 16172 36966
rect 16196 36964 16252 36966
rect 16394 37032 16450 37088
rect 16118 36352 16174 36408
rect 16210 36216 16266 36272
rect 16578 37712 16634 37768
rect 16854 37984 16910 38040
rect 15956 35930 16012 35932
rect 16036 35930 16092 35932
rect 16116 35930 16172 35932
rect 16196 35930 16252 35932
rect 15956 35878 15982 35930
rect 15982 35878 16012 35930
rect 16036 35878 16046 35930
rect 16046 35878 16092 35930
rect 16116 35878 16162 35930
rect 16162 35878 16172 35930
rect 16196 35878 16226 35930
rect 16226 35878 16252 35930
rect 15956 35876 16012 35878
rect 16036 35876 16092 35878
rect 16116 35876 16172 35878
rect 16196 35876 16252 35878
rect 16394 35808 16450 35864
rect 15934 35692 15990 35728
rect 15934 35672 15936 35692
rect 15936 35672 15988 35692
rect 15988 35672 15990 35692
rect 16026 35572 16028 35592
rect 16028 35572 16080 35592
rect 16080 35572 16082 35592
rect 16026 35536 16082 35572
rect 15956 34842 16012 34844
rect 16036 34842 16092 34844
rect 16116 34842 16172 34844
rect 16196 34842 16252 34844
rect 15956 34790 15982 34842
rect 15982 34790 16012 34842
rect 16036 34790 16046 34842
rect 16046 34790 16092 34842
rect 16116 34790 16162 34842
rect 16162 34790 16172 34842
rect 16196 34790 16226 34842
rect 16226 34790 16252 34842
rect 15956 34788 16012 34790
rect 16036 34788 16092 34790
rect 16116 34788 16172 34790
rect 16196 34788 16252 34790
rect 15956 33754 16012 33756
rect 16036 33754 16092 33756
rect 16116 33754 16172 33756
rect 16196 33754 16252 33756
rect 15956 33702 15982 33754
rect 15982 33702 16012 33754
rect 16036 33702 16046 33754
rect 16046 33702 16092 33754
rect 16116 33702 16162 33754
rect 16162 33702 16172 33754
rect 16196 33702 16226 33754
rect 16226 33702 16252 33754
rect 15956 33700 16012 33702
rect 16036 33700 16092 33702
rect 16116 33700 16172 33702
rect 16196 33700 16252 33702
rect 16210 33360 16266 33416
rect 16026 33224 16082 33280
rect 15934 32972 15990 33008
rect 15934 32952 15936 32972
rect 15936 32952 15988 32972
rect 15988 32952 15990 32972
rect 16762 35944 16818 36000
rect 16854 35128 16910 35184
rect 16486 33804 16488 33824
rect 16488 33804 16540 33824
rect 16540 33804 16542 33824
rect 16486 33768 16542 33804
rect 15956 32666 16012 32668
rect 16036 32666 16092 32668
rect 16116 32666 16172 32668
rect 16196 32666 16252 32668
rect 15956 32614 15982 32666
rect 15982 32614 16012 32666
rect 16036 32614 16046 32666
rect 16046 32614 16092 32666
rect 16116 32614 16162 32666
rect 16162 32614 16172 32666
rect 16196 32614 16226 32666
rect 16226 32614 16252 32666
rect 15956 32612 16012 32614
rect 16036 32612 16092 32614
rect 16116 32612 16172 32614
rect 16196 32612 16252 32614
rect 15750 31592 15806 31648
rect 15956 31578 16012 31580
rect 16036 31578 16092 31580
rect 16116 31578 16172 31580
rect 16196 31578 16252 31580
rect 15956 31526 15982 31578
rect 15982 31526 16012 31578
rect 16036 31526 16046 31578
rect 16046 31526 16092 31578
rect 16116 31526 16162 31578
rect 16162 31526 16172 31578
rect 16196 31526 16226 31578
rect 16226 31526 16252 31578
rect 15956 31524 16012 31526
rect 16036 31524 16092 31526
rect 16116 31524 16172 31526
rect 16196 31524 16252 31526
rect 15658 31320 15714 31376
rect 16394 31476 16450 31512
rect 16394 31456 16396 31476
rect 16396 31456 16448 31476
rect 16448 31456 16450 31476
rect 15750 29452 15752 29472
rect 15752 29452 15804 29472
rect 15804 29452 15806 29472
rect 15750 29416 15806 29452
rect 15750 29280 15806 29336
rect 15290 23160 15346 23216
rect 15566 27240 15622 27296
rect 15566 25064 15622 25120
rect 16762 33904 16818 33960
rect 16670 32136 16726 32192
rect 16578 31220 16580 31240
rect 16580 31220 16632 31240
rect 16632 31220 16634 31240
rect 16578 31184 16634 31220
rect 16394 30912 16450 30968
rect 16762 32000 16818 32056
rect 15956 30490 16012 30492
rect 16036 30490 16092 30492
rect 16116 30490 16172 30492
rect 16196 30490 16252 30492
rect 15956 30438 15982 30490
rect 15982 30438 16012 30490
rect 16036 30438 16046 30490
rect 16046 30438 16092 30490
rect 16116 30438 16162 30490
rect 16162 30438 16172 30490
rect 16196 30438 16226 30490
rect 16226 30438 16252 30490
rect 15956 30436 16012 30438
rect 16036 30436 16092 30438
rect 16116 30436 16172 30438
rect 16196 30436 16252 30438
rect 15934 30132 15936 30152
rect 15936 30132 15988 30152
rect 15988 30132 15990 30152
rect 15934 30096 15990 30132
rect 16210 29552 16266 29608
rect 15956 29402 16012 29404
rect 16036 29402 16092 29404
rect 16116 29402 16172 29404
rect 16196 29402 16252 29404
rect 15956 29350 15982 29402
rect 15982 29350 16012 29402
rect 16036 29350 16046 29402
rect 16046 29350 16092 29402
rect 16116 29350 16162 29402
rect 16162 29350 16172 29402
rect 16196 29350 16226 29402
rect 16226 29350 16252 29402
rect 15956 29348 16012 29350
rect 16036 29348 16092 29350
rect 16116 29348 16172 29350
rect 16196 29348 16252 29350
rect 16026 28736 16082 28792
rect 15934 28600 15990 28656
rect 16762 30776 16818 30832
rect 16670 30676 16672 30696
rect 16672 30676 16724 30696
rect 16724 30676 16726 30696
rect 16486 30232 16542 30288
rect 16670 30640 16726 30676
rect 16670 30504 16726 30560
rect 16394 28736 16450 28792
rect 16578 29280 16634 29336
rect 15956 28314 16012 28316
rect 16036 28314 16092 28316
rect 16116 28314 16172 28316
rect 16196 28314 16252 28316
rect 15956 28262 15982 28314
rect 15982 28262 16012 28314
rect 16036 28262 16046 28314
rect 16046 28262 16092 28314
rect 16116 28262 16162 28314
rect 16162 28262 16172 28314
rect 16196 28262 16226 28314
rect 16226 28262 16252 28314
rect 15956 28260 16012 28262
rect 16036 28260 16092 28262
rect 16116 28260 16172 28262
rect 16196 28260 16252 28262
rect 15934 28056 15990 28112
rect 16394 27648 16450 27704
rect 16210 27376 16266 27432
rect 15956 27226 16012 27228
rect 16036 27226 16092 27228
rect 16116 27226 16172 27228
rect 16196 27226 16252 27228
rect 15956 27174 15982 27226
rect 15982 27174 16012 27226
rect 16036 27174 16046 27226
rect 16046 27174 16092 27226
rect 16116 27174 16162 27226
rect 16162 27174 16172 27226
rect 16196 27174 16226 27226
rect 16226 27174 16252 27226
rect 15956 27172 16012 27174
rect 16036 27172 16092 27174
rect 16116 27172 16172 27174
rect 16196 27172 16252 27174
rect 15658 24928 15714 24984
rect 15382 22616 15438 22672
rect 15290 21936 15346 21992
rect 15658 21528 15714 21584
rect 15566 21120 15622 21176
rect 15382 19488 15438 19544
rect 15566 17876 15622 17912
rect 15566 17856 15568 17876
rect 15568 17856 15620 17876
rect 15620 17856 15622 17876
rect 16394 27124 16450 27160
rect 16394 27104 16396 27124
rect 16396 27104 16448 27124
rect 16448 27104 16450 27124
rect 16854 29824 16910 29880
rect 16854 29008 16910 29064
rect 16762 28872 16818 28928
rect 16670 28192 16726 28248
rect 16762 27920 16818 27976
rect 16670 27532 16726 27568
rect 16670 27512 16672 27532
rect 16672 27512 16724 27532
rect 16724 27512 16726 27532
rect 16670 27376 16726 27432
rect 15956 26138 16012 26140
rect 16036 26138 16092 26140
rect 16116 26138 16172 26140
rect 16196 26138 16252 26140
rect 15956 26086 15982 26138
rect 15982 26086 16012 26138
rect 16036 26086 16046 26138
rect 16046 26086 16092 26138
rect 16116 26086 16162 26138
rect 16162 26086 16172 26138
rect 16196 26086 16226 26138
rect 16226 26086 16252 26138
rect 15956 26084 16012 26086
rect 16036 26084 16092 26086
rect 16116 26084 16172 26086
rect 16196 26084 16252 26086
rect 16210 25644 16212 25664
rect 16212 25644 16264 25664
rect 16264 25644 16266 25664
rect 16210 25608 16266 25644
rect 15956 25050 16012 25052
rect 16036 25050 16092 25052
rect 16116 25050 16172 25052
rect 16196 25050 16252 25052
rect 15956 24998 15982 25050
rect 15982 24998 16012 25050
rect 16036 24998 16046 25050
rect 16046 24998 16092 25050
rect 16116 24998 16162 25050
rect 16162 24998 16172 25050
rect 16196 24998 16226 25050
rect 16226 24998 16252 25050
rect 15956 24996 16012 24998
rect 16036 24996 16092 24998
rect 16116 24996 16172 24998
rect 16196 24996 16252 24998
rect 15842 24656 15898 24712
rect 17038 28872 17094 28928
rect 15956 23962 16012 23964
rect 16036 23962 16092 23964
rect 16116 23962 16172 23964
rect 16196 23962 16252 23964
rect 15956 23910 15982 23962
rect 15982 23910 16012 23962
rect 16036 23910 16046 23962
rect 16046 23910 16092 23962
rect 16116 23910 16162 23962
rect 16162 23910 16172 23962
rect 16196 23910 16226 23962
rect 16226 23910 16252 23962
rect 15956 23908 16012 23910
rect 16036 23908 16092 23910
rect 16116 23908 16172 23910
rect 16196 23908 16252 23910
rect 15956 22874 16012 22876
rect 16036 22874 16092 22876
rect 16116 22874 16172 22876
rect 16196 22874 16252 22876
rect 15956 22822 15982 22874
rect 15982 22822 16012 22874
rect 16036 22822 16046 22874
rect 16046 22822 16092 22874
rect 16116 22822 16162 22874
rect 16162 22822 16172 22874
rect 16196 22822 16226 22874
rect 16226 22822 16252 22874
rect 15956 22820 16012 22822
rect 16036 22820 16092 22822
rect 16116 22820 16172 22822
rect 16196 22820 16252 22822
rect 15566 17332 15622 17368
rect 15566 17312 15568 17332
rect 15568 17312 15620 17332
rect 15620 17312 15622 17332
rect 15382 15952 15438 16008
rect 15956 21786 16012 21788
rect 16036 21786 16092 21788
rect 16116 21786 16172 21788
rect 16196 21786 16252 21788
rect 15956 21734 15982 21786
rect 15982 21734 16012 21786
rect 16036 21734 16046 21786
rect 16046 21734 16092 21786
rect 16116 21734 16162 21786
rect 16162 21734 16172 21786
rect 16196 21734 16226 21786
rect 16226 21734 16252 21786
rect 15956 21732 16012 21734
rect 16036 21732 16092 21734
rect 16116 21732 16172 21734
rect 16196 21732 16252 21734
rect 16486 23740 16488 23760
rect 16488 23740 16540 23760
rect 16540 23740 16542 23760
rect 16486 23704 16542 23740
rect 16670 23704 16726 23760
rect 16486 23568 16542 23624
rect 16578 22380 16580 22400
rect 16580 22380 16632 22400
rect 16632 22380 16634 22400
rect 16578 22344 16634 22380
rect 16210 21392 16266 21448
rect 15956 20698 16012 20700
rect 16036 20698 16092 20700
rect 16116 20698 16172 20700
rect 16196 20698 16252 20700
rect 15956 20646 15982 20698
rect 15982 20646 16012 20698
rect 16036 20646 16046 20698
rect 16046 20646 16092 20698
rect 16116 20646 16162 20698
rect 16162 20646 16172 20698
rect 16196 20646 16226 20698
rect 16226 20646 16252 20698
rect 15956 20644 16012 20646
rect 16036 20644 16092 20646
rect 16116 20644 16172 20646
rect 16196 20644 16252 20646
rect 15956 19610 16012 19612
rect 16036 19610 16092 19612
rect 16116 19610 16172 19612
rect 16196 19610 16252 19612
rect 15956 19558 15982 19610
rect 15982 19558 16012 19610
rect 16036 19558 16046 19610
rect 16046 19558 16092 19610
rect 16116 19558 16162 19610
rect 16162 19558 16172 19610
rect 16196 19558 16226 19610
rect 16226 19558 16252 19610
rect 15956 19556 16012 19558
rect 16036 19556 16092 19558
rect 16116 19556 16172 19558
rect 16196 19556 16252 19558
rect 15956 18522 16012 18524
rect 16036 18522 16092 18524
rect 16116 18522 16172 18524
rect 16196 18522 16252 18524
rect 15956 18470 15982 18522
rect 15982 18470 16012 18522
rect 16036 18470 16046 18522
rect 16046 18470 16092 18522
rect 16116 18470 16162 18522
rect 16162 18470 16172 18522
rect 16196 18470 16226 18522
rect 16226 18470 16252 18522
rect 15956 18468 16012 18470
rect 16036 18468 16092 18470
rect 16116 18468 16172 18470
rect 16196 18468 16252 18470
rect 15956 17434 16012 17436
rect 16036 17434 16092 17436
rect 16116 17434 16172 17436
rect 16196 17434 16252 17436
rect 15956 17382 15982 17434
rect 15982 17382 16012 17434
rect 16036 17382 16046 17434
rect 16046 17382 16092 17434
rect 16116 17382 16162 17434
rect 16162 17382 16172 17434
rect 16196 17382 16226 17434
rect 16226 17382 16252 17434
rect 15956 17380 16012 17382
rect 16036 17380 16092 17382
rect 16116 17380 16172 17382
rect 16196 17380 16252 17382
rect 15956 16346 16012 16348
rect 16036 16346 16092 16348
rect 16116 16346 16172 16348
rect 16196 16346 16252 16348
rect 15956 16294 15982 16346
rect 15982 16294 16012 16346
rect 16036 16294 16046 16346
rect 16046 16294 16092 16346
rect 16116 16294 16162 16346
rect 16162 16294 16172 16346
rect 16196 16294 16226 16346
rect 16226 16294 16252 16346
rect 15956 16292 16012 16294
rect 16036 16292 16092 16294
rect 16116 16292 16172 16294
rect 16196 16292 16252 16294
rect 16210 16088 16266 16144
rect 15474 15580 15476 15600
rect 15476 15580 15528 15600
rect 15528 15580 15530 15600
rect 15474 15544 15530 15580
rect 15956 15258 16012 15260
rect 16036 15258 16092 15260
rect 16116 15258 16172 15260
rect 16196 15258 16252 15260
rect 15956 15206 15982 15258
rect 15982 15206 16012 15258
rect 16036 15206 16046 15258
rect 16046 15206 16092 15258
rect 16116 15206 16162 15258
rect 16162 15206 16172 15258
rect 16196 15206 16226 15258
rect 16226 15206 16252 15258
rect 15956 15204 16012 15206
rect 16036 15204 16092 15206
rect 16116 15204 16172 15206
rect 16196 15204 16252 15206
rect 15566 13932 15622 13968
rect 15566 13912 15568 13932
rect 15568 13912 15620 13932
rect 15620 13912 15622 13932
rect 15382 12144 15438 12200
rect 15956 14170 16012 14172
rect 16036 14170 16092 14172
rect 16116 14170 16172 14172
rect 16196 14170 16252 14172
rect 15956 14118 15982 14170
rect 15982 14118 16012 14170
rect 16036 14118 16046 14170
rect 16046 14118 16092 14170
rect 16116 14118 16162 14170
rect 16162 14118 16172 14170
rect 16196 14118 16226 14170
rect 16226 14118 16252 14170
rect 15956 14116 16012 14118
rect 16036 14116 16092 14118
rect 16116 14116 16172 14118
rect 16196 14116 16252 14118
rect 15956 13082 16012 13084
rect 16036 13082 16092 13084
rect 16116 13082 16172 13084
rect 16196 13082 16252 13084
rect 15956 13030 15982 13082
rect 15982 13030 16012 13082
rect 16036 13030 16046 13082
rect 16046 13030 16092 13082
rect 16116 13030 16162 13082
rect 16162 13030 16172 13082
rect 16196 13030 16226 13082
rect 16226 13030 16252 13082
rect 15956 13028 16012 13030
rect 16036 13028 16092 13030
rect 16116 13028 16172 13030
rect 16196 13028 16252 13030
rect 15956 11994 16012 11996
rect 16036 11994 16092 11996
rect 16116 11994 16172 11996
rect 16196 11994 16252 11996
rect 15956 11942 15982 11994
rect 15982 11942 16012 11994
rect 16036 11942 16046 11994
rect 16046 11942 16092 11994
rect 16116 11942 16162 11994
rect 16162 11942 16172 11994
rect 16196 11942 16226 11994
rect 16226 11942 16252 11994
rect 15956 11940 16012 11942
rect 16036 11940 16092 11942
rect 16116 11940 16172 11942
rect 16196 11940 16252 11942
rect 15198 8200 15254 8256
rect 15956 10906 16012 10908
rect 16036 10906 16092 10908
rect 16116 10906 16172 10908
rect 16196 10906 16252 10908
rect 15956 10854 15982 10906
rect 15982 10854 16012 10906
rect 16036 10854 16046 10906
rect 16046 10854 16092 10906
rect 16116 10854 16162 10906
rect 16162 10854 16172 10906
rect 16196 10854 16226 10906
rect 16226 10854 16252 10906
rect 15956 10852 16012 10854
rect 16036 10852 16092 10854
rect 16116 10852 16172 10854
rect 16196 10852 16252 10854
rect 16670 20884 16672 20904
rect 16672 20884 16724 20904
rect 16724 20884 16726 20904
rect 16670 20848 16726 20884
rect 17314 47912 17370 47968
rect 17590 71032 17646 71088
rect 17682 67768 17738 67824
rect 18786 71440 18842 71496
rect 18602 67496 18658 67552
rect 17774 66020 17830 66056
rect 17774 66000 17776 66020
rect 17776 66000 17828 66020
rect 17828 66000 17830 66020
rect 18694 65456 18750 65512
rect 18234 64932 18290 64968
rect 18234 64912 18236 64932
rect 18236 64912 18288 64932
rect 18288 64912 18290 64932
rect 18602 63980 18658 64016
rect 18602 63960 18604 63980
rect 18604 63960 18656 63980
rect 18656 63960 18658 63980
rect 19706 72664 19762 72720
rect 18878 70352 18934 70408
rect 19062 68856 19118 68912
rect 18878 63960 18934 64016
rect 18786 63416 18842 63472
rect 17958 62736 18014 62792
rect 17590 59100 17592 59120
rect 17592 59100 17644 59120
rect 17644 59100 17646 59120
rect 17590 59064 17646 59100
rect 17774 58928 17830 58984
rect 17498 57704 17554 57760
rect 17774 55836 17776 55856
rect 17776 55836 17828 55856
rect 17828 55836 17830 55856
rect 17774 55800 17830 55836
rect 17774 55392 17830 55448
rect 17590 52128 17646 52184
rect 17682 50768 17738 50824
rect 17498 48320 17554 48376
rect 17590 47540 17592 47560
rect 17592 47540 17644 47560
rect 17644 47540 17646 47560
rect 17590 47504 17646 47540
rect 17682 47232 17738 47288
rect 17222 44648 17278 44704
rect 17222 43832 17278 43888
rect 17222 43560 17278 43616
rect 17774 45736 17830 45792
rect 17498 44396 17554 44432
rect 17498 44376 17500 44396
rect 17500 44376 17552 44396
rect 17552 44376 17554 44396
rect 17682 44140 17684 44160
rect 17684 44140 17736 44160
rect 17736 44140 17738 44160
rect 17682 44104 17738 44140
rect 17590 43868 17592 43888
rect 17592 43868 17644 43888
rect 17644 43868 17646 43888
rect 17590 43832 17646 43868
rect 17222 37304 17278 37360
rect 17222 34448 17278 34504
rect 17222 31728 17278 31784
rect 17222 30252 17278 30288
rect 17222 30232 17224 30252
rect 17224 30232 17276 30252
rect 17276 30232 17278 30252
rect 17222 28500 17224 28520
rect 17224 28500 17276 28520
rect 17276 28500 17278 28520
rect 17222 28464 17278 28500
rect 16946 21120 17002 21176
rect 16670 20440 16726 20496
rect 16762 19216 16818 19272
rect 17038 19896 17094 19952
rect 17130 19352 17186 19408
rect 17038 19216 17094 19272
rect 16854 15680 16910 15736
rect 17682 36760 17738 36816
rect 17590 35264 17646 35320
rect 17498 31592 17554 31648
rect 17498 30268 17500 30288
rect 17500 30268 17552 30288
rect 17552 30268 17554 30288
rect 17498 30232 17554 30268
rect 17774 35128 17830 35184
rect 17774 32680 17830 32736
rect 17682 31728 17738 31784
rect 17590 28600 17646 28656
rect 17590 27668 17646 27704
rect 17590 27648 17592 27668
rect 17592 27648 17644 27668
rect 17644 27648 17646 27668
rect 17590 26696 17646 26752
rect 17406 17076 17408 17096
rect 17408 17076 17460 17096
rect 17460 17076 17462 17096
rect 17406 17040 17462 17076
rect 17406 14592 17462 14648
rect 17682 21548 17738 21584
rect 17682 21528 17684 21548
rect 17684 21528 17736 21548
rect 17736 21528 17738 21548
rect 17498 13640 17554 13696
rect 17222 11736 17278 11792
rect 15474 8064 15530 8120
rect 15956 9818 16012 9820
rect 16036 9818 16092 9820
rect 16116 9818 16172 9820
rect 16196 9818 16252 9820
rect 15956 9766 15982 9818
rect 15982 9766 16012 9818
rect 16036 9766 16046 9818
rect 16046 9766 16092 9818
rect 16116 9766 16162 9818
rect 16162 9766 16172 9818
rect 16196 9766 16226 9818
rect 16226 9766 16252 9818
rect 15956 9764 16012 9766
rect 16036 9764 16092 9766
rect 16116 9764 16172 9766
rect 16196 9764 16252 9766
rect 16302 9424 16358 9480
rect 17038 9036 17094 9072
rect 17038 9016 17040 9036
rect 17040 9016 17092 9036
rect 17092 9016 17094 9036
rect 15956 8730 16012 8732
rect 16036 8730 16092 8732
rect 16116 8730 16172 8732
rect 16196 8730 16252 8732
rect 15956 8678 15982 8730
rect 15982 8678 16012 8730
rect 16036 8678 16046 8730
rect 16046 8678 16092 8730
rect 16116 8678 16162 8730
rect 16162 8678 16172 8730
rect 16196 8678 16226 8730
rect 16226 8678 16252 8730
rect 15956 8676 16012 8678
rect 16036 8676 16092 8678
rect 16116 8676 16172 8678
rect 16196 8676 16252 8678
rect 16854 8880 16910 8936
rect 16486 8472 16542 8528
rect 17038 8336 17094 8392
rect 15956 7642 16012 7644
rect 16036 7642 16092 7644
rect 16116 7642 16172 7644
rect 16196 7642 16252 7644
rect 15956 7590 15982 7642
rect 15982 7590 16012 7642
rect 16036 7590 16046 7642
rect 16046 7590 16092 7642
rect 16116 7590 16162 7642
rect 16162 7590 16172 7642
rect 16196 7590 16226 7642
rect 16226 7590 16252 7642
rect 15956 7588 16012 7590
rect 16036 7588 16092 7590
rect 16116 7588 16172 7590
rect 16196 7588 16252 7590
rect 15956 6554 16012 6556
rect 16036 6554 16092 6556
rect 16116 6554 16172 6556
rect 16196 6554 16252 6556
rect 15956 6502 15982 6554
rect 15982 6502 16012 6554
rect 16036 6502 16046 6554
rect 16046 6502 16092 6554
rect 16116 6502 16162 6554
rect 16162 6502 16172 6554
rect 16196 6502 16226 6554
rect 16226 6502 16252 6554
rect 15956 6500 16012 6502
rect 16036 6500 16092 6502
rect 16116 6500 16172 6502
rect 16196 6500 16252 6502
rect 15198 3984 15254 4040
rect 15956 5466 16012 5468
rect 16036 5466 16092 5468
rect 16116 5466 16172 5468
rect 16196 5466 16252 5468
rect 15956 5414 15982 5466
rect 15982 5414 16012 5466
rect 16036 5414 16046 5466
rect 16046 5414 16092 5466
rect 16116 5414 16162 5466
rect 16162 5414 16172 5466
rect 16196 5414 16226 5466
rect 16226 5414 16252 5466
rect 15956 5412 16012 5414
rect 16036 5412 16092 5414
rect 16116 5412 16172 5414
rect 16196 5412 16252 5414
rect 15956 4378 16012 4380
rect 16036 4378 16092 4380
rect 16116 4378 16172 4380
rect 16196 4378 16252 4380
rect 15956 4326 15982 4378
rect 15982 4326 16012 4378
rect 16036 4326 16046 4378
rect 16046 4326 16092 4378
rect 16116 4326 16162 4378
rect 16162 4326 16172 4378
rect 16196 4326 16226 4378
rect 16226 4326 16252 4378
rect 15956 4324 16012 4326
rect 16036 4324 16092 4326
rect 16116 4324 16172 4326
rect 16196 4324 16252 4326
rect 16302 3984 16358 4040
rect 15566 3440 15622 3496
rect 15956 3290 16012 3292
rect 16036 3290 16092 3292
rect 16116 3290 16172 3292
rect 16196 3290 16252 3292
rect 15956 3238 15982 3290
rect 15982 3238 16012 3290
rect 16036 3238 16046 3290
rect 16046 3238 16092 3290
rect 16116 3238 16162 3290
rect 16162 3238 16172 3290
rect 16196 3238 16226 3290
rect 16226 3238 16252 3290
rect 15956 3236 16012 3238
rect 16036 3236 16092 3238
rect 16116 3236 16172 3238
rect 16196 3236 16252 3238
rect 15956 2202 16012 2204
rect 16036 2202 16092 2204
rect 16116 2202 16172 2204
rect 16196 2202 16252 2204
rect 15956 2150 15982 2202
rect 15982 2150 16012 2202
rect 16036 2150 16046 2202
rect 16046 2150 16092 2202
rect 16116 2150 16162 2202
rect 16162 2150 16172 2202
rect 16196 2150 16226 2202
rect 16226 2150 16252 2202
rect 15956 2148 16012 2150
rect 16036 2148 16092 2150
rect 16116 2148 16172 2150
rect 16196 2148 16252 2150
rect 18878 60732 18880 60752
rect 18880 60732 18932 60752
rect 18932 60732 18934 60752
rect 18878 60696 18934 60732
rect 18234 59472 18290 59528
rect 17958 58520 18014 58576
rect 17958 55528 18014 55584
rect 18970 58792 19026 58848
rect 19154 59200 19210 59256
rect 18510 57704 18566 57760
rect 18694 57704 18750 57760
rect 18050 52672 18106 52728
rect 18234 53488 18290 53544
rect 17958 50380 18014 50416
rect 17958 50360 17960 50380
rect 17960 50360 18012 50380
rect 18012 50360 18014 50380
rect 18050 48628 18052 48648
rect 18052 48628 18104 48648
rect 18104 48628 18106 48648
rect 18050 48592 18106 48628
rect 18050 48048 18106 48104
rect 18786 56208 18842 56264
rect 18694 55256 18750 55312
rect 18602 54576 18658 54632
rect 18510 52944 18566 53000
rect 18786 53760 18842 53816
rect 18694 53644 18750 53680
rect 18694 53624 18696 53644
rect 18696 53624 18748 53644
rect 18748 53624 18750 53644
rect 18694 50088 18750 50144
rect 19062 56480 19118 56536
rect 18878 50632 18934 50688
rect 18694 49716 18696 49736
rect 18696 49716 18748 49736
rect 18748 49716 18750 49736
rect 18694 49680 18750 49716
rect 19154 51312 19210 51368
rect 18970 48320 19026 48376
rect 18142 47640 18198 47696
rect 19062 48184 19118 48240
rect 18234 47368 18290 47424
rect 18142 46280 18198 46336
rect 18878 45872 18934 45928
rect 18510 44276 18512 44296
rect 18512 44276 18564 44296
rect 18564 44276 18566 44296
rect 18510 44240 18566 44276
rect 18050 43424 18106 43480
rect 18878 44376 18934 44432
rect 18142 40840 18198 40896
rect 17958 36216 18014 36272
rect 18142 35828 18198 35864
rect 18142 35808 18144 35828
rect 18144 35808 18196 35828
rect 18196 35808 18198 35828
rect 18234 35708 18236 35728
rect 18236 35708 18288 35728
rect 18288 35708 18290 35728
rect 18234 35672 18290 35708
rect 17958 34720 18014 34776
rect 18142 30504 18198 30560
rect 18050 29688 18106 29744
rect 18050 27920 18106 27976
rect 18142 27104 18198 27160
rect 18234 26968 18290 27024
rect 18142 26560 18198 26616
rect 18050 24112 18106 24168
rect 18050 21664 18106 21720
rect 18050 21392 18106 21448
rect 17866 12144 17922 12200
rect 18142 8200 18198 8256
rect 17774 7248 17830 7304
rect 18510 38004 18566 38040
rect 18510 37984 18512 38004
rect 18512 37984 18564 38004
rect 18564 37984 18566 38004
rect 19062 42744 19118 42800
rect 18970 40976 19026 41032
rect 18694 39208 18750 39264
rect 18786 34312 18842 34368
rect 18786 33768 18842 33824
rect 18878 33632 18934 33688
rect 18418 26988 18474 27024
rect 18418 26968 18420 26988
rect 18420 26968 18472 26988
rect 18472 26968 18474 26988
rect 18418 26036 18474 26072
rect 18418 26016 18420 26036
rect 18420 26016 18472 26036
rect 18472 26016 18474 26036
rect 18418 25744 18474 25800
rect 18510 23568 18566 23624
rect 18786 31320 18842 31376
rect 19154 35672 19210 35728
rect 19062 34720 19118 34776
rect 19062 34604 19118 34640
rect 19062 34584 19064 34604
rect 19064 34584 19116 34604
rect 19116 34584 19118 34604
rect 19338 57996 19394 58032
rect 19338 57976 19340 57996
rect 19340 57976 19392 57996
rect 19392 57976 19394 57996
rect 19338 57024 19394 57080
rect 19338 54576 19394 54632
rect 20956 77818 21012 77820
rect 21036 77818 21092 77820
rect 21116 77818 21172 77820
rect 21196 77818 21252 77820
rect 20956 77766 20982 77818
rect 20982 77766 21012 77818
rect 21036 77766 21046 77818
rect 21046 77766 21092 77818
rect 21116 77766 21162 77818
rect 21162 77766 21172 77818
rect 21196 77766 21226 77818
rect 21226 77766 21252 77818
rect 20956 77764 21012 77766
rect 21036 77764 21092 77766
rect 21116 77764 21172 77766
rect 21196 77764 21252 77766
rect 20956 76730 21012 76732
rect 21036 76730 21092 76732
rect 21116 76730 21172 76732
rect 21196 76730 21252 76732
rect 20956 76678 20982 76730
rect 20982 76678 21012 76730
rect 21036 76678 21046 76730
rect 21046 76678 21092 76730
rect 21116 76678 21162 76730
rect 21162 76678 21172 76730
rect 21196 76678 21226 76730
rect 21226 76678 21252 76730
rect 20956 76676 21012 76678
rect 21036 76676 21092 76678
rect 21116 76676 21172 76678
rect 21196 76676 21252 76678
rect 21270 76336 21326 76392
rect 20810 75656 20866 75712
rect 20956 75642 21012 75644
rect 21036 75642 21092 75644
rect 21116 75642 21172 75644
rect 21196 75642 21252 75644
rect 20956 75590 20982 75642
rect 20982 75590 21012 75642
rect 21036 75590 21046 75642
rect 21046 75590 21092 75642
rect 21116 75590 21162 75642
rect 21162 75590 21172 75642
rect 21196 75590 21226 75642
rect 21226 75590 21252 75642
rect 20956 75588 21012 75590
rect 21036 75588 21092 75590
rect 21116 75588 21172 75590
rect 21196 75588 21252 75590
rect 20810 75248 20866 75304
rect 20956 74554 21012 74556
rect 21036 74554 21092 74556
rect 21116 74554 21172 74556
rect 21196 74554 21252 74556
rect 20956 74502 20982 74554
rect 20982 74502 21012 74554
rect 21036 74502 21046 74554
rect 21046 74502 21092 74554
rect 21116 74502 21162 74554
rect 21162 74502 21172 74554
rect 21196 74502 21226 74554
rect 21226 74502 21252 74554
rect 20956 74500 21012 74502
rect 21036 74500 21092 74502
rect 21116 74500 21172 74502
rect 21196 74500 21252 74502
rect 20956 73466 21012 73468
rect 21036 73466 21092 73468
rect 21116 73466 21172 73468
rect 21196 73466 21252 73468
rect 20956 73414 20982 73466
rect 20982 73414 21012 73466
rect 21036 73414 21046 73466
rect 21046 73414 21092 73466
rect 21116 73414 21162 73466
rect 21162 73414 21172 73466
rect 21196 73414 21226 73466
rect 21226 73414 21252 73466
rect 20956 73412 21012 73414
rect 21036 73412 21092 73414
rect 21116 73412 21172 73414
rect 21196 73412 21252 73414
rect 20810 73344 20866 73400
rect 20956 72378 21012 72380
rect 21036 72378 21092 72380
rect 21116 72378 21172 72380
rect 21196 72378 21252 72380
rect 20956 72326 20982 72378
rect 20982 72326 21012 72378
rect 21036 72326 21046 72378
rect 21046 72326 21092 72378
rect 21116 72326 21162 72378
rect 21162 72326 21172 72378
rect 21196 72326 21226 72378
rect 21226 72326 21252 72378
rect 20956 72324 21012 72326
rect 21036 72324 21092 72326
rect 21116 72324 21172 72326
rect 21196 72324 21252 72326
rect 20718 68992 20774 69048
rect 20350 62328 20406 62384
rect 20166 62192 20222 62248
rect 19614 58928 19670 58984
rect 19522 51992 19578 52048
rect 19338 48728 19394 48784
rect 19430 48456 19486 48512
rect 19430 47096 19486 47152
rect 19430 43968 19486 44024
rect 19338 43152 19394 43208
rect 19430 39888 19486 39944
rect 20258 58792 20314 58848
rect 20074 50768 20130 50824
rect 19982 48864 20038 48920
rect 19890 48592 19946 48648
rect 20074 48456 20130 48512
rect 19982 47776 20038 47832
rect 19522 38800 19578 38856
rect 19706 44648 19762 44704
rect 20074 45772 20076 45792
rect 20076 45772 20128 45792
rect 20128 45772 20130 45792
rect 20074 45736 20130 45772
rect 19890 44104 19946 44160
rect 19890 42336 19946 42392
rect 20074 41928 20130 41984
rect 19798 41112 19854 41168
rect 19614 36760 19670 36816
rect 19614 36624 19670 36680
rect 19430 35536 19486 35592
rect 19338 35400 19394 35456
rect 19430 34992 19486 35048
rect 19430 33260 19432 33280
rect 19432 33260 19484 33280
rect 19484 33260 19486 33280
rect 19430 33224 19486 33260
rect 19706 33224 19762 33280
rect 18970 31184 19026 31240
rect 18694 29960 18750 30016
rect 18878 28756 18934 28792
rect 18878 28736 18880 28756
rect 18880 28736 18932 28756
rect 18932 28736 18934 28756
rect 18694 27512 18750 27568
rect 19246 30268 19248 30288
rect 19248 30268 19300 30288
rect 19300 30268 19302 30288
rect 19246 30232 19302 30268
rect 19430 30116 19486 30152
rect 19430 30096 19432 30116
rect 19432 30096 19484 30116
rect 19484 30096 19486 30116
rect 19062 29416 19118 29472
rect 19338 28872 19394 28928
rect 19614 28192 19670 28248
rect 19430 28056 19486 28112
rect 19246 25200 19302 25256
rect 19154 24792 19210 24848
rect 19062 21256 19118 21312
rect 18418 11600 18474 11656
rect 19062 10532 19118 10568
rect 19062 10512 19064 10532
rect 19064 10512 19116 10532
rect 19116 10512 19118 10532
rect 18326 5480 18382 5536
rect 19246 20748 19248 20768
rect 19248 20748 19300 20768
rect 19300 20748 19302 20768
rect 19246 20712 19302 20748
rect 19522 20304 19578 20360
rect 19430 5480 19486 5536
rect 19154 5208 19210 5264
rect 17682 1944 17738 2000
rect 19982 36488 20038 36544
rect 19890 34448 19946 34504
rect 19982 32716 19984 32736
rect 19984 32716 20036 32736
rect 20036 32716 20038 32736
rect 19982 32680 20038 32716
rect 20074 31592 20130 31648
rect 19982 31084 19984 31104
rect 19984 31084 20036 31104
rect 20036 31084 20038 31104
rect 19982 31048 20038 31084
rect 19890 29300 19946 29336
rect 19890 29280 19892 29300
rect 19892 29280 19944 29300
rect 19944 29280 19946 29300
rect 20074 27820 20076 27840
rect 20076 27820 20128 27840
rect 20128 27820 20130 27840
rect 20074 27784 20130 27820
rect 20074 27532 20130 27568
rect 20074 27512 20076 27532
rect 20076 27512 20128 27532
rect 20128 27512 20130 27532
rect 19890 21392 19946 21448
rect 20718 63960 20774 64016
rect 20956 71290 21012 71292
rect 21036 71290 21092 71292
rect 21116 71290 21172 71292
rect 21196 71290 21252 71292
rect 20956 71238 20982 71290
rect 20982 71238 21012 71290
rect 21036 71238 21046 71290
rect 21046 71238 21092 71290
rect 21116 71238 21162 71290
rect 21162 71238 21172 71290
rect 21196 71238 21226 71290
rect 21226 71238 21252 71290
rect 20956 71236 21012 71238
rect 21036 71236 21092 71238
rect 21116 71236 21172 71238
rect 21196 71236 21252 71238
rect 20902 70524 20904 70544
rect 20904 70524 20956 70544
rect 20956 70524 20958 70544
rect 20902 70488 20958 70524
rect 20956 70202 21012 70204
rect 21036 70202 21092 70204
rect 21116 70202 21172 70204
rect 21196 70202 21252 70204
rect 20956 70150 20982 70202
rect 20982 70150 21012 70202
rect 21036 70150 21046 70202
rect 21046 70150 21092 70202
rect 21116 70150 21162 70202
rect 21162 70150 21172 70202
rect 21196 70150 21226 70202
rect 21226 70150 21252 70202
rect 20956 70148 21012 70150
rect 21036 70148 21092 70150
rect 21116 70148 21172 70150
rect 21196 70148 21252 70150
rect 21270 69672 21326 69728
rect 20956 69114 21012 69116
rect 21036 69114 21092 69116
rect 21116 69114 21172 69116
rect 21196 69114 21252 69116
rect 20956 69062 20982 69114
rect 20982 69062 21012 69114
rect 21036 69062 21046 69114
rect 21046 69062 21092 69114
rect 21116 69062 21162 69114
rect 21162 69062 21172 69114
rect 21196 69062 21226 69114
rect 21226 69062 21252 69114
rect 20956 69060 21012 69062
rect 21036 69060 21092 69062
rect 21116 69060 21172 69062
rect 21196 69060 21252 69062
rect 20956 68026 21012 68028
rect 21036 68026 21092 68028
rect 21116 68026 21172 68028
rect 21196 68026 21252 68028
rect 20956 67974 20982 68026
rect 20982 67974 21012 68026
rect 21036 67974 21046 68026
rect 21046 67974 21092 68026
rect 21116 67974 21162 68026
rect 21162 67974 21172 68026
rect 21196 67974 21226 68026
rect 21226 67974 21252 68026
rect 20956 67972 21012 67974
rect 21036 67972 21092 67974
rect 21116 67972 21172 67974
rect 21196 67972 21252 67974
rect 21454 67632 21510 67688
rect 20956 66938 21012 66940
rect 21036 66938 21092 66940
rect 21116 66938 21172 66940
rect 21196 66938 21252 66940
rect 20956 66886 20982 66938
rect 20982 66886 21012 66938
rect 21036 66886 21046 66938
rect 21046 66886 21092 66938
rect 21116 66886 21162 66938
rect 21162 66886 21172 66938
rect 21196 66886 21226 66938
rect 21226 66886 21252 66938
rect 20956 66884 21012 66886
rect 21036 66884 21092 66886
rect 21116 66884 21172 66886
rect 21196 66884 21252 66886
rect 20956 65850 21012 65852
rect 21036 65850 21092 65852
rect 21116 65850 21172 65852
rect 21196 65850 21252 65852
rect 20956 65798 20982 65850
rect 20982 65798 21012 65850
rect 21036 65798 21046 65850
rect 21046 65798 21092 65850
rect 21116 65798 21162 65850
rect 21162 65798 21172 65850
rect 21196 65798 21226 65850
rect 21226 65798 21252 65850
rect 20956 65796 21012 65798
rect 21036 65796 21092 65798
rect 21116 65796 21172 65798
rect 21196 65796 21252 65798
rect 20956 64762 21012 64764
rect 21036 64762 21092 64764
rect 21116 64762 21172 64764
rect 21196 64762 21252 64764
rect 20956 64710 20982 64762
rect 20982 64710 21012 64762
rect 21036 64710 21046 64762
rect 21046 64710 21092 64762
rect 21116 64710 21162 64762
rect 21162 64710 21172 64762
rect 21196 64710 21226 64762
rect 21226 64710 21252 64762
rect 20956 64708 21012 64710
rect 21036 64708 21092 64710
rect 21116 64708 21172 64710
rect 21196 64708 21252 64710
rect 20956 63674 21012 63676
rect 21036 63674 21092 63676
rect 21116 63674 21172 63676
rect 21196 63674 21252 63676
rect 20956 63622 20982 63674
rect 20982 63622 21012 63674
rect 21036 63622 21046 63674
rect 21046 63622 21092 63674
rect 21116 63622 21162 63674
rect 21162 63622 21172 63674
rect 21196 63622 21226 63674
rect 21226 63622 21252 63674
rect 20956 63620 21012 63622
rect 21036 63620 21092 63622
rect 21116 63620 21172 63622
rect 21196 63620 21252 63622
rect 20956 62586 21012 62588
rect 21036 62586 21092 62588
rect 21116 62586 21172 62588
rect 21196 62586 21252 62588
rect 20956 62534 20982 62586
rect 20982 62534 21012 62586
rect 21036 62534 21046 62586
rect 21046 62534 21092 62586
rect 21116 62534 21162 62586
rect 21162 62534 21172 62586
rect 21196 62534 21226 62586
rect 21226 62534 21252 62586
rect 20956 62532 21012 62534
rect 21036 62532 21092 62534
rect 21116 62532 21172 62534
rect 21196 62532 21252 62534
rect 20956 61498 21012 61500
rect 21036 61498 21092 61500
rect 21116 61498 21172 61500
rect 21196 61498 21252 61500
rect 20956 61446 20982 61498
rect 20982 61446 21012 61498
rect 21036 61446 21046 61498
rect 21046 61446 21092 61498
rect 21116 61446 21162 61498
rect 21162 61446 21172 61498
rect 21196 61446 21226 61498
rect 21226 61446 21252 61498
rect 20956 61444 21012 61446
rect 21036 61444 21092 61446
rect 21116 61444 21172 61446
rect 21196 61444 21252 61446
rect 21914 69808 21970 69864
rect 21638 63960 21694 64016
rect 21822 63552 21878 63608
rect 20956 60410 21012 60412
rect 21036 60410 21092 60412
rect 21116 60410 21172 60412
rect 21196 60410 21252 60412
rect 20956 60358 20982 60410
rect 20982 60358 21012 60410
rect 21036 60358 21046 60410
rect 21046 60358 21092 60410
rect 21116 60358 21162 60410
rect 21162 60358 21172 60410
rect 21196 60358 21226 60410
rect 21226 60358 21252 60410
rect 20956 60356 21012 60358
rect 21036 60356 21092 60358
rect 21116 60356 21172 60358
rect 21196 60356 21252 60358
rect 20956 59322 21012 59324
rect 21036 59322 21092 59324
rect 21116 59322 21172 59324
rect 21196 59322 21252 59324
rect 20956 59270 20982 59322
rect 20982 59270 21012 59322
rect 21036 59270 21046 59322
rect 21046 59270 21092 59322
rect 21116 59270 21162 59322
rect 21162 59270 21172 59322
rect 21196 59270 21226 59322
rect 21226 59270 21252 59322
rect 20956 59268 21012 59270
rect 21036 59268 21092 59270
rect 21116 59268 21172 59270
rect 21196 59268 21252 59270
rect 21270 58384 21326 58440
rect 20956 58234 21012 58236
rect 21036 58234 21092 58236
rect 21116 58234 21172 58236
rect 21196 58234 21252 58236
rect 20956 58182 20982 58234
rect 20982 58182 21012 58234
rect 21036 58182 21046 58234
rect 21046 58182 21092 58234
rect 21116 58182 21162 58234
rect 21162 58182 21172 58234
rect 21196 58182 21226 58234
rect 21226 58182 21252 58234
rect 20956 58180 21012 58182
rect 21036 58180 21092 58182
rect 21116 58180 21172 58182
rect 21196 58180 21252 58182
rect 20718 57876 20720 57896
rect 20720 57876 20772 57896
rect 20772 57876 20774 57896
rect 20718 57840 20774 57876
rect 20718 56500 20774 56536
rect 20718 56480 20720 56500
rect 20720 56480 20772 56500
rect 20772 56480 20774 56500
rect 20718 56244 20720 56264
rect 20720 56244 20772 56264
rect 20772 56244 20774 56264
rect 20718 56208 20774 56244
rect 20626 55528 20682 55584
rect 20626 52536 20682 52592
rect 20350 49816 20406 49872
rect 20350 44820 20352 44840
rect 20352 44820 20404 44840
rect 20404 44820 20406 44840
rect 20350 44784 20406 44820
rect 20442 42628 20498 42664
rect 20442 42608 20444 42628
rect 20444 42608 20496 42628
rect 20496 42608 20498 42628
rect 20258 41384 20314 41440
rect 20350 37732 20406 37768
rect 20350 37712 20352 37732
rect 20352 37712 20404 37732
rect 20404 37712 20406 37732
rect 20534 41248 20590 41304
rect 20534 41112 20590 41168
rect 20534 38120 20590 38176
rect 20258 36100 20314 36136
rect 20258 36080 20260 36100
rect 20260 36080 20312 36100
rect 20312 36080 20314 36100
rect 20994 57296 21050 57352
rect 20956 57146 21012 57148
rect 21036 57146 21092 57148
rect 21116 57146 21172 57148
rect 21196 57146 21252 57148
rect 20956 57094 20982 57146
rect 20982 57094 21012 57146
rect 21036 57094 21046 57146
rect 21046 57094 21092 57146
rect 21116 57094 21162 57146
rect 21162 57094 21172 57146
rect 21196 57094 21226 57146
rect 21226 57094 21252 57146
rect 20956 57092 21012 57094
rect 21036 57092 21092 57094
rect 21116 57092 21172 57094
rect 21196 57092 21252 57094
rect 20994 56344 21050 56400
rect 20956 56058 21012 56060
rect 21036 56058 21092 56060
rect 21116 56058 21172 56060
rect 21196 56058 21252 56060
rect 20956 56006 20982 56058
rect 20982 56006 21012 56058
rect 21036 56006 21046 56058
rect 21046 56006 21092 56058
rect 21116 56006 21162 56058
rect 21162 56006 21172 56058
rect 21196 56006 21226 56058
rect 21226 56006 21252 56058
rect 20956 56004 21012 56006
rect 21036 56004 21092 56006
rect 21116 56004 21172 56006
rect 21196 56004 21252 56006
rect 20902 55820 20958 55856
rect 20902 55800 20904 55820
rect 20904 55800 20956 55820
rect 20956 55800 20958 55820
rect 21362 55392 21418 55448
rect 21086 55256 21142 55312
rect 21270 55256 21326 55312
rect 21362 54984 21418 55040
rect 20956 54970 21012 54972
rect 21036 54970 21092 54972
rect 21116 54970 21172 54972
rect 21196 54970 21252 54972
rect 20956 54918 20982 54970
rect 20982 54918 21012 54970
rect 21036 54918 21046 54970
rect 21046 54918 21092 54970
rect 21116 54918 21162 54970
rect 21162 54918 21172 54970
rect 21196 54918 21226 54970
rect 21226 54918 21252 54970
rect 20956 54916 21012 54918
rect 21036 54916 21092 54918
rect 21116 54916 21172 54918
rect 21196 54916 21252 54918
rect 21086 54732 21142 54768
rect 21086 54712 21088 54732
rect 21088 54712 21140 54732
rect 21140 54712 21142 54732
rect 20956 53882 21012 53884
rect 21036 53882 21092 53884
rect 21116 53882 21172 53884
rect 21196 53882 21252 53884
rect 20956 53830 20982 53882
rect 20982 53830 21012 53882
rect 21036 53830 21046 53882
rect 21046 53830 21092 53882
rect 21116 53830 21162 53882
rect 21162 53830 21172 53882
rect 21196 53830 21226 53882
rect 21226 53830 21252 53882
rect 20956 53828 21012 53830
rect 21036 53828 21092 53830
rect 21116 53828 21172 53830
rect 21196 53828 21252 53830
rect 21086 52964 21142 53000
rect 21086 52944 21088 52964
rect 21088 52944 21140 52964
rect 21140 52944 21142 52964
rect 20956 52794 21012 52796
rect 21036 52794 21092 52796
rect 21116 52794 21172 52796
rect 21196 52794 21252 52796
rect 20956 52742 20982 52794
rect 20982 52742 21012 52794
rect 21036 52742 21046 52794
rect 21046 52742 21092 52794
rect 21116 52742 21162 52794
rect 21162 52742 21172 52794
rect 21196 52742 21226 52794
rect 21226 52742 21252 52794
rect 20956 52740 21012 52742
rect 21036 52740 21092 52742
rect 21116 52740 21172 52742
rect 21196 52740 21252 52742
rect 20956 51706 21012 51708
rect 21036 51706 21092 51708
rect 21116 51706 21172 51708
rect 21196 51706 21252 51708
rect 20956 51654 20982 51706
rect 20982 51654 21012 51706
rect 21036 51654 21046 51706
rect 21046 51654 21092 51706
rect 21116 51654 21162 51706
rect 21162 51654 21172 51706
rect 21196 51654 21226 51706
rect 21226 51654 21252 51706
rect 20956 51652 21012 51654
rect 21036 51652 21092 51654
rect 21116 51652 21172 51654
rect 21196 51652 21252 51654
rect 21178 51448 21234 51504
rect 20956 50618 21012 50620
rect 21036 50618 21092 50620
rect 21116 50618 21172 50620
rect 21196 50618 21252 50620
rect 20956 50566 20982 50618
rect 20982 50566 21012 50618
rect 21036 50566 21046 50618
rect 21046 50566 21092 50618
rect 21116 50566 21162 50618
rect 21162 50566 21172 50618
rect 21196 50566 21226 50618
rect 21226 50566 21252 50618
rect 20956 50564 21012 50566
rect 21036 50564 21092 50566
rect 21116 50564 21172 50566
rect 21196 50564 21252 50566
rect 22558 73480 22614 73536
rect 22282 69672 22338 69728
rect 22190 62192 22246 62248
rect 21546 58520 21602 58576
rect 21822 57160 21878 57216
rect 21546 53080 21602 53136
rect 20902 49852 20904 49872
rect 20904 49852 20956 49872
rect 20956 49852 20958 49872
rect 20902 49816 20958 49852
rect 20718 49408 20774 49464
rect 20956 49530 21012 49532
rect 21036 49530 21092 49532
rect 21116 49530 21172 49532
rect 21196 49530 21252 49532
rect 20956 49478 20982 49530
rect 20982 49478 21012 49530
rect 21036 49478 21046 49530
rect 21046 49478 21092 49530
rect 21116 49478 21162 49530
rect 21162 49478 21172 49530
rect 21196 49478 21226 49530
rect 21226 49478 21252 49530
rect 20956 49476 21012 49478
rect 21036 49476 21092 49478
rect 21116 49476 21172 49478
rect 21196 49476 21252 49478
rect 20810 49136 20866 49192
rect 20956 48442 21012 48444
rect 21036 48442 21092 48444
rect 21116 48442 21172 48444
rect 21196 48442 21252 48444
rect 20956 48390 20982 48442
rect 20982 48390 21012 48442
rect 21036 48390 21046 48442
rect 21046 48390 21092 48442
rect 21116 48390 21162 48442
rect 21162 48390 21172 48442
rect 21196 48390 21226 48442
rect 21226 48390 21252 48442
rect 20956 48388 21012 48390
rect 21036 48388 21092 48390
rect 21116 48388 21172 48390
rect 21196 48388 21252 48390
rect 20718 41692 20720 41712
rect 20720 41692 20772 41712
rect 20772 41692 20774 41712
rect 20718 41656 20774 41692
rect 20718 41520 20774 41576
rect 20956 47354 21012 47356
rect 21036 47354 21092 47356
rect 21116 47354 21172 47356
rect 21196 47354 21252 47356
rect 20956 47302 20982 47354
rect 20982 47302 21012 47354
rect 21036 47302 21046 47354
rect 21046 47302 21092 47354
rect 21116 47302 21162 47354
rect 21162 47302 21172 47354
rect 21196 47302 21226 47354
rect 21226 47302 21252 47354
rect 20956 47300 21012 47302
rect 21036 47300 21092 47302
rect 21116 47300 21172 47302
rect 21196 47300 21252 47302
rect 20956 46266 21012 46268
rect 21036 46266 21092 46268
rect 21116 46266 21172 46268
rect 21196 46266 21252 46268
rect 20956 46214 20982 46266
rect 20982 46214 21012 46266
rect 21036 46214 21046 46266
rect 21046 46214 21092 46266
rect 21116 46214 21162 46266
rect 21162 46214 21172 46266
rect 21196 46214 21226 46266
rect 21226 46214 21252 46266
rect 20956 46212 21012 46214
rect 21036 46212 21092 46214
rect 21116 46212 21172 46214
rect 21196 46212 21252 46214
rect 20956 45178 21012 45180
rect 21036 45178 21092 45180
rect 21116 45178 21172 45180
rect 21196 45178 21252 45180
rect 20956 45126 20982 45178
rect 20982 45126 21012 45178
rect 21036 45126 21046 45178
rect 21046 45126 21092 45178
rect 21116 45126 21162 45178
rect 21162 45126 21172 45178
rect 21196 45126 21226 45178
rect 21226 45126 21252 45178
rect 20956 45124 21012 45126
rect 21036 45124 21092 45126
rect 21116 45124 21172 45126
rect 21196 45124 21252 45126
rect 21178 44820 21180 44840
rect 21180 44820 21232 44840
rect 21232 44820 21234 44840
rect 21178 44784 21234 44820
rect 20956 44090 21012 44092
rect 21036 44090 21092 44092
rect 21116 44090 21172 44092
rect 21196 44090 21252 44092
rect 20956 44038 20982 44090
rect 20982 44038 21012 44090
rect 21036 44038 21046 44090
rect 21046 44038 21092 44090
rect 21116 44038 21162 44090
rect 21162 44038 21172 44090
rect 21196 44038 21226 44090
rect 21226 44038 21252 44090
rect 20956 44036 21012 44038
rect 21036 44036 21092 44038
rect 21116 44036 21172 44038
rect 21196 44036 21252 44038
rect 21086 43852 21142 43888
rect 21086 43832 21088 43852
rect 21088 43832 21140 43852
rect 21140 43832 21142 43852
rect 20956 43002 21012 43004
rect 21036 43002 21092 43004
rect 21116 43002 21172 43004
rect 21196 43002 21252 43004
rect 20956 42950 20982 43002
rect 20982 42950 21012 43002
rect 21036 42950 21046 43002
rect 21046 42950 21092 43002
rect 21116 42950 21162 43002
rect 21162 42950 21172 43002
rect 21196 42950 21226 43002
rect 21226 42950 21252 43002
rect 20956 42948 21012 42950
rect 21036 42948 21092 42950
rect 21116 42948 21172 42950
rect 21196 42948 21252 42950
rect 20956 41914 21012 41916
rect 21036 41914 21092 41916
rect 21116 41914 21172 41916
rect 21196 41914 21252 41916
rect 20956 41862 20982 41914
rect 20982 41862 21012 41914
rect 21036 41862 21046 41914
rect 21046 41862 21092 41914
rect 21116 41862 21162 41914
rect 21162 41862 21172 41914
rect 21196 41862 21226 41914
rect 21226 41862 21252 41914
rect 20956 41860 21012 41862
rect 21036 41860 21092 41862
rect 21116 41860 21172 41862
rect 21196 41860 21252 41862
rect 21178 41132 21234 41168
rect 21178 41112 21180 41132
rect 21180 41112 21232 41132
rect 21232 41112 21234 41132
rect 20810 40840 20866 40896
rect 20956 40826 21012 40828
rect 21036 40826 21092 40828
rect 21116 40826 21172 40828
rect 21196 40826 21252 40828
rect 20956 40774 20982 40826
rect 20982 40774 21012 40826
rect 21036 40774 21046 40826
rect 21046 40774 21092 40826
rect 21116 40774 21162 40826
rect 21162 40774 21172 40826
rect 21196 40774 21226 40826
rect 21226 40774 21252 40826
rect 20956 40772 21012 40774
rect 21036 40772 21092 40774
rect 21116 40772 21172 40774
rect 21196 40772 21252 40774
rect 20956 39738 21012 39740
rect 21036 39738 21092 39740
rect 21116 39738 21172 39740
rect 21196 39738 21252 39740
rect 20956 39686 20982 39738
rect 20982 39686 21012 39738
rect 21036 39686 21046 39738
rect 21046 39686 21092 39738
rect 21116 39686 21162 39738
rect 21162 39686 21172 39738
rect 21196 39686 21226 39738
rect 21226 39686 21252 39738
rect 20956 39684 21012 39686
rect 21036 39684 21092 39686
rect 21116 39684 21172 39686
rect 21196 39684 21252 39686
rect 21178 39480 21234 39536
rect 20956 38650 21012 38652
rect 21036 38650 21092 38652
rect 21116 38650 21172 38652
rect 21196 38650 21252 38652
rect 20956 38598 20982 38650
rect 20982 38598 21012 38650
rect 21036 38598 21046 38650
rect 21046 38598 21092 38650
rect 21116 38598 21162 38650
rect 21162 38598 21172 38650
rect 21196 38598 21226 38650
rect 21226 38598 21252 38650
rect 20956 38596 21012 38598
rect 21036 38596 21092 38598
rect 21116 38596 21172 38598
rect 21196 38596 21252 38598
rect 21546 50224 21602 50280
rect 21546 50124 21548 50144
rect 21548 50124 21600 50144
rect 21600 50124 21602 50144
rect 21546 50088 21602 50124
rect 21454 49952 21510 50008
rect 22098 55528 22154 55584
rect 21638 49000 21694 49056
rect 21546 48084 21548 48104
rect 21548 48084 21600 48104
rect 21600 48084 21602 48104
rect 21546 48048 21602 48084
rect 21546 47948 21548 47968
rect 21548 47948 21600 47968
rect 21600 47948 21602 47968
rect 21546 47912 21602 47948
rect 20626 35672 20682 35728
rect 20956 37562 21012 37564
rect 21036 37562 21092 37564
rect 21116 37562 21172 37564
rect 21196 37562 21252 37564
rect 20956 37510 20982 37562
rect 20982 37510 21012 37562
rect 21036 37510 21046 37562
rect 21046 37510 21092 37562
rect 21116 37510 21162 37562
rect 21162 37510 21172 37562
rect 21196 37510 21226 37562
rect 21226 37510 21252 37562
rect 20956 37508 21012 37510
rect 21036 37508 21092 37510
rect 21116 37508 21172 37510
rect 21196 37508 21252 37510
rect 20956 36474 21012 36476
rect 21036 36474 21092 36476
rect 21116 36474 21172 36476
rect 21196 36474 21252 36476
rect 20956 36422 20982 36474
rect 20982 36422 21012 36474
rect 21036 36422 21046 36474
rect 21046 36422 21092 36474
rect 21116 36422 21162 36474
rect 21162 36422 21172 36474
rect 21196 36422 21226 36474
rect 21226 36422 21252 36474
rect 20956 36420 21012 36422
rect 21036 36420 21092 36422
rect 21116 36420 21172 36422
rect 21196 36420 21252 36422
rect 21178 35672 21234 35728
rect 20956 35386 21012 35388
rect 21036 35386 21092 35388
rect 21116 35386 21172 35388
rect 21196 35386 21252 35388
rect 20956 35334 20982 35386
rect 20982 35334 21012 35386
rect 21036 35334 21046 35386
rect 21046 35334 21092 35386
rect 21116 35334 21162 35386
rect 21162 35334 21172 35386
rect 21196 35334 21226 35386
rect 21226 35334 21252 35386
rect 20956 35332 21012 35334
rect 21036 35332 21092 35334
rect 21116 35332 21172 35334
rect 21196 35332 21252 35334
rect 20902 35128 20958 35184
rect 20956 34298 21012 34300
rect 21036 34298 21092 34300
rect 21116 34298 21172 34300
rect 21196 34298 21252 34300
rect 20956 34246 20982 34298
rect 20982 34246 21012 34298
rect 21036 34246 21046 34298
rect 21046 34246 21092 34298
rect 21116 34246 21162 34298
rect 21162 34246 21172 34298
rect 21196 34246 21226 34298
rect 21226 34246 21252 34298
rect 20956 34244 21012 34246
rect 21036 34244 21092 34246
rect 21116 34244 21172 34246
rect 21196 34244 21252 34246
rect 20810 34040 20866 34096
rect 20258 32680 20314 32736
rect 20258 32408 20314 32464
rect 20442 33224 20498 33280
rect 20442 33088 20498 33144
rect 20534 31456 20590 31512
rect 20258 24792 20314 24848
rect 20166 19488 20222 19544
rect 20956 33210 21012 33212
rect 21036 33210 21092 33212
rect 21116 33210 21172 33212
rect 21196 33210 21252 33212
rect 20956 33158 20982 33210
rect 20982 33158 21012 33210
rect 21036 33158 21046 33210
rect 21046 33158 21092 33210
rect 21116 33158 21162 33210
rect 21162 33158 21172 33210
rect 21196 33158 21226 33210
rect 21226 33158 21252 33210
rect 20956 33156 21012 33158
rect 21036 33156 21092 33158
rect 21116 33156 21172 33158
rect 21196 33156 21252 33158
rect 20956 32122 21012 32124
rect 21036 32122 21092 32124
rect 21116 32122 21172 32124
rect 21196 32122 21252 32124
rect 20956 32070 20982 32122
rect 20982 32070 21012 32122
rect 21036 32070 21046 32122
rect 21046 32070 21092 32122
rect 21116 32070 21162 32122
rect 21162 32070 21172 32122
rect 21196 32070 21226 32122
rect 21226 32070 21252 32122
rect 20956 32068 21012 32070
rect 21036 32068 21092 32070
rect 21116 32068 21172 32070
rect 21196 32068 21252 32070
rect 20902 31320 20958 31376
rect 21178 31184 21234 31240
rect 20810 31048 20866 31104
rect 20718 28600 20774 28656
rect 20956 31034 21012 31036
rect 21036 31034 21092 31036
rect 21116 31034 21172 31036
rect 21196 31034 21252 31036
rect 20956 30982 20982 31034
rect 20982 30982 21012 31034
rect 21036 30982 21046 31034
rect 21046 30982 21092 31034
rect 21116 30982 21162 31034
rect 21162 30982 21172 31034
rect 21196 30982 21226 31034
rect 21226 30982 21252 31034
rect 20956 30980 21012 30982
rect 21036 30980 21092 30982
rect 21116 30980 21172 30982
rect 21196 30980 21252 30982
rect 20902 30796 20958 30832
rect 20902 30776 20904 30796
rect 20904 30776 20956 30796
rect 20956 30776 20958 30796
rect 21086 30660 21142 30696
rect 21086 30640 21088 30660
rect 21088 30640 21140 30660
rect 21140 30640 21142 30660
rect 20956 29946 21012 29948
rect 21036 29946 21092 29948
rect 21116 29946 21172 29948
rect 21196 29946 21252 29948
rect 20956 29894 20982 29946
rect 20982 29894 21012 29946
rect 21036 29894 21046 29946
rect 21046 29894 21092 29946
rect 21116 29894 21162 29946
rect 21162 29894 21172 29946
rect 21196 29894 21226 29946
rect 21226 29894 21252 29946
rect 20956 29892 21012 29894
rect 21036 29892 21092 29894
rect 21116 29892 21172 29894
rect 21196 29892 21252 29894
rect 20994 29416 21050 29472
rect 20956 28858 21012 28860
rect 21036 28858 21092 28860
rect 21116 28858 21172 28860
rect 21196 28858 21252 28860
rect 20956 28806 20982 28858
rect 20982 28806 21012 28858
rect 21036 28806 21046 28858
rect 21046 28806 21092 28858
rect 21116 28806 21162 28858
rect 21162 28806 21172 28858
rect 21196 28806 21226 28858
rect 21226 28806 21252 28858
rect 20956 28804 21012 28806
rect 21036 28804 21092 28806
rect 21116 28804 21172 28806
rect 21196 28804 21252 28806
rect 20956 27770 21012 27772
rect 21036 27770 21092 27772
rect 21116 27770 21172 27772
rect 21196 27770 21252 27772
rect 20956 27718 20982 27770
rect 20982 27718 21012 27770
rect 21036 27718 21046 27770
rect 21046 27718 21092 27770
rect 21116 27718 21162 27770
rect 21162 27718 21172 27770
rect 21196 27718 21226 27770
rect 21226 27718 21252 27770
rect 20956 27716 21012 27718
rect 21036 27716 21092 27718
rect 21116 27716 21172 27718
rect 21196 27716 21252 27718
rect 18602 1944 18658 2000
rect 20956 26682 21012 26684
rect 21036 26682 21092 26684
rect 21116 26682 21172 26684
rect 21196 26682 21252 26684
rect 20956 26630 20982 26682
rect 20982 26630 21012 26682
rect 21036 26630 21046 26682
rect 21046 26630 21092 26682
rect 21116 26630 21162 26682
rect 21162 26630 21172 26682
rect 21196 26630 21226 26682
rect 21226 26630 21252 26682
rect 20956 26628 21012 26630
rect 21036 26628 21092 26630
rect 21116 26628 21172 26630
rect 21196 26628 21252 26630
rect 20956 25594 21012 25596
rect 21036 25594 21092 25596
rect 21116 25594 21172 25596
rect 21196 25594 21252 25596
rect 20956 25542 20982 25594
rect 20982 25542 21012 25594
rect 21036 25542 21046 25594
rect 21046 25542 21092 25594
rect 21116 25542 21162 25594
rect 21162 25542 21172 25594
rect 21196 25542 21226 25594
rect 21226 25542 21252 25594
rect 20956 25540 21012 25542
rect 21036 25540 21092 25542
rect 21116 25540 21172 25542
rect 21196 25540 21252 25542
rect 20956 24506 21012 24508
rect 21036 24506 21092 24508
rect 21116 24506 21172 24508
rect 21196 24506 21252 24508
rect 20956 24454 20982 24506
rect 20982 24454 21012 24506
rect 21036 24454 21046 24506
rect 21046 24454 21092 24506
rect 21116 24454 21162 24506
rect 21162 24454 21172 24506
rect 21196 24454 21226 24506
rect 21226 24454 21252 24506
rect 20956 24452 21012 24454
rect 21036 24452 21092 24454
rect 21116 24452 21172 24454
rect 21196 24452 21252 24454
rect 20956 23418 21012 23420
rect 21036 23418 21092 23420
rect 21116 23418 21172 23420
rect 21196 23418 21252 23420
rect 20956 23366 20982 23418
rect 20982 23366 21012 23418
rect 21036 23366 21046 23418
rect 21046 23366 21092 23418
rect 21116 23366 21162 23418
rect 21162 23366 21172 23418
rect 21196 23366 21226 23418
rect 21226 23366 21252 23418
rect 20956 23364 21012 23366
rect 21036 23364 21092 23366
rect 21116 23364 21172 23366
rect 21196 23364 21252 23366
rect 20956 22330 21012 22332
rect 21036 22330 21092 22332
rect 21116 22330 21172 22332
rect 21196 22330 21252 22332
rect 20956 22278 20982 22330
rect 20982 22278 21012 22330
rect 21036 22278 21046 22330
rect 21046 22278 21092 22330
rect 21116 22278 21162 22330
rect 21162 22278 21172 22330
rect 21196 22278 21226 22330
rect 21226 22278 21252 22330
rect 20956 22276 21012 22278
rect 21036 22276 21092 22278
rect 21116 22276 21172 22278
rect 21196 22276 21252 22278
rect 20956 21242 21012 21244
rect 21036 21242 21092 21244
rect 21116 21242 21172 21244
rect 21196 21242 21252 21244
rect 20956 21190 20982 21242
rect 20982 21190 21012 21242
rect 21036 21190 21046 21242
rect 21046 21190 21092 21242
rect 21116 21190 21162 21242
rect 21162 21190 21172 21242
rect 21196 21190 21226 21242
rect 21226 21190 21252 21242
rect 20956 21188 21012 21190
rect 21036 21188 21092 21190
rect 21116 21188 21172 21190
rect 21196 21188 21252 21190
rect 20956 20154 21012 20156
rect 21036 20154 21092 20156
rect 21116 20154 21172 20156
rect 21196 20154 21252 20156
rect 20956 20102 20982 20154
rect 20982 20102 21012 20154
rect 21036 20102 21046 20154
rect 21046 20102 21092 20154
rect 21116 20102 21162 20154
rect 21162 20102 21172 20154
rect 21196 20102 21226 20154
rect 21226 20102 21252 20154
rect 20956 20100 21012 20102
rect 21036 20100 21092 20102
rect 21116 20100 21172 20102
rect 21196 20100 21252 20102
rect 21178 19488 21234 19544
rect 20956 19066 21012 19068
rect 21036 19066 21092 19068
rect 21116 19066 21172 19068
rect 21196 19066 21252 19068
rect 20956 19014 20982 19066
rect 20982 19014 21012 19066
rect 21036 19014 21046 19066
rect 21046 19014 21092 19066
rect 21116 19014 21162 19066
rect 21162 19014 21172 19066
rect 21196 19014 21226 19066
rect 21226 19014 21252 19066
rect 20956 19012 21012 19014
rect 21036 19012 21092 19014
rect 21116 19012 21172 19014
rect 21196 19012 21252 19014
rect 20956 17978 21012 17980
rect 21036 17978 21092 17980
rect 21116 17978 21172 17980
rect 21196 17978 21252 17980
rect 20956 17926 20982 17978
rect 20982 17926 21012 17978
rect 21036 17926 21046 17978
rect 21046 17926 21092 17978
rect 21116 17926 21162 17978
rect 21162 17926 21172 17978
rect 21196 17926 21226 17978
rect 21226 17926 21252 17978
rect 20956 17924 21012 17926
rect 21036 17924 21092 17926
rect 21116 17924 21172 17926
rect 21196 17924 21252 17926
rect 20956 16890 21012 16892
rect 21036 16890 21092 16892
rect 21116 16890 21172 16892
rect 21196 16890 21252 16892
rect 20956 16838 20982 16890
rect 20982 16838 21012 16890
rect 21036 16838 21046 16890
rect 21046 16838 21092 16890
rect 21116 16838 21162 16890
rect 21162 16838 21172 16890
rect 21196 16838 21226 16890
rect 21226 16838 21252 16890
rect 20956 16836 21012 16838
rect 21036 16836 21092 16838
rect 21116 16836 21172 16838
rect 21196 16836 21252 16838
rect 20956 15802 21012 15804
rect 21036 15802 21092 15804
rect 21116 15802 21172 15804
rect 21196 15802 21252 15804
rect 20956 15750 20982 15802
rect 20982 15750 21012 15802
rect 21036 15750 21046 15802
rect 21046 15750 21092 15802
rect 21116 15750 21162 15802
rect 21162 15750 21172 15802
rect 21196 15750 21226 15802
rect 21226 15750 21252 15802
rect 20956 15748 21012 15750
rect 21036 15748 21092 15750
rect 21116 15748 21172 15750
rect 21196 15748 21252 15750
rect 20956 14714 21012 14716
rect 21036 14714 21092 14716
rect 21116 14714 21172 14716
rect 21196 14714 21252 14716
rect 20956 14662 20982 14714
rect 20982 14662 21012 14714
rect 21036 14662 21046 14714
rect 21046 14662 21092 14714
rect 21116 14662 21162 14714
rect 21162 14662 21172 14714
rect 21196 14662 21226 14714
rect 21226 14662 21252 14714
rect 20956 14660 21012 14662
rect 21036 14660 21092 14662
rect 21116 14660 21172 14662
rect 21196 14660 21252 14662
rect 20956 13626 21012 13628
rect 21036 13626 21092 13628
rect 21116 13626 21172 13628
rect 21196 13626 21252 13628
rect 20956 13574 20982 13626
rect 20982 13574 21012 13626
rect 21036 13574 21046 13626
rect 21046 13574 21092 13626
rect 21116 13574 21162 13626
rect 21162 13574 21172 13626
rect 21196 13574 21226 13626
rect 21226 13574 21252 13626
rect 20956 13572 21012 13574
rect 21036 13572 21092 13574
rect 21116 13572 21172 13574
rect 21196 13572 21252 13574
rect 20956 12538 21012 12540
rect 21036 12538 21092 12540
rect 21116 12538 21172 12540
rect 21196 12538 21252 12540
rect 20956 12486 20982 12538
rect 20982 12486 21012 12538
rect 21036 12486 21046 12538
rect 21046 12486 21092 12538
rect 21116 12486 21162 12538
rect 21162 12486 21172 12538
rect 21196 12486 21226 12538
rect 21226 12486 21252 12538
rect 20956 12484 21012 12486
rect 21036 12484 21092 12486
rect 21116 12484 21172 12486
rect 21196 12484 21252 12486
rect 20956 11450 21012 11452
rect 21036 11450 21092 11452
rect 21116 11450 21172 11452
rect 21196 11450 21252 11452
rect 20956 11398 20982 11450
rect 20982 11398 21012 11450
rect 21036 11398 21046 11450
rect 21046 11398 21092 11450
rect 21116 11398 21162 11450
rect 21162 11398 21172 11450
rect 21196 11398 21226 11450
rect 21226 11398 21252 11450
rect 20956 11396 21012 11398
rect 21036 11396 21092 11398
rect 21116 11396 21172 11398
rect 21196 11396 21252 11398
rect 22190 54068 22192 54088
rect 22192 54068 22244 54088
rect 22244 54068 22246 54088
rect 22190 54032 22246 54068
rect 22006 50788 22062 50824
rect 22006 50768 22008 50788
rect 22008 50768 22060 50788
rect 22060 50768 22062 50788
rect 23662 74704 23718 74760
rect 23110 74296 23166 74352
rect 23202 73752 23258 73808
rect 22926 62328 22982 62384
rect 22742 61784 22798 61840
rect 22650 59064 22706 59120
rect 22558 57740 22560 57760
rect 22560 57740 22612 57760
rect 22612 57740 22614 57760
rect 22558 57704 22614 57740
rect 22466 56480 22522 56536
rect 22742 54984 22798 55040
rect 22466 53624 22522 53680
rect 22006 50396 22008 50416
rect 22008 50396 22060 50416
rect 22060 50396 22062 50416
rect 22006 50360 22062 50396
rect 22006 50260 22008 50280
rect 22008 50260 22060 50280
rect 22060 50260 22062 50280
rect 22006 50224 22062 50260
rect 22006 49680 22062 49736
rect 22190 49816 22246 49872
rect 22006 49000 22062 49056
rect 21822 48456 21878 48512
rect 21730 46588 21732 46608
rect 21732 46588 21784 46608
rect 21784 46588 21786 46608
rect 21730 46552 21786 46588
rect 21822 46144 21878 46200
rect 21730 46008 21786 46064
rect 21546 41112 21602 41168
rect 21546 39888 21602 39944
rect 22926 51176 22982 51232
rect 22282 48184 22338 48240
rect 22190 48048 22246 48104
rect 22650 48204 22706 48240
rect 22650 48184 22652 48204
rect 22652 48184 22704 48204
rect 22704 48184 22706 48204
rect 22742 47912 22798 47968
rect 22374 46824 22430 46880
rect 22190 46144 22246 46200
rect 22190 43424 22246 43480
rect 22650 44512 22706 44568
rect 22282 42764 22338 42800
rect 22282 42744 22284 42764
rect 22284 42744 22336 42764
rect 22336 42744 22338 42764
rect 21914 41248 21970 41304
rect 21822 40704 21878 40760
rect 21546 37304 21602 37360
rect 21730 38800 21786 38856
rect 21546 35808 21602 35864
rect 21914 38664 21970 38720
rect 21638 34176 21694 34232
rect 21638 33360 21694 33416
rect 21822 36352 21878 36408
rect 23202 51312 23258 51368
rect 23294 50768 23350 50824
rect 23110 47796 23166 47832
rect 23110 47776 23112 47796
rect 23112 47776 23164 47796
rect 23164 47776 23166 47796
rect 23018 46688 23074 46744
rect 23294 47232 23350 47288
rect 22926 43560 22982 43616
rect 22834 43016 22890 43072
rect 23110 45872 23166 45928
rect 23294 45328 23350 45384
rect 23294 45076 23350 45112
rect 23294 45056 23296 45076
rect 23296 45056 23348 45076
rect 23348 45056 23350 45076
rect 23110 43968 23166 44024
rect 22926 41656 22982 41712
rect 22374 37032 22430 37088
rect 22006 35148 22062 35184
rect 22006 35128 22008 35148
rect 22008 35128 22060 35148
rect 22060 35128 22062 35148
rect 22190 34584 22246 34640
rect 21822 33632 21878 33688
rect 21822 33224 21878 33280
rect 21730 32680 21786 32736
rect 22006 32408 22062 32464
rect 21638 28872 21694 28928
rect 21638 25744 21694 25800
rect 21730 23704 21786 23760
rect 21730 20576 21786 20632
rect 21454 20168 21510 20224
rect 21638 13640 21694 13696
rect 20956 10362 21012 10364
rect 21036 10362 21092 10364
rect 21116 10362 21172 10364
rect 21196 10362 21252 10364
rect 20956 10310 20982 10362
rect 20982 10310 21012 10362
rect 21036 10310 21046 10362
rect 21046 10310 21092 10362
rect 21116 10310 21162 10362
rect 21162 10310 21172 10362
rect 21196 10310 21226 10362
rect 21226 10310 21252 10362
rect 20956 10308 21012 10310
rect 21036 10308 21092 10310
rect 21116 10308 21172 10310
rect 21196 10308 21252 10310
rect 20956 9274 21012 9276
rect 21036 9274 21092 9276
rect 21116 9274 21172 9276
rect 21196 9274 21252 9276
rect 20956 9222 20982 9274
rect 20982 9222 21012 9274
rect 21036 9222 21046 9274
rect 21046 9222 21092 9274
rect 21116 9222 21162 9274
rect 21162 9222 21172 9274
rect 21196 9222 21226 9274
rect 21226 9222 21252 9274
rect 20956 9220 21012 9222
rect 21036 9220 21092 9222
rect 21116 9220 21172 9222
rect 21196 9220 21252 9222
rect 20956 8186 21012 8188
rect 21036 8186 21092 8188
rect 21116 8186 21172 8188
rect 21196 8186 21252 8188
rect 20956 8134 20982 8186
rect 20982 8134 21012 8186
rect 21036 8134 21046 8186
rect 21046 8134 21092 8186
rect 21116 8134 21162 8186
rect 21162 8134 21172 8186
rect 21196 8134 21226 8186
rect 21226 8134 21252 8186
rect 20956 8132 21012 8134
rect 21036 8132 21092 8134
rect 21116 8132 21172 8134
rect 21196 8132 21252 8134
rect 20956 7098 21012 7100
rect 21036 7098 21092 7100
rect 21116 7098 21172 7100
rect 21196 7098 21252 7100
rect 20956 7046 20982 7098
rect 20982 7046 21012 7098
rect 21036 7046 21046 7098
rect 21046 7046 21092 7098
rect 21116 7046 21162 7098
rect 21162 7046 21172 7098
rect 21196 7046 21226 7098
rect 21226 7046 21252 7098
rect 20956 7044 21012 7046
rect 21036 7044 21092 7046
rect 21116 7044 21172 7046
rect 21196 7044 21252 7046
rect 20956 6010 21012 6012
rect 21036 6010 21092 6012
rect 21116 6010 21172 6012
rect 21196 6010 21252 6012
rect 20956 5958 20982 6010
rect 20982 5958 21012 6010
rect 21036 5958 21046 6010
rect 21046 5958 21092 6010
rect 21116 5958 21162 6010
rect 21162 5958 21172 6010
rect 21196 5958 21226 6010
rect 21226 5958 21252 6010
rect 20956 5956 21012 5958
rect 21036 5956 21092 5958
rect 21116 5956 21172 5958
rect 21196 5956 21252 5958
rect 20956 4922 21012 4924
rect 21036 4922 21092 4924
rect 21116 4922 21172 4924
rect 21196 4922 21252 4924
rect 20956 4870 20982 4922
rect 20982 4870 21012 4922
rect 21036 4870 21046 4922
rect 21046 4870 21092 4922
rect 21116 4870 21162 4922
rect 21162 4870 21172 4922
rect 21196 4870 21226 4922
rect 21226 4870 21252 4922
rect 20956 4868 21012 4870
rect 21036 4868 21092 4870
rect 21116 4868 21172 4870
rect 21196 4868 21252 4870
rect 21454 4800 21510 4856
rect 20956 3834 21012 3836
rect 21036 3834 21092 3836
rect 21116 3834 21172 3836
rect 21196 3834 21252 3836
rect 20956 3782 20982 3834
rect 20982 3782 21012 3834
rect 21036 3782 21046 3834
rect 21046 3782 21092 3834
rect 21116 3782 21162 3834
rect 21162 3782 21172 3834
rect 21196 3782 21226 3834
rect 21226 3782 21252 3834
rect 20956 3780 21012 3782
rect 21036 3780 21092 3782
rect 21116 3780 21172 3782
rect 21196 3780 21252 3782
rect 21730 10240 21786 10296
rect 21914 19216 21970 19272
rect 21822 8336 21878 8392
rect 21638 3576 21694 3632
rect 22558 35536 22614 35592
rect 22466 34720 22522 34776
rect 22374 33768 22430 33824
rect 22558 33516 22614 33552
rect 22558 33496 22560 33516
rect 22560 33496 22612 33516
rect 22612 33496 22614 33516
rect 22282 32852 22284 32872
rect 22284 32852 22336 32872
rect 22336 32852 22338 32872
rect 22282 32816 22338 32852
rect 22742 37324 22798 37360
rect 22742 37304 22744 37324
rect 22744 37304 22796 37324
rect 22796 37304 22798 37324
rect 22834 35436 22836 35456
rect 22836 35436 22888 35456
rect 22888 35436 22890 35456
rect 22834 35400 22890 35436
rect 22742 32952 22798 33008
rect 22650 29960 22706 30016
rect 22282 20576 22338 20632
rect 22006 13912 22062 13968
rect 22006 6160 22062 6216
rect 22466 15272 22522 15328
rect 22558 14320 22614 14376
rect 22742 13640 22798 13696
rect 22558 11736 22614 11792
rect 22374 3984 22430 4040
rect 20956 2746 21012 2748
rect 21036 2746 21092 2748
rect 21116 2746 21172 2748
rect 21196 2746 21252 2748
rect 20956 2694 20982 2746
rect 20982 2694 21012 2746
rect 21036 2694 21046 2746
rect 21046 2694 21092 2746
rect 21116 2694 21162 2746
rect 21162 2694 21172 2746
rect 21196 2694 21226 2746
rect 21226 2694 21252 2746
rect 20956 2692 21012 2694
rect 21036 2692 21092 2694
rect 21116 2692 21172 2694
rect 21196 2692 21252 2694
rect 20902 2372 20958 2408
rect 20902 2352 20904 2372
rect 20904 2352 20956 2372
rect 20956 2352 20958 2372
rect 20534 856 20590 912
rect 20718 856 20774 912
rect 23202 41656 23258 41712
rect 23202 41384 23258 41440
rect 23478 59084 23534 59120
rect 23478 59064 23480 59084
rect 23480 59064 23532 59084
rect 23532 59064 23534 59084
rect 23938 74432 23994 74488
rect 24398 74296 24454 74352
rect 24490 68992 24546 69048
rect 23938 58384 23994 58440
rect 23478 54032 23534 54088
rect 23754 52420 23810 52456
rect 23754 52400 23756 52420
rect 23756 52400 23808 52420
rect 23808 52400 23810 52420
rect 23662 51448 23718 51504
rect 23570 50904 23626 50960
rect 23570 50632 23626 50688
rect 23754 50632 23810 50688
rect 23570 48048 23626 48104
rect 23478 46588 23480 46608
rect 23480 46588 23532 46608
rect 23532 46588 23534 46608
rect 23478 46552 23534 46588
rect 24214 52264 24270 52320
rect 24030 48456 24086 48512
rect 23570 44376 23626 44432
rect 23478 43324 23480 43344
rect 23480 43324 23532 43344
rect 23532 43324 23534 43344
rect 23478 43288 23534 43324
rect 23662 42200 23718 42256
rect 23478 39908 23534 39944
rect 23478 39888 23480 39908
rect 23480 39888 23532 39908
rect 23532 39888 23534 39908
rect 23846 44920 23902 44976
rect 24122 47640 24178 47696
rect 24122 46028 24178 46064
rect 24122 46008 24124 46028
rect 24124 46008 24176 46028
rect 24176 46008 24178 46028
rect 23662 38412 23718 38448
rect 23662 38392 23664 38412
rect 23664 38392 23716 38412
rect 23716 38392 23718 38412
rect 24582 59336 24638 59392
rect 25870 78240 25926 78296
rect 25956 77274 26012 77276
rect 26036 77274 26092 77276
rect 26116 77274 26172 77276
rect 26196 77274 26252 77276
rect 25956 77222 25982 77274
rect 25982 77222 26012 77274
rect 26036 77222 26046 77274
rect 26046 77222 26092 77274
rect 26116 77222 26162 77274
rect 26162 77222 26172 77274
rect 26196 77222 26226 77274
rect 26226 77222 26252 77274
rect 25956 77220 26012 77222
rect 26036 77220 26092 77222
rect 26116 77220 26172 77222
rect 26196 77220 26252 77222
rect 25134 76336 25190 76392
rect 25042 75928 25098 75984
rect 24858 74568 24914 74624
rect 25226 74840 25282 74896
rect 25778 76880 25834 76936
rect 25686 74704 25742 74760
rect 25502 70080 25558 70136
rect 25226 68992 25282 69048
rect 25134 68856 25190 68912
rect 25502 67768 25558 67824
rect 25502 66680 25558 66736
rect 25956 76186 26012 76188
rect 26036 76186 26092 76188
rect 26116 76186 26172 76188
rect 26196 76186 26252 76188
rect 25956 76134 25982 76186
rect 25982 76134 26012 76186
rect 26036 76134 26046 76186
rect 26046 76134 26092 76186
rect 26116 76134 26162 76186
rect 26162 76134 26172 76186
rect 26196 76134 26226 76186
rect 26226 76134 26252 76186
rect 25956 76132 26012 76134
rect 26036 76132 26092 76134
rect 26116 76132 26172 76134
rect 26196 76132 26252 76134
rect 26698 75248 26754 75304
rect 25956 75098 26012 75100
rect 26036 75098 26092 75100
rect 26116 75098 26172 75100
rect 26196 75098 26252 75100
rect 25956 75046 25982 75098
rect 25982 75046 26012 75098
rect 26036 75046 26046 75098
rect 26046 75046 26092 75098
rect 26116 75046 26162 75098
rect 26162 75046 26172 75098
rect 26196 75046 26226 75098
rect 26226 75046 26252 75098
rect 25956 75044 26012 75046
rect 26036 75044 26092 75046
rect 26116 75044 26172 75046
rect 26196 75044 26252 75046
rect 25956 74010 26012 74012
rect 26036 74010 26092 74012
rect 26116 74010 26172 74012
rect 26196 74010 26252 74012
rect 25956 73958 25982 74010
rect 25982 73958 26012 74010
rect 26036 73958 26046 74010
rect 26046 73958 26092 74010
rect 26116 73958 26162 74010
rect 26162 73958 26172 74010
rect 26196 73958 26226 74010
rect 26226 73958 26252 74010
rect 25956 73956 26012 73958
rect 26036 73956 26092 73958
rect 26116 73956 26172 73958
rect 26196 73956 26252 73958
rect 25956 72922 26012 72924
rect 26036 72922 26092 72924
rect 26116 72922 26172 72924
rect 26196 72922 26252 72924
rect 25956 72870 25982 72922
rect 25982 72870 26012 72922
rect 26036 72870 26046 72922
rect 26046 72870 26092 72922
rect 26116 72870 26162 72922
rect 26162 72870 26172 72922
rect 26196 72870 26226 72922
rect 26226 72870 26252 72922
rect 25956 72868 26012 72870
rect 26036 72868 26092 72870
rect 26116 72868 26172 72870
rect 26196 72868 26252 72870
rect 25956 71834 26012 71836
rect 26036 71834 26092 71836
rect 26116 71834 26172 71836
rect 26196 71834 26252 71836
rect 25956 71782 25982 71834
rect 25982 71782 26012 71834
rect 26036 71782 26046 71834
rect 26046 71782 26092 71834
rect 26116 71782 26162 71834
rect 26162 71782 26172 71834
rect 26196 71782 26226 71834
rect 26226 71782 26252 71834
rect 25956 71780 26012 71782
rect 26036 71780 26092 71782
rect 26116 71780 26172 71782
rect 26196 71780 26252 71782
rect 26422 71712 26478 71768
rect 25956 70746 26012 70748
rect 26036 70746 26092 70748
rect 26116 70746 26172 70748
rect 26196 70746 26252 70748
rect 25956 70694 25982 70746
rect 25982 70694 26012 70746
rect 26036 70694 26046 70746
rect 26046 70694 26092 70746
rect 26116 70694 26162 70746
rect 26162 70694 26172 70746
rect 26196 70694 26226 70746
rect 26226 70694 26252 70746
rect 25956 70692 26012 70694
rect 26036 70692 26092 70694
rect 26116 70692 26172 70694
rect 26196 70692 26252 70694
rect 25956 69658 26012 69660
rect 26036 69658 26092 69660
rect 26116 69658 26172 69660
rect 26196 69658 26252 69660
rect 25956 69606 25982 69658
rect 25982 69606 26012 69658
rect 26036 69606 26046 69658
rect 26046 69606 26092 69658
rect 26116 69606 26162 69658
rect 26162 69606 26172 69658
rect 26196 69606 26226 69658
rect 26226 69606 26252 69658
rect 25956 69604 26012 69606
rect 26036 69604 26092 69606
rect 26116 69604 26172 69606
rect 26196 69604 26252 69606
rect 25956 68570 26012 68572
rect 26036 68570 26092 68572
rect 26116 68570 26172 68572
rect 26196 68570 26252 68572
rect 25956 68518 25982 68570
rect 25982 68518 26012 68570
rect 26036 68518 26046 68570
rect 26046 68518 26092 68570
rect 26116 68518 26162 68570
rect 26162 68518 26172 68570
rect 26196 68518 26226 68570
rect 26226 68518 26252 68570
rect 25956 68516 26012 68518
rect 26036 68516 26092 68518
rect 26116 68516 26172 68518
rect 26196 68516 26252 68518
rect 25956 67482 26012 67484
rect 26036 67482 26092 67484
rect 26116 67482 26172 67484
rect 26196 67482 26252 67484
rect 25956 67430 25982 67482
rect 25982 67430 26012 67482
rect 26036 67430 26046 67482
rect 26046 67430 26092 67482
rect 26116 67430 26162 67482
rect 26162 67430 26172 67482
rect 26196 67430 26226 67482
rect 26226 67430 26252 67482
rect 25956 67428 26012 67430
rect 26036 67428 26092 67430
rect 26116 67428 26172 67430
rect 26196 67428 26252 67430
rect 25956 66394 26012 66396
rect 26036 66394 26092 66396
rect 26116 66394 26172 66396
rect 26196 66394 26252 66396
rect 25956 66342 25982 66394
rect 25982 66342 26012 66394
rect 26036 66342 26046 66394
rect 26046 66342 26092 66394
rect 26116 66342 26162 66394
rect 26162 66342 26172 66394
rect 26196 66342 26226 66394
rect 26226 66342 26252 66394
rect 25956 66340 26012 66342
rect 26036 66340 26092 66342
rect 26116 66340 26172 66342
rect 26196 66340 26252 66342
rect 25956 65306 26012 65308
rect 26036 65306 26092 65308
rect 26116 65306 26172 65308
rect 26196 65306 26252 65308
rect 25956 65254 25982 65306
rect 25982 65254 26012 65306
rect 26036 65254 26046 65306
rect 26046 65254 26092 65306
rect 26116 65254 26162 65306
rect 26162 65254 26172 65306
rect 26196 65254 26226 65306
rect 26226 65254 26252 65306
rect 25956 65252 26012 65254
rect 26036 65252 26092 65254
rect 26116 65252 26172 65254
rect 26196 65252 26252 65254
rect 25594 65048 25650 65104
rect 25870 64640 25926 64696
rect 25778 63280 25834 63336
rect 25594 62872 25650 62928
rect 25594 61784 25650 61840
rect 24950 61240 25006 61296
rect 24490 53100 24546 53136
rect 24490 53080 24492 53100
rect 24492 53080 24544 53100
rect 24544 53080 24546 53100
rect 24306 47232 24362 47288
rect 24490 47096 24546 47152
rect 23570 34176 23626 34232
rect 23386 34060 23442 34096
rect 23386 34040 23388 34060
rect 23388 34040 23440 34060
rect 23440 34040 23442 34060
rect 22926 31220 22928 31240
rect 22928 31220 22980 31240
rect 22980 31220 22982 31240
rect 22926 31184 22982 31220
rect 23754 33224 23810 33280
rect 22926 21120 22982 21176
rect 23938 37032 23994 37088
rect 23938 36080 23994 36136
rect 23938 31340 23994 31376
rect 23938 31320 23940 31340
rect 23940 31320 23992 31340
rect 23992 31320 23994 31340
rect 23846 23160 23902 23216
rect 24122 28600 24178 28656
rect 23754 20748 23756 20768
rect 23756 20748 23808 20768
rect 23808 20748 23810 20768
rect 23754 20712 23810 20748
rect 24030 20712 24086 20768
rect 24490 43696 24546 43752
rect 24858 47948 24860 47968
rect 24860 47948 24912 47968
rect 24912 47948 24914 47968
rect 24858 47912 24914 47948
rect 24674 43832 24730 43888
rect 24306 41792 24362 41848
rect 24674 41792 24730 41848
rect 24306 40840 24362 40896
rect 24306 35128 24362 35184
rect 24306 34720 24362 34776
rect 24214 19216 24270 19272
rect 22834 10648 22890 10704
rect 24582 41384 24638 41440
rect 24490 39092 24546 39128
rect 24490 39072 24492 39092
rect 24492 39072 24544 39092
rect 24544 39072 24546 39092
rect 24766 38256 24822 38312
rect 24398 6840 24454 6896
rect 25042 55120 25098 55176
rect 25410 53760 25466 53816
rect 25318 52400 25374 52456
rect 25226 51584 25282 51640
rect 25226 50360 25282 50416
rect 25226 48728 25282 48784
rect 25134 48220 25136 48240
rect 25136 48220 25188 48240
rect 25188 48220 25190 48240
rect 25134 48184 25190 48220
rect 25410 50224 25466 50280
rect 25134 45600 25190 45656
rect 25134 45348 25190 45384
rect 25134 45328 25136 45348
rect 25136 45328 25188 45348
rect 25188 45328 25190 45348
rect 25042 44512 25098 44568
rect 25134 43696 25190 43752
rect 25042 41792 25098 41848
rect 25134 35400 25190 35456
rect 25042 34040 25098 34096
rect 24950 32000 25006 32056
rect 24950 30232 25006 30288
rect 25134 27614 25190 27670
rect 25042 26016 25098 26072
rect 25410 44784 25466 44840
rect 25318 44512 25374 44568
rect 25410 43016 25466 43072
rect 25410 41928 25466 41984
rect 25956 64218 26012 64220
rect 26036 64218 26092 64220
rect 26116 64218 26172 64220
rect 26196 64218 26252 64220
rect 25956 64166 25982 64218
rect 25982 64166 26012 64218
rect 26036 64166 26046 64218
rect 26046 64166 26092 64218
rect 26116 64166 26162 64218
rect 26162 64166 26172 64218
rect 26196 64166 26226 64218
rect 26226 64166 26252 64218
rect 25956 64164 26012 64166
rect 26036 64164 26092 64166
rect 26116 64164 26172 64166
rect 26196 64164 26252 64166
rect 27526 63552 27582 63608
rect 25956 63130 26012 63132
rect 26036 63130 26092 63132
rect 26116 63130 26172 63132
rect 26196 63130 26252 63132
rect 25956 63078 25982 63130
rect 25982 63078 26012 63130
rect 26036 63078 26046 63130
rect 26046 63078 26092 63130
rect 26116 63078 26162 63130
rect 26162 63078 26172 63130
rect 26196 63078 26226 63130
rect 26226 63078 26252 63130
rect 25956 63076 26012 63078
rect 26036 63076 26092 63078
rect 26116 63076 26172 63078
rect 26196 63076 26252 63078
rect 29918 72528 29974 72584
rect 25956 62042 26012 62044
rect 26036 62042 26092 62044
rect 26116 62042 26172 62044
rect 26196 62042 26252 62044
rect 25956 61990 25982 62042
rect 25982 61990 26012 62042
rect 26036 61990 26046 62042
rect 26046 61990 26092 62042
rect 26116 61990 26162 62042
rect 26162 61990 26172 62042
rect 26196 61990 26226 62042
rect 26226 61990 26252 62042
rect 25956 61988 26012 61990
rect 26036 61988 26092 61990
rect 26116 61988 26172 61990
rect 26196 61988 26252 61990
rect 26698 61920 26754 61976
rect 25778 59608 25834 59664
rect 25956 60954 26012 60956
rect 26036 60954 26092 60956
rect 26116 60954 26172 60956
rect 26196 60954 26252 60956
rect 25956 60902 25982 60954
rect 25982 60902 26012 60954
rect 26036 60902 26046 60954
rect 26046 60902 26092 60954
rect 26116 60902 26162 60954
rect 26162 60902 26172 60954
rect 26196 60902 26226 60954
rect 26226 60902 26252 60954
rect 25956 60900 26012 60902
rect 26036 60900 26092 60902
rect 26116 60900 26172 60902
rect 26196 60900 26252 60902
rect 25956 59866 26012 59868
rect 26036 59866 26092 59868
rect 26116 59866 26172 59868
rect 26196 59866 26252 59868
rect 25956 59814 25982 59866
rect 25982 59814 26012 59866
rect 26036 59814 26046 59866
rect 26046 59814 26092 59866
rect 26116 59814 26162 59866
rect 26162 59814 26172 59866
rect 26196 59814 26226 59866
rect 26226 59814 26252 59866
rect 25956 59812 26012 59814
rect 26036 59812 26092 59814
rect 26116 59812 26172 59814
rect 26196 59812 26252 59814
rect 26514 59336 26570 59392
rect 25956 58778 26012 58780
rect 26036 58778 26092 58780
rect 26116 58778 26172 58780
rect 26196 58778 26252 58780
rect 25956 58726 25982 58778
rect 25982 58726 26012 58778
rect 26036 58726 26046 58778
rect 26046 58726 26092 58778
rect 26116 58726 26162 58778
rect 26162 58726 26172 58778
rect 26196 58726 26226 58778
rect 26226 58726 26252 58778
rect 25956 58724 26012 58726
rect 26036 58724 26092 58726
rect 26116 58724 26172 58726
rect 26196 58724 26252 58726
rect 25956 57690 26012 57692
rect 26036 57690 26092 57692
rect 26116 57690 26172 57692
rect 26196 57690 26252 57692
rect 25956 57638 25982 57690
rect 25982 57638 26012 57690
rect 26036 57638 26046 57690
rect 26046 57638 26092 57690
rect 26116 57638 26162 57690
rect 26162 57638 26172 57690
rect 26196 57638 26226 57690
rect 26226 57638 26252 57690
rect 25956 57636 26012 57638
rect 26036 57636 26092 57638
rect 26116 57636 26172 57638
rect 26196 57636 26252 57638
rect 25956 56602 26012 56604
rect 26036 56602 26092 56604
rect 26116 56602 26172 56604
rect 26196 56602 26252 56604
rect 25956 56550 25982 56602
rect 25982 56550 26012 56602
rect 26036 56550 26046 56602
rect 26046 56550 26092 56602
rect 26116 56550 26162 56602
rect 26162 56550 26172 56602
rect 26196 56550 26226 56602
rect 26226 56550 26252 56602
rect 25956 56548 26012 56550
rect 26036 56548 26092 56550
rect 26116 56548 26172 56550
rect 26196 56548 26252 56550
rect 25962 56344 26018 56400
rect 25956 55514 26012 55516
rect 26036 55514 26092 55516
rect 26116 55514 26172 55516
rect 26196 55514 26252 55516
rect 25956 55462 25982 55514
rect 25982 55462 26012 55514
rect 26036 55462 26046 55514
rect 26046 55462 26092 55514
rect 26116 55462 26162 55514
rect 26162 55462 26172 55514
rect 26196 55462 26226 55514
rect 26226 55462 26252 55514
rect 25956 55460 26012 55462
rect 26036 55460 26092 55462
rect 26116 55460 26172 55462
rect 26196 55460 26252 55462
rect 26606 54984 26662 55040
rect 25956 54426 26012 54428
rect 26036 54426 26092 54428
rect 26116 54426 26172 54428
rect 26196 54426 26252 54428
rect 25956 54374 25982 54426
rect 25982 54374 26012 54426
rect 26036 54374 26046 54426
rect 26046 54374 26092 54426
rect 26116 54374 26162 54426
rect 26162 54374 26172 54426
rect 26196 54374 26226 54426
rect 26226 54374 26252 54426
rect 25956 54372 26012 54374
rect 26036 54372 26092 54374
rect 26116 54372 26172 54374
rect 26196 54372 26252 54374
rect 25956 53338 26012 53340
rect 26036 53338 26092 53340
rect 26116 53338 26172 53340
rect 26196 53338 26252 53340
rect 25956 53286 25982 53338
rect 25982 53286 26012 53338
rect 26036 53286 26046 53338
rect 26046 53286 26092 53338
rect 26116 53286 26162 53338
rect 26162 53286 26172 53338
rect 26196 53286 26226 53338
rect 26226 53286 26252 53338
rect 25956 53284 26012 53286
rect 26036 53284 26092 53286
rect 26116 53284 26172 53286
rect 26196 53284 26252 53286
rect 25686 52536 25742 52592
rect 25778 52264 25834 52320
rect 25956 52250 26012 52252
rect 26036 52250 26092 52252
rect 26116 52250 26172 52252
rect 26196 52250 26252 52252
rect 25956 52198 25982 52250
rect 25982 52198 26012 52250
rect 26036 52198 26046 52250
rect 26046 52198 26092 52250
rect 26116 52198 26162 52250
rect 26162 52198 26172 52250
rect 26196 52198 26226 52250
rect 26226 52198 26252 52250
rect 25956 52196 26012 52198
rect 26036 52196 26092 52198
rect 26116 52196 26172 52198
rect 26196 52196 26252 52198
rect 25686 51720 25742 51776
rect 25956 51162 26012 51164
rect 26036 51162 26092 51164
rect 26116 51162 26172 51164
rect 26196 51162 26252 51164
rect 25956 51110 25982 51162
rect 25982 51110 26012 51162
rect 26036 51110 26046 51162
rect 26046 51110 26092 51162
rect 26116 51110 26162 51162
rect 26162 51110 26172 51162
rect 26196 51110 26226 51162
rect 26226 51110 26252 51162
rect 25956 51108 26012 51110
rect 26036 51108 26092 51110
rect 26116 51108 26172 51110
rect 26196 51108 26252 51110
rect 25956 50074 26012 50076
rect 26036 50074 26092 50076
rect 26116 50074 26172 50076
rect 26196 50074 26252 50076
rect 25956 50022 25982 50074
rect 25982 50022 26012 50074
rect 26036 50022 26046 50074
rect 26046 50022 26092 50074
rect 26116 50022 26162 50074
rect 26162 50022 26172 50074
rect 26196 50022 26226 50074
rect 26226 50022 26252 50074
rect 25956 50020 26012 50022
rect 26036 50020 26092 50022
rect 26116 50020 26172 50022
rect 26196 50020 26252 50022
rect 25956 48986 26012 48988
rect 26036 48986 26092 48988
rect 26116 48986 26172 48988
rect 26196 48986 26252 48988
rect 25956 48934 25982 48986
rect 25982 48934 26012 48986
rect 26036 48934 26046 48986
rect 26046 48934 26092 48986
rect 26116 48934 26162 48986
rect 26162 48934 26172 48986
rect 26196 48934 26226 48986
rect 26226 48934 26252 48986
rect 25956 48932 26012 48934
rect 26036 48932 26092 48934
rect 26116 48932 26172 48934
rect 26196 48932 26252 48934
rect 25956 47898 26012 47900
rect 26036 47898 26092 47900
rect 26116 47898 26172 47900
rect 26196 47898 26252 47900
rect 25956 47846 25982 47898
rect 25982 47846 26012 47898
rect 26036 47846 26046 47898
rect 26046 47846 26092 47898
rect 26116 47846 26162 47898
rect 26162 47846 26172 47898
rect 26196 47846 26226 47898
rect 26226 47846 26252 47898
rect 25956 47844 26012 47846
rect 26036 47844 26092 47846
rect 26116 47844 26172 47846
rect 26196 47844 26252 47846
rect 26698 47640 26754 47696
rect 25870 47232 25926 47288
rect 25686 46960 25742 47016
rect 25502 41520 25558 41576
rect 25502 38528 25558 38584
rect 25594 38120 25650 38176
rect 25318 34584 25374 34640
rect 26514 47116 26570 47152
rect 26514 47096 26516 47116
rect 26516 47096 26568 47116
rect 26568 47096 26570 47116
rect 25956 46810 26012 46812
rect 26036 46810 26092 46812
rect 26116 46810 26172 46812
rect 26196 46810 26252 46812
rect 25956 46758 25982 46810
rect 25982 46758 26012 46810
rect 26036 46758 26046 46810
rect 26046 46758 26092 46810
rect 26116 46758 26162 46810
rect 26162 46758 26172 46810
rect 26196 46758 26226 46810
rect 26226 46758 26252 46810
rect 25956 46756 26012 46758
rect 26036 46756 26092 46758
rect 26116 46756 26172 46758
rect 26196 46756 26252 46758
rect 25956 45722 26012 45724
rect 26036 45722 26092 45724
rect 26116 45722 26172 45724
rect 26196 45722 26252 45724
rect 25956 45670 25982 45722
rect 25982 45670 26012 45722
rect 26036 45670 26046 45722
rect 26046 45670 26092 45722
rect 26116 45670 26162 45722
rect 26162 45670 26172 45722
rect 26196 45670 26226 45722
rect 26226 45670 26252 45722
rect 25956 45668 26012 45670
rect 26036 45668 26092 45670
rect 26116 45668 26172 45670
rect 26196 45668 26252 45670
rect 26514 45872 26570 45928
rect 26422 45464 26478 45520
rect 26330 45056 26386 45112
rect 25956 44634 26012 44636
rect 26036 44634 26092 44636
rect 26116 44634 26172 44636
rect 26196 44634 26252 44636
rect 25956 44582 25982 44634
rect 25982 44582 26012 44634
rect 26036 44582 26046 44634
rect 26046 44582 26092 44634
rect 26116 44582 26162 44634
rect 26162 44582 26172 44634
rect 26196 44582 26226 44634
rect 26226 44582 26252 44634
rect 25956 44580 26012 44582
rect 26036 44580 26092 44582
rect 26116 44580 26172 44582
rect 26196 44580 26252 44582
rect 25956 43546 26012 43548
rect 26036 43546 26092 43548
rect 26116 43546 26172 43548
rect 26196 43546 26252 43548
rect 25956 43494 25982 43546
rect 25982 43494 26012 43546
rect 26036 43494 26046 43546
rect 26046 43494 26092 43546
rect 26116 43494 26162 43546
rect 26162 43494 26172 43546
rect 26196 43494 26226 43546
rect 26226 43494 26252 43546
rect 25956 43492 26012 43494
rect 26036 43492 26092 43494
rect 26116 43492 26172 43494
rect 26196 43492 26252 43494
rect 26606 44784 26662 44840
rect 26882 43868 26884 43888
rect 26884 43868 26936 43888
rect 26936 43868 26938 43888
rect 26882 43832 26938 43868
rect 25956 42458 26012 42460
rect 26036 42458 26092 42460
rect 26116 42458 26172 42460
rect 26196 42458 26252 42460
rect 25956 42406 25982 42458
rect 25982 42406 26012 42458
rect 26036 42406 26046 42458
rect 26046 42406 26092 42458
rect 26116 42406 26162 42458
rect 26162 42406 26172 42458
rect 26196 42406 26226 42458
rect 26226 42406 26252 42458
rect 25956 42404 26012 42406
rect 26036 42404 26092 42406
rect 26116 42404 26172 42406
rect 26196 42404 26252 42406
rect 25962 42236 25964 42256
rect 25964 42236 26016 42256
rect 26016 42236 26018 42256
rect 25962 42200 26018 42236
rect 26606 42200 26662 42256
rect 26514 42064 26570 42120
rect 25956 41370 26012 41372
rect 26036 41370 26092 41372
rect 26116 41370 26172 41372
rect 26196 41370 26252 41372
rect 25956 41318 25982 41370
rect 25982 41318 26012 41370
rect 26036 41318 26046 41370
rect 26046 41318 26092 41370
rect 26116 41318 26162 41370
rect 26162 41318 26172 41370
rect 26196 41318 26226 41370
rect 26226 41318 26252 41370
rect 25956 41316 26012 41318
rect 26036 41316 26092 41318
rect 26116 41316 26172 41318
rect 26196 41316 26252 41318
rect 25956 40282 26012 40284
rect 26036 40282 26092 40284
rect 26116 40282 26172 40284
rect 26196 40282 26252 40284
rect 25956 40230 25982 40282
rect 25982 40230 26012 40282
rect 26036 40230 26046 40282
rect 26046 40230 26092 40282
rect 26116 40230 26162 40282
rect 26162 40230 26172 40282
rect 26196 40230 26226 40282
rect 26226 40230 26252 40282
rect 25956 40228 26012 40230
rect 26036 40228 26092 40230
rect 26116 40228 26172 40230
rect 26196 40228 26252 40230
rect 25870 40024 25926 40080
rect 25956 39194 26012 39196
rect 26036 39194 26092 39196
rect 26116 39194 26172 39196
rect 26196 39194 26252 39196
rect 25956 39142 25982 39194
rect 25982 39142 26012 39194
rect 26036 39142 26046 39194
rect 26046 39142 26092 39194
rect 26116 39142 26162 39194
rect 26162 39142 26172 39194
rect 26196 39142 26226 39194
rect 26226 39142 26252 39194
rect 25956 39140 26012 39142
rect 26036 39140 26092 39142
rect 26116 39140 26172 39142
rect 26196 39140 26252 39142
rect 26422 38836 26424 38856
rect 26424 38836 26476 38856
rect 26476 38836 26478 38856
rect 26422 38800 26478 38836
rect 25956 38106 26012 38108
rect 26036 38106 26092 38108
rect 26116 38106 26172 38108
rect 26196 38106 26252 38108
rect 25956 38054 25982 38106
rect 25982 38054 26012 38106
rect 26036 38054 26046 38106
rect 26046 38054 26092 38106
rect 26116 38054 26162 38106
rect 26162 38054 26172 38106
rect 26196 38054 26226 38106
rect 26226 38054 26252 38106
rect 25956 38052 26012 38054
rect 26036 38052 26092 38054
rect 26116 38052 26172 38054
rect 26196 38052 26252 38054
rect 25956 37018 26012 37020
rect 26036 37018 26092 37020
rect 26116 37018 26172 37020
rect 26196 37018 26252 37020
rect 25956 36966 25982 37018
rect 25982 36966 26012 37018
rect 26036 36966 26046 37018
rect 26046 36966 26092 37018
rect 26116 36966 26162 37018
rect 26162 36966 26172 37018
rect 26196 36966 26226 37018
rect 26226 36966 26252 37018
rect 25956 36964 26012 36966
rect 26036 36964 26092 36966
rect 26116 36964 26172 36966
rect 26196 36964 26252 36966
rect 25956 35930 26012 35932
rect 26036 35930 26092 35932
rect 26116 35930 26172 35932
rect 26196 35930 26252 35932
rect 25956 35878 25982 35930
rect 25982 35878 26012 35930
rect 26036 35878 26046 35930
rect 26046 35878 26092 35930
rect 26116 35878 26162 35930
rect 26162 35878 26172 35930
rect 26196 35878 26226 35930
rect 26226 35878 26252 35930
rect 25956 35876 26012 35878
rect 26036 35876 26092 35878
rect 26116 35876 26172 35878
rect 26196 35876 26252 35878
rect 25956 34842 26012 34844
rect 26036 34842 26092 34844
rect 26116 34842 26172 34844
rect 26196 34842 26252 34844
rect 25956 34790 25982 34842
rect 25982 34790 26012 34842
rect 26036 34790 26046 34842
rect 26046 34790 26092 34842
rect 26116 34790 26162 34842
rect 26162 34790 26172 34842
rect 26196 34790 26226 34842
rect 26226 34790 26252 34842
rect 25956 34788 26012 34790
rect 26036 34788 26092 34790
rect 26116 34788 26172 34790
rect 26196 34788 26252 34790
rect 25594 33360 25650 33416
rect 25686 30640 25742 30696
rect 25410 27648 25466 27704
rect 25502 26560 25558 26616
rect 25686 26152 25742 26208
rect 25956 33754 26012 33756
rect 26036 33754 26092 33756
rect 26116 33754 26172 33756
rect 26196 33754 26252 33756
rect 25956 33702 25982 33754
rect 25982 33702 26012 33754
rect 26036 33702 26046 33754
rect 26046 33702 26092 33754
rect 26116 33702 26162 33754
rect 26162 33702 26172 33754
rect 26196 33702 26226 33754
rect 26226 33702 26252 33754
rect 25956 33700 26012 33702
rect 26036 33700 26092 33702
rect 26116 33700 26172 33702
rect 26196 33700 26252 33702
rect 25956 32666 26012 32668
rect 26036 32666 26092 32668
rect 26116 32666 26172 32668
rect 26196 32666 26252 32668
rect 25956 32614 25982 32666
rect 25982 32614 26012 32666
rect 26036 32614 26046 32666
rect 26046 32614 26092 32666
rect 26116 32614 26162 32666
rect 26162 32614 26172 32666
rect 26196 32614 26226 32666
rect 26226 32614 26252 32666
rect 25956 32612 26012 32614
rect 26036 32612 26092 32614
rect 26116 32612 26172 32614
rect 26196 32612 26252 32614
rect 25956 31578 26012 31580
rect 26036 31578 26092 31580
rect 26116 31578 26172 31580
rect 26196 31578 26252 31580
rect 25956 31526 25982 31578
rect 25982 31526 26012 31578
rect 26036 31526 26046 31578
rect 26046 31526 26092 31578
rect 26116 31526 26162 31578
rect 26162 31526 26172 31578
rect 26196 31526 26226 31578
rect 26226 31526 26252 31578
rect 25956 31524 26012 31526
rect 26036 31524 26092 31526
rect 26116 31524 26172 31526
rect 26196 31524 26252 31526
rect 25956 30490 26012 30492
rect 26036 30490 26092 30492
rect 26116 30490 26172 30492
rect 26196 30490 26252 30492
rect 25956 30438 25982 30490
rect 25982 30438 26012 30490
rect 26036 30438 26046 30490
rect 26046 30438 26092 30490
rect 26116 30438 26162 30490
rect 26162 30438 26172 30490
rect 26196 30438 26226 30490
rect 26226 30438 26252 30490
rect 25956 30436 26012 30438
rect 26036 30436 26092 30438
rect 26116 30436 26172 30438
rect 26196 30436 26252 30438
rect 25956 29402 26012 29404
rect 26036 29402 26092 29404
rect 26116 29402 26172 29404
rect 26196 29402 26252 29404
rect 25956 29350 25982 29402
rect 25982 29350 26012 29402
rect 26036 29350 26046 29402
rect 26046 29350 26092 29402
rect 26116 29350 26162 29402
rect 26162 29350 26172 29402
rect 26196 29350 26226 29402
rect 26226 29350 26252 29402
rect 25956 29348 26012 29350
rect 26036 29348 26092 29350
rect 26116 29348 26172 29350
rect 26196 29348 26252 29350
rect 25870 28872 25926 28928
rect 25956 28314 26012 28316
rect 26036 28314 26092 28316
rect 26116 28314 26172 28316
rect 26196 28314 26252 28316
rect 25956 28262 25982 28314
rect 25982 28262 26012 28314
rect 26036 28262 26046 28314
rect 26046 28262 26092 28314
rect 26116 28262 26162 28314
rect 26162 28262 26172 28314
rect 26196 28262 26226 28314
rect 26226 28262 26252 28314
rect 25956 28260 26012 28262
rect 26036 28260 26092 28262
rect 26116 28260 26172 28262
rect 26196 28260 26252 28262
rect 25956 27226 26012 27228
rect 26036 27226 26092 27228
rect 26116 27226 26172 27228
rect 26196 27226 26252 27228
rect 25956 27174 25982 27226
rect 25982 27174 26012 27226
rect 26036 27174 26046 27226
rect 26046 27174 26092 27226
rect 26116 27174 26162 27226
rect 26162 27174 26172 27226
rect 26196 27174 26226 27226
rect 26226 27174 26252 27226
rect 25956 27172 26012 27174
rect 26036 27172 26092 27174
rect 26116 27172 26172 27174
rect 26196 27172 26252 27174
rect 25956 26138 26012 26140
rect 26036 26138 26092 26140
rect 26116 26138 26172 26140
rect 26196 26138 26252 26140
rect 25956 26086 25982 26138
rect 25982 26086 26012 26138
rect 26036 26086 26046 26138
rect 26046 26086 26092 26138
rect 26116 26086 26162 26138
rect 26162 26086 26172 26138
rect 26196 26086 26226 26138
rect 26226 26086 26252 26138
rect 25956 26084 26012 26086
rect 26036 26084 26092 26086
rect 26116 26084 26172 26086
rect 26196 26084 26252 26086
rect 25870 25200 25926 25256
rect 25956 25050 26012 25052
rect 26036 25050 26092 25052
rect 26116 25050 26172 25052
rect 26196 25050 26252 25052
rect 25956 24998 25982 25050
rect 25982 24998 26012 25050
rect 26036 24998 26046 25050
rect 26046 24998 26092 25050
rect 26116 24998 26162 25050
rect 26162 24998 26172 25050
rect 26196 24998 26226 25050
rect 26226 24998 26252 25050
rect 25956 24996 26012 24998
rect 26036 24996 26092 24998
rect 26116 24996 26172 24998
rect 26196 24996 26252 24998
rect 25956 23962 26012 23964
rect 26036 23962 26092 23964
rect 26116 23962 26172 23964
rect 26196 23962 26252 23964
rect 25956 23910 25982 23962
rect 25982 23910 26012 23962
rect 26036 23910 26046 23962
rect 26046 23910 26092 23962
rect 26116 23910 26162 23962
rect 26162 23910 26172 23962
rect 26196 23910 26226 23962
rect 26226 23910 26252 23962
rect 25956 23908 26012 23910
rect 26036 23908 26092 23910
rect 26116 23908 26172 23910
rect 26196 23908 26252 23910
rect 25956 22874 26012 22876
rect 26036 22874 26092 22876
rect 26116 22874 26172 22876
rect 26196 22874 26252 22876
rect 25956 22822 25982 22874
rect 25982 22822 26012 22874
rect 26036 22822 26046 22874
rect 26046 22822 26092 22874
rect 26116 22822 26162 22874
rect 26162 22822 26172 22874
rect 26196 22822 26226 22874
rect 26226 22822 26252 22874
rect 25956 22820 26012 22822
rect 26036 22820 26092 22822
rect 26116 22820 26172 22822
rect 26196 22820 26252 22822
rect 26330 21800 26386 21856
rect 25956 21786 26012 21788
rect 26036 21786 26092 21788
rect 26116 21786 26172 21788
rect 26196 21786 26252 21788
rect 25956 21734 25982 21786
rect 25982 21734 26012 21786
rect 26036 21734 26046 21786
rect 26046 21734 26092 21786
rect 26116 21734 26162 21786
rect 26162 21734 26172 21786
rect 26196 21734 26226 21786
rect 26226 21734 26252 21786
rect 25956 21732 26012 21734
rect 26036 21732 26092 21734
rect 26116 21732 26172 21734
rect 26196 21732 26252 21734
rect 25778 21120 25834 21176
rect 26330 20984 26386 21040
rect 25956 20698 26012 20700
rect 26036 20698 26092 20700
rect 26116 20698 26172 20700
rect 26196 20698 26252 20700
rect 25956 20646 25982 20698
rect 25982 20646 26012 20698
rect 26036 20646 26046 20698
rect 26046 20646 26092 20698
rect 26116 20646 26162 20698
rect 26162 20646 26172 20698
rect 26196 20646 26226 20698
rect 26226 20646 26252 20698
rect 25956 20644 26012 20646
rect 26036 20644 26092 20646
rect 26116 20644 26172 20646
rect 26196 20644 26252 20646
rect 25594 20168 25650 20224
rect 25956 19610 26012 19612
rect 26036 19610 26092 19612
rect 26116 19610 26172 19612
rect 26196 19610 26252 19612
rect 25956 19558 25982 19610
rect 25982 19558 26012 19610
rect 26036 19558 26046 19610
rect 26046 19558 26092 19610
rect 26116 19558 26162 19610
rect 26162 19558 26172 19610
rect 26196 19558 26226 19610
rect 26226 19558 26252 19610
rect 25956 19556 26012 19558
rect 26036 19556 26092 19558
rect 26116 19556 26172 19558
rect 26196 19556 26252 19558
rect 25594 18672 25650 18728
rect 25956 18522 26012 18524
rect 26036 18522 26092 18524
rect 26116 18522 26172 18524
rect 26196 18522 26252 18524
rect 25956 18470 25982 18522
rect 25982 18470 26012 18522
rect 26036 18470 26046 18522
rect 26046 18470 26092 18522
rect 26116 18470 26162 18522
rect 26162 18470 26172 18522
rect 26196 18470 26226 18522
rect 26226 18470 26252 18522
rect 25956 18468 26012 18470
rect 26036 18468 26092 18470
rect 26116 18468 26172 18470
rect 26196 18468 26252 18470
rect 25502 17720 25558 17776
rect 25410 13368 25466 13424
rect 25226 11600 25282 11656
rect 24950 7384 25006 7440
rect 24858 5208 24914 5264
rect 23938 3984 23994 4040
rect 23018 3712 23074 3768
rect 3146 720 3202 776
rect 25318 6840 25374 6896
rect 25318 4120 25374 4176
rect 25318 2624 25374 2680
rect 24950 720 25006 776
rect 25956 17434 26012 17436
rect 26036 17434 26092 17436
rect 26116 17434 26172 17436
rect 26196 17434 26252 17436
rect 25956 17382 25982 17434
rect 25982 17382 26012 17434
rect 26036 17382 26046 17434
rect 26046 17382 26092 17434
rect 26116 17382 26162 17434
rect 26162 17382 26172 17434
rect 26196 17382 26226 17434
rect 26226 17382 26252 17434
rect 25956 17380 26012 17382
rect 26036 17380 26092 17382
rect 26116 17380 26172 17382
rect 26196 17380 26252 17382
rect 25956 16346 26012 16348
rect 26036 16346 26092 16348
rect 26116 16346 26172 16348
rect 26196 16346 26252 16348
rect 25956 16294 25982 16346
rect 25982 16294 26012 16346
rect 26036 16294 26046 16346
rect 26046 16294 26092 16346
rect 26116 16294 26162 16346
rect 26162 16294 26172 16346
rect 26196 16294 26226 16346
rect 26226 16294 26252 16346
rect 25956 16292 26012 16294
rect 26036 16292 26092 16294
rect 26116 16292 26172 16294
rect 26196 16292 26252 16294
rect 25956 15258 26012 15260
rect 26036 15258 26092 15260
rect 26116 15258 26172 15260
rect 26196 15258 26252 15260
rect 25956 15206 25982 15258
rect 25982 15206 26012 15258
rect 26036 15206 26046 15258
rect 26046 15206 26092 15258
rect 26116 15206 26162 15258
rect 26162 15206 26172 15258
rect 26196 15206 26226 15258
rect 26226 15206 26252 15258
rect 25956 15204 26012 15206
rect 26036 15204 26092 15206
rect 26116 15204 26172 15206
rect 26196 15204 26252 15206
rect 25956 14170 26012 14172
rect 26036 14170 26092 14172
rect 26116 14170 26172 14172
rect 26196 14170 26252 14172
rect 25956 14118 25982 14170
rect 25982 14118 26012 14170
rect 26036 14118 26046 14170
rect 26046 14118 26092 14170
rect 26116 14118 26162 14170
rect 26162 14118 26172 14170
rect 26196 14118 26226 14170
rect 26226 14118 26252 14170
rect 25956 14116 26012 14118
rect 26036 14116 26092 14118
rect 26116 14116 26172 14118
rect 26196 14116 26252 14118
rect 26238 13796 26294 13832
rect 26238 13776 26240 13796
rect 26240 13776 26292 13796
rect 26292 13776 26294 13796
rect 25956 13082 26012 13084
rect 26036 13082 26092 13084
rect 26116 13082 26172 13084
rect 26196 13082 26252 13084
rect 25956 13030 25982 13082
rect 25982 13030 26012 13082
rect 26036 13030 26046 13082
rect 26046 13030 26092 13082
rect 26116 13030 26162 13082
rect 26162 13030 26172 13082
rect 26196 13030 26226 13082
rect 26226 13030 26252 13082
rect 25956 13028 26012 13030
rect 26036 13028 26092 13030
rect 26116 13028 26172 13030
rect 26196 13028 26252 13030
rect 25956 11994 26012 11996
rect 26036 11994 26092 11996
rect 26116 11994 26172 11996
rect 26196 11994 26252 11996
rect 25956 11942 25982 11994
rect 25982 11942 26012 11994
rect 26036 11942 26046 11994
rect 26046 11942 26092 11994
rect 26116 11942 26162 11994
rect 26162 11942 26172 11994
rect 26196 11942 26226 11994
rect 26226 11942 26252 11994
rect 25956 11940 26012 11942
rect 26036 11940 26092 11942
rect 26116 11940 26172 11942
rect 26196 11940 26252 11942
rect 26330 11464 26386 11520
rect 25956 10906 26012 10908
rect 26036 10906 26092 10908
rect 26116 10906 26172 10908
rect 26196 10906 26252 10908
rect 25956 10854 25982 10906
rect 25982 10854 26012 10906
rect 26036 10854 26046 10906
rect 26046 10854 26092 10906
rect 26116 10854 26162 10906
rect 26162 10854 26172 10906
rect 26196 10854 26226 10906
rect 26226 10854 26252 10906
rect 25956 10852 26012 10854
rect 26036 10852 26092 10854
rect 26116 10852 26172 10854
rect 26196 10852 26252 10854
rect 25956 9818 26012 9820
rect 26036 9818 26092 9820
rect 26116 9818 26172 9820
rect 26196 9818 26252 9820
rect 25956 9766 25982 9818
rect 25982 9766 26012 9818
rect 26036 9766 26046 9818
rect 26046 9766 26092 9818
rect 26116 9766 26162 9818
rect 26162 9766 26172 9818
rect 26196 9766 26226 9818
rect 26226 9766 26252 9818
rect 25956 9764 26012 9766
rect 26036 9764 26092 9766
rect 26116 9764 26172 9766
rect 26196 9764 26252 9766
rect 25956 8730 26012 8732
rect 26036 8730 26092 8732
rect 26116 8730 26172 8732
rect 26196 8730 26252 8732
rect 25956 8678 25982 8730
rect 25982 8678 26012 8730
rect 26036 8678 26046 8730
rect 26046 8678 26092 8730
rect 26116 8678 26162 8730
rect 26162 8678 26172 8730
rect 26196 8678 26226 8730
rect 26226 8678 26252 8730
rect 25956 8676 26012 8678
rect 26036 8676 26092 8678
rect 26116 8676 26172 8678
rect 26196 8676 26252 8678
rect 25956 7642 26012 7644
rect 26036 7642 26092 7644
rect 26116 7642 26172 7644
rect 26196 7642 26252 7644
rect 25956 7590 25982 7642
rect 25982 7590 26012 7642
rect 26036 7590 26046 7642
rect 26046 7590 26092 7642
rect 26116 7590 26162 7642
rect 26162 7590 26172 7642
rect 26196 7590 26226 7642
rect 26226 7590 26252 7642
rect 25956 7588 26012 7590
rect 26036 7588 26092 7590
rect 26116 7588 26172 7590
rect 26196 7588 26252 7590
rect 25956 6554 26012 6556
rect 26036 6554 26092 6556
rect 26116 6554 26172 6556
rect 26196 6554 26252 6556
rect 25956 6502 25982 6554
rect 25982 6502 26012 6554
rect 26036 6502 26046 6554
rect 26046 6502 26092 6554
rect 26116 6502 26162 6554
rect 26162 6502 26172 6554
rect 26196 6502 26226 6554
rect 26226 6502 26252 6554
rect 25956 6500 26012 6502
rect 26036 6500 26092 6502
rect 26116 6500 26172 6502
rect 26196 6500 26252 6502
rect 25956 5466 26012 5468
rect 26036 5466 26092 5468
rect 26116 5466 26172 5468
rect 26196 5466 26252 5468
rect 25956 5414 25982 5466
rect 25982 5414 26012 5466
rect 26036 5414 26046 5466
rect 26046 5414 26092 5466
rect 26116 5414 26162 5466
rect 26162 5414 26172 5466
rect 26196 5414 26226 5466
rect 26226 5414 26252 5466
rect 25956 5412 26012 5414
rect 26036 5412 26092 5414
rect 26116 5412 26172 5414
rect 26196 5412 26252 5414
rect 25956 4378 26012 4380
rect 26036 4378 26092 4380
rect 26116 4378 26172 4380
rect 26196 4378 26252 4380
rect 25956 4326 25982 4378
rect 25982 4326 26012 4378
rect 26036 4326 26046 4378
rect 26046 4326 26092 4378
rect 26116 4326 26162 4378
rect 26162 4326 26172 4378
rect 26196 4326 26226 4378
rect 26226 4326 26252 4378
rect 25956 4324 26012 4326
rect 26036 4324 26092 4326
rect 26116 4324 26172 4326
rect 26196 4324 26252 4326
rect 25956 3290 26012 3292
rect 26036 3290 26092 3292
rect 26116 3290 26172 3292
rect 26196 3290 26252 3292
rect 25956 3238 25982 3290
rect 25982 3238 26012 3290
rect 26036 3238 26046 3290
rect 26046 3238 26092 3290
rect 26116 3238 26162 3290
rect 26162 3238 26172 3290
rect 26196 3238 26226 3290
rect 26226 3238 26252 3290
rect 25956 3236 26012 3238
rect 26036 3236 26092 3238
rect 26116 3236 26172 3238
rect 26196 3236 26252 3238
rect 25956 2202 26012 2204
rect 26036 2202 26092 2204
rect 26116 2202 26172 2204
rect 26196 2202 26252 2204
rect 25956 2150 25982 2202
rect 25982 2150 26012 2202
rect 26036 2150 26046 2202
rect 26046 2150 26092 2202
rect 26116 2150 26162 2202
rect 26162 2150 26172 2202
rect 26196 2150 26226 2202
rect 26226 2150 26252 2202
rect 25956 2148 26012 2150
rect 26036 2148 26092 2150
rect 26116 2148 26172 2150
rect 26196 2148 26252 2150
rect 27986 66136 28042 66192
rect 27986 56616 28042 56672
rect 27894 52944 27950 53000
rect 27342 52400 27398 52456
rect 27710 49544 27766 49600
rect 27526 43968 27582 44024
rect 27250 43288 27306 43344
rect 27342 42744 27398 42800
rect 27710 42608 27766 42664
rect 27066 41656 27122 41712
rect 27710 36080 27766 36136
rect 27710 35672 27766 35728
rect 28078 48456 28134 48512
rect 27802 33224 27858 33280
rect 27618 31184 27674 31240
rect 26974 23840 27030 23896
rect 27710 20304 27766 20360
rect 27618 13932 27674 13968
rect 27618 13912 27620 13932
rect 27620 13912 27672 13932
rect 27672 13912 27674 13932
rect 26514 13812 26516 13832
rect 26516 13812 26568 13832
rect 26568 13812 26570 13832
rect 26514 13776 26570 13812
rect 29458 8472 29514 8528
rect 28538 4800 28594 4856
rect 26514 2080 26570 2136
rect 28078 1944 28134 2000
rect 25502 40 25558 96
<< metal3 >>
rect 0 79658 800 79688
rect 4061 79658 4127 79661
rect 0 79656 4127 79658
rect 0 79600 4066 79656
rect 4122 79600 4127 79656
rect 0 79598 4127 79600
rect 0 79568 800 79598
rect 4061 79595 4127 79598
rect 24669 79658 24735 79661
rect 29200 79658 30000 79688
rect 24669 79656 30000 79658
rect 24669 79600 24674 79656
rect 24730 79600 30000 79656
rect 24669 79598 30000 79600
rect 24669 79595 24735 79598
rect 29200 79568 30000 79598
rect 0 78298 800 78328
rect 3325 78298 3391 78301
rect 0 78296 3391 78298
rect 0 78240 3330 78296
rect 3386 78240 3391 78296
rect 0 78238 3391 78240
rect 0 78208 800 78238
rect 3325 78235 3391 78238
rect 25865 78298 25931 78301
rect 29200 78298 30000 78328
rect 25865 78296 30000 78298
rect 25865 78240 25870 78296
rect 25926 78240 30000 78296
rect 25865 78238 30000 78240
rect 25865 78235 25931 78238
rect 29200 78208 30000 78238
rect 10944 77824 11264 77825
rect 10944 77760 10952 77824
rect 11016 77760 11032 77824
rect 11096 77760 11112 77824
rect 11176 77760 11192 77824
rect 11256 77760 11264 77824
rect 10944 77759 11264 77760
rect 20944 77824 21264 77825
rect 20944 77760 20952 77824
rect 21016 77760 21032 77824
rect 21096 77760 21112 77824
rect 21176 77760 21192 77824
rect 21256 77760 21264 77824
rect 20944 77759 21264 77760
rect 4061 77482 4127 77485
rect 20662 77482 20668 77484
rect 4061 77480 20668 77482
rect 4061 77424 4066 77480
rect 4122 77424 20668 77480
rect 4061 77422 20668 77424
rect 4061 77419 4127 77422
rect 20662 77420 20668 77422
rect 20732 77420 20738 77484
rect 5944 77280 6264 77281
rect 5944 77216 5952 77280
rect 6016 77216 6032 77280
rect 6096 77216 6112 77280
rect 6176 77216 6192 77280
rect 6256 77216 6264 77280
rect 5944 77215 6264 77216
rect 15944 77280 16264 77281
rect 15944 77216 15952 77280
rect 16016 77216 16032 77280
rect 16096 77216 16112 77280
rect 16176 77216 16192 77280
rect 16256 77216 16264 77280
rect 15944 77215 16264 77216
rect 25944 77280 26264 77281
rect 25944 77216 25952 77280
rect 26016 77216 26032 77280
rect 26096 77216 26112 77280
rect 26176 77216 26192 77280
rect 26256 77216 26264 77280
rect 25944 77215 26264 77216
rect 9581 77074 9647 77077
rect 798 77072 9647 77074
rect 798 77016 9586 77072
rect 9642 77016 9647 77072
rect 798 77014 9647 77016
rect 798 76968 858 77014
rect 9581 77011 9647 77014
rect 0 76878 858 76968
rect 25773 76938 25839 76941
rect 29200 76938 30000 76968
rect 25773 76936 30000 76938
rect 25773 76880 25778 76936
rect 25834 76880 30000 76936
rect 25773 76878 30000 76880
rect 0 76848 800 76878
rect 25773 76875 25839 76878
rect 29200 76848 30000 76878
rect 10944 76736 11264 76737
rect 10944 76672 10952 76736
rect 11016 76672 11032 76736
rect 11096 76672 11112 76736
rect 11176 76672 11192 76736
rect 11256 76672 11264 76736
rect 10944 76671 11264 76672
rect 20944 76736 21264 76737
rect 20944 76672 20952 76736
rect 21016 76672 21032 76736
rect 21096 76672 21112 76736
rect 21176 76672 21192 76736
rect 21256 76672 21264 76736
rect 20944 76671 21264 76672
rect 9581 76394 9647 76397
rect 13721 76394 13787 76397
rect 21265 76394 21331 76397
rect 9581 76392 11714 76394
rect 9581 76336 9586 76392
rect 9642 76336 11714 76392
rect 9581 76334 11714 76336
rect 9581 76331 9647 76334
rect 5944 76192 6264 76193
rect 5944 76128 5952 76192
rect 6016 76128 6032 76192
rect 6096 76128 6112 76192
rect 6176 76128 6192 76192
rect 6256 76128 6264 76192
rect 5944 76127 6264 76128
rect 11654 75986 11714 76334
rect 13721 76392 21331 76394
rect 13721 76336 13726 76392
rect 13782 76336 21270 76392
rect 21326 76336 21331 76392
rect 13721 76334 21331 76336
rect 13721 76331 13787 76334
rect 21265 76331 21331 76334
rect 25129 76394 25195 76397
rect 25129 76392 26618 76394
rect 25129 76336 25134 76392
rect 25190 76336 26618 76392
rect 25129 76334 26618 76336
rect 25129 76331 25195 76334
rect 26558 76258 26618 76334
rect 29200 76258 30000 76288
rect 26558 76198 30000 76258
rect 15944 76192 16264 76193
rect 15944 76128 15952 76192
rect 16016 76128 16032 76192
rect 16096 76128 16112 76192
rect 16176 76128 16192 76192
rect 16256 76128 16264 76192
rect 15944 76127 16264 76128
rect 25944 76192 26264 76193
rect 25944 76128 25952 76192
rect 26016 76128 26032 76192
rect 26096 76128 26112 76192
rect 26176 76128 26192 76192
rect 26256 76128 26264 76192
rect 29200 76168 30000 76198
rect 25944 76127 26264 76128
rect 25037 75986 25103 75989
rect 11654 75984 25103 75986
rect 11654 75928 25042 75984
rect 25098 75928 25103 75984
rect 11654 75926 25103 75928
rect 25037 75923 25103 75926
rect 2313 75850 2379 75853
rect 5349 75850 5415 75853
rect 2313 75848 5415 75850
rect 2313 75792 2318 75848
rect 2374 75792 5354 75848
rect 5410 75792 5415 75848
rect 2313 75790 5415 75792
rect 2313 75787 2379 75790
rect 5349 75787 5415 75790
rect 10133 75850 10199 75853
rect 12157 75850 12223 75853
rect 10133 75848 12223 75850
rect 10133 75792 10138 75848
rect 10194 75792 12162 75848
rect 12218 75792 12223 75848
rect 10133 75790 12223 75792
rect 10133 75787 10199 75790
rect 12157 75787 12223 75790
rect 13353 75850 13419 75853
rect 15101 75850 15167 75853
rect 16573 75850 16639 75853
rect 13353 75848 15026 75850
rect 13353 75792 13358 75848
rect 13414 75792 15026 75848
rect 13353 75790 15026 75792
rect 13353 75787 13419 75790
rect 11830 75652 11836 75716
rect 11900 75714 11906 75716
rect 13353 75714 13419 75717
rect 11900 75712 13419 75714
rect 11900 75656 13358 75712
rect 13414 75656 13419 75712
rect 11900 75654 13419 75656
rect 14966 75714 15026 75790
rect 15101 75848 16639 75850
rect 15101 75792 15106 75848
rect 15162 75792 16578 75848
rect 16634 75792 16639 75848
rect 15101 75790 16639 75792
rect 15101 75787 15167 75790
rect 16573 75787 16639 75790
rect 20805 75714 20871 75717
rect 14966 75712 20871 75714
rect 14966 75656 20810 75712
rect 20866 75656 20871 75712
rect 14966 75654 20871 75656
rect 11900 75652 11906 75654
rect 13353 75651 13419 75654
rect 20805 75651 20871 75654
rect 10944 75648 11264 75649
rect 0 75578 800 75608
rect 10944 75584 10952 75648
rect 11016 75584 11032 75648
rect 11096 75584 11112 75648
rect 11176 75584 11192 75648
rect 11256 75584 11264 75648
rect 10944 75583 11264 75584
rect 20944 75648 21264 75649
rect 20944 75584 20952 75648
rect 21016 75584 21032 75648
rect 21096 75584 21112 75648
rect 21176 75584 21192 75648
rect 21256 75584 21264 75648
rect 20944 75583 21264 75584
rect 2957 75578 3023 75581
rect 0 75576 3023 75578
rect 0 75520 2962 75576
rect 3018 75520 3023 75576
rect 0 75518 3023 75520
rect 0 75488 800 75518
rect 2957 75515 3023 75518
rect 6913 75306 6979 75309
rect 18597 75306 18663 75309
rect 6913 75304 18663 75306
rect 6913 75248 6918 75304
rect 6974 75248 18602 75304
rect 18658 75248 18663 75304
rect 6913 75246 18663 75248
rect 6913 75243 6979 75246
rect 18597 75243 18663 75246
rect 20805 75306 20871 75309
rect 26693 75306 26759 75309
rect 20805 75304 26759 75306
rect 20805 75248 20810 75304
rect 20866 75248 26698 75304
rect 26754 75248 26759 75304
rect 20805 75246 26759 75248
rect 20805 75243 20871 75246
rect 26693 75243 26759 75246
rect 5944 75104 6264 75105
rect 5944 75040 5952 75104
rect 6016 75040 6032 75104
rect 6096 75040 6112 75104
rect 6176 75040 6192 75104
rect 6256 75040 6264 75104
rect 5944 75039 6264 75040
rect 15944 75104 16264 75105
rect 15944 75040 15952 75104
rect 16016 75040 16032 75104
rect 16096 75040 16112 75104
rect 16176 75040 16192 75104
rect 16256 75040 16264 75104
rect 15944 75039 16264 75040
rect 25944 75104 26264 75105
rect 25944 75040 25952 75104
rect 26016 75040 26032 75104
rect 26096 75040 26112 75104
rect 26176 75040 26192 75104
rect 26256 75040 26264 75104
rect 25944 75039 26264 75040
rect 0 74898 800 74928
rect 3233 74898 3299 74901
rect 5625 74898 5691 74901
rect 0 74808 858 74898
rect 3233 74896 5691 74898
rect 3233 74840 3238 74896
rect 3294 74840 5630 74896
rect 5686 74840 5691 74896
rect 3233 74838 5691 74840
rect 3233 74835 3299 74838
rect 5625 74835 5691 74838
rect 25221 74898 25287 74901
rect 29200 74898 30000 74928
rect 25221 74896 30000 74898
rect 25221 74840 25226 74896
rect 25282 74840 30000 74896
rect 25221 74838 30000 74840
rect 25221 74835 25287 74838
rect 29200 74808 30000 74838
rect 798 74762 858 74808
rect 3417 74762 3483 74765
rect 798 74760 3483 74762
rect 798 74704 3422 74760
rect 3478 74704 3483 74760
rect 798 74702 3483 74704
rect 3417 74699 3483 74702
rect 5533 74762 5599 74765
rect 7465 74762 7531 74765
rect 5533 74760 7531 74762
rect 5533 74704 5538 74760
rect 5594 74704 7470 74760
rect 7526 74704 7531 74760
rect 5533 74702 7531 74704
rect 5533 74699 5599 74702
rect 7465 74699 7531 74702
rect 9673 74762 9739 74765
rect 9990 74762 9996 74764
rect 9673 74760 9996 74762
rect 9673 74704 9678 74760
rect 9734 74704 9996 74760
rect 9673 74702 9996 74704
rect 9673 74699 9739 74702
rect 9990 74700 9996 74702
rect 10060 74700 10066 74764
rect 23657 74762 23723 74765
rect 25681 74762 25747 74765
rect 23657 74760 25747 74762
rect 23657 74704 23662 74760
rect 23718 74704 25686 74760
rect 25742 74704 25747 74760
rect 23657 74702 25747 74704
rect 23657 74699 23723 74702
rect 25681 74699 25747 74702
rect 24853 74626 24919 74629
rect 25078 74626 25084 74628
rect 24853 74624 25084 74626
rect 24853 74568 24858 74624
rect 24914 74568 25084 74624
rect 24853 74566 25084 74568
rect 24853 74563 24919 74566
rect 25078 74564 25084 74566
rect 25148 74564 25154 74628
rect 10944 74560 11264 74561
rect 10944 74496 10952 74560
rect 11016 74496 11032 74560
rect 11096 74496 11112 74560
rect 11176 74496 11192 74560
rect 11256 74496 11264 74560
rect 10944 74495 11264 74496
rect 20944 74560 21264 74561
rect 20944 74496 20952 74560
rect 21016 74496 21032 74560
rect 21096 74496 21112 74560
rect 21176 74496 21192 74560
rect 21256 74496 21264 74560
rect 20944 74495 21264 74496
rect 23933 74490 23999 74493
rect 24894 74490 24900 74492
rect 23933 74488 24900 74490
rect 23933 74432 23938 74488
rect 23994 74432 24900 74488
rect 23933 74430 24900 74432
rect 23933 74427 23999 74430
rect 24894 74428 24900 74430
rect 24964 74428 24970 74492
rect 23105 74354 23171 74357
rect 24393 74354 24459 74357
rect 23105 74352 24459 74354
rect 23105 74296 23110 74352
rect 23166 74296 24398 74352
rect 24454 74296 24459 74352
rect 23105 74294 24459 74296
rect 23105 74291 23171 74294
rect 24393 74291 24459 74294
rect 5944 74016 6264 74017
rect 5944 73952 5952 74016
rect 6016 73952 6032 74016
rect 6096 73952 6112 74016
rect 6176 73952 6192 74016
rect 6256 73952 6264 74016
rect 5944 73951 6264 73952
rect 15944 74016 16264 74017
rect 15944 73952 15952 74016
rect 16016 73952 16032 74016
rect 16096 73952 16112 74016
rect 16176 73952 16192 74016
rect 16256 73952 16264 74016
rect 15944 73951 16264 73952
rect 25944 74016 26264 74017
rect 25944 73952 25952 74016
rect 26016 73952 26032 74016
rect 26096 73952 26112 74016
rect 26176 73952 26192 74016
rect 26256 73952 26264 74016
rect 25944 73951 26264 73952
rect 6913 73810 6979 73813
rect 23197 73810 23263 73813
rect 6913 73808 23263 73810
rect 6913 73752 6918 73808
rect 6974 73752 23202 73808
rect 23258 73752 23263 73808
rect 6913 73750 23263 73752
rect 6913 73747 6979 73750
rect 23197 73747 23263 73750
rect 1393 73674 1459 73677
rect 7741 73674 7807 73677
rect 1393 73672 7807 73674
rect 1393 73616 1398 73672
rect 1454 73616 7746 73672
rect 7802 73616 7807 73672
rect 1393 73614 7807 73616
rect 1393 73611 1459 73614
rect 7741 73611 7807 73614
rect 0 73538 800 73568
rect 22553 73538 22619 73541
rect 29200 73538 30000 73568
rect 0 73448 858 73538
rect 22553 73536 30000 73538
rect 22553 73480 22558 73536
rect 22614 73480 30000 73536
rect 22553 73478 30000 73480
rect 22553 73475 22619 73478
rect 798 73266 858 73448
rect 10944 73472 11264 73473
rect 10944 73408 10952 73472
rect 11016 73408 11032 73472
rect 11096 73408 11112 73472
rect 11176 73408 11192 73472
rect 11256 73408 11264 73472
rect 10944 73407 11264 73408
rect 20944 73472 21264 73473
rect 20944 73408 20952 73472
rect 21016 73408 21032 73472
rect 21096 73408 21112 73472
rect 21176 73408 21192 73472
rect 21256 73408 21264 73472
rect 29200 73448 30000 73478
rect 20944 73407 21264 73408
rect 17033 73402 17099 73405
rect 20805 73402 20871 73405
rect 17033 73400 20871 73402
rect 17033 73344 17038 73400
rect 17094 73344 20810 73400
rect 20866 73344 20871 73400
rect 17033 73342 20871 73344
rect 17033 73339 17099 73342
rect 20805 73339 20871 73342
rect 11513 73266 11579 73269
rect 798 73264 11579 73266
rect 798 73208 11518 73264
rect 11574 73208 11579 73264
rect 798 73206 11579 73208
rect 11513 73203 11579 73206
rect 14365 73266 14431 73269
rect 17401 73266 17467 73269
rect 14365 73264 17467 73266
rect 14365 73208 14370 73264
rect 14426 73208 17406 73264
rect 17462 73208 17467 73264
rect 14365 73206 17467 73208
rect 14365 73203 14431 73206
rect 17401 73203 17467 73206
rect 5349 73130 5415 73133
rect 7557 73130 7623 73133
rect 5349 73128 7623 73130
rect 5349 73072 5354 73128
rect 5410 73072 7562 73128
rect 7618 73072 7623 73128
rect 5349 73070 7623 73072
rect 5349 73067 5415 73070
rect 7557 73067 7623 73070
rect 5944 72928 6264 72929
rect 5944 72864 5952 72928
rect 6016 72864 6032 72928
rect 6096 72864 6112 72928
rect 6176 72864 6192 72928
rect 6256 72864 6264 72928
rect 5944 72863 6264 72864
rect 15944 72928 16264 72929
rect 15944 72864 15952 72928
rect 16016 72864 16032 72928
rect 16096 72864 16112 72928
rect 16176 72864 16192 72928
rect 16256 72864 16264 72928
rect 15944 72863 16264 72864
rect 25944 72928 26264 72929
rect 25944 72864 25952 72928
rect 26016 72864 26032 72928
rect 26096 72864 26112 72928
rect 26176 72864 26192 72928
rect 26256 72864 26264 72928
rect 25944 72863 26264 72864
rect 105 72722 171 72725
rect 19701 72722 19767 72725
rect 105 72720 19767 72722
rect 105 72664 110 72720
rect 166 72664 19706 72720
rect 19762 72664 19767 72720
rect 105 72662 19767 72664
rect 105 72659 171 72662
rect 19701 72659 19767 72662
rect 7281 72586 7347 72589
rect 29913 72586 29979 72589
rect 7281 72584 29979 72586
rect 7281 72528 7286 72584
rect 7342 72528 29918 72584
rect 29974 72528 29979 72584
rect 7281 72526 29979 72528
rect 7281 72523 7347 72526
rect 29913 72523 29979 72526
rect 10944 72384 11264 72385
rect 10944 72320 10952 72384
rect 11016 72320 11032 72384
rect 11096 72320 11112 72384
rect 11176 72320 11192 72384
rect 11256 72320 11264 72384
rect 10944 72319 11264 72320
rect 20944 72384 21264 72385
rect 20944 72320 20952 72384
rect 21016 72320 21032 72384
rect 21096 72320 21112 72384
rect 21176 72320 21192 72384
rect 21256 72320 21264 72384
rect 20944 72319 21264 72320
rect 0 72178 800 72208
rect 1761 72178 1827 72181
rect 29200 72178 30000 72208
rect 0 72176 1827 72178
rect 0 72120 1766 72176
rect 1822 72120 1827 72176
rect 0 72118 1827 72120
rect 0 72088 800 72118
rect 1761 72115 1827 72118
rect 26558 72118 30000 72178
rect 5944 71840 6264 71841
rect 5944 71776 5952 71840
rect 6016 71776 6032 71840
rect 6096 71776 6112 71840
rect 6176 71776 6192 71840
rect 6256 71776 6264 71840
rect 5944 71775 6264 71776
rect 15944 71840 16264 71841
rect 15944 71776 15952 71840
rect 16016 71776 16032 71840
rect 16096 71776 16112 71840
rect 16176 71776 16192 71840
rect 16256 71776 16264 71840
rect 15944 71775 16264 71776
rect 25944 71840 26264 71841
rect 25944 71776 25952 71840
rect 26016 71776 26032 71840
rect 26096 71776 26112 71840
rect 26176 71776 26192 71840
rect 26256 71776 26264 71840
rect 25944 71775 26264 71776
rect 26417 71770 26483 71773
rect 26558 71770 26618 72118
rect 29200 72088 30000 72118
rect 26417 71768 26618 71770
rect 26417 71712 26422 71768
rect 26478 71712 26618 71768
rect 26417 71710 26618 71712
rect 26417 71707 26483 71710
rect 0 71498 800 71528
rect 2773 71498 2839 71501
rect 0 71496 2839 71498
rect 0 71440 2778 71496
rect 2834 71440 2839 71496
rect 0 71438 2839 71440
rect 0 71408 800 71438
rect 2773 71435 2839 71438
rect 18781 71498 18847 71501
rect 29200 71498 30000 71528
rect 18781 71496 30000 71498
rect 18781 71440 18786 71496
rect 18842 71440 30000 71496
rect 18781 71438 30000 71440
rect 18781 71435 18847 71438
rect 29200 71408 30000 71438
rect 10944 71296 11264 71297
rect 10944 71232 10952 71296
rect 11016 71232 11032 71296
rect 11096 71232 11112 71296
rect 11176 71232 11192 71296
rect 11256 71232 11264 71296
rect 10944 71231 11264 71232
rect 20944 71296 21264 71297
rect 20944 71232 20952 71296
rect 21016 71232 21032 71296
rect 21096 71232 21112 71296
rect 21176 71232 21192 71296
rect 21256 71232 21264 71296
rect 20944 71231 21264 71232
rect 5533 71090 5599 71093
rect 17585 71090 17651 71093
rect 5533 71088 17651 71090
rect 5533 71032 5538 71088
rect 5594 71032 17590 71088
rect 17646 71032 17651 71088
rect 5533 71030 17651 71032
rect 5533 71027 5599 71030
rect 17585 71027 17651 71030
rect 5944 70752 6264 70753
rect 5944 70688 5952 70752
rect 6016 70688 6032 70752
rect 6096 70688 6112 70752
rect 6176 70688 6192 70752
rect 6256 70688 6264 70752
rect 5944 70687 6264 70688
rect 15944 70752 16264 70753
rect 15944 70688 15952 70752
rect 16016 70688 16032 70752
rect 16096 70688 16112 70752
rect 16176 70688 16192 70752
rect 16256 70688 16264 70752
rect 15944 70687 16264 70688
rect 25944 70752 26264 70753
rect 25944 70688 25952 70752
rect 26016 70688 26032 70752
rect 26096 70688 26112 70752
rect 26176 70688 26192 70752
rect 26256 70688 26264 70752
rect 25944 70687 26264 70688
rect 20897 70546 20963 70549
rect 3374 70544 20963 70546
rect 3374 70488 20902 70544
rect 20958 70488 20963 70544
rect 3374 70486 20963 70488
rect 0 70138 800 70168
rect 3374 70138 3434 70486
rect 20897 70483 20963 70486
rect 12617 70410 12683 70413
rect 18873 70410 18939 70413
rect 12617 70408 18939 70410
rect 12617 70352 12622 70408
rect 12678 70352 18878 70408
rect 18934 70352 18939 70408
rect 12617 70350 18939 70352
rect 12617 70347 12683 70350
rect 18873 70347 18939 70350
rect 10944 70208 11264 70209
rect 10944 70144 10952 70208
rect 11016 70144 11032 70208
rect 11096 70144 11112 70208
rect 11176 70144 11192 70208
rect 11256 70144 11264 70208
rect 10944 70143 11264 70144
rect 20944 70208 21264 70209
rect 20944 70144 20952 70208
rect 21016 70144 21032 70208
rect 21096 70144 21112 70208
rect 21176 70144 21192 70208
rect 21256 70144 21264 70208
rect 20944 70143 21264 70144
rect 0 70078 3434 70138
rect 25497 70138 25563 70141
rect 29200 70138 30000 70168
rect 25497 70136 30000 70138
rect 25497 70080 25502 70136
rect 25558 70080 30000 70136
rect 25497 70078 30000 70080
rect 0 70048 800 70078
rect 25497 70075 25563 70078
rect 29200 70048 30000 70078
rect 5625 69866 5691 69869
rect 21909 69866 21975 69869
rect 5625 69864 21975 69866
rect 5625 69808 5630 69864
rect 5686 69808 21914 69864
rect 21970 69808 21975 69864
rect 5625 69806 21975 69808
rect 5625 69803 5691 69806
rect 21909 69803 21975 69806
rect 21265 69730 21331 69733
rect 22277 69730 22343 69733
rect 21265 69728 22343 69730
rect 21265 69672 21270 69728
rect 21326 69672 22282 69728
rect 22338 69672 22343 69728
rect 21265 69670 22343 69672
rect 21265 69667 21331 69670
rect 22277 69667 22343 69670
rect 5944 69664 6264 69665
rect 5944 69600 5952 69664
rect 6016 69600 6032 69664
rect 6096 69600 6112 69664
rect 6176 69600 6192 69664
rect 6256 69600 6264 69664
rect 5944 69599 6264 69600
rect 15944 69664 16264 69665
rect 15944 69600 15952 69664
rect 16016 69600 16032 69664
rect 16096 69600 16112 69664
rect 16176 69600 16192 69664
rect 16256 69600 16264 69664
rect 15944 69599 16264 69600
rect 25944 69664 26264 69665
rect 25944 69600 25952 69664
rect 26016 69600 26032 69664
rect 26096 69600 26112 69664
rect 26176 69600 26192 69664
rect 26256 69600 26264 69664
rect 25944 69599 26264 69600
rect 2037 69458 2103 69461
rect 9121 69458 9187 69461
rect 10777 69458 10843 69461
rect 2037 69456 10843 69458
rect 2037 69400 2042 69456
rect 2098 69400 9126 69456
rect 9182 69400 10782 69456
rect 10838 69400 10843 69456
rect 2037 69398 10843 69400
rect 2037 69395 2103 69398
rect 9121 69395 9187 69398
rect 10777 69395 10843 69398
rect 1669 69322 1735 69325
rect 17166 69322 17172 69324
rect 1669 69320 17172 69322
rect 1669 69264 1674 69320
rect 1730 69264 17172 69320
rect 1669 69262 17172 69264
rect 1669 69259 1735 69262
rect 17166 69260 17172 69262
rect 17236 69260 17242 69324
rect 10944 69120 11264 69121
rect 10944 69056 10952 69120
rect 11016 69056 11032 69120
rect 11096 69056 11112 69120
rect 11176 69056 11192 69120
rect 11256 69056 11264 69120
rect 10944 69055 11264 69056
rect 20944 69120 21264 69121
rect 20944 69056 20952 69120
rect 21016 69056 21032 69120
rect 21096 69056 21112 69120
rect 21176 69056 21192 69120
rect 21256 69056 21264 69120
rect 20944 69055 21264 69056
rect 16573 69050 16639 69053
rect 20713 69050 20779 69053
rect 16573 69048 20779 69050
rect 16573 68992 16578 69048
rect 16634 68992 20718 69048
rect 20774 68992 20779 69048
rect 16573 68990 20779 68992
rect 16573 68987 16639 68990
rect 20713 68987 20779 68990
rect 24485 69050 24551 69053
rect 25221 69050 25287 69053
rect 24485 69048 25287 69050
rect 24485 68992 24490 69048
rect 24546 68992 25226 69048
rect 25282 68992 25287 69048
rect 24485 68990 25287 68992
rect 24485 68987 24551 68990
rect 25221 68987 25287 68990
rect 11513 68914 11579 68917
rect 15193 68914 15259 68917
rect 11513 68912 15259 68914
rect 11513 68856 11518 68912
rect 11574 68856 15198 68912
rect 15254 68856 15259 68912
rect 11513 68854 15259 68856
rect 11513 68851 11579 68854
rect 15193 68851 15259 68854
rect 19057 68914 19123 68917
rect 25129 68914 25195 68917
rect 19057 68912 25195 68914
rect 19057 68856 19062 68912
rect 19118 68856 25134 68912
rect 25190 68856 25195 68912
rect 19057 68854 25195 68856
rect 19057 68851 19123 68854
rect 25129 68851 25195 68854
rect 0 68778 800 68808
rect 3233 68778 3299 68781
rect 0 68776 3299 68778
rect 0 68720 3238 68776
rect 3294 68720 3299 68776
rect 0 68718 3299 68720
rect 0 68688 800 68718
rect 3233 68715 3299 68718
rect 25630 68716 25636 68780
rect 25700 68778 25706 68780
rect 29200 68778 30000 68808
rect 25700 68718 30000 68778
rect 25700 68716 25706 68718
rect 29200 68688 30000 68718
rect 5944 68576 6264 68577
rect 5944 68512 5952 68576
rect 6016 68512 6032 68576
rect 6096 68512 6112 68576
rect 6176 68512 6192 68576
rect 6256 68512 6264 68576
rect 5944 68511 6264 68512
rect 15944 68576 16264 68577
rect 15944 68512 15952 68576
rect 16016 68512 16032 68576
rect 16096 68512 16112 68576
rect 16176 68512 16192 68576
rect 16256 68512 16264 68576
rect 15944 68511 16264 68512
rect 25944 68576 26264 68577
rect 25944 68512 25952 68576
rect 26016 68512 26032 68576
rect 26096 68512 26112 68576
rect 26176 68512 26192 68576
rect 26256 68512 26264 68576
rect 25944 68511 26264 68512
rect 0 68098 800 68128
rect 29200 68098 30000 68128
rect 0 68008 858 68098
rect 25638 68038 30000 68098
rect 798 67690 858 68008
rect 10944 68032 11264 68033
rect 10944 67968 10952 68032
rect 11016 67968 11032 68032
rect 11096 67968 11112 68032
rect 11176 67968 11192 68032
rect 11256 67968 11264 68032
rect 10944 67967 11264 67968
rect 20944 68032 21264 68033
rect 20944 67968 20952 68032
rect 21016 67968 21032 68032
rect 21096 67968 21112 68032
rect 21176 67968 21192 68032
rect 21256 67968 21264 68032
rect 20944 67967 21264 67968
rect 17677 67826 17743 67829
rect 25497 67826 25563 67829
rect 17677 67824 25563 67826
rect 17677 67768 17682 67824
rect 17738 67768 25502 67824
rect 25558 67768 25563 67824
rect 17677 67766 25563 67768
rect 17677 67763 17743 67766
rect 25497 67763 25563 67766
rect 11237 67690 11303 67693
rect 798 67688 11303 67690
rect 798 67632 11242 67688
rect 11298 67632 11303 67688
rect 798 67630 11303 67632
rect 11237 67627 11303 67630
rect 11605 67690 11671 67693
rect 11973 67690 12039 67693
rect 21449 67690 21515 67693
rect 11605 67688 11714 67690
rect 11605 67632 11610 67688
rect 11666 67632 11714 67688
rect 11605 67627 11714 67632
rect 11973 67688 21515 67690
rect 11973 67632 11978 67688
rect 12034 67632 21454 67688
rect 21510 67632 21515 67688
rect 11973 67630 21515 67632
rect 11973 67627 12039 67630
rect 21449 67627 21515 67630
rect 5944 67488 6264 67489
rect 5944 67424 5952 67488
rect 6016 67424 6032 67488
rect 6096 67424 6112 67488
rect 6176 67424 6192 67488
rect 6256 67424 6264 67488
rect 5944 67423 6264 67424
rect 11513 67418 11579 67421
rect 11654 67418 11714 67627
rect 12249 67554 12315 67557
rect 15377 67554 15443 67557
rect 12249 67552 15443 67554
rect 12249 67496 12254 67552
rect 12310 67496 15382 67552
rect 15438 67496 15443 67552
rect 12249 67494 15443 67496
rect 12249 67491 12315 67494
rect 15377 67491 15443 67494
rect 18597 67554 18663 67557
rect 25638 67554 25698 68038
rect 29200 68008 30000 68038
rect 18597 67552 25698 67554
rect 18597 67496 18602 67552
rect 18658 67496 25698 67552
rect 18597 67494 25698 67496
rect 18597 67491 18663 67494
rect 15944 67488 16264 67489
rect 15944 67424 15952 67488
rect 16016 67424 16032 67488
rect 16096 67424 16112 67488
rect 16176 67424 16192 67488
rect 16256 67424 16264 67488
rect 15944 67423 16264 67424
rect 25944 67488 26264 67489
rect 25944 67424 25952 67488
rect 26016 67424 26032 67488
rect 26096 67424 26112 67488
rect 26176 67424 26192 67488
rect 26256 67424 26264 67488
rect 25944 67423 26264 67424
rect 11513 67416 11714 67418
rect 11513 67360 11518 67416
rect 11574 67360 11714 67416
rect 11513 67358 11714 67360
rect 11513 67355 11579 67358
rect 10944 66944 11264 66945
rect 10944 66880 10952 66944
rect 11016 66880 11032 66944
rect 11096 66880 11112 66944
rect 11176 66880 11192 66944
rect 11256 66880 11264 66944
rect 10944 66879 11264 66880
rect 20944 66944 21264 66945
rect 20944 66880 20952 66944
rect 21016 66880 21032 66944
rect 21096 66880 21112 66944
rect 21176 66880 21192 66944
rect 21256 66880 21264 66944
rect 20944 66879 21264 66880
rect 0 66738 800 66768
rect 4061 66738 4127 66741
rect 0 66736 4127 66738
rect 0 66680 4066 66736
rect 4122 66680 4127 66736
rect 0 66678 4127 66680
rect 0 66648 800 66678
rect 4061 66675 4127 66678
rect 25497 66738 25563 66741
rect 29200 66738 30000 66768
rect 25497 66736 30000 66738
rect 25497 66680 25502 66736
rect 25558 66680 30000 66736
rect 25497 66678 30000 66680
rect 25497 66675 25563 66678
rect 29200 66648 30000 66678
rect 5944 66400 6264 66401
rect 5944 66336 5952 66400
rect 6016 66336 6032 66400
rect 6096 66336 6112 66400
rect 6176 66336 6192 66400
rect 6256 66336 6264 66400
rect 5944 66335 6264 66336
rect 15944 66400 16264 66401
rect 15944 66336 15952 66400
rect 16016 66336 16032 66400
rect 16096 66336 16112 66400
rect 16176 66336 16192 66400
rect 16256 66336 16264 66400
rect 15944 66335 16264 66336
rect 25944 66400 26264 66401
rect 25944 66336 25952 66400
rect 26016 66336 26032 66400
rect 26096 66336 26112 66400
rect 26176 66336 26192 66400
rect 26256 66336 26264 66400
rect 25944 66335 26264 66336
rect 8201 66194 8267 66197
rect 15101 66194 15167 66197
rect 8201 66192 15167 66194
rect 8201 66136 8206 66192
rect 8262 66136 15106 66192
rect 15162 66136 15167 66192
rect 8201 66134 15167 66136
rect 8201 66131 8267 66134
rect 15101 66131 15167 66134
rect 27838 66132 27844 66196
rect 27908 66194 27914 66196
rect 27981 66194 28047 66197
rect 27908 66192 28047 66194
rect 27908 66136 27986 66192
rect 28042 66136 28047 66192
rect 27908 66134 28047 66136
rect 27908 66132 27914 66134
rect 27981 66131 28047 66134
rect 4061 66058 4127 66061
rect 17769 66058 17835 66061
rect 4061 66056 17835 66058
rect 4061 66000 4066 66056
rect 4122 66000 17774 66056
rect 17830 66000 17835 66056
rect 4061 65998 17835 66000
rect 4061 65995 4127 65998
rect 17769 65995 17835 65998
rect 10944 65856 11264 65857
rect 10944 65792 10952 65856
rect 11016 65792 11032 65856
rect 11096 65792 11112 65856
rect 11176 65792 11192 65856
rect 11256 65792 11264 65856
rect 10944 65791 11264 65792
rect 20944 65856 21264 65857
rect 20944 65792 20952 65856
rect 21016 65792 21032 65856
rect 21096 65792 21112 65856
rect 21176 65792 21192 65856
rect 21256 65792 21264 65856
rect 20944 65791 21264 65792
rect 18689 65514 18755 65517
rect 21950 65514 21956 65516
rect 18689 65512 21956 65514
rect 18689 65456 18694 65512
rect 18750 65456 21956 65512
rect 18689 65454 21956 65456
rect 18689 65451 18755 65454
rect 21950 65452 21956 65454
rect 22020 65452 22026 65516
rect 0 65378 800 65408
rect 29200 65378 30000 65408
rect 0 65288 858 65378
rect 26374 65318 30000 65378
rect 798 65242 858 65288
rect 5944 65312 6264 65313
rect 5944 65248 5952 65312
rect 6016 65248 6032 65312
rect 6096 65248 6112 65312
rect 6176 65248 6192 65312
rect 6256 65248 6264 65312
rect 5944 65247 6264 65248
rect 15944 65312 16264 65313
rect 15944 65248 15952 65312
rect 16016 65248 16032 65312
rect 16096 65248 16112 65312
rect 16176 65248 16192 65312
rect 16256 65248 16264 65312
rect 15944 65247 16264 65248
rect 25944 65312 26264 65313
rect 25944 65248 25952 65312
rect 26016 65248 26032 65312
rect 26096 65248 26112 65312
rect 26176 65248 26192 65312
rect 26256 65248 26264 65312
rect 25944 65247 26264 65248
rect 4797 65242 4863 65245
rect 798 65240 4863 65242
rect 798 65184 4802 65240
rect 4858 65184 4863 65240
rect 798 65182 4863 65184
rect 4797 65179 4863 65182
rect 25589 65106 25655 65109
rect 26374 65106 26434 65318
rect 29200 65288 30000 65318
rect 25589 65104 26434 65106
rect 25589 65048 25594 65104
rect 25650 65048 26434 65104
rect 25589 65046 26434 65048
rect 25589 65043 25655 65046
rect 15469 64970 15535 64973
rect 18229 64970 18295 64973
rect 15469 64968 18295 64970
rect 15469 64912 15474 64968
rect 15530 64912 18234 64968
rect 18290 64912 18295 64968
rect 15469 64910 18295 64912
rect 15469 64907 15535 64910
rect 18229 64907 18295 64910
rect 10944 64768 11264 64769
rect 10944 64704 10952 64768
rect 11016 64704 11032 64768
rect 11096 64704 11112 64768
rect 11176 64704 11192 64768
rect 11256 64704 11264 64768
rect 10944 64703 11264 64704
rect 20944 64768 21264 64769
rect 20944 64704 20952 64768
rect 21016 64704 21032 64768
rect 21096 64704 21112 64768
rect 21176 64704 21192 64768
rect 21256 64704 21264 64768
rect 20944 64703 21264 64704
rect 25865 64698 25931 64701
rect 29200 64698 30000 64728
rect 25865 64696 30000 64698
rect 25865 64640 25870 64696
rect 25926 64640 30000 64696
rect 25865 64638 30000 64640
rect 25865 64635 25931 64638
rect 29200 64608 30000 64638
rect 4797 64562 4863 64565
rect 21582 64562 21588 64564
rect 4797 64560 21588 64562
rect 4797 64504 4802 64560
rect 4858 64504 21588 64560
rect 4797 64502 21588 64504
rect 4797 64499 4863 64502
rect 21582 64500 21588 64502
rect 21652 64500 21658 64564
rect 5944 64224 6264 64225
rect 5944 64160 5952 64224
rect 6016 64160 6032 64224
rect 6096 64160 6112 64224
rect 6176 64160 6192 64224
rect 6256 64160 6264 64224
rect 5944 64159 6264 64160
rect 15944 64224 16264 64225
rect 15944 64160 15952 64224
rect 16016 64160 16032 64224
rect 16096 64160 16112 64224
rect 16176 64160 16192 64224
rect 16256 64160 16264 64224
rect 15944 64159 16264 64160
rect 25944 64224 26264 64225
rect 25944 64160 25952 64224
rect 26016 64160 26032 64224
rect 26096 64160 26112 64224
rect 26176 64160 26192 64224
rect 26256 64160 26264 64224
rect 25944 64159 26264 64160
rect 0 64018 800 64048
rect 18597 64018 18663 64021
rect 0 64016 18663 64018
rect 0 63960 18602 64016
rect 18658 63960 18663 64016
rect 0 63958 18663 63960
rect 0 63928 800 63958
rect 18597 63955 18663 63958
rect 18873 64018 18939 64021
rect 20713 64018 20779 64021
rect 21633 64018 21699 64021
rect 18873 64016 21699 64018
rect 18873 63960 18878 64016
rect 18934 63960 20718 64016
rect 20774 63960 21638 64016
rect 21694 63960 21699 64016
rect 18873 63958 21699 63960
rect 18873 63955 18939 63958
rect 20713 63955 20779 63958
rect 21633 63955 21699 63958
rect 10944 63680 11264 63681
rect 10944 63616 10952 63680
rect 11016 63616 11032 63680
rect 11096 63616 11112 63680
rect 11176 63616 11192 63680
rect 11256 63616 11264 63680
rect 10944 63615 11264 63616
rect 20944 63680 21264 63681
rect 20944 63616 20952 63680
rect 21016 63616 21032 63680
rect 21096 63616 21112 63680
rect 21176 63616 21192 63680
rect 21256 63616 21264 63680
rect 20944 63615 21264 63616
rect 21817 63610 21883 63613
rect 27521 63610 27587 63613
rect 21817 63608 27587 63610
rect 21817 63552 21822 63608
rect 21878 63552 27526 63608
rect 27582 63552 27587 63608
rect 21817 63550 27587 63552
rect 21817 63547 21883 63550
rect 27521 63547 27587 63550
rect 16757 63474 16823 63477
rect 18781 63474 18847 63477
rect 16757 63472 18847 63474
rect 16757 63416 16762 63472
rect 16818 63416 18786 63472
rect 18842 63416 18847 63472
rect 16757 63414 18847 63416
rect 16757 63411 16823 63414
rect 18781 63411 18847 63414
rect 0 63338 800 63368
rect 3785 63338 3851 63341
rect 0 63336 3851 63338
rect 0 63280 3790 63336
rect 3846 63280 3851 63336
rect 0 63278 3851 63280
rect 0 63248 800 63278
rect 3785 63275 3851 63278
rect 25773 63338 25839 63341
rect 29200 63338 30000 63368
rect 25773 63336 30000 63338
rect 25773 63280 25778 63336
rect 25834 63280 30000 63336
rect 25773 63278 30000 63280
rect 25773 63275 25839 63278
rect 29200 63248 30000 63278
rect 5944 63136 6264 63137
rect 5944 63072 5952 63136
rect 6016 63072 6032 63136
rect 6096 63072 6112 63136
rect 6176 63072 6192 63136
rect 6256 63072 6264 63136
rect 5944 63071 6264 63072
rect 15944 63136 16264 63137
rect 15944 63072 15952 63136
rect 16016 63072 16032 63136
rect 16096 63072 16112 63136
rect 16176 63072 16192 63136
rect 16256 63072 16264 63136
rect 15944 63071 16264 63072
rect 25944 63136 26264 63137
rect 25944 63072 25952 63136
rect 26016 63072 26032 63136
rect 26096 63072 26112 63136
rect 26176 63072 26192 63136
rect 26256 63072 26264 63136
rect 25944 63071 26264 63072
rect 18086 62868 18092 62932
rect 18156 62930 18162 62932
rect 25589 62930 25655 62933
rect 18156 62928 25655 62930
rect 18156 62872 25594 62928
rect 25650 62872 25655 62928
rect 18156 62870 25655 62872
rect 18156 62868 18162 62870
rect 25589 62867 25655 62870
rect 3417 62794 3483 62797
rect 17953 62794 18019 62797
rect 3417 62792 18019 62794
rect 3417 62736 3422 62792
rect 3478 62736 17958 62792
rect 18014 62736 18019 62792
rect 3417 62734 18019 62736
rect 3417 62731 3483 62734
rect 17953 62731 18019 62734
rect 10944 62592 11264 62593
rect 10944 62528 10952 62592
rect 11016 62528 11032 62592
rect 11096 62528 11112 62592
rect 11176 62528 11192 62592
rect 11256 62528 11264 62592
rect 10944 62527 11264 62528
rect 20944 62592 21264 62593
rect 20944 62528 20952 62592
rect 21016 62528 21032 62592
rect 21096 62528 21112 62592
rect 21176 62528 21192 62592
rect 21256 62528 21264 62592
rect 20944 62527 21264 62528
rect 20345 62386 20411 62389
rect 22921 62386 22987 62389
rect 20345 62384 22987 62386
rect 20345 62328 20350 62384
rect 20406 62328 22926 62384
rect 22982 62328 22987 62384
rect 20345 62326 22987 62328
rect 20345 62323 20411 62326
rect 22921 62323 22987 62326
rect 20161 62250 20227 62253
rect 22185 62250 22251 62253
rect 20161 62248 22251 62250
rect 20161 62192 20166 62248
rect 20222 62192 22190 62248
rect 22246 62192 22251 62248
rect 20161 62190 22251 62192
rect 20161 62187 20227 62190
rect 22185 62187 22251 62190
rect 5944 62048 6264 62049
rect 0 61978 800 62008
rect 5944 61984 5952 62048
rect 6016 61984 6032 62048
rect 6096 61984 6112 62048
rect 6176 61984 6192 62048
rect 6256 61984 6264 62048
rect 5944 61983 6264 61984
rect 15944 62048 16264 62049
rect 15944 61984 15952 62048
rect 16016 61984 16032 62048
rect 16096 61984 16112 62048
rect 16176 61984 16192 62048
rect 16256 61984 16264 62048
rect 15944 61983 16264 61984
rect 25944 62048 26264 62049
rect 25944 61984 25952 62048
rect 26016 61984 26032 62048
rect 26096 61984 26112 62048
rect 26176 61984 26192 62048
rect 26256 61984 26264 62048
rect 25944 61983 26264 61984
rect 2773 61978 2839 61981
rect 0 61976 2839 61978
rect 0 61920 2778 61976
rect 2834 61920 2839 61976
rect 0 61918 2839 61920
rect 0 61888 800 61918
rect 2773 61915 2839 61918
rect 26693 61978 26759 61981
rect 29200 61978 30000 62008
rect 26693 61976 30000 61978
rect 26693 61920 26698 61976
rect 26754 61920 30000 61976
rect 26693 61918 30000 61920
rect 26693 61915 26759 61918
rect 29200 61888 30000 61918
rect 22737 61842 22803 61845
rect 25589 61842 25655 61845
rect 22737 61840 25655 61842
rect 22737 61784 22742 61840
rect 22798 61784 25594 61840
rect 25650 61784 25655 61840
rect 22737 61782 25655 61784
rect 22737 61779 22803 61782
rect 25589 61779 25655 61782
rect 10944 61504 11264 61505
rect 10944 61440 10952 61504
rect 11016 61440 11032 61504
rect 11096 61440 11112 61504
rect 11176 61440 11192 61504
rect 11256 61440 11264 61504
rect 10944 61439 11264 61440
rect 20944 61504 21264 61505
rect 20944 61440 20952 61504
rect 21016 61440 21032 61504
rect 21096 61440 21112 61504
rect 21176 61440 21192 61504
rect 21256 61440 21264 61504
rect 20944 61439 21264 61440
rect 24945 61298 25011 61301
rect 29200 61298 30000 61328
rect 24945 61296 30000 61298
rect 24945 61240 24950 61296
rect 25006 61240 30000 61296
rect 24945 61238 30000 61240
rect 24945 61235 25011 61238
rect 29200 61208 30000 61238
rect 5944 60960 6264 60961
rect 5944 60896 5952 60960
rect 6016 60896 6032 60960
rect 6096 60896 6112 60960
rect 6176 60896 6192 60960
rect 6256 60896 6264 60960
rect 5944 60895 6264 60896
rect 15944 60960 16264 60961
rect 15944 60896 15952 60960
rect 16016 60896 16032 60960
rect 16096 60896 16112 60960
rect 16176 60896 16192 60960
rect 16256 60896 16264 60960
rect 15944 60895 16264 60896
rect 25944 60960 26264 60961
rect 25944 60896 25952 60960
rect 26016 60896 26032 60960
rect 26096 60896 26112 60960
rect 26176 60896 26192 60960
rect 26256 60896 26264 60960
rect 25944 60895 26264 60896
rect 5441 60754 5507 60757
rect 18873 60754 18939 60757
rect 5441 60752 18939 60754
rect 5441 60696 5446 60752
rect 5502 60696 18878 60752
rect 18934 60696 18939 60752
rect 5441 60694 18939 60696
rect 5441 60691 5507 60694
rect 18873 60691 18939 60694
rect 0 60618 800 60648
rect 7925 60618 7991 60621
rect 0 60616 7991 60618
rect 0 60560 7930 60616
rect 7986 60560 7991 60616
rect 0 60558 7991 60560
rect 0 60528 800 60558
rect 7925 60555 7991 60558
rect 10944 60416 11264 60417
rect 10944 60352 10952 60416
rect 11016 60352 11032 60416
rect 11096 60352 11112 60416
rect 11176 60352 11192 60416
rect 11256 60352 11264 60416
rect 10944 60351 11264 60352
rect 20944 60416 21264 60417
rect 20944 60352 20952 60416
rect 21016 60352 21032 60416
rect 21096 60352 21112 60416
rect 21176 60352 21192 60416
rect 21256 60352 21264 60416
rect 20944 60351 21264 60352
rect 0 59938 800 59968
rect 2865 59938 2931 59941
rect 29200 59938 30000 59968
rect 0 59936 2931 59938
rect 0 59880 2870 59936
rect 2926 59880 2931 59936
rect 0 59878 2931 59880
rect 0 59848 800 59878
rect 2865 59875 2931 59878
rect 26374 59878 30000 59938
rect 5944 59872 6264 59873
rect 5944 59808 5952 59872
rect 6016 59808 6032 59872
rect 6096 59808 6112 59872
rect 6176 59808 6192 59872
rect 6256 59808 6264 59872
rect 5944 59807 6264 59808
rect 15944 59872 16264 59873
rect 15944 59808 15952 59872
rect 16016 59808 16032 59872
rect 16096 59808 16112 59872
rect 16176 59808 16192 59872
rect 16256 59808 16264 59872
rect 15944 59807 16264 59808
rect 25944 59872 26264 59873
rect 25944 59808 25952 59872
rect 26016 59808 26032 59872
rect 26096 59808 26112 59872
rect 26176 59808 26192 59872
rect 26256 59808 26264 59872
rect 25944 59807 26264 59808
rect 25773 59666 25839 59669
rect 26374 59666 26434 59878
rect 29200 59848 30000 59878
rect 25773 59664 26434 59666
rect 25773 59608 25778 59664
rect 25834 59608 26434 59664
rect 25773 59606 26434 59608
rect 25773 59603 25839 59606
rect 16205 59530 16271 59533
rect 16665 59530 16731 59533
rect 18229 59530 18295 59533
rect 16205 59528 18295 59530
rect 16205 59472 16210 59528
rect 16266 59472 16670 59528
rect 16726 59472 18234 59528
rect 18290 59472 18295 59528
rect 16205 59470 18295 59472
rect 16205 59467 16271 59470
rect 16665 59467 16731 59470
rect 18229 59467 18295 59470
rect 14457 59394 14523 59397
rect 17033 59394 17099 59397
rect 14457 59392 17099 59394
rect 14457 59336 14462 59392
rect 14518 59336 17038 59392
rect 17094 59336 17099 59392
rect 14457 59334 17099 59336
rect 14457 59331 14523 59334
rect 17033 59331 17099 59334
rect 24577 59394 24643 59397
rect 26509 59394 26575 59397
rect 24577 59392 26575 59394
rect 24577 59336 24582 59392
rect 24638 59336 26514 59392
rect 26570 59336 26575 59392
rect 24577 59334 26575 59336
rect 24577 59331 24643 59334
rect 26509 59331 26575 59334
rect 10944 59328 11264 59329
rect 10944 59264 10952 59328
rect 11016 59264 11032 59328
rect 11096 59264 11112 59328
rect 11176 59264 11192 59328
rect 11256 59264 11264 59328
rect 10944 59263 11264 59264
rect 20944 59328 21264 59329
rect 20944 59264 20952 59328
rect 21016 59264 21032 59328
rect 21096 59264 21112 59328
rect 21176 59264 21192 59328
rect 21256 59264 21264 59328
rect 20944 59263 21264 59264
rect 16573 59258 16639 59261
rect 19149 59258 19215 59261
rect 16573 59256 19215 59258
rect 16573 59200 16578 59256
rect 16634 59200 19154 59256
rect 19210 59200 19215 59256
rect 16573 59198 19215 59200
rect 16573 59195 16639 59198
rect 19149 59195 19215 59198
rect 14365 59122 14431 59125
rect 17585 59122 17651 59125
rect 14365 59120 17651 59122
rect 14365 59064 14370 59120
rect 14426 59064 17590 59120
rect 17646 59064 17651 59120
rect 14365 59062 17651 59064
rect 14365 59059 14431 59062
rect 17585 59059 17651 59062
rect 22645 59122 22711 59125
rect 23473 59122 23539 59125
rect 22645 59120 23539 59122
rect 22645 59064 22650 59120
rect 22706 59064 23478 59120
rect 23534 59064 23539 59120
rect 22645 59062 23539 59064
rect 22645 59059 22711 59062
rect 23473 59059 23539 59062
rect 17769 58986 17835 58989
rect 19609 58986 19675 58989
rect 17769 58984 19675 58986
rect 17769 58928 17774 58984
rect 17830 58928 19614 58984
rect 19670 58928 19675 58984
rect 17769 58926 19675 58928
rect 17769 58923 17835 58926
rect 19609 58923 19675 58926
rect 18965 58850 19031 58853
rect 20253 58850 20319 58853
rect 18965 58848 20319 58850
rect 18965 58792 18970 58848
rect 19026 58792 20258 58848
rect 20314 58792 20319 58848
rect 18965 58790 20319 58792
rect 18965 58787 19031 58790
rect 20253 58787 20319 58790
rect 5944 58784 6264 58785
rect 5944 58720 5952 58784
rect 6016 58720 6032 58784
rect 6096 58720 6112 58784
rect 6176 58720 6192 58784
rect 6256 58720 6264 58784
rect 5944 58719 6264 58720
rect 15944 58784 16264 58785
rect 15944 58720 15952 58784
rect 16016 58720 16032 58784
rect 16096 58720 16112 58784
rect 16176 58720 16192 58784
rect 16256 58720 16264 58784
rect 15944 58719 16264 58720
rect 25944 58784 26264 58785
rect 25944 58720 25952 58784
rect 26016 58720 26032 58784
rect 26096 58720 26112 58784
rect 26176 58720 26192 58784
rect 26256 58720 26264 58784
rect 25944 58719 26264 58720
rect 0 58578 800 58608
rect 3049 58578 3115 58581
rect 0 58576 3115 58578
rect 0 58520 3054 58576
rect 3110 58520 3115 58576
rect 0 58518 3115 58520
rect 0 58488 800 58518
rect 3049 58515 3115 58518
rect 14641 58578 14707 58581
rect 16205 58578 16271 58581
rect 17953 58578 18019 58581
rect 14641 58576 18019 58578
rect 14641 58520 14646 58576
rect 14702 58520 16210 58576
rect 16266 58520 17958 58576
rect 18014 58520 18019 58576
rect 14641 58518 18019 58520
rect 14641 58515 14707 58518
rect 16205 58515 16271 58518
rect 17953 58515 18019 58518
rect 21541 58578 21607 58581
rect 29200 58578 30000 58608
rect 21541 58576 30000 58578
rect 21541 58520 21546 58576
rect 21602 58520 30000 58576
rect 21541 58518 30000 58520
rect 21541 58515 21607 58518
rect 29200 58488 30000 58518
rect 21265 58442 21331 58445
rect 23933 58442 23999 58445
rect 21265 58440 23999 58442
rect 21265 58384 21270 58440
rect 21326 58384 23938 58440
rect 23994 58384 23999 58440
rect 21265 58382 23999 58384
rect 21265 58379 21331 58382
rect 23933 58379 23999 58382
rect 14825 58306 14891 58309
rect 16573 58306 16639 58309
rect 14825 58304 16639 58306
rect 14825 58248 14830 58304
rect 14886 58248 16578 58304
rect 16634 58248 16639 58304
rect 14825 58246 16639 58248
rect 14825 58243 14891 58246
rect 16573 58243 16639 58246
rect 10944 58240 11264 58241
rect 10944 58176 10952 58240
rect 11016 58176 11032 58240
rect 11096 58176 11112 58240
rect 11176 58176 11192 58240
rect 11256 58176 11264 58240
rect 10944 58175 11264 58176
rect 20944 58240 21264 58241
rect 20944 58176 20952 58240
rect 21016 58176 21032 58240
rect 21096 58176 21112 58240
rect 21176 58176 21192 58240
rect 21256 58176 21264 58240
rect 20944 58175 21264 58176
rect 11513 58036 11579 58037
rect 11462 58034 11468 58036
rect 11422 57974 11468 58034
rect 11532 58032 11579 58036
rect 11574 57976 11579 58032
rect 11462 57972 11468 57974
rect 11532 57972 11579 57976
rect 11513 57971 11579 57972
rect 19333 58032 19399 58037
rect 19333 57976 19338 58032
rect 19394 57976 19399 58032
rect 19333 57971 19399 57976
rect 3325 57898 3391 57901
rect 7005 57898 7071 57901
rect 3325 57896 7071 57898
rect 3325 57840 3330 57896
rect 3386 57840 7010 57896
rect 7066 57840 7071 57896
rect 3325 57838 7071 57840
rect 3325 57835 3391 57838
rect 7005 57835 7071 57838
rect 15377 57898 15443 57901
rect 19336 57898 19396 57971
rect 20713 57898 20779 57901
rect 15377 57896 20779 57898
rect 15377 57840 15382 57896
rect 15438 57840 20718 57896
rect 20774 57840 20779 57896
rect 15377 57838 20779 57840
rect 15377 57835 15443 57838
rect 20713 57835 20779 57838
rect 17493 57762 17559 57765
rect 18505 57762 18571 57765
rect 17493 57760 18571 57762
rect 17493 57704 17498 57760
rect 17554 57704 18510 57760
rect 18566 57704 18571 57760
rect 17493 57702 18571 57704
rect 17493 57699 17559 57702
rect 18505 57699 18571 57702
rect 18689 57762 18755 57765
rect 22553 57762 22619 57765
rect 18689 57760 22619 57762
rect 18689 57704 18694 57760
rect 18750 57704 22558 57760
rect 22614 57704 22619 57760
rect 18689 57702 22619 57704
rect 18689 57699 18755 57702
rect 22553 57699 22619 57702
rect 5944 57696 6264 57697
rect 5944 57632 5952 57696
rect 6016 57632 6032 57696
rect 6096 57632 6112 57696
rect 6176 57632 6192 57696
rect 6256 57632 6264 57696
rect 5944 57631 6264 57632
rect 15944 57696 16264 57697
rect 15944 57632 15952 57696
rect 16016 57632 16032 57696
rect 16096 57632 16112 57696
rect 16176 57632 16192 57696
rect 16256 57632 16264 57696
rect 15944 57631 16264 57632
rect 25944 57696 26264 57697
rect 25944 57632 25952 57696
rect 26016 57632 26032 57696
rect 26096 57632 26112 57696
rect 26176 57632 26192 57696
rect 26256 57632 26264 57696
rect 25944 57631 26264 57632
rect 2681 57490 2747 57493
rect 2681 57488 11530 57490
rect 2681 57432 2686 57488
rect 2742 57432 11530 57488
rect 2681 57430 11530 57432
rect 2681 57427 2747 57430
rect 0 57218 800 57248
rect 1669 57218 1735 57221
rect 0 57216 1735 57218
rect 0 57160 1674 57216
rect 1730 57160 1735 57216
rect 0 57158 1735 57160
rect 0 57128 800 57158
rect 1669 57155 1735 57158
rect 2221 57218 2287 57221
rect 3325 57218 3391 57221
rect 2221 57216 3391 57218
rect 2221 57160 2226 57216
rect 2282 57160 3330 57216
rect 3386 57160 3391 57216
rect 2221 57158 3391 57160
rect 2221 57155 2287 57158
rect 3325 57155 3391 57158
rect 3601 57218 3667 57221
rect 8753 57218 8819 57221
rect 3601 57216 8819 57218
rect 3601 57160 3606 57216
rect 3662 57160 8758 57216
rect 8814 57160 8819 57216
rect 3601 57158 8819 57160
rect 11470 57218 11530 57430
rect 20478 57292 20484 57356
rect 20548 57354 20554 57356
rect 20989 57354 21055 57357
rect 20548 57352 21055 57354
rect 20548 57296 20994 57352
rect 21050 57296 21055 57352
rect 20548 57294 21055 57296
rect 20548 57292 20554 57294
rect 20989 57291 21055 57294
rect 17309 57218 17375 57221
rect 11470 57216 17375 57218
rect 11470 57160 17314 57216
rect 17370 57160 17375 57216
rect 11470 57158 17375 57160
rect 3601 57155 3667 57158
rect 8753 57155 8819 57158
rect 17309 57155 17375 57158
rect 21817 57218 21883 57221
rect 29200 57218 30000 57248
rect 21817 57216 30000 57218
rect 21817 57160 21822 57216
rect 21878 57160 30000 57216
rect 21817 57158 30000 57160
rect 21817 57155 21883 57158
rect 10944 57152 11264 57153
rect 10944 57088 10952 57152
rect 11016 57088 11032 57152
rect 11096 57088 11112 57152
rect 11176 57088 11192 57152
rect 11256 57088 11264 57152
rect 10944 57087 11264 57088
rect 20944 57152 21264 57153
rect 20944 57088 20952 57152
rect 21016 57088 21032 57152
rect 21096 57088 21112 57152
rect 21176 57088 21192 57152
rect 21256 57088 21264 57152
rect 29200 57128 30000 57158
rect 20944 57087 21264 57088
rect 14641 57082 14707 57085
rect 19333 57082 19399 57085
rect 14641 57080 19399 57082
rect 14641 57024 14646 57080
rect 14702 57024 19338 57080
rect 19394 57024 19399 57080
rect 14641 57022 19399 57024
rect 14641 57019 14707 57022
rect 19333 57019 19399 57022
rect 16665 56946 16731 56949
rect 3558 56944 16731 56946
rect 3558 56888 16670 56944
rect 16726 56888 16731 56944
rect 3558 56886 16731 56888
rect 0 56538 800 56568
rect 3558 56538 3618 56886
rect 16665 56883 16731 56886
rect 12065 56810 12131 56813
rect 12065 56808 17786 56810
rect 12065 56752 12070 56808
rect 12126 56752 17786 56808
rect 12065 56750 17786 56752
rect 12065 56747 12131 56750
rect 15745 56676 15811 56677
rect 15694 56674 15700 56676
rect 15654 56614 15700 56674
rect 15764 56672 15811 56676
rect 15806 56616 15811 56672
rect 15694 56612 15700 56614
rect 15764 56612 15811 56616
rect 15745 56611 15811 56612
rect 5944 56608 6264 56609
rect 5944 56544 5952 56608
rect 6016 56544 6032 56608
rect 6096 56544 6112 56608
rect 6176 56544 6192 56608
rect 6256 56544 6264 56608
rect 5944 56543 6264 56544
rect 15944 56608 16264 56609
rect 15944 56544 15952 56608
rect 16016 56544 16032 56608
rect 16096 56544 16112 56608
rect 16176 56544 16192 56608
rect 16256 56544 16264 56608
rect 15944 56543 16264 56544
rect 0 56478 3618 56538
rect 15469 56538 15535 56541
rect 15745 56538 15811 56541
rect 17726 56540 17786 56750
rect 27838 56612 27844 56676
rect 27908 56674 27914 56676
rect 27981 56674 28047 56677
rect 27908 56672 28047 56674
rect 27908 56616 27986 56672
rect 28042 56616 28047 56672
rect 27908 56614 28047 56616
rect 27908 56612 27914 56614
rect 27981 56611 28047 56614
rect 25944 56608 26264 56609
rect 25944 56544 25952 56608
rect 26016 56544 26032 56608
rect 26096 56544 26112 56608
rect 26176 56544 26192 56608
rect 26256 56544 26264 56608
rect 25944 56543 26264 56544
rect 17718 56538 17724 56540
rect 15469 56536 15811 56538
rect 15469 56480 15474 56536
rect 15530 56480 15750 56536
rect 15806 56480 15811 56536
rect 15469 56478 15811 56480
rect 17596 56478 17724 56538
rect 0 56448 800 56478
rect 15469 56475 15535 56478
rect 15745 56475 15811 56478
rect 17718 56476 17724 56478
rect 17788 56538 17794 56540
rect 19057 56538 19123 56541
rect 17788 56536 19123 56538
rect 17788 56480 19062 56536
rect 19118 56480 19123 56536
rect 17788 56478 19123 56480
rect 17788 56476 17794 56478
rect 19057 56475 19123 56478
rect 20713 56538 20779 56541
rect 22461 56538 22527 56541
rect 29200 56538 30000 56568
rect 20713 56536 22527 56538
rect 20713 56480 20718 56536
rect 20774 56480 22466 56536
rect 22522 56480 22527 56536
rect 20713 56478 22527 56480
rect 20713 56475 20779 56478
rect 22461 56475 22527 56478
rect 26374 56478 30000 56538
rect 13721 56402 13787 56405
rect 14181 56402 14247 56405
rect 16573 56402 16639 56405
rect 20989 56402 21055 56405
rect 13721 56400 16639 56402
rect 13721 56344 13726 56400
rect 13782 56344 14186 56400
rect 14242 56344 16578 56400
rect 16634 56344 16639 56400
rect 13721 56342 16639 56344
rect 13721 56339 13787 56342
rect 14181 56339 14247 56342
rect 16573 56339 16639 56342
rect 18646 56400 21055 56402
rect 18646 56344 20994 56400
rect 21050 56344 21055 56400
rect 18646 56342 21055 56344
rect 13537 56266 13603 56269
rect 14181 56266 14247 56269
rect 18646 56266 18706 56342
rect 20989 56339 21055 56342
rect 25957 56402 26023 56405
rect 26374 56402 26434 56478
rect 29200 56448 30000 56478
rect 25957 56400 26434 56402
rect 25957 56344 25962 56400
rect 26018 56344 26434 56400
rect 25957 56342 26434 56344
rect 25957 56339 26023 56342
rect 13537 56264 18706 56266
rect 13537 56208 13542 56264
rect 13598 56208 14186 56264
rect 14242 56208 18706 56264
rect 13537 56206 18706 56208
rect 18781 56266 18847 56269
rect 20713 56266 20779 56269
rect 18781 56264 20779 56266
rect 18781 56208 18786 56264
rect 18842 56208 20718 56264
rect 20774 56208 20779 56264
rect 18781 56206 20779 56208
rect 13537 56203 13603 56206
rect 14181 56203 14247 56206
rect 18781 56203 18847 56206
rect 20713 56203 20779 56206
rect 13261 56130 13327 56133
rect 16665 56130 16731 56133
rect 13261 56128 16731 56130
rect 13261 56072 13266 56128
rect 13322 56072 16670 56128
rect 16726 56072 16731 56128
rect 13261 56070 16731 56072
rect 13261 56067 13327 56070
rect 16665 56067 16731 56070
rect 10944 56064 11264 56065
rect 10944 56000 10952 56064
rect 11016 56000 11032 56064
rect 11096 56000 11112 56064
rect 11176 56000 11192 56064
rect 11256 56000 11264 56064
rect 10944 55999 11264 56000
rect 20944 56064 21264 56065
rect 20944 56000 20952 56064
rect 21016 56000 21032 56064
rect 21096 56000 21112 56064
rect 21176 56000 21192 56064
rect 21256 56000 21264 56064
rect 20944 55999 21264 56000
rect 3417 55858 3483 55861
rect 12157 55858 12223 55861
rect 3417 55856 12223 55858
rect 3417 55800 3422 55856
rect 3478 55800 12162 55856
rect 12218 55800 12223 55856
rect 3417 55798 12223 55800
rect 3417 55795 3483 55798
rect 12157 55795 12223 55798
rect 14273 55858 14339 55861
rect 16941 55858 17007 55861
rect 14273 55856 17007 55858
rect 14273 55800 14278 55856
rect 14334 55800 16946 55856
rect 17002 55800 17007 55856
rect 14273 55798 17007 55800
rect 14273 55795 14339 55798
rect 16941 55795 17007 55798
rect 17769 55858 17835 55861
rect 20897 55858 20963 55861
rect 17769 55856 20963 55858
rect 17769 55800 17774 55856
rect 17830 55800 20902 55856
rect 20958 55800 20963 55856
rect 17769 55798 20963 55800
rect 17769 55795 17835 55798
rect 20897 55795 20963 55798
rect 11789 55722 11855 55725
rect 17033 55722 17099 55725
rect 11789 55720 17099 55722
rect 11789 55664 11794 55720
rect 11850 55664 17038 55720
rect 17094 55664 17099 55720
rect 11789 55662 17099 55664
rect 11789 55659 11855 55662
rect 17033 55659 17099 55662
rect 16481 55586 16547 55589
rect 17217 55586 17283 55589
rect 17953 55586 18019 55589
rect 16481 55584 18019 55586
rect 16481 55528 16486 55584
rect 16542 55528 17222 55584
rect 17278 55528 17958 55584
rect 18014 55528 18019 55584
rect 16481 55526 18019 55528
rect 16481 55523 16547 55526
rect 17217 55523 17283 55526
rect 17953 55523 18019 55526
rect 20621 55586 20687 55589
rect 22093 55586 22159 55589
rect 20621 55584 22159 55586
rect 20621 55528 20626 55584
rect 20682 55528 22098 55584
rect 22154 55528 22159 55584
rect 20621 55526 22159 55528
rect 20621 55523 20687 55526
rect 22093 55523 22159 55526
rect 5944 55520 6264 55521
rect 5944 55456 5952 55520
rect 6016 55456 6032 55520
rect 6096 55456 6112 55520
rect 6176 55456 6192 55520
rect 6256 55456 6264 55520
rect 5944 55455 6264 55456
rect 15944 55520 16264 55521
rect 15944 55456 15952 55520
rect 16016 55456 16032 55520
rect 16096 55456 16112 55520
rect 16176 55456 16192 55520
rect 16256 55456 16264 55520
rect 15944 55455 16264 55456
rect 25944 55520 26264 55521
rect 25944 55456 25952 55520
rect 26016 55456 26032 55520
rect 26096 55456 26112 55520
rect 26176 55456 26192 55520
rect 26256 55456 26264 55520
rect 25944 55455 26264 55456
rect 12065 55450 12131 55453
rect 14549 55450 14615 55453
rect 12065 55448 14615 55450
rect 12065 55392 12070 55448
rect 12126 55392 14554 55448
rect 14610 55392 14615 55448
rect 12065 55390 14615 55392
rect 12065 55387 12131 55390
rect 14549 55387 14615 55390
rect 17769 55450 17835 55453
rect 21357 55450 21423 55453
rect 17769 55448 21423 55450
rect 17769 55392 17774 55448
rect 17830 55392 21362 55448
rect 21418 55392 21423 55448
rect 17769 55390 21423 55392
rect 17769 55387 17835 55390
rect 21357 55387 21423 55390
rect 15101 55314 15167 55317
rect 18689 55314 18755 55317
rect 21081 55314 21147 55317
rect 15101 55312 21147 55314
rect 15101 55256 15106 55312
rect 15162 55256 18694 55312
rect 18750 55256 21086 55312
rect 21142 55256 21147 55312
rect 15101 55254 21147 55256
rect 15101 55251 15167 55254
rect 18689 55251 18755 55254
rect 21081 55251 21147 55254
rect 21265 55314 21331 55317
rect 21398 55314 21404 55316
rect 21265 55312 21404 55314
rect 21265 55256 21270 55312
rect 21326 55256 21404 55312
rect 21265 55254 21404 55256
rect 21265 55251 21331 55254
rect 21398 55252 21404 55254
rect 21468 55252 21474 55316
rect 0 55178 800 55208
rect 25037 55178 25103 55181
rect 29200 55178 30000 55208
rect 0 55088 858 55178
rect 25037 55176 30000 55178
rect 25037 55120 25042 55176
rect 25098 55120 30000 55176
rect 25037 55118 30000 55120
rect 25037 55115 25103 55118
rect 29200 55088 30000 55118
rect 798 54770 858 55088
rect 21357 55042 21423 55045
rect 22737 55042 22803 55045
rect 26601 55042 26667 55045
rect 21357 55040 26667 55042
rect 21357 54984 21362 55040
rect 21418 54984 22742 55040
rect 22798 54984 26606 55040
rect 26662 54984 26667 55040
rect 21357 54982 26667 54984
rect 21357 54979 21423 54982
rect 22737 54979 22803 54982
rect 26601 54979 26667 54982
rect 10944 54976 11264 54977
rect 10944 54912 10952 54976
rect 11016 54912 11032 54976
rect 11096 54912 11112 54976
rect 11176 54912 11192 54976
rect 11256 54912 11264 54976
rect 10944 54911 11264 54912
rect 20944 54976 21264 54977
rect 20944 54912 20952 54976
rect 21016 54912 21032 54976
rect 21096 54912 21112 54976
rect 21176 54912 21192 54976
rect 21256 54912 21264 54976
rect 20944 54911 21264 54912
rect 14917 54906 14983 54909
rect 16665 54906 16731 54909
rect 14917 54904 16731 54906
rect 14917 54848 14922 54904
rect 14978 54848 16670 54904
rect 16726 54848 16731 54904
rect 14917 54846 16731 54848
rect 14917 54843 14983 54846
rect 16665 54843 16731 54846
rect 21081 54770 21147 54773
rect 798 54768 21147 54770
rect 798 54712 21086 54768
rect 21142 54712 21147 54768
rect 798 54710 21147 54712
rect 21081 54707 21147 54710
rect 13169 54634 13235 54637
rect 18597 54634 18663 54637
rect 19333 54634 19399 54637
rect 13169 54632 19399 54634
rect 13169 54576 13174 54632
rect 13230 54576 18602 54632
rect 18658 54576 19338 54632
rect 19394 54576 19399 54632
rect 13169 54574 19399 54576
rect 13169 54571 13235 54574
rect 18597 54571 18663 54574
rect 19333 54571 19399 54574
rect 5944 54432 6264 54433
rect 5944 54368 5952 54432
rect 6016 54368 6032 54432
rect 6096 54368 6112 54432
rect 6176 54368 6192 54432
rect 6256 54368 6264 54432
rect 5944 54367 6264 54368
rect 15944 54432 16264 54433
rect 15944 54368 15952 54432
rect 16016 54368 16032 54432
rect 16096 54368 16112 54432
rect 16176 54368 16192 54432
rect 16256 54368 16264 54432
rect 15944 54367 16264 54368
rect 25944 54432 26264 54433
rect 25944 54368 25952 54432
rect 26016 54368 26032 54432
rect 26096 54368 26112 54432
rect 26176 54368 26192 54432
rect 26256 54368 26264 54432
rect 25944 54367 26264 54368
rect 11881 54226 11947 54229
rect 16021 54226 16087 54229
rect 11881 54224 16087 54226
rect 11881 54168 11886 54224
rect 11942 54168 16026 54224
rect 16082 54168 16087 54224
rect 11881 54166 16087 54168
rect 11881 54163 11947 54166
rect 16021 54163 16087 54166
rect 11513 54090 11579 54093
rect 13169 54090 13235 54093
rect 11513 54088 13235 54090
rect 11513 54032 11518 54088
rect 11574 54032 13174 54088
rect 13230 54032 13235 54088
rect 11513 54030 13235 54032
rect 11513 54027 11579 54030
rect 13169 54027 13235 54030
rect 13445 54090 13511 54093
rect 15193 54090 15259 54093
rect 13445 54088 15259 54090
rect 13445 54032 13450 54088
rect 13506 54032 15198 54088
rect 15254 54032 15259 54088
rect 13445 54030 15259 54032
rect 13445 54027 13511 54030
rect 15193 54027 15259 54030
rect 22185 54090 22251 54093
rect 23473 54090 23539 54093
rect 22185 54088 23539 54090
rect 22185 54032 22190 54088
rect 22246 54032 23478 54088
rect 23534 54032 23539 54088
rect 22185 54030 23539 54032
rect 22185 54027 22251 54030
rect 23473 54027 23539 54030
rect 11881 53954 11947 53957
rect 13997 53954 14063 53957
rect 11881 53952 14063 53954
rect 11881 53896 11886 53952
rect 11942 53896 14002 53952
rect 14058 53896 14063 53952
rect 11881 53894 14063 53896
rect 11881 53891 11947 53894
rect 13997 53891 14063 53894
rect 10944 53888 11264 53889
rect 0 53818 800 53848
rect 10944 53824 10952 53888
rect 11016 53824 11032 53888
rect 11096 53824 11112 53888
rect 11176 53824 11192 53888
rect 11256 53824 11264 53888
rect 10944 53823 11264 53824
rect 20944 53888 21264 53889
rect 20944 53824 20952 53888
rect 21016 53824 21032 53888
rect 21096 53824 21112 53888
rect 21176 53824 21192 53888
rect 21256 53824 21264 53888
rect 20944 53823 21264 53824
rect 1669 53818 1735 53821
rect 0 53816 1735 53818
rect 0 53760 1674 53816
rect 1730 53760 1735 53816
rect 0 53758 1735 53760
rect 0 53728 800 53758
rect 1669 53755 1735 53758
rect 18781 53818 18847 53821
rect 25405 53818 25471 53821
rect 29200 53818 30000 53848
rect 18781 53816 18890 53818
rect 18781 53760 18786 53816
rect 18842 53760 18890 53816
rect 18781 53755 18890 53760
rect 25405 53816 30000 53818
rect 25405 53760 25410 53816
rect 25466 53760 30000 53816
rect 25405 53758 30000 53760
rect 25405 53755 25471 53758
rect 11605 53682 11671 53685
rect 982 53680 11671 53682
rect 982 53624 11610 53680
rect 11666 53624 11671 53680
rect 982 53622 11671 53624
rect 982 53274 1042 53622
rect 11605 53619 11671 53622
rect 14733 53682 14799 53685
rect 18689 53682 18755 53685
rect 14733 53680 18755 53682
rect 14733 53624 14738 53680
rect 14794 53624 18694 53680
rect 18750 53624 18755 53680
rect 14733 53622 18755 53624
rect 18830 53682 18890 53755
rect 29200 53728 30000 53758
rect 22461 53682 22527 53685
rect 18830 53680 22527 53682
rect 18830 53624 22466 53680
rect 22522 53624 22527 53680
rect 18830 53622 22527 53624
rect 14733 53619 14799 53622
rect 18689 53619 18755 53622
rect 22461 53619 22527 53622
rect 14457 53546 14523 53549
rect 18229 53546 18295 53549
rect 14457 53544 18295 53546
rect 14457 53488 14462 53544
rect 14518 53488 18234 53544
rect 18290 53488 18295 53544
rect 14457 53486 18295 53488
rect 14457 53483 14523 53486
rect 18229 53483 18295 53486
rect 11421 53410 11487 53413
rect 14641 53410 14707 53413
rect 15101 53410 15167 53413
rect 11421 53408 15167 53410
rect 11421 53352 11426 53408
rect 11482 53352 14646 53408
rect 14702 53352 15106 53408
rect 15162 53352 15167 53408
rect 11421 53350 15167 53352
rect 11421 53347 11487 53350
rect 14641 53347 14707 53350
rect 15101 53347 15167 53350
rect 5944 53344 6264 53345
rect 5944 53280 5952 53344
rect 6016 53280 6032 53344
rect 6096 53280 6112 53344
rect 6176 53280 6192 53344
rect 6256 53280 6264 53344
rect 5944 53279 6264 53280
rect 15944 53344 16264 53345
rect 15944 53280 15952 53344
rect 16016 53280 16032 53344
rect 16096 53280 16112 53344
rect 16176 53280 16192 53344
rect 16256 53280 16264 53344
rect 15944 53279 16264 53280
rect 25944 53344 26264 53345
rect 25944 53280 25952 53344
rect 26016 53280 26032 53344
rect 26096 53280 26112 53344
rect 26176 53280 26192 53344
rect 26256 53280 26264 53344
rect 25944 53279 26264 53280
rect 798 53214 1042 53274
rect 16573 53274 16639 53277
rect 16941 53274 17007 53277
rect 16573 53272 17007 53274
rect 16573 53216 16578 53272
rect 16634 53216 16946 53272
rect 17002 53216 17007 53272
rect 16573 53214 17007 53216
rect 798 53168 858 53214
rect 16573 53211 16639 53214
rect 16941 53211 17007 53214
rect 0 53078 858 53168
rect 21541 53138 21607 53141
rect 21766 53138 21772 53140
rect 21541 53136 21772 53138
rect 21541 53080 21546 53136
rect 21602 53080 21772 53136
rect 21541 53078 21772 53080
rect 0 53048 800 53078
rect 21541 53075 21607 53078
rect 21766 53076 21772 53078
rect 21836 53076 21842 53140
rect 24485 53138 24551 53141
rect 29200 53138 30000 53168
rect 24485 53136 30000 53138
rect 24485 53080 24490 53136
rect 24546 53080 30000 53136
rect 24485 53078 30000 53080
rect 24485 53075 24551 53078
rect 29200 53048 30000 53078
rect 14825 53002 14891 53005
rect 16941 53002 17007 53005
rect 14825 53000 17007 53002
rect 14825 52944 14830 53000
rect 14886 52944 16946 53000
rect 17002 52944 17007 53000
rect 14825 52942 17007 52944
rect 14825 52939 14891 52942
rect 16941 52939 17007 52942
rect 18505 53002 18571 53005
rect 21081 53002 21147 53005
rect 18505 53000 21147 53002
rect 18505 52944 18510 53000
rect 18566 52944 21086 53000
rect 21142 52944 21147 53000
rect 18505 52942 21147 52944
rect 18505 52939 18571 52942
rect 21081 52939 21147 52942
rect 25446 52940 25452 53004
rect 25516 53002 25522 53004
rect 27889 53002 27955 53005
rect 25516 53000 27955 53002
rect 25516 52944 27894 53000
rect 27950 52944 27955 53000
rect 25516 52942 27955 52944
rect 25516 52940 25522 52942
rect 27889 52939 27955 52942
rect 14273 52866 14339 52869
rect 17217 52866 17283 52869
rect 14273 52864 17283 52866
rect 14273 52808 14278 52864
rect 14334 52808 17222 52864
rect 17278 52808 17283 52864
rect 14273 52806 17283 52808
rect 14273 52803 14339 52806
rect 17217 52803 17283 52806
rect 10944 52800 11264 52801
rect 10944 52736 10952 52800
rect 11016 52736 11032 52800
rect 11096 52736 11112 52800
rect 11176 52736 11192 52800
rect 11256 52736 11264 52800
rect 10944 52735 11264 52736
rect 20944 52800 21264 52801
rect 20944 52736 20952 52800
rect 21016 52736 21032 52800
rect 21096 52736 21112 52800
rect 21176 52736 21192 52800
rect 21256 52736 21264 52800
rect 20944 52735 21264 52736
rect 11329 52730 11395 52733
rect 13997 52730 14063 52733
rect 11329 52728 14063 52730
rect 11329 52672 11334 52728
rect 11390 52672 14002 52728
rect 14058 52672 14063 52728
rect 11329 52670 14063 52672
rect 11329 52667 11395 52670
rect 13997 52667 14063 52670
rect 15009 52730 15075 52733
rect 18045 52730 18111 52733
rect 15009 52728 18111 52730
rect 15009 52672 15014 52728
rect 15070 52672 18050 52728
rect 18106 52672 18111 52728
rect 15009 52670 18111 52672
rect 15009 52667 15075 52670
rect 18045 52667 18111 52670
rect 4061 52594 4127 52597
rect 12014 52594 12020 52596
rect 4061 52592 12020 52594
rect 4061 52536 4066 52592
rect 4122 52536 12020 52592
rect 4061 52534 12020 52536
rect 4061 52531 4127 52534
rect 12014 52532 12020 52534
rect 12084 52532 12090 52596
rect 12249 52594 12315 52597
rect 15193 52594 15259 52597
rect 16481 52596 16547 52597
rect 16430 52594 16436 52596
rect 12249 52592 15259 52594
rect 12249 52536 12254 52592
rect 12310 52536 15198 52592
rect 15254 52536 15259 52592
rect 12249 52534 15259 52536
rect 16390 52534 16436 52594
rect 16500 52592 16547 52596
rect 16542 52536 16547 52592
rect 12249 52531 12315 52534
rect 15193 52531 15259 52534
rect 16430 52532 16436 52534
rect 16500 52532 16547 52536
rect 16481 52531 16547 52532
rect 20621 52594 20687 52597
rect 25681 52594 25747 52597
rect 20621 52592 25747 52594
rect 20621 52536 20626 52592
rect 20682 52536 25686 52592
rect 25742 52536 25747 52592
rect 20621 52534 25747 52536
rect 20621 52531 20687 52534
rect 25681 52531 25747 52534
rect 11605 52458 11671 52461
rect 23749 52458 23815 52461
rect 11605 52456 23815 52458
rect 11605 52400 11610 52456
rect 11666 52400 23754 52456
rect 23810 52400 23815 52456
rect 11605 52398 23815 52400
rect 11605 52395 11671 52398
rect 23749 52395 23815 52398
rect 25313 52458 25379 52461
rect 27337 52458 27403 52461
rect 25313 52456 27403 52458
rect 25313 52400 25318 52456
rect 25374 52400 27342 52456
rect 27398 52400 27403 52456
rect 25313 52398 27403 52400
rect 25313 52395 25379 52398
rect 27337 52395 27403 52398
rect 10961 52322 11027 52325
rect 12617 52322 12683 52325
rect 10961 52320 12683 52322
rect 10961 52264 10966 52320
rect 11022 52264 12622 52320
rect 12678 52264 12683 52320
rect 10961 52262 12683 52264
rect 10961 52259 11027 52262
rect 12617 52259 12683 52262
rect 24209 52322 24275 52325
rect 25773 52322 25839 52325
rect 24209 52320 25839 52322
rect 24209 52264 24214 52320
rect 24270 52264 25778 52320
rect 25834 52264 25839 52320
rect 24209 52262 25839 52264
rect 24209 52259 24275 52262
rect 25773 52259 25839 52262
rect 5944 52256 6264 52257
rect 5944 52192 5952 52256
rect 6016 52192 6032 52256
rect 6096 52192 6112 52256
rect 6176 52192 6192 52256
rect 6256 52192 6264 52256
rect 5944 52191 6264 52192
rect 15944 52256 16264 52257
rect 15944 52192 15952 52256
rect 16016 52192 16032 52256
rect 16096 52192 16112 52256
rect 16176 52192 16192 52256
rect 16256 52192 16264 52256
rect 15944 52191 16264 52192
rect 25944 52256 26264 52257
rect 25944 52192 25952 52256
rect 26016 52192 26032 52256
rect 26096 52192 26112 52256
rect 26176 52192 26192 52256
rect 26256 52192 26264 52256
rect 25944 52191 26264 52192
rect 8385 52186 8451 52189
rect 11697 52186 11763 52189
rect 8385 52184 11763 52186
rect 8385 52128 8390 52184
rect 8446 52128 11702 52184
rect 11758 52128 11763 52184
rect 8385 52126 11763 52128
rect 8385 52123 8451 52126
rect 11697 52123 11763 52126
rect 17585 52186 17651 52189
rect 17718 52186 17724 52188
rect 17585 52184 17724 52186
rect 17585 52128 17590 52184
rect 17646 52128 17724 52184
rect 17585 52126 17724 52128
rect 17585 52123 17651 52126
rect 17718 52124 17724 52126
rect 17788 52124 17794 52188
rect 13537 52050 13603 52053
rect 15285 52050 15351 52053
rect 13537 52048 15351 52050
rect 13537 51992 13542 52048
rect 13598 51992 15290 52048
rect 15346 51992 15351 52048
rect 13537 51990 15351 51992
rect 13537 51987 13603 51990
rect 15285 51987 15351 51990
rect 19517 52050 19583 52053
rect 19517 52048 21466 52050
rect 19517 51992 19522 52048
rect 19578 51992 21466 52048
rect 19517 51990 21466 51992
rect 19517 51987 19583 51990
rect 0 51778 800 51808
rect 16941 51778 17007 51781
rect 0 51688 858 51778
rect 16941 51776 17050 51778
rect 16941 51720 16946 51776
rect 17002 51720 17050 51776
rect 16941 51715 17050 51720
rect 798 51506 858 51688
rect 10944 51712 11264 51713
rect 10944 51648 10952 51712
rect 11016 51648 11032 51712
rect 11096 51648 11112 51712
rect 11176 51648 11192 51712
rect 11256 51648 11264 51712
rect 10944 51647 11264 51648
rect 12433 51506 12499 51509
rect 798 51504 12499 51506
rect 798 51448 12438 51504
rect 12494 51448 12499 51504
rect 798 51446 12499 51448
rect 12433 51443 12499 51446
rect 12709 51506 12775 51509
rect 16665 51506 16731 51509
rect 12709 51504 16731 51506
rect 12709 51448 12714 51504
rect 12770 51448 16670 51504
rect 16726 51448 16731 51504
rect 12709 51446 16731 51448
rect 12709 51443 12775 51446
rect 16665 51443 16731 51446
rect 6269 51370 6335 51373
rect 7833 51370 7899 51373
rect 10409 51370 10475 51373
rect 6269 51368 10475 51370
rect 6269 51312 6274 51368
rect 6330 51312 7838 51368
rect 7894 51312 10414 51368
rect 10470 51312 10475 51368
rect 6269 51310 10475 51312
rect 6269 51307 6335 51310
rect 7833 51307 7899 51310
rect 10409 51307 10475 51310
rect 15510 51308 15516 51372
rect 15580 51370 15586 51372
rect 15837 51370 15903 51373
rect 15580 51368 15903 51370
rect 15580 51312 15842 51368
rect 15898 51312 15903 51368
rect 15580 51310 15903 51312
rect 15580 51308 15586 51310
rect 15837 51307 15903 51310
rect 16990 51234 17050 51715
rect 20944 51712 21264 51713
rect 20944 51648 20952 51712
rect 21016 51648 21032 51712
rect 21096 51648 21112 51712
rect 21176 51648 21192 51712
rect 21256 51648 21264 51712
rect 20944 51647 21264 51648
rect 21406 51642 21466 51990
rect 25681 51778 25747 51781
rect 29200 51778 30000 51808
rect 25681 51776 30000 51778
rect 25681 51720 25686 51776
rect 25742 51720 30000 51776
rect 25681 51718 30000 51720
rect 25681 51715 25747 51718
rect 29200 51688 30000 51718
rect 25221 51642 25287 51645
rect 21406 51640 25287 51642
rect 21406 51584 25226 51640
rect 25282 51584 25287 51640
rect 21406 51582 25287 51584
rect 25221 51579 25287 51582
rect 21173 51506 21239 51509
rect 23657 51506 23723 51509
rect 21173 51504 23723 51506
rect 21173 51448 21178 51504
rect 21234 51448 23662 51504
rect 23718 51448 23723 51504
rect 21173 51446 23723 51448
rect 21173 51443 21239 51446
rect 23657 51443 23723 51446
rect 19149 51370 19215 51373
rect 23197 51370 23263 51373
rect 19149 51368 23263 51370
rect 19149 51312 19154 51368
rect 19210 51312 23202 51368
rect 23258 51312 23263 51368
rect 19149 51310 23263 51312
rect 19149 51307 19215 51310
rect 23197 51307 23263 51310
rect 22921 51234 22987 51237
rect 16990 51232 22987 51234
rect 16990 51176 22926 51232
rect 22982 51176 22987 51232
rect 16990 51174 22987 51176
rect 22921 51171 22987 51174
rect 5944 51168 6264 51169
rect 5944 51104 5952 51168
rect 6016 51104 6032 51168
rect 6096 51104 6112 51168
rect 6176 51104 6192 51168
rect 6256 51104 6264 51168
rect 5944 51103 6264 51104
rect 15944 51168 16264 51169
rect 15944 51104 15952 51168
rect 16016 51104 16032 51168
rect 16096 51104 16112 51168
rect 16176 51104 16192 51168
rect 16256 51104 16264 51168
rect 15944 51103 16264 51104
rect 25944 51168 26264 51169
rect 25944 51104 25952 51168
rect 26016 51104 26032 51168
rect 26096 51104 26112 51168
rect 26176 51104 26192 51168
rect 26256 51104 26264 51168
rect 25944 51103 26264 51104
rect 15009 51098 15075 51101
rect 15193 51098 15259 51101
rect 15009 51096 15259 51098
rect 15009 51040 15014 51096
rect 15070 51040 15198 51096
rect 15254 51040 15259 51096
rect 15009 51038 15259 51040
rect 15009 51035 15075 51038
rect 15193 51035 15259 51038
rect 1577 50962 1643 50965
rect 5809 50962 5875 50965
rect 7373 50962 7439 50965
rect 1577 50960 7439 50962
rect 1577 50904 1582 50960
rect 1638 50904 5814 50960
rect 5870 50904 7378 50960
rect 7434 50904 7439 50960
rect 1577 50902 7439 50904
rect 1577 50899 1643 50902
rect 5809 50899 5875 50902
rect 7373 50899 7439 50902
rect 11513 50962 11579 50965
rect 13813 50962 13879 50965
rect 11513 50960 13879 50962
rect 11513 50904 11518 50960
rect 11574 50904 13818 50960
rect 13874 50904 13879 50960
rect 11513 50902 13879 50904
rect 11513 50899 11579 50902
rect 13813 50899 13879 50902
rect 14457 50962 14523 50965
rect 23565 50962 23631 50965
rect 14457 50960 16130 50962
rect 14457 50904 14462 50960
rect 14518 50904 16130 50960
rect 14457 50902 16130 50904
rect 14457 50899 14523 50902
rect 13997 50826 14063 50829
rect 15510 50826 15516 50828
rect 13997 50824 15516 50826
rect 13997 50768 14002 50824
rect 14058 50768 15516 50824
rect 13997 50766 15516 50768
rect 13997 50763 14063 50766
rect 15510 50764 15516 50766
rect 15580 50764 15586 50828
rect 16070 50826 16130 50902
rect 23565 50960 23812 50962
rect 23565 50904 23570 50960
rect 23626 50904 23812 50960
rect 23565 50902 23812 50904
rect 23565 50899 23631 50902
rect 17677 50826 17743 50829
rect 16070 50824 17743 50826
rect 16070 50768 17682 50824
rect 17738 50768 17743 50824
rect 16070 50766 17743 50768
rect 17677 50763 17743 50766
rect 20069 50826 20135 50829
rect 22001 50826 22067 50829
rect 23289 50826 23355 50829
rect 20069 50824 21466 50826
rect 20069 50768 20074 50824
rect 20130 50768 21466 50824
rect 20069 50766 21466 50768
rect 20069 50763 20135 50766
rect 12249 50690 12315 50693
rect 13077 50690 13143 50693
rect 12249 50688 13143 50690
rect 12249 50632 12254 50688
rect 12310 50632 13082 50688
rect 13138 50632 13143 50688
rect 12249 50630 13143 50632
rect 12249 50627 12315 50630
rect 13077 50627 13143 50630
rect 15561 50690 15627 50693
rect 18873 50690 18939 50693
rect 15561 50688 18939 50690
rect 15561 50632 15566 50688
rect 15622 50632 18878 50688
rect 18934 50632 18939 50688
rect 15561 50630 18939 50632
rect 21406 50690 21466 50766
rect 22001 50824 23355 50826
rect 22001 50768 22006 50824
rect 22062 50768 23294 50824
rect 23350 50768 23355 50824
rect 22001 50766 23355 50768
rect 22001 50763 22067 50766
rect 23289 50763 23355 50766
rect 23752 50693 23812 50902
rect 23565 50690 23631 50693
rect 21406 50688 23631 50690
rect 21406 50632 23570 50688
rect 23626 50632 23631 50688
rect 21406 50630 23631 50632
rect 15561 50627 15627 50630
rect 18873 50627 18939 50630
rect 23565 50627 23631 50630
rect 23749 50688 23815 50693
rect 23749 50632 23754 50688
rect 23810 50632 23815 50688
rect 23749 50627 23815 50632
rect 10944 50624 11264 50625
rect 10944 50560 10952 50624
rect 11016 50560 11032 50624
rect 11096 50560 11112 50624
rect 11176 50560 11192 50624
rect 11256 50560 11264 50624
rect 10944 50559 11264 50560
rect 20944 50624 21264 50625
rect 20944 50560 20952 50624
rect 21016 50560 21032 50624
rect 21096 50560 21112 50624
rect 21176 50560 21192 50624
rect 21256 50560 21264 50624
rect 20944 50559 21264 50560
rect 17309 50554 17375 50557
rect 17309 50552 20730 50554
rect 17309 50496 17314 50552
rect 17370 50496 20730 50552
rect 17309 50494 20730 50496
rect 17309 50491 17375 50494
rect 0 50418 800 50448
rect 4061 50418 4127 50421
rect 0 50416 4127 50418
rect 0 50360 4066 50416
rect 4122 50360 4127 50416
rect 0 50358 4127 50360
rect 0 50328 800 50358
rect 4061 50355 4127 50358
rect 13077 50418 13143 50421
rect 14181 50418 14247 50421
rect 17953 50418 18019 50421
rect 13077 50416 18019 50418
rect 13077 50360 13082 50416
rect 13138 50360 14186 50416
rect 14242 50360 17958 50416
rect 18014 50360 18019 50416
rect 13077 50358 18019 50360
rect 20670 50418 20730 50494
rect 22001 50418 22067 50421
rect 20670 50416 22067 50418
rect 20670 50360 22006 50416
rect 22062 50360 22067 50416
rect 20670 50358 22067 50360
rect 13077 50355 13143 50358
rect 14181 50355 14247 50358
rect 17953 50355 18019 50358
rect 22001 50355 22067 50358
rect 25221 50418 25287 50421
rect 29200 50418 30000 50448
rect 25221 50416 30000 50418
rect 25221 50360 25226 50416
rect 25282 50360 30000 50416
rect 25221 50358 30000 50360
rect 25221 50355 25287 50358
rect 29200 50328 30000 50358
rect 8937 50282 9003 50285
rect 21541 50282 21607 50285
rect 8937 50280 21607 50282
rect 8937 50224 8942 50280
rect 8998 50224 21546 50280
rect 21602 50224 21607 50280
rect 8937 50222 21607 50224
rect 8937 50219 9003 50222
rect 21541 50219 21607 50222
rect 22001 50282 22067 50285
rect 25405 50282 25471 50285
rect 22001 50280 25471 50282
rect 22001 50224 22006 50280
rect 22062 50224 25410 50280
rect 25466 50224 25471 50280
rect 22001 50222 25471 50224
rect 22001 50219 22067 50222
rect 25405 50219 25471 50222
rect 18689 50146 18755 50149
rect 21541 50146 21607 50149
rect 18689 50144 21607 50146
rect 18689 50088 18694 50144
rect 18750 50088 21546 50144
rect 21602 50088 21607 50144
rect 18689 50086 21607 50088
rect 18689 50083 18755 50086
rect 21541 50083 21607 50086
rect 5944 50080 6264 50081
rect 5944 50016 5952 50080
rect 6016 50016 6032 50080
rect 6096 50016 6112 50080
rect 6176 50016 6192 50080
rect 6256 50016 6264 50080
rect 5944 50015 6264 50016
rect 15944 50080 16264 50081
rect 15944 50016 15952 50080
rect 16016 50016 16032 50080
rect 16096 50016 16112 50080
rect 16176 50016 16192 50080
rect 16256 50016 16264 50080
rect 15944 50015 16264 50016
rect 25944 50080 26264 50081
rect 25944 50016 25952 50080
rect 26016 50016 26032 50080
rect 26096 50016 26112 50080
rect 26176 50016 26192 50080
rect 26256 50016 26264 50080
rect 25944 50015 26264 50016
rect 20294 49948 20300 50012
rect 20364 50010 20370 50012
rect 21449 50010 21515 50013
rect 20364 50008 21515 50010
rect 20364 49952 21454 50008
rect 21510 49952 21515 50008
rect 20364 49950 21515 49952
rect 20364 49948 20370 49950
rect 21449 49947 21515 49950
rect 10501 49874 10567 49877
rect 16849 49874 16915 49877
rect 20345 49874 20411 49877
rect 10501 49872 16915 49874
rect 10501 49816 10506 49872
rect 10562 49816 16854 49872
rect 16910 49816 16915 49872
rect 10501 49814 16915 49816
rect 10501 49811 10567 49814
rect 16849 49811 16915 49814
rect 16990 49872 20411 49874
rect 16990 49816 20350 49872
rect 20406 49816 20411 49872
rect 16990 49814 20411 49816
rect 4061 49738 4127 49741
rect 12617 49738 12683 49741
rect 4061 49736 12683 49738
rect 4061 49680 4066 49736
rect 4122 49680 12622 49736
rect 12678 49680 12683 49736
rect 4061 49678 12683 49680
rect 4061 49675 4127 49678
rect 12617 49675 12683 49678
rect 15285 49738 15351 49741
rect 16990 49738 17050 49814
rect 20345 49811 20411 49814
rect 20897 49874 20963 49877
rect 22185 49874 22251 49877
rect 20897 49872 22251 49874
rect 20897 49816 20902 49872
rect 20958 49816 22190 49872
rect 22246 49816 22251 49872
rect 20897 49814 22251 49816
rect 20897 49811 20963 49814
rect 22185 49811 22251 49814
rect 15285 49736 17050 49738
rect 15285 49680 15290 49736
rect 15346 49680 17050 49736
rect 15285 49678 17050 49680
rect 18689 49738 18755 49741
rect 22001 49738 22067 49741
rect 29200 49738 30000 49768
rect 18689 49736 22067 49738
rect 18689 49680 18694 49736
rect 18750 49680 22006 49736
rect 22062 49680 22067 49736
rect 18689 49678 22067 49680
rect 15285 49675 15351 49678
rect 18689 49675 18755 49678
rect 22001 49675 22067 49678
rect 27846 49678 30000 49738
rect 11973 49602 12039 49605
rect 15745 49602 15811 49605
rect 11973 49600 15811 49602
rect 11973 49544 11978 49600
rect 12034 49544 15750 49600
rect 15806 49544 15811 49600
rect 11973 49542 15811 49544
rect 11973 49539 12039 49542
rect 15745 49539 15811 49542
rect 16021 49602 16087 49605
rect 16430 49602 16436 49604
rect 16021 49600 16436 49602
rect 16021 49544 16026 49600
rect 16082 49544 16436 49600
rect 16021 49542 16436 49544
rect 16021 49539 16087 49542
rect 16430 49540 16436 49542
rect 16500 49540 16506 49604
rect 27705 49602 27771 49605
rect 27846 49602 27906 49678
rect 29200 49648 30000 49678
rect 27705 49600 27906 49602
rect 27705 49544 27710 49600
rect 27766 49544 27906 49600
rect 27705 49542 27906 49544
rect 27705 49539 27771 49542
rect 10944 49536 11264 49537
rect 10944 49472 10952 49536
rect 11016 49472 11032 49536
rect 11096 49472 11112 49536
rect 11176 49472 11192 49536
rect 11256 49472 11264 49536
rect 10944 49471 11264 49472
rect 20944 49536 21264 49537
rect 20944 49472 20952 49536
rect 21016 49472 21032 49536
rect 21096 49472 21112 49536
rect 21176 49472 21192 49536
rect 21256 49472 21264 49536
rect 20944 49471 21264 49472
rect 20478 49404 20484 49468
rect 20548 49466 20554 49468
rect 20713 49466 20779 49469
rect 20548 49464 20779 49466
rect 20548 49408 20718 49464
rect 20774 49408 20779 49464
rect 20548 49406 20779 49408
rect 20548 49404 20554 49406
rect 20713 49403 20779 49406
rect 13537 49194 13603 49197
rect 14273 49194 14339 49197
rect 15285 49194 15351 49197
rect 13537 49192 15351 49194
rect 13537 49136 13542 49192
rect 13598 49136 14278 49192
rect 14334 49136 15290 49192
rect 15346 49136 15351 49192
rect 13537 49134 15351 49136
rect 13537 49131 13603 49134
rect 14273 49131 14339 49134
rect 15285 49131 15351 49134
rect 20294 49132 20300 49196
rect 20364 49194 20370 49196
rect 20805 49194 20871 49197
rect 20364 49192 20871 49194
rect 20364 49136 20810 49192
rect 20866 49136 20871 49192
rect 20364 49134 20871 49136
rect 20364 49132 20370 49134
rect 20805 49131 20871 49134
rect 0 49058 800 49088
rect 3693 49058 3759 49061
rect 0 49056 3759 49058
rect 0 49000 3698 49056
rect 3754 49000 3759 49056
rect 0 48998 3759 49000
rect 0 48968 800 48998
rect 3693 48995 3759 48998
rect 21633 49058 21699 49061
rect 22001 49058 22067 49061
rect 21633 49056 22067 49058
rect 21633 49000 21638 49056
rect 21694 49000 22006 49056
rect 22062 49000 22067 49056
rect 21633 48998 22067 49000
rect 21633 48995 21699 48998
rect 22001 48995 22067 48998
rect 5944 48992 6264 48993
rect 5944 48928 5952 48992
rect 6016 48928 6032 48992
rect 6096 48928 6112 48992
rect 6176 48928 6192 48992
rect 6256 48928 6264 48992
rect 5944 48927 6264 48928
rect 15944 48992 16264 48993
rect 15944 48928 15952 48992
rect 16016 48928 16032 48992
rect 16096 48928 16112 48992
rect 16176 48928 16192 48992
rect 16256 48928 16264 48992
rect 15944 48927 16264 48928
rect 25944 48992 26264 48993
rect 25944 48928 25952 48992
rect 26016 48928 26032 48992
rect 26096 48928 26112 48992
rect 26176 48928 26192 48992
rect 26256 48928 26264 48992
rect 25944 48927 26264 48928
rect 13629 48922 13695 48925
rect 15469 48922 15535 48925
rect 13629 48920 15535 48922
rect 13629 48864 13634 48920
rect 13690 48864 15474 48920
rect 15530 48864 15535 48920
rect 13629 48862 15535 48864
rect 13629 48859 13695 48862
rect 15469 48859 15535 48862
rect 17125 48922 17191 48925
rect 19977 48922 20043 48925
rect 17125 48920 20043 48922
rect 17125 48864 17130 48920
rect 17186 48864 19982 48920
rect 20038 48864 20043 48920
rect 17125 48862 20043 48864
rect 17125 48859 17191 48862
rect 19977 48859 20043 48862
rect 19333 48786 19399 48789
rect 25221 48786 25287 48789
rect 19333 48784 25287 48786
rect 19333 48728 19338 48784
rect 19394 48728 25226 48784
rect 25282 48728 25287 48784
rect 19333 48726 25287 48728
rect 19333 48723 19399 48726
rect 25221 48723 25287 48726
rect 3509 48650 3575 48653
rect 12065 48650 12131 48653
rect 3509 48648 12131 48650
rect 3509 48592 3514 48648
rect 3570 48592 12070 48648
rect 12126 48592 12131 48648
rect 3509 48590 12131 48592
rect 3509 48587 3575 48590
rect 12065 48587 12131 48590
rect 13169 48650 13235 48653
rect 18045 48650 18111 48653
rect 13169 48648 18111 48650
rect 13169 48592 13174 48648
rect 13230 48592 18050 48648
rect 18106 48592 18111 48648
rect 13169 48590 18111 48592
rect 13169 48587 13235 48590
rect 18045 48587 18111 48590
rect 19885 48650 19951 48653
rect 19885 48648 21420 48650
rect 19885 48592 19890 48648
rect 19946 48592 21420 48648
rect 19885 48590 21420 48592
rect 19885 48587 19951 48590
rect 12801 48514 12867 48517
rect 16941 48514 17007 48517
rect 12801 48512 17007 48514
rect 12801 48456 12806 48512
rect 12862 48456 16946 48512
rect 17002 48456 17007 48512
rect 12801 48454 17007 48456
rect 12801 48451 12867 48454
rect 16941 48451 17007 48454
rect 19425 48514 19491 48517
rect 20069 48514 20135 48517
rect 19425 48512 20135 48514
rect 19425 48456 19430 48512
rect 19486 48456 20074 48512
rect 20130 48456 20135 48512
rect 19425 48454 20135 48456
rect 19425 48451 19491 48454
rect 20069 48451 20135 48454
rect 10944 48448 11264 48449
rect 0 48378 800 48408
rect 10944 48384 10952 48448
rect 11016 48384 11032 48448
rect 11096 48384 11112 48448
rect 11176 48384 11192 48448
rect 11256 48384 11264 48448
rect 10944 48383 11264 48384
rect 20944 48448 21264 48449
rect 20944 48384 20952 48448
rect 21016 48384 21032 48448
rect 21096 48384 21112 48448
rect 21176 48384 21192 48448
rect 21256 48384 21264 48448
rect 20944 48383 21264 48384
rect 4061 48378 4127 48381
rect 0 48376 4127 48378
rect 0 48320 4066 48376
rect 4122 48320 4127 48376
rect 0 48318 4127 48320
rect 0 48288 800 48318
rect 4061 48315 4127 48318
rect 15326 48316 15332 48380
rect 15396 48378 15402 48380
rect 15469 48378 15535 48381
rect 15396 48376 15535 48378
rect 15396 48320 15474 48376
rect 15530 48320 15535 48376
rect 15396 48318 15535 48320
rect 15396 48316 15402 48318
rect 15469 48315 15535 48318
rect 17493 48378 17559 48381
rect 18965 48378 19031 48381
rect 17493 48376 19031 48378
rect 17493 48320 17498 48376
rect 17554 48320 18970 48376
rect 19026 48320 19031 48376
rect 17493 48318 19031 48320
rect 21360 48378 21420 48590
rect 21817 48516 21883 48517
rect 21766 48514 21772 48516
rect 21726 48454 21772 48514
rect 21836 48512 21883 48516
rect 21878 48456 21883 48512
rect 21766 48452 21772 48454
rect 21836 48452 21883 48456
rect 21817 48451 21883 48452
rect 24025 48514 24091 48517
rect 28073 48514 28139 48517
rect 24025 48512 28139 48514
rect 24025 48456 24030 48512
rect 24086 48456 28078 48512
rect 28134 48456 28139 48512
rect 24025 48454 28139 48456
rect 24025 48451 24091 48454
rect 28073 48451 28139 48454
rect 29200 48378 30000 48408
rect 21360 48318 30000 48378
rect 17493 48315 17559 48318
rect 18965 48315 19031 48318
rect 29200 48288 30000 48318
rect 3601 48242 3667 48245
rect 7189 48242 7255 48245
rect 3601 48240 7255 48242
rect 3601 48184 3606 48240
rect 3662 48184 7194 48240
rect 7250 48184 7255 48240
rect 3601 48182 7255 48184
rect 3601 48179 3667 48182
rect 7189 48179 7255 48182
rect 8201 48242 8267 48245
rect 11421 48242 11487 48245
rect 8201 48240 11487 48242
rect 8201 48184 8206 48240
rect 8262 48184 11426 48240
rect 11482 48184 11487 48240
rect 8201 48182 11487 48184
rect 8201 48179 8267 48182
rect 11421 48179 11487 48182
rect 19057 48242 19123 48245
rect 22277 48242 22343 48245
rect 19057 48240 22343 48242
rect 19057 48184 19062 48240
rect 19118 48184 22282 48240
rect 22338 48184 22343 48240
rect 19057 48182 22343 48184
rect 19057 48179 19123 48182
rect 22277 48179 22343 48182
rect 22645 48242 22711 48245
rect 25129 48242 25195 48245
rect 22645 48240 25195 48242
rect 22645 48184 22650 48240
rect 22706 48184 25134 48240
rect 25190 48184 25195 48240
rect 22645 48182 25195 48184
rect 22645 48179 22711 48182
rect 25129 48179 25195 48182
rect 3785 48106 3851 48109
rect 7833 48106 7899 48109
rect 3785 48104 7899 48106
rect 3785 48048 3790 48104
rect 3846 48048 7838 48104
rect 7894 48048 7899 48104
rect 3785 48046 7899 48048
rect 3785 48043 3851 48046
rect 7833 48043 7899 48046
rect 9397 48106 9463 48109
rect 12893 48106 12959 48109
rect 9397 48104 12959 48106
rect 9397 48048 9402 48104
rect 9458 48048 12898 48104
rect 12954 48048 12959 48104
rect 9397 48046 12959 48048
rect 9397 48043 9463 48046
rect 12893 48043 12959 48046
rect 13077 48106 13143 48109
rect 18045 48106 18111 48109
rect 21541 48106 21607 48109
rect 13077 48104 21607 48106
rect 13077 48048 13082 48104
rect 13138 48048 18050 48104
rect 18106 48048 21546 48104
rect 21602 48048 21607 48104
rect 13077 48046 21607 48048
rect 13077 48043 13143 48046
rect 18045 48043 18111 48046
rect 21541 48043 21607 48046
rect 22185 48106 22251 48109
rect 23565 48106 23631 48109
rect 22185 48104 23631 48106
rect 22185 48048 22190 48104
rect 22246 48048 23570 48104
rect 23626 48048 23631 48104
rect 22185 48046 23631 48048
rect 22185 48043 22251 48046
rect 23565 48043 23631 48046
rect 17309 47970 17375 47973
rect 19926 47970 19932 47972
rect 17309 47968 19932 47970
rect 17309 47912 17314 47968
rect 17370 47912 19932 47968
rect 17309 47910 19932 47912
rect 17309 47907 17375 47910
rect 19926 47908 19932 47910
rect 19996 47970 20002 47972
rect 21541 47970 21607 47973
rect 19996 47968 21607 47970
rect 19996 47912 21546 47968
rect 21602 47912 21607 47968
rect 19996 47910 21607 47912
rect 19996 47908 20002 47910
rect 21541 47907 21607 47910
rect 22737 47970 22803 47973
rect 24853 47970 24919 47973
rect 22737 47968 24919 47970
rect 22737 47912 22742 47968
rect 22798 47912 24858 47968
rect 24914 47912 24919 47968
rect 22737 47910 24919 47912
rect 22737 47907 22803 47910
rect 24853 47907 24919 47910
rect 5944 47904 6264 47905
rect 5944 47840 5952 47904
rect 6016 47840 6032 47904
rect 6096 47840 6112 47904
rect 6176 47840 6192 47904
rect 6256 47840 6264 47904
rect 5944 47839 6264 47840
rect 15944 47904 16264 47905
rect 15944 47840 15952 47904
rect 16016 47840 16032 47904
rect 16096 47840 16112 47904
rect 16176 47840 16192 47904
rect 16256 47840 16264 47904
rect 15944 47839 16264 47840
rect 25944 47904 26264 47905
rect 25944 47840 25952 47904
rect 26016 47840 26032 47904
rect 26096 47840 26112 47904
rect 26176 47840 26192 47904
rect 26256 47840 26264 47904
rect 25944 47839 26264 47840
rect 19977 47834 20043 47837
rect 23105 47834 23171 47837
rect 19977 47832 23171 47834
rect 19977 47776 19982 47832
rect 20038 47776 23110 47832
rect 23166 47776 23171 47832
rect 19977 47774 23171 47776
rect 19977 47771 20043 47774
rect 23105 47771 23171 47774
rect 16297 47698 16363 47701
rect 18137 47698 18203 47701
rect 16297 47696 18203 47698
rect 16297 47640 16302 47696
rect 16358 47640 18142 47696
rect 18198 47640 18203 47696
rect 16297 47638 18203 47640
rect 16297 47635 16363 47638
rect 18137 47635 18203 47638
rect 23974 47636 23980 47700
rect 24044 47698 24050 47700
rect 24117 47698 24183 47701
rect 26693 47698 26759 47701
rect 24044 47696 26759 47698
rect 24044 47640 24122 47696
rect 24178 47640 26698 47696
rect 26754 47640 26759 47696
rect 24044 47638 26759 47640
rect 24044 47636 24050 47638
rect 24117 47635 24183 47638
rect 26693 47635 26759 47638
rect 11973 47562 12039 47565
rect 17585 47562 17651 47565
rect 11973 47560 17651 47562
rect 11973 47504 11978 47560
rect 12034 47504 17590 47560
rect 17646 47504 17651 47560
rect 11973 47502 17651 47504
rect 11973 47499 12039 47502
rect 17585 47499 17651 47502
rect 14733 47426 14799 47429
rect 18229 47426 18295 47429
rect 14733 47424 18295 47426
rect 14733 47368 14738 47424
rect 14794 47368 18234 47424
rect 18290 47368 18295 47424
rect 14733 47366 18295 47368
rect 14733 47363 14799 47366
rect 18229 47363 18295 47366
rect 10944 47360 11264 47361
rect 10944 47296 10952 47360
rect 11016 47296 11032 47360
rect 11096 47296 11112 47360
rect 11176 47296 11192 47360
rect 11256 47296 11264 47360
rect 10944 47295 11264 47296
rect 20944 47360 21264 47361
rect 20944 47296 20952 47360
rect 21016 47296 21032 47360
rect 21096 47296 21112 47360
rect 21176 47296 21192 47360
rect 21256 47296 21264 47360
rect 20944 47295 21264 47296
rect 13997 47290 14063 47293
rect 17677 47290 17743 47293
rect 13997 47288 17743 47290
rect 13997 47232 14002 47288
rect 14058 47232 17682 47288
rect 17738 47232 17743 47288
rect 13997 47230 17743 47232
rect 13997 47227 14063 47230
rect 17677 47227 17743 47230
rect 23289 47290 23355 47293
rect 24301 47290 24367 47293
rect 25865 47290 25931 47293
rect 23289 47288 25931 47290
rect 23289 47232 23294 47288
rect 23350 47232 24306 47288
rect 24362 47232 25870 47288
rect 25926 47232 25931 47288
rect 23289 47230 25931 47232
rect 23289 47227 23355 47230
rect 24301 47227 24367 47230
rect 25865 47227 25931 47230
rect 15009 47154 15075 47157
rect 19425 47154 19491 47157
rect 15009 47152 19491 47154
rect 15009 47096 15014 47152
rect 15070 47096 19430 47152
rect 19486 47096 19491 47152
rect 15009 47094 19491 47096
rect 15009 47091 15075 47094
rect 19425 47091 19491 47094
rect 24485 47154 24551 47157
rect 26509 47154 26575 47157
rect 24485 47152 26575 47154
rect 24485 47096 24490 47152
rect 24546 47096 26514 47152
rect 26570 47096 26575 47152
rect 24485 47094 26575 47096
rect 24485 47091 24551 47094
rect 26509 47091 26575 47094
rect 0 47018 800 47048
rect 7373 47018 7439 47021
rect 0 47016 7439 47018
rect 0 46960 7378 47016
rect 7434 46960 7439 47016
rect 0 46958 7439 46960
rect 0 46928 800 46958
rect 7373 46955 7439 46958
rect 9622 46956 9628 47020
rect 9692 47018 9698 47020
rect 9765 47018 9831 47021
rect 9692 47016 9831 47018
rect 9692 46960 9770 47016
rect 9826 46960 9831 47016
rect 9692 46958 9831 46960
rect 9692 46956 9698 46958
rect 9765 46955 9831 46958
rect 15510 46956 15516 47020
rect 15580 47018 15586 47020
rect 16113 47018 16179 47021
rect 16481 47020 16547 47021
rect 16430 47018 16436 47020
rect 15580 47016 16179 47018
rect 15580 46960 16118 47016
rect 16174 46960 16179 47016
rect 15580 46958 16179 46960
rect 16390 46958 16436 47018
rect 16500 47016 16547 47020
rect 16542 46960 16547 47016
rect 15580 46956 15586 46958
rect 16113 46955 16179 46958
rect 16430 46956 16436 46958
rect 16500 46956 16547 46960
rect 16481 46955 16547 46956
rect 25681 47018 25747 47021
rect 29200 47018 30000 47048
rect 25681 47016 30000 47018
rect 25681 46960 25686 47016
rect 25742 46960 30000 47016
rect 25681 46958 30000 46960
rect 25681 46955 25747 46958
rect 29200 46928 30000 46958
rect 22369 46882 22435 46885
rect 17174 46880 22435 46882
rect 17174 46824 22374 46880
rect 22430 46824 22435 46880
rect 17174 46822 22435 46824
rect 5944 46816 6264 46817
rect 5944 46752 5952 46816
rect 6016 46752 6032 46816
rect 6096 46752 6112 46816
rect 6176 46752 6192 46816
rect 6256 46752 6264 46816
rect 5944 46751 6264 46752
rect 15944 46816 16264 46817
rect 15944 46752 15952 46816
rect 16016 46752 16032 46816
rect 16096 46752 16112 46816
rect 16176 46752 16192 46816
rect 16256 46752 16264 46816
rect 15944 46751 16264 46752
rect 8293 46610 8359 46613
rect 17174 46610 17234 46822
rect 22369 46819 22435 46822
rect 25944 46816 26264 46817
rect 25944 46752 25952 46816
rect 26016 46752 26032 46816
rect 26096 46752 26112 46816
rect 26176 46752 26192 46816
rect 26256 46752 26264 46816
rect 25944 46751 26264 46752
rect 20110 46684 20116 46748
rect 20180 46746 20186 46748
rect 23013 46746 23079 46749
rect 20180 46744 23079 46746
rect 20180 46688 23018 46744
rect 23074 46688 23079 46744
rect 20180 46686 23079 46688
rect 20180 46684 20186 46686
rect 23013 46683 23079 46686
rect 8293 46608 17234 46610
rect 8293 46552 8298 46608
rect 8354 46552 17234 46608
rect 8293 46550 17234 46552
rect 21725 46610 21791 46613
rect 23473 46610 23539 46613
rect 21725 46608 23539 46610
rect 21725 46552 21730 46608
rect 21786 46552 23478 46608
rect 23534 46552 23539 46608
rect 21725 46550 23539 46552
rect 8293 46547 8359 46550
rect 21725 46547 21791 46550
rect 23473 46547 23539 46550
rect 4061 46474 4127 46477
rect 9489 46474 9555 46477
rect 4061 46472 9555 46474
rect 4061 46416 4066 46472
rect 4122 46416 9494 46472
rect 9550 46416 9555 46472
rect 4061 46414 9555 46416
rect 4061 46411 4127 46414
rect 9489 46411 9555 46414
rect 15561 46338 15627 46341
rect 18137 46338 18203 46341
rect 15561 46336 18203 46338
rect 15561 46280 15566 46336
rect 15622 46280 18142 46336
rect 18198 46280 18203 46336
rect 15561 46278 18203 46280
rect 15561 46275 15627 46278
rect 18137 46275 18203 46278
rect 10944 46272 11264 46273
rect 10944 46208 10952 46272
rect 11016 46208 11032 46272
rect 11096 46208 11112 46272
rect 11176 46208 11192 46272
rect 11256 46208 11264 46272
rect 10944 46207 11264 46208
rect 20944 46272 21264 46273
rect 20944 46208 20952 46272
rect 21016 46208 21032 46272
rect 21096 46208 21112 46272
rect 21176 46208 21192 46272
rect 21256 46208 21264 46272
rect 20944 46207 21264 46208
rect 21817 46202 21883 46205
rect 22185 46202 22251 46205
rect 21817 46200 22251 46202
rect 21817 46144 21822 46200
rect 21878 46144 22190 46200
rect 22246 46144 22251 46200
rect 21817 46142 22251 46144
rect 21817 46139 21883 46142
rect 22185 46139 22251 46142
rect 21725 46066 21791 46069
rect 24117 46066 24183 46069
rect 21725 46064 24183 46066
rect 21725 46008 21730 46064
rect 21786 46008 24122 46064
rect 24178 46008 24183 46064
rect 21725 46006 24183 46008
rect 21725 46003 21791 46006
rect 24117 46003 24183 46006
rect 6269 45930 6335 45933
rect 16113 45930 16179 45933
rect 6269 45928 16179 45930
rect 6269 45872 6274 45928
rect 6330 45872 16118 45928
rect 16174 45872 16179 45928
rect 6269 45870 16179 45872
rect 6269 45867 6335 45870
rect 16113 45867 16179 45870
rect 16481 45930 16547 45933
rect 18873 45930 18939 45933
rect 16481 45928 18939 45930
rect 16481 45872 16486 45928
rect 16542 45872 18878 45928
rect 18934 45872 18939 45928
rect 16481 45870 18939 45872
rect 16481 45867 16547 45870
rect 18873 45867 18939 45870
rect 23105 45930 23171 45933
rect 26509 45930 26575 45933
rect 23105 45928 26575 45930
rect 23105 45872 23110 45928
rect 23166 45872 26514 45928
rect 26570 45872 26575 45928
rect 23105 45870 26575 45872
rect 23105 45867 23171 45870
rect 26509 45867 26575 45870
rect 17769 45794 17835 45797
rect 20069 45794 20135 45797
rect 17769 45792 20135 45794
rect 17769 45736 17774 45792
rect 17830 45736 20074 45792
rect 20130 45736 20135 45792
rect 17769 45734 20135 45736
rect 17769 45731 17835 45734
rect 20069 45731 20135 45734
rect 5944 45728 6264 45729
rect 0 45658 800 45688
rect 5944 45664 5952 45728
rect 6016 45664 6032 45728
rect 6096 45664 6112 45728
rect 6176 45664 6192 45728
rect 6256 45664 6264 45728
rect 5944 45663 6264 45664
rect 15944 45728 16264 45729
rect 15944 45664 15952 45728
rect 16016 45664 16032 45728
rect 16096 45664 16112 45728
rect 16176 45664 16192 45728
rect 16256 45664 16264 45728
rect 15944 45663 16264 45664
rect 25944 45728 26264 45729
rect 25944 45664 25952 45728
rect 26016 45664 26032 45728
rect 26096 45664 26112 45728
rect 26176 45664 26192 45728
rect 26256 45664 26264 45728
rect 25944 45663 26264 45664
rect 1945 45658 2011 45661
rect 0 45656 2011 45658
rect 0 45600 1950 45656
rect 2006 45600 2011 45656
rect 0 45598 2011 45600
rect 0 45568 800 45598
rect 1945 45595 2011 45598
rect 16849 45658 16915 45661
rect 20110 45658 20116 45660
rect 16849 45656 20116 45658
rect 16849 45600 16854 45656
rect 16910 45600 20116 45656
rect 16849 45598 20116 45600
rect 16849 45595 16915 45598
rect 20110 45596 20116 45598
rect 20180 45596 20186 45660
rect 25129 45658 25195 45661
rect 25262 45658 25268 45660
rect 25129 45656 25268 45658
rect 25129 45600 25134 45656
rect 25190 45600 25268 45656
rect 25129 45598 25268 45600
rect 25129 45595 25195 45598
rect 25262 45596 25268 45598
rect 25332 45596 25338 45660
rect 29200 45658 30000 45688
rect 26558 45598 30000 45658
rect 26417 45522 26483 45525
rect 26558 45522 26618 45598
rect 29200 45568 30000 45598
rect 26417 45520 26618 45522
rect 26417 45464 26422 45520
rect 26478 45464 26618 45520
rect 26417 45462 26618 45464
rect 26417 45459 26483 45462
rect 23289 45386 23355 45389
rect 25129 45386 25195 45389
rect 23289 45384 25195 45386
rect 23289 45328 23294 45384
rect 23350 45328 25134 45384
rect 25190 45328 25195 45384
rect 23289 45326 25195 45328
rect 23289 45323 23355 45326
rect 25129 45323 25195 45326
rect 10944 45184 11264 45185
rect 10944 45120 10952 45184
rect 11016 45120 11032 45184
rect 11096 45120 11112 45184
rect 11176 45120 11192 45184
rect 11256 45120 11264 45184
rect 10944 45119 11264 45120
rect 20944 45184 21264 45185
rect 20944 45120 20952 45184
rect 21016 45120 21032 45184
rect 21096 45120 21112 45184
rect 21176 45120 21192 45184
rect 21256 45120 21264 45184
rect 20944 45119 21264 45120
rect 23289 45114 23355 45117
rect 26325 45114 26391 45117
rect 23289 45112 26391 45114
rect 23289 45056 23294 45112
rect 23350 45056 26330 45112
rect 26386 45056 26391 45112
rect 23289 45054 26391 45056
rect 23289 45051 23355 45054
rect 26325 45051 26391 45054
rect 0 44978 800 45008
rect 1761 44978 1827 44981
rect 0 44976 1827 44978
rect 0 44920 1766 44976
rect 1822 44920 1827 44976
rect 0 44918 1827 44920
rect 0 44888 800 44918
rect 1761 44915 1827 44918
rect 23841 44978 23907 44981
rect 29200 44978 30000 45008
rect 23841 44976 30000 44978
rect 23841 44920 23846 44976
rect 23902 44920 30000 44976
rect 23841 44918 30000 44920
rect 23841 44915 23907 44918
rect 29200 44888 30000 44918
rect 6729 44842 6795 44845
rect 15653 44842 15719 44845
rect 20345 44844 20411 44845
rect 6729 44840 15719 44842
rect 6729 44784 6734 44840
rect 6790 44784 15658 44840
rect 15714 44784 15719 44840
rect 6729 44782 15719 44784
rect 6729 44779 6795 44782
rect 15653 44779 15719 44782
rect 20294 44780 20300 44844
rect 20364 44842 20411 44844
rect 21173 44842 21239 44845
rect 25405 44842 25471 44845
rect 26601 44842 26667 44845
rect 20364 44840 20456 44842
rect 20406 44784 20456 44840
rect 20364 44782 20456 44784
rect 21173 44840 25471 44842
rect 21173 44784 21178 44840
rect 21234 44784 25410 44840
rect 25466 44784 25471 44840
rect 21173 44782 25471 44784
rect 20364 44780 20411 44782
rect 20302 44779 20411 44780
rect 21173 44779 21239 44782
rect 25405 44779 25471 44782
rect 25822 44840 26667 44842
rect 25822 44784 26606 44840
rect 26662 44784 26667 44840
rect 25822 44782 26667 44784
rect 17217 44706 17283 44709
rect 19701 44706 19767 44709
rect 20302 44706 20362 44779
rect 17217 44704 20362 44706
rect 17217 44648 17222 44704
rect 17278 44648 19706 44704
rect 19762 44648 20362 44704
rect 17217 44646 20362 44648
rect 17217 44643 17283 44646
rect 19701 44643 19767 44646
rect 23054 44644 23060 44708
rect 23124 44706 23130 44708
rect 25822 44706 25882 44782
rect 26601 44779 26667 44782
rect 23124 44646 25882 44706
rect 23124 44644 23130 44646
rect 5944 44640 6264 44641
rect 5944 44576 5952 44640
rect 6016 44576 6032 44640
rect 6096 44576 6112 44640
rect 6176 44576 6192 44640
rect 6256 44576 6264 44640
rect 5944 44575 6264 44576
rect 15944 44640 16264 44641
rect 15944 44576 15952 44640
rect 16016 44576 16032 44640
rect 16096 44576 16112 44640
rect 16176 44576 16192 44640
rect 16256 44576 16264 44640
rect 15944 44575 16264 44576
rect 25944 44640 26264 44641
rect 25944 44576 25952 44640
rect 26016 44576 26032 44640
rect 26096 44576 26112 44640
rect 26176 44576 26192 44640
rect 26256 44576 26264 44640
rect 25944 44575 26264 44576
rect 2957 44570 3023 44573
rect 3182 44570 3188 44572
rect 2957 44568 3188 44570
rect 2957 44512 2962 44568
rect 3018 44512 3188 44568
rect 2957 44510 3188 44512
rect 2957 44507 3023 44510
rect 3182 44508 3188 44510
rect 3252 44508 3258 44572
rect 22645 44570 22711 44573
rect 17174 44568 22711 44570
rect 17174 44512 22650 44568
rect 22706 44512 22711 44568
rect 17174 44510 22711 44512
rect 7741 44434 7807 44437
rect 17174 44434 17234 44510
rect 22645 44507 22711 44510
rect 25037 44570 25103 44573
rect 25313 44570 25379 44573
rect 25037 44568 25379 44570
rect 25037 44512 25042 44568
rect 25098 44512 25318 44568
rect 25374 44512 25379 44568
rect 25037 44510 25379 44512
rect 25037 44507 25103 44510
rect 25313 44507 25379 44510
rect 7741 44432 17234 44434
rect 7741 44376 7746 44432
rect 7802 44376 17234 44432
rect 7741 44374 17234 44376
rect 17493 44434 17559 44437
rect 18873 44434 18939 44437
rect 23565 44434 23631 44437
rect 17493 44432 23631 44434
rect 17493 44376 17498 44432
rect 17554 44376 18878 44432
rect 18934 44376 23570 44432
rect 23626 44376 23631 44432
rect 17493 44374 23631 44376
rect 7741 44371 7807 44374
rect 17493 44371 17559 44374
rect 18873 44371 18939 44374
rect 23565 44371 23631 44374
rect 16113 44298 16179 44301
rect 18505 44298 18571 44301
rect 16113 44296 18571 44298
rect 16113 44240 16118 44296
rect 16174 44240 18510 44296
rect 18566 44240 18571 44296
rect 16113 44238 18571 44240
rect 16113 44235 16179 44238
rect 18505 44235 18571 44238
rect 17677 44162 17743 44165
rect 19885 44162 19951 44165
rect 17677 44160 19951 44162
rect 17677 44104 17682 44160
rect 17738 44104 19890 44160
rect 19946 44104 19951 44160
rect 17677 44102 19951 44104
rect 17677 44099 17743 44102
rect 19885 44099 19951 44102
rect 10944 44096 11264 44097
rect 10944 44032 10952 44096
rect 11016 44032 11032 44096
rect 11096 44032 11112 44096
rect 11176 44032 11192 44096
rect 11256 44032 11264 44096
rect 10944 44031 11264 44032
rect 20944 44096 21264 44097
rect 20944 44032 20952 44096
rect 21016 44032 21032 44096
rect 21096 44032 21112 44096
rect 21176 44032 21192 44096
rect 21256 44032 21264 44096
rect 20944 44031 21264 44032
rect 13997 44026 14063 44029
rect 19425 44026 19491 44029
rect 13997 44024 19491 44026
rect 13997 43968 14002 44024
rect 14058 43968 19430 44024
rect 19486 43968 19491 44024
rect 13997 43966 19491 43968
rect 13997 43963 14063 43966
rect 19425 43963 19491 43966
rect 23105 44026 23171 44029
rect 27521 44026 27587 44029
rect 23105 44024 27587 44026
rect 23105 43968 23110 44024
rect 23166 43968 27526 44024
rect 27582 43968 27587 44024
rect 23105 43966 27587 43968
rect 23105 43963 23171 43966
rect 27521 43963 27587 43966
rect 4061 43890 4127 43893
rect 8569 43890 8635 43893
rect 4061 43888 8635 43890
rect 4061 43832 4066 43888
rect 4122 43832 8574 43888
rect 8630 43832 8635 43888
rect 4061 43830 8635 43832
rect 4061 43827 4127 43830
rect 8569 43827 8635 43830
rect 8753 43890 8819 43893
rect 17217 43890 17283 43893
rect 8753 43888 17283 43890
rect 8753 43832 8758 43888
rect 8814 43832 17222 43888
rect 17278 43832 17283 43888
rect 8753 43830 17283 43832
rect 8753 43827 8819 43830
rect 17217 43827 17283 43830
rect 17585 43890 17651 43893
rect 21081 43890 21147 43893
rect 17585 43888 21147 43890
rect 17585 43832 17590 43888
rect 17646 43832 21086 43888
rect 21142 43832 21147 43888
rect 17585 43830 21147 43832
rect 17585 43827 17651 43830
rect 21081 43827 21147 43830
rect 24669 43890 24735 43893
rect 26877 43890 26943 43893
rect 24669 43888 26943 43890
rect 24669 43832 24674 43888
rect 24730 43832 26882 43888
rect 26938 43832 26943 43888
rect 24669 43830 26943 43832
rect 24669 43827 24735 43830
rect 26877 43827 26943 43830
rect 3141 43754 3207 43757
rect 24485 43754 24551 43757
rect 3141 43752 24551 43754
rect 3141 43696 3146 43752
rect 3202 43696 24490 43752
rect 24546 43696 24551 43752
rect 3141 43694 24551 43696
rect 3141 43691 3207 43694
rect 24485 43691 24551 43694
rect 25129 43754 25195 43757
rect 25129 43752 26434 43754
rect 25129 43696 25134 43752
rect 25190 43696 26434 43752
rect 25129 43694 26434 43696
rect 25129 43691 25195 43694
rect 0 43618 800 43648
rect 3417 43618 3483 43621
rect 0 43616 3483 43618
rect 0 43560 3422 43616
rect 3478 43560 3483 43616
rect 0 43558 3483 43560
rect 0 43528 800 43558
rect 3417 43555 3483 43558
rect 17217 43618 17283 43621
rect 22921 43618 22987 43621
rect 17217 43616 22987 43618
rect 17217 43560 17222 43616
rect 17278 43560 22926 43616
rect 22982 43560 22987 43616
rect 17217 43558 22987 43560
rect 26374 43618 26434 43694
rect 29200 43618 30000 43648
rect 26374 43558 30000 43618
rect 17217 43555 17283 43558
rect 22921 43555 22987 43558
rect 5944 43552 6264 43553
rect 5944 43488 5952 43552
rect 6016 43488 6032 43552
rect 6096 43488 6112 43552
rect 6176 43488 6192 43552
rect 6256 43488 6264 43552
rect 5944 43487 6264 43488
rect 15944 43552 16264 43553
rect 15944 43488 15952 43552
rect 16016 43488 16032 43552
rect 16096 43488 16112 43552
rect 16176 43488 16192 43552
rect 16256 43488 16264 43552
rect 15944 43487 16264 43488
rect 25944 43552 26264 43553
rect 25944 43488 25952 43552
rect 26016 43488 26032 43552
rect 26096 43488 26112 43552
rect 26176 43488 26192 43552
rect 26256 43488 26264 43552
rect 29200 43528 30000 43558
rect 25944 43487 26264 43488
rect 18045 43482 18111 43485
rect 22185 43482 22251 43485
rect 18045 43480 22251 43482
rect 18045 43424 18050 43480
rect 18106 43424 22190 43480
rect 22246 43424 22251 43480
rect 18045 43422 22251 43424
rect 18045 43419 18111 43422
rect 22185 43419 22251 43422
rect 23473 43346 23539 43349
rect 27245 43346 27311 43349
rect 23473 43344 27311 43346
rect 23473 43288 23478 43344
rect 23534 43288 27250 43344
rect 27306 43288 27311 43344
rect 23473 43286 27311 43288
rect 23473 43283 23539 43286
rect 27245 43283 27311 43286
rect 3141 43210 3207 43213
rect 19333 43210 19399 43213
rect 3141 43208 19399 43210
rect 3141 43152 3146 43208
rect 3202 43152 19338 43208
rect 19394 43152 19399 43208
rect 3141 43150 19399 43152
rect 3141 43147 3207 43150
rect 19333 43147 19399 43150
rect 3325 43074 3391 43077
rect 10593 43074 10659 43077
rect 3325 43072 10659 43074
rect 3325 43016 3330 43072
rect 3386 43016 10598 43072
rect 10654 43016 10659 43072
rect 3325 43014 10659 43016
rect 3325 43011 3391 43014
rect 10593 43011 10659 43014
rect 22829 43074 22895 43077
rect 25405 43074 25471 43077
rect 22829 43072 25471 43074
rect 22829 43016 22834 43072
rect 22890 43016 25410 43072
rect 25466 43016 25471 43072
rect 22829 43014 25471 43016
rect 22829 43011 22895 43014
rect 25405 43011 25471 43014
rect 10944 43008 11264 43009
rect 10944 42944 10952 43008
rect 11016 42944 11032 43008
rect 11096 42944 11112 43008
rect 11176 42944 11192 43008
rect 11256 42944 11264 43008
rect 10944 42943 11264 42944
rect 20944 43008 21264 43009
rect 20944 42944 20952 43008
rect 21016 42944 21032 43008
rect 21096 42944 21112 43008
rect 21176 42944 21192 43008
rect 21256 42944 21264 43008
rect 20944 42943 21264 42944
rect 13261 42938 13327 42941
rect 13670 42938 13676 42940
rect 13261 42936 13676 42938
rect 13261 42880 13266 42936
rect 13322 42880 13676 42936
rect 13261 42878 13676 42880
rect 13261 42875 13327 42878
rect 13670 42876 13676 42878
rect 13740 42876 13746 42940
rect 14641 42802 14707 42805
rect 19057 42802 19123 42805
rect 14641 42800 19123 42802
rect 14641 42744 14646 42800
rect 14702 42744 19062 42800
rect 19118 42744 19123 42800
rect 14641 42742 19123 42744
rect 14641 42739 14707 42742
rect 19057 42739 19123 42742
rect 22277 42802 22343 42805
rect 27337 42802 27403 42805
rect 22277 42800 27403 42802
rect 22277 42744 22282 42800
rect 22338 42744 27342 42800
rect 27398 42744 27403 42800
rect 22277 42742 27403 42744
rect 22277 42739 22343 42742
rect 27337 42739 27403 42742
rect 20437 42666 20503 42669
rect 27705 42666 27771 42669
rect 20437 42664 27771 42666
rect 20437 42608 20442 42664
rect 20498 42608 27710 42664
rect 27766 42608 27771 42664
rect 20437 42606 27771 42608
rect 20437 42603 20503 42606
rect 27705 42603 27771 42606
rect 5944 42464 6264 42465
rect 5944 42400 5952 42464
rect 6016 42400 6032 42464
rect 6096 42400 6112 42464
rect 6176 42400 6192 42464
rect 6256 42400 6264 42464
rect 5944 42399 6264 42400
rect 15944 42464 16264 42465
rect 15944 42400 15952 42464
rect 16016 42400 16032 42464
rect 16096 42400 16112 42464
rect 16176 42400 16192 42464
rect 16256 42400 16264 42464
rect 15944 42399 16264 42400
rect 25944 42464 26264 42465
rect 25944 42400 25952 42464
rect 26016 42400 26032 42464
rect 26096 42400 26112 42464
rect 26176 42400 26192 42464
rect 26256 42400 26264 42464
rect 25944 42399 26264 42400
rect 19885 42396 19951 42397
rect 19885 42394 19932 42396
rect 19840 42392 19932 42394
rect 19840 42336 19890 42392
rect 19840 42334 19932 42336
rect 19885 42332 19932 42334
rect 19996 42332 20002 42396
rect 19885 42331 19951 42332
rect 0 42258 800 42288
rect 14825 42258 14891 42261
rect 0 42256 14891 42258
rect 0 42200 14830 42256
rect 14886 42200 14891 42256
rect 0 42198 14891 42200
rect 0 42168 800 42198
rect 14825 42195 14891 42198
rect 23657 42258 23723 42261
rect 25957 42258 26023 42261
rect 26601 42258 26667 42261
rect 29200 42258 30000 42288
rect 23657 42256 26667 42258
rect 23657 42200 23662 42256
rect 23718 42200 25962 42256
rect 26018 42200 26606 42256
rect 26662 42200 26667 42256
rect 23657 42198 26667 42200
rect 23657 42195 23723 42198
rect 25957 42195 26023 42198
rect 26601 42195 26667 42198
rect 26742 42198 30000 42258
rect 9213 42122 9279 42125
rect 10777 42122 10843 42125
rect 9213 42120 10843 42122
rect 9213 42064 9218 42120
rect 9274 42064 10782 42120
rect 10838 42064 10843 42120
rect 9213 42062 10843 42064
rect 9213 42059 9279 42062
rect 10777 42059 10843 42062
rect 12382 42060 12388 42124
rect 12452 42122 12458 42124
rect 15101 42122 15167 42125
rect 26509 42122 26575 42125
rect 12452 42120 26575 42122
rect 12452 42064 15106 42120
rect 15162 42064 26514 42120
rect 26570 42064 26575 42120
rect 12452 42062 26575 42064
rect 12452 42060 12458 42062
rect 15101 42059 15167 42062
rect 26509 42059 26575 42062
rect 20069 41988 20135 41989
rect 20069 41986 20116 41988
rect 20024 41984 20116 41986
rect 20024 41928 20074 41984
rect 20024 41926 20116 41928
rect 20069 41924 20116 41926
rect 20180 41924 20186 41988
rect 25405 41986 25471 41989
rect 26742 41986 26802 42198
rect 29200 42168 30000 42198
rect 25405 41984 26802 41986
rect 25405 41928 25410 41984
rect 25466 41928 26802 41984
rect 25405 41926 26802 41928
rect 20069 41923 20135 41924
rect 25405 41923 25471 41926
rect 10944 41920 11264 41921
rect 10944 41856 10952 41920
rect 11016 41856 11032 41920
rect 11096 41856 11112 41920
rect 11176 41856 11192 41920
rect 11256 41856 11264 41920
rect 10944 41855 11264 41856
rect 20944 41920 21264 41921
rect 20944 41856 20952 41920
rect 21016 41856 21032 41920
rect 21096 41856 21112 41920
rect 21176 41856 21192 41920
rect 21256 41856 21264 41920
rect 20944 41855 21264 41856
rect 12934 41788 12940 41852
rect 13004 41850 13010 41852
rect 13997 41850 14063 41853
rect 13004 41848 14063 41850
rect 13004 41792 14002 41848
rect 14058 41792 14063 41848
rect 13004 41790 14063 41792
rect 13004 41788 13010 41790
rect 13997 41787 14063 41790
rect 24301 41850 24367 41853
rect 24669 41850 24735 41853
rect 24301 41848 24735 41850
rect 24301 41792 24306 41848
rect 24362 41792 24674 41848
rect 24730 41792 24735 41848
rect 24301 41790 24735 41792
rect 24301 41787 24367 41790
rect 24669 41787 24735 41790
rect 25037 41850 25103 41853
rect 25037 41848 27354 41850
rect 25037 41792 25042 41848
rect 25098 41792 27354 41848
rect 25037 41790 27354 41792
rect 25037 41787 25103 41790
rect 20713 41714 20779 41717
rect 22921 41714 22987 41717
rect 20713 41712 22987 41714
rect 20713 41656 20718 41712
rect 20774 41656 22926 41712
rect 22982 41656 22987 41712
rect 20713 41654 22987 41656
rect 20713 41651 20779 41654
rect 22921 41651 22987 41654
rect 23197 41714 23263 41717
rect 27061 41714 27127 41717
rect 23197 41712 27127 41714
rect 23197 41656 23202 41712
rect 23258 41656 27066 41712
rect 27122 41656 27127 41712
rect 23197 41654 27127 41656
rect 23197 41651 23263 41654
rect 27061 41651 27127 41654
rect 0 41578 800 41608
rect 1761 41578 1827 41581
rect 0 41576 1827 41578
rect 0 41520 1766 41576
rect 1822 41520 1827 41576
rect 0 41518 1827 41520
rect 0 41488 800 41518
rect 1761 41515 1827 41518
rect 20478 41516 20484 41580
rect 20548 41578 20554 41580
rect 20713 41578 20779 41581
rect 20548 41576 20779 41578
rect 20548 41520 20718 41576
rect 20774 41520 20779 41576
rect 20548 41518 20779 41520
rect 20548 41516 20554 41518
rect 20713 41515 20779 41518
rect 24710 41516 24716 41580
rect 24780 41578 24786 41580
rect 25497 41578 25563 41581
rect 24780 41576 25563 41578
rect 24780 41520 25502 41576
rect 25558 41520 25563 41576
rect 24780 41518 25563 41520
rect 27294 41578 27354 41790
rect 29200 41578 30000 41608
rect 27294 41518 30000 41578
rect 24780 41516 24786 41518
rect 25497 41515 25563 41518
rect 29200 41488 30000 41518
rect 2313 41442 2379 41445
rect 3233 41442 3299 41445
rect 2313 41440 3299 41442
rect 2313 41384 2318 41440
rect 2374 41384 3238 41440
rect 3294 41384 3299 41440
rect 2313 41382 3299 41384
rect 2313 41379 2379 41382
rect 3233 41379 3299 41382
rect 9029 41442 9095 41445
rect 10409 41442 10475 41445
rect 9029 41440 10475 41442
rect 9029 41384 9034 41440
rect 9090 41384 10414 41440
rect 10470 41384 10475 41440
rect 9029 41382 10475 41384
rect 9029 41379 9095 41382
rect 10409 41379 10475 41382
rect 20253 41442 20319 41445
rect 20478 41442 20484 41444
rect 20253 41440 20484 41442
rect 20253 41384 20258 41440
rect 20314 41384 20484 41440
rect 20253 41382 20484 41384
rect 20253 41379 20319 41382
rect 20478 41380 20484 41382
rect 20548 41380 20554 41444
rect 23054 41380 23060 41444
rect 23124 41442 23130 41444
rect 23197 41442 23263 41445
rect 24577 41442 24643 41445
rect 23124 41440 24643 41442
rect 23124 41384 23202 41440
rect 23258 41384 24582 41440
rect 24638 41384 24643 41440
rect 23124 41382 24643 41384
rect 23124 41380 23130 41382
rect 23197 41379 23263 41382
rect 24577 41379 24643 41382
rect 5944 41376 6264 41377
rect 5944 41312 5952 41376
rect 6016 41312 6032 41376
rect 6096 41312 6112 41376
rect 6176 41312 6192 41376
rect 6256 41312 6264 41376
rect 5944 41311 6264 41312
rect 15944 41376 16264 41377
rect 15944 41312 15952 41376
rect 16016 41312 16032 41376
rect 16096 41312 16112 41376
rect 16176 41312 16192 41376
rect 16256 41312 16264 41376
rect 15944 41311 16264 41312
rect 25944 41376 26264 41377
rect 25944 41312 25952 41376
rect 26016 41312 26032 41376
rect 26096 41312 26112 41376
rect 26176 41312 26192 41376
rect 26256 41312 26264 41376
rect 25944 41311 26264 41312
rect 11697 41306 11763 41309
rect 15745 41306 15811 41309
rect 20529 41306 20595 41309
rect 21909 41306 21975 41309
rect 11697 41304 15811 41306
rect 11697 41248 11702 41304
rect 11758 41248 15750 41304
rect 15806 41248 15811 41304
rect 11697 41246 15811 41248
rect 11697 41243 11763 41246
rect 15745 41243 15811 41246
rect 19796 41304 20595 41306
rect 19796 41248 20534 41304
rect 20590 41248 20595 41304
rect 19796 41246 20595 41248
rect 19796 41173 19856 41246
rect 20529 41243 20595 41246
rect 21774 41304 21975 41306
rect 21774 41248 21914 41304
rect 21970 41248 21975 41304
rect 21774 41246 21975 41248
rect 11881 41170 11947 41173
rect 15101 41170 15167 41173
rect 11881 41168 15167 41170
rect 11881 41112 11886 41168
rect 11942 41112 15106 41168
rect 15162 41112 15167 41168
rect 11881 41110 15167 41112
rect 11881 41107 11947 41110
rect 15101 41107 15167 41110
rect 19793 41168 19859 41173
rect 20529 41172 20595 41173
rect 20478 41170 20484 41172
rect 19793 41112 19798 41168
rect 19854 41112 19859 41168
rect 19793 41107 19859 41112
rect 20438 41110 20484 41170
rect 20548 41168 20595 41172
rect 20590 41112 20595 41168
rect 20478 41108 20484 41110
rect 20548 41108 20595 41112
rect 20662 41108 20668 41172
rect 20732 41170 20738 41172
rect 21173 41170 21239 41173
rect 21541 41170 21607 41173
rect 20732 41168 21239 41170
rect 20732 41112 21178 41168
rect 21234 41112 21239 41168
rect 20732 41110 21239 41112
rect 20732 41108 20738 41110
rect 20529 41107 20595 41108
rect 21173 41107 21239 41110
rect 21406 41168 21607 41170
rect 21406 41112 21546 41168
rect 21602 41112 21607 41168
rect 21406 41110 21607 41112
rect 18965 41034 19031 41037
rect 21406 41034 21466 41110
rect 21541 41107 21607 41110
rect 18965 41032 21466 41034
rect 18965 40976 18970 41032
rect 19026 40976 21466 41032
rect 18965 40974 21466 40976
rect 18965 40971 19031 40974
rect 13077 40898 13143 40901
rect 18137 40898 18203 40901
rect 13077 40896 18203 40898
rect 13077 40840 13082 40896
rect 13138 40840 18142 40896
rect 18198 40840 18203 40896
rect 13077 40838 18203 40840
rect 13077 40835 13143 40838
rect 18137 40835 18203 40838
rect 20478 40836 20484 40900
rect 20548 40898 20554 40900
rect 20805 40898 20871 40901
rect 20548 40896 20871 40898
rect 20548 40840 20810 40896
rect 20866 40840 20871 40896
rect 20548 40838 20871 40840
rect 20548 40836 20554 40838
rect 20805 40835 20871 40838
rect 10944 40832 11264 40833
rect 10944 40768 10952 40832
rect 11016 40768 11032 40832
rect 11096 40768 11112 40832
rect 11176 40768 11192 40832
rect 11256 40768 11264 40832
rect 10944 40767 11264 40768
rect 20944 40832 21264 40833
rect 20944 40768 20952 40832
rect 21016 40768 21032 40832
rect 21096 40768 21112 40832
rect 21176 40768 21192 40832
rect 21256 40768 21264 40832
rect 20944 40767 21264 40768
rect 21774 40765 21834 41246
rect 21909 41243 21975 41246
rect 23974 40836 23980 40900
rect 24044 40898 24050 40900
rect 24301 40898 24367 40901
rect 24044 40896 24367 40898
rect 24044 40840 24306 40896
rect 24362 40840 24367 40896
rect 24044 40838 24367 40840
rect 24044 40836 24050 40838
rect 24301 40835 24367 40838
rect 21774 40760 21883 40765
rect 21774 40704 21822 40760
rect 21878 40704 21883 40760
rect 21774 40702 21883 40704
rect 21817 40699 21883 40702
rect 5944 40288 6264 40289
rect 0 40218 800 40248
rect 5944 40224 5952 40288
rect 6016 40224 6032 40288
rect 6096 40224 6112 40288
rect 6176 40224 6192 40288
rect 6256 40224 6264 40288
rect 5944 40223 6264 40224
rect 15944 40288 16264 40289
rect 15944 40224 15952 40288
rect 16016 40224 16032 40288
rect 16096 40224 16112 40288
rect 16176 40224 16192 40288
rect 16256 40224 16264 40288
rect 15944 40223 16264 40224
rect 25944 40288 26264 40289
rect 25944 40224 25952 40288
rect 26016 40224 26032 40288
rect 26096 40224 26112 40288
rect 26176 40224 26192 40288
rect 26256 40224 26264 40288
rect 25944 40223 26264 40224
rect 2129 40218 2195 40221
rect 29200 40218 30000 40248
rect 0 40216 2195 40218
rect 0 40160 2134 40216
rect 2190 40160 2195 40216
rect 0 40158 2195 40160
rect 0 40128 800 40158
rect 2129 40155 2195 40158
rect 26604 40158 30000 40218
rect 9949 40082 10015 40085
rect 15653 40082 15719 40085
rect 15929 40082 15995 40085
rect 9949 40080 15995 40082
rect 9949 40024 9954 40080
rect 10010 40024 15658 40080
rect 15714 40024 15934 40080
rect 15990 40024 15995 40080
rect 9949 40022 15995 40024
rect 9949 40019 10015 40022
rect 15653 40019 15719 40022
rect 15929 40019 15995 40022
rect 25865 40082 25931 40085
rect 26604 40082 26664 40158
rect 29200 40128 30000 40158
rect 25865 40080 26664 40082
rect 25865 40024 25870 40080
rect 25926 40024 26664 40080
rect 25865 40022 26664 40024
rect 25865 40019 25931 40022
rect 13445 39946 13511 39949
rect 19425 39946 19491 39949
rect 13445 39944 19491 39946
rect 13445 39888 13450 39944
rect 13506 39888 19430 39944
rect 19486 39888 19491 39944
rect 13445 39886 19491 39888
rect 13445 39883 13511 39886
rect 19425 39883 19491 39886
rect 21541 39946 21607 39949
rect 23473 39946 23539 39949
rect 21541 39944 23539 39946
rect 21541 39888 21546 39944
rect 21602 39888 23478 39944
rect 23534 39888 23539 39944
rect 21541 39886 23539 39888
rect 21541 39883 21607 39886
rect 23473 39883 23539 39886
rect 13486 39748 13492 39812
rect 13556 39810 13562 39812
rect 13629 39810 13695 39813
rect 13556 39808 13695 39810
rect 13556 39752 13634 39808
rect 13690 39752 13695 39808
rect 13556 39750 13695 39752
rect 13556 39748 13562 39750
rect 13629 39747 13695 39750
rect 10944 39744 11264 39745
rect 10944 39680 10952 39744
rect 11016 39680 11032 39744
rect 11096 39680 11112 39744
rect 11176 39680 11192 39744
rect 11256 39680 11264 39744
rect 10944 39679 11264 39680
rect 20944 39744 21264 39745
rect 20944 39680 20952 39744
rect 21016 39680 21032 39744
rect 21096 39680 21112 39744
rect 21176 39680 21192 39744
rect 21256 39680 21264 39744
rect 20944 39679 21264 39680
rect 11421 39674 11487 39677
rect 12750 39674 12756 39676
rect 11421 39672 12756 39674
rect 11421 39616 11426 39672
rect 11482 39616 12756 39672
rect 11421 39614 12756 39616
rect 11421 39611 11487 39614
rect 12750 39612 12756 39614
rect 12820 39674 12826 39676
rect 13302 39674 13308 39676
rect 12820 39614 13308 39674
rect 12820 39612 12826 39614
rect 13302 39612 13308 39614
rect 13372 39612 13378 39676
rect 3141 39538 3207 39541
rect 21173 39538 21239 39541
rect 3141 39536 21239 39538
rect 3141 39480 3146 39536
rect 3202 39480 21178 39536
rect 21234 39480 21239 39536
rect 3141 39478 21239 39480
rect 3141 39475 3207 39478
rect 21173 39475 21239 39478
rect 13302 39340 13308 39404
rect 13372 39402 13378 39404
rect 13372 39342 16498 39402
rect 13372 39340 13378 39342
rect 5944 39200 6264 39201
rect 5944 39136 5952 39200
rect 6016 39136 6032 39200
rect 6096 39136 6112 39200
rect 6176 39136 6192 39200
rect 6256 39136 6264 39200
rect 5944 39135 6264 39136
rect 15944 39200 16264 39201
rect 15944 39136 15952 39200
rect 16016 39136 16032 39200
rect 16096 39136 16112 39200
rect 16176 39136 16192 39200
rect 16256 39136 16264 39200
rect 15944 39135 16264 39136
rect 16438 39130 16498 39342
rect 18689 39266 18755 39269
rect 24710 39266 24716 39268
rect 18689 39264 24716 39266
rect 18689 39208 18694 39264
rect 18750 39208 24716 39264
rect 18689 39206 24716 39208
rect 18689 39203 18755 39206
rect 24710 39204 24716 39206
rect 24780 39204 24786 39268
rect 25944 39200 26264 39201
rect 25944 39136 25952 39200
rect 26016 39136 26032 39200
rect 26096 39136 26112 39200
rect 26176 39136 26192 39200
rect 26256 39136 26264 39200
rect 25944 39135 26264 39136
rect 24485 39130 24551 39133
rect 16438 39128 24551 39130
rect 16438 39072 24490 39128
rect 24546 39072 24551 39128
rect 16438 39070 24551 39072
rect 24485 39067 24551 39070
rect 3141 38994 3207 38997
rect 3141 38992 17970 38994
rect 3141 38936 3146 38992
rect 3202 38936 17970 38992
rect 3141 38934 17970 38936
rect 3141 38931 3207 38934
rect 0 38858 800 38888
rect 8293 38858 8359 38861
rect 0 38856 8359 38858
rect 0 38800 8298 38856
rect 8354 38800 8359 38856
rect 0 38798 8359 38800
rect 0 38768 800 38798
rect 8293 38795 8359 38798
rect 13537 38858 13603 38861
rect 16481 38858 16547 38861
rect 13537 38856 16547 38858
rect 13537 38800 13542 38856
rect 13598 38800 16486 38856
rect 16542 38800 16547 38856
rect 13537 38798 16547 38800
rect 13537 38795 13603 38798
rect 16481 38795 16547 38798
rect 10944 38656 11264 38657
rect 10944 38592 10952 38656
rect 11016 38592 11032 38656
rect 11096 38592 11112 38656
rect 11176 38592 11192 38656
rect 11256 38592 11264 38656
rect 10944 38591 11264 38592
rect 11973 38586 12039 38589
rect 12985 38586 13051 38589
rect 11973 38584 13051 38586
rect 11973 38528 11978 38584
rect 12034 38528 12990 38584
rect 13046 38528 13051 38584
rect 11973 38526 13051 38528
rect 11973 38523 12039 38526
rect 12985 38523 13051 38526
rect 8661 38450 8727 38453
rect 10869 38450 10935 38453
rect 13118 38450 13124 38452
rect 8661 38448 13124 38450
rect 8661 38392 8666 38448
rect 8722 38392 10874 38448
rect 10930 38392 13124 38448
rect 8661 38390 13124 38392
rect 8661 38387 8727 38390
rect 10869 38387 10935 38390
rect 13118 38388 13124 38390
rect 13188 38450 13194 38452
rect 13721 38450 13787 38453
rect 13188 38448 13787 38450
rect 13188 38392 13726 38448
rect 13782 38392 13787 38448
rect 13188 38390 13787 38392
rect 17910 38450 17970 38934
rect 19517 38858 19583 38861
rect 21725 38858 21791 38861
rect 19517 38856 21791 38858
rect 19517 38800 19522 38856
rect 19578 38800 21730 38856
rect 21786 38800 21791 38856
rect 19517 38798 21791 38800
rect 19517 38795 19583 38798
rect 21725 38795 21791 38798
rect 26417 38858 26483 38861
rect 29200 38858 30000 38888
rect 26417 38856 30000 38858
rect 26417 38800 26422 38856
rect 26478 38800 30000 38856
rect 26417 38798 30000 38800
rect 26417 38795 26483 38798
rect 29200 38768 30000 38798
rect 21766 38660 21772 38724
rect 21836 38722 21842 38724
rect 21909 38722 21975 38725
rect 21836 38720 21975 38722
rect 21836 38664 21914 38720
rect 21970 38664 21975 38720
rect 21836 38662 21975 38664
rect 21836 38660 21842 38662
rect 21909 38659 21975 38662
rect 20944 38656 21264 38657
rect 20944 38592 20952 38656
rect 21016 38592 21032 38656
rect 21096 38592 21112 38656
rect 21176 38592 21192 38656
rect 21256 38592 21264 38656
rect 20944 38591 21264 38592
rect 25497 38588 25563 38589
rect 25446 38586 25452 38588
rect 25406 38526 25452 38586
rect 25516 38584 25563 38588
rect 25558 38528 25563 38584
rect 25446 38524 25452 38526
rect 25516 38524 25563 38528
rect 25497 38523 25563 38524
rect 23657 38450 23723 38453
rect 17910 38448 23723 38450
rect 17910 38392 23662 38448
rect 23718 38392 23723 38448
rect 17910 38390 23723 38392
rect 13188 38388 13194 38390
rect 13721 38387 13787 38390
rect 23657 38387 23723 38390
rect 24342 38388 24348 38452
rect 24412 38450 24418 38452
rect 25446 38450 25452 38452
rect 24412 38390 25452 38450
rect 24412 38388 24418 38390
rect 25446 38388 25452 38390
rect 25516 38388 25522 38452
rect 24761 38314 24827 38317
rect 24761 38312 26434 38314
rect 24761 38256 24766 38312
rect 24822 38256 26434 38312
rect 24761 38254 26434 38256
rect 24761 38251 24827 38254
rect 9029 38178 9095 38181
rect 12525 38178 12591 38181
rect 9029 38176 12591 38178
rect 9029 38120 9034 38176
rect 9090 38120 12530 38176
rect 12586 38120 12591 38176
rect 9029 38118 12591 38120
rect 9029 38115 9095 38118
rect 12525 38115 12591 38118
rect 20529 38178 20595 38181
rect 25589 38178 25655 38181
rect 20529 38176 25655 38178
rect 20529 38120 20534 38176
rect 20590 38120 25594 38176
rect 25650 38120 25655 38176
rect 20529 38118 25655 38120
rect 26374 38178 26434 38254
rect 29200 38178 30000 38208
rect 26374 38118 30000 38178
rect 20529 38115 20595 38118
rect 25589 38115 25655 38118
rect 5944 38112 6264 38113
rect 5944 38048 5952 38112
rect 6016 38048 6032 38112
rect 6096 38048 6112 38112
rect 6176 38048 6192 38112
rect 6256 38048 6264 38112
rect 5944 38047 6264 38048
rect 15944 38112 16264 38113
rect 15944 38048 15952 38112
rect 16016 38048 16032 38112
rect 16096 38048 16112 38112
rect 16176 38048 16192 38112
rect 16256 38048 16264 38112
rect 15944 38047 16264 38048
rect 25944 38112 26264 38113
rect 25944 38048 25952 38112
rect 26016 38048 26032 38112
rect 26096 38048 26112 38112
rect 26176 38048 26192 38112
rect 26256 38048 26264 38112
rect 29200 38088 30000 38118
rect 25944 38047 26264 38048
rect 9397 38042 9463 38045
rect 11329 38042 11395 38045
rect 9397 38040 11395 38042
rect 9397 37984 9402 38040
rect 9458 37984 11334 38040
rect 11390 37984 11395 38040
rect 9397 37982 11395 37984
rect 9397 37979 9463 37982
rect 11329 37979 11395 37982
rect 16849 38042 16915 38045
rect 18505 38042 18571 38045
rect 16849 38040 18571 38042
rect 16849 37984 16854 38040
rect 16910 37984 18510 38040
rect 18566 37984 18571 38040
rect 16849 37982 18571 37984
rect 16849 37979 16915 37982
rect 18505 37979 18571 37982
rect 13169 37906 13235 37909
rect 15469 37906 15535 37909
rect 13169 37904 15535 37906
rect 13169 37848 13174 37904
rect 13230 37848 15474 37904
rect 15530 37848 15535 37904
rect 13169 37846 15535 37848
rect 13169 37843 13235 37846
rect 15469 37843 15535 37846
rect 8201 37770 8267 37773
rect 10225 37770 10291 37773
rect 8201 37768 10291 37770
rect 8201 37712 8206 37768
rect 8262 37712 10230 37768
rect 10286 37712 10291 37768
rect 8201 37710 10291 37712
rect 8201 37707 8267 37710
rect 10225 37707 10291 37710
rect 10358 37708 10364 37772
rect 10428 37770 10434 37772
rect 13077 37770 13143 37773
rect 13537 37770 13603 37773
rect 16573 37770 16639 37773
rect 10428 37710 11484 37770
rect 10428 37708 10434 37710
rect 9857 37636 9923 37637
rect 9806 37572 9812 37636
rect 9876 37634 9923 37636
rect 11424 37634 11484 37710
rect 13077 37768 16639 37770
rect 13077 37712 13082 37768
rect 13138 37712 13542 37768
rect 13598 37712 16578 37768
rect 16634 37712 16639 37768
rect 13077 37710 16639 37712
rect 13077 37707 13143 37710
rect 13537 37707 13603 37710
rect 16573 37707 16639 37710
rect 19374 37708 19380 37772
rect 19444 37770 19450 37772
rect 20345 37770 20411 37773
rect 19444 37768 20411 37770
rect 19444 37712 20350 37768
rect 20406 37712 20411 37768
rect 19444 37710 20411 37712
rect 19444 37708 19450 37710
rect 20345 37707 20411 37710
rect 14273 37634 14339 37637
rect 9876 37632 9968 37634
rect 9918 37576 9968 37632
rect 9876 37574 9968 37576
rect 11424 37632 14339 37634
rect 11424 37576 14278 37632
rect 14334 37576 14339 37632
rect 11424 37574 14339 37576
rect 9876 37572 9923 37574
rect 9857 37571 9923 37572
rect 14273 37571 14339 37574
rect 14457 37634 14523 37637
rect 14590 37634 14596 37636
rect 14457 37632 14596 37634
rect 14457 37576 14462 37632
rect 14518 37576 14596 37632
rect 14457 37574 14596 37576
rect 14457 37571 14523 37574
rect 14590 37572 14596 37574
rect 14660 37572 14666 37636
rect 10944 37568 11264 37569
rect 0 37498 800 37528
rect 10944 37504 10952 37568
rect 11016 37504 11032 37568
rect 11096 37504 11112 37568
rect 11176 37504 11192 37568
rect 11256 37504 11264 37568
rect 10944 37503 11264 37504
rect 20944 37568 21264 37569
rect 20944 37504 20952 37568
rect 21016 37504 21032 37568
rect 21096 37504 21112 37568
rect 21176 37504 21192 37568
rect 21256 37504 21264 37568
rect 20944 37503 21264 37504
rect 1669 37498 1735 37501
rect 0 37496 1735 37498
rect 0 37440 1674 37496
rect 1730 37440 1735 37496
rect 0 37438 1735 37440
rect 0 37408 800 37438
rect 1669 37435 1735 37438
rect 14917 37498 14983 37501
rect 16798 37498 16804 37500
rect 14917 37496 16804 37498
rect 14917 37440 14922 37496
rect 14978 37440 16804 37496
rect 14917 37438 16804 37440
rect 14917 37435 14983 37438
rect 16798 37436 16804 37438
rect 16868 37436 16874 37500
rect 8477 37362 8543 37365
rect 9622 37362 9628 37364
rect 8477 37360 9628 37362
rect 8477 37304 8482 37360
rect 8538 37304 9628 37360
rect 8477 37302 9628 37304
rect 8477 37299 8543 37302
rect 9622 37300 9628 37302
rect 9692 37362 9698 37364
rect 10174 37362 10180 37364
rect 9692 37302 10180 37362
rect 9692 37300 9698 37302
rect 10174 37300 10180 37302
rect 10244 37300 10250 37364
rect 10869 37362 10935 37365
rect 14641 37362 14707 37365
rect 10869 37360 14707 37362
rect 10869 37304 10874 37360
rect 10930 37304 14646 37360
rect 14702 37304 14707 37360
rect 10869 37302 14707 37304
rect 10869 37299 10935 37302
rect 14641 37299 14707 37302
rect 15745 37362 15811 37365
rect 17217 37362 17283 37365
rect 15745 37360 17283 37362
rect 15745 37304 15750 37360
rect 15806 37304 17222 37360
rect 17278 37304 17283 37360
rect 15745 37302 17283 37304
rect 15745 37299 15811 37302
rect 17217 37299 17283 37302
rect 21541 37362 21607 37365
rect 22737 37362 22803 37365
rect 21541 37360 22803 37362
rect 21541 37304 21546 37360
rect 21602 37304 22742 37360
rect 22798 37304 22803 37360
rect 21541 37302 22803 37304
rect 21541 37299 21607 37302
rect 22737 37299 22803 37302
rect 5073 37226 5139 37229
rect 11237 37226 11303 37229
rect 5073 37224 11303 37226
rect 5073 37168 5078 37224
rect 5134 37168 11242 37224
rect 11298 37168 11303 37224
rect 5073 37166 11303 37168
rect 5073 37163 5139 37166
rect 11237 37163 11303 37166
rect 13445 37226 13511 37229
rect 15929 37226 15995 37229
rect 13445 37224 15995 37226
rect 13445 37168 13450 37224
rect 13506 37168 15934 37224
rect 15990 37168 15995 37224
rect 13445 37166 15995 37168
rect 13445 37163 13511 37166
rect 15929 37163 15995 37166
rect 16113 37226 16179 37229
rect 16614 37226 16620 37228
rect 16113 37224 16620 37226
rect 16113 37168 16118 37224
rect 16174 37168 16620 37224
rect 16113 37166 16620 37168
rect 16113 37163 16179 37166
rect 16614 37164 16620 37166
rect 16684 37164 16690 37228
rect 8293 37090 8359 37093
rect 10542 37090 10548 37092
rect 8293 37088 10548 37090
rect 8293 37032 8298 37088
rect 8354 37032 10548 37088
rect 8293 37030 10548 37032
rect 8293 37027 8359 37030
rect 10542 37028 10548 37030
rect 10612 37028 10618 37092
rect 14733 37090 14799 37093
rect 15745 37090 15811 37093
rect 14733 37088 15811 37090
rect 14733 37032 14738 37088
rect 14794 37032 15750 37088
rect 15806 37032 15811 37088
rect 14733 37030 15811 37032
rect 14733 37027 14799 37030
rect 15745 37027 15811 37030
rect 16389 37090 16455 37093
rect 22369 37090 22435 37093
rect 16389 37088 22435 37090
rect 16389 37032 16394 37088
rect 16450 37032 22374 37088
rect 22430 37032 22435 37088
rect 16389 37030 22435 37032
rect 16389 37027 16455 37030
rect 22369 37027 22435 37030
rect 23790 37028 23796 37092
rect 23860 37090 23866 37092
rect 23933 37090 23999 37093
rect 23860 37088 23999 37090
rect 23860 37032 23938 37088
rect 23994 37032 23999 37088
rect 23860 37030 23999 37032
rect 23860 37028 23866 37030
rect 23933 37027 23999 37030
rect 5944 37024 6264 37025
rect 5944 36960 5952 37024
rect 6016 36960 6032 37024
rect 6096 36960 6112 37024
rect 6176 36960 6192 37024
rect 6256 36960 6264 37024
rect 5944 36959 6264 36960
rect 15944 37024 16264 37025
rect 15944 36960 15952 37024
rect 16016 36960 16032 37024
rect 16096 36960 16112 37024
rect 16176 36960 16192 37024
rect 16256 36960 16264 37024
rect 15944 36959 16264 36960
rect 25944 37024 26264 37025
rect 25944 36960 25952 37024
rect 26016 36960 26032 37024
rect 26096 36960 26112 37024
rect 26176 36960 26192 37024
rect 26256 36960 26264 37024
rect 25944 36959 26264 36960
rect 6821 36954 6887 36957
rect 11053 36954 11119 36957
rect 6821 36952 11119 36954
rect 6821 36896 6826 36952
rect 6882 36896 11058 36952
rect 11114 36896 11119 36952
rect 6821 36894 11119 36896
rect 6821 36891 6887 36894
rect 11053 36891 11119 36894
rect 13261 36954 13327 36957
rect 13261 36952 15762 36954
rect 13261 36896 13266 36952
rect 13322 36896 15762 36952
rect 13261 36894 15762 36896
rect 13261 36891 13327 36894
rect 0 36818 800 36848
rect 6545 36818 6611 36821
rect 0 36816 6611 36818
rect 0 36760 6550 36816
rect 6606 36760 6611 36816
rect 0 36758 6611 36760
rect 0 36728 800 36758
rect 6545 36755 6611 36758
rect 8201 36818 8267 36821
rect 11145 36818 11211 36821
rect 8201 36816 11211 36818
rect 8201 36760 8206 36816
rect 8262 36760 11150 36816
rect 11206 36760 11211 36816
rect 8201 36758 11211 36760
rect 8201 36755 8267 36758
rect 11145 36755 11211 36758
rect 12985 36818 13051 36821
rect 15702 36818 15762 36894
rect 17677 36818 17743 36821
rect 12985 36816 15578 36818
rect 12985 36760 12990 36816
rect 13046 36760 15578 36816
rect 12985 36758 15578 36760
rect 15702 36816 17743 36818
rect 15702 36760 17682 36816
rect 17738 36760 17743 36816
rect 15702 36758 17743 36760
rect 12985 36755 13051 36758
rect 15518 36682 15578 36758
rect 17677 36755 17743 36758
rect 19609 36818 19675 36821
rect 29200 36818 30000 36848
rect 19609 36816 30000 36818
rect 19609 36760 19614 36816
rect 19670 36760 30000 36816
rect 19609 36758 30000 36760
rect 19609 36755 19675 36758
rect 29200 36728 30000 36758
rect 19609 36682 19675 36685
rect 15518 36680 19675 36682
rect 15518 36624 19614 36680
rect 19670 36624 19675 36680
rect 15518 36622 19675 36624
rect 19609 36619 19675 36622
rect 15009 36546 15075 36549
rect 19977 36546 20043 36549
rect 15009 36544 20043 36546
rect 15009 36488 15014 36544
rect 15070 36488 19982 36544
rect 20038 36488 20043 36544
rect 15009 36486 20043 36488
rect 15009 36483 15075 36486
rect 19977 36483 20043 36486
rect 10944 36480 11264 36481
rect 10944 36416 10952 36480
rect 11016 36416 11032 36480
rect 11096 36416 11112 36480
rect 11176 36416 11192 36480
rect 11256 36416 11264 36480
rect 10944 36415 11264 36416
rect 20944 36480 21264 36481
rect 20944 36416 20952 36480
rect 21016 36416 21032 36480
rect 21096 36416 21112 36480
rect 21176 36416 21192 36480
rect 21256 36416 21264 36480
rect 20944 36415 21264 36416
rect 4613 36410 4679 36413
rect 8569 36410 8635 36413
rect 4613 36408 8635 36410
rect 4613 36352 4618 36408
rect 4674 36352 8574 36408
rect 8630 36352 8635 36408
rect 4613 36350 8635 36352
rect 4613 36347 4679 36350
rect 8569 36347 8635 36350
rect 13353 36410 13419 36413
rect 15653 36410 15719 36413
rect 13353 36408 15719 36410
rect 13353 36352 13358 36408
rect 13414 36352 15658 36408
rect 15714 36352 15719 36408
rect 13353 36350 15719 36352
rect 13353 36347 13419 36350
rect 15653 36347 15719 36350
rect 16113 36410 16179 36413
rect 16614 36410 16620 36412
rect 16113 36408 16620 36410
rect 16113 36352 16118 36408
rect 16174 36352 16620 36408
rect 16113 36350 16620 36352
rect 16113 36347 16179 36350
rect 16614 36348 16620 36350
rect 16684 36348 16690 36412
rect 21817 36410 21883 36413
rect 21950 36410 21956 36412
rect 21817 36408 21956 36410
rect 21817 36352 21822 36408
rect 21878 36352 21956 36408
rect 21817 36350 21956 36352
rect 21817 36347 21883 36350
rect 21950 36348 21956 36350
rect 22020 36348 22026 36412
rect 8845 36274 8911 36277
rect 13813 36274 13879 36277
rect 8845 36272 13879 36274
rect 8845 36216 8850 36272
rect 8906 36216 13818 36272
rect 13874 36216 13879 36272
rect 8845 36214 13879 36216
rect 8845 36211 8911 36214
rect 13813 36211 13879 36214
rect 16205 36274 16271 36277
rect 17953 36274 18019 36277
rect 16205 36272 18019 36274
rect 16205 36216 16210 36272
rect 16266 36216 17958 36272
rect 18014 36216 18019 36272
rect 16205 36214 18019 36216
rect 16205 36211 16271 36214
rect 17953 36211 18019 36214
rect 5441 36138 5507 36141
rect 15561 36138 15627 36141
rect 20253 36138 20319 36141
rect 5441 36136 10978 36138
rect 5441 36080 5446 36136
rect 5502 36080 10978 36136
rect 5441 36078 10978 36080
rect 5441 36075 5507 36078
rect 9673 36004 9739 36005
rect 9622 36002 9628 36004
rect 9582 35942 9628 36002
rect 9692 36000 9739 36004
rect 9734 35944 9739 36000
rect 9622 35940 9628 35942
rect 9692 35940 9739 35944
rect 9673 35939 9739 35940
rect 5944 35936 6264 35937
rect 5944 35872 5952 35936
rect 6016 35872 6032 35936
rect 6096 35872 6112 35936
rect 6176 35872 6192 35936
rect 6256 35872 6264 35936
rect 5944 35871 6264 35872
rect 10918 35866 10978 36078
rect 15561 36136 20319 36138
rect 15561 36080 15566 36136
rect 15622 36080 20258 36136
rect 20314 36080 20319 36136
rect 15561 36078 20319 36080
rect 15561 36075 15627 36078
rect 20253 36075 20319 36078
rect 23933 36138 23999 36141
rect 27705 36138 27771 36141
rect 23933 36136 27771 36138
rect 23933 36080 23938 36136
rect 23994 36080 27710 36136
rect 27766 36080 27771 36136
rect 23933 36078 27771 36080
rect 23933 36075 23999 36078
rect 27705 36075 27771 36078
rect 11646 35940 11652 36004
rect 11716 36002 11722 36004
rect 12709 36002 12775 36005
rect 11716 36000 12775 36002
rect 11716 35944 12714 36000
rect 12770 35944 12775 36000
rect 11716 35942 12775 35944
rect 11716 35940 11722 35942
rect 12709 35939 12775 35942
rect 16757 36002 16823 36005
rect 16982 36002 16988 36004
rect 16757 36000 16988 36002
rect 16757 35944 16762 36000
rect 16818 35944 16988 36000
rect 16757 35942 16988 35944
rect 16757 35939 16823 35942
rect 16982 35940 16988 35942
rect 17052 35940 17058 36004
rect 15944 35936 16264 35937
rect 15944 35872 15952 35936
rect 16016 35872 16032 35936
rect 16096 35872 16112 35936
rect 16176 35872 16192 35936
rect 16256 35872 16264 35936
rect 15944 35871 16264 35872
rect 25944 35936 26264 35937
rect 25944 35872 25952 35936
rect 26016 35872 26032 35936
rect 26096 35872 26112 35936
rect 26176 35872 26192 35936
rect 26256 35872 26264 35936
rect 25944 35871 26264 35872
rect 11421 35866 11487 35869
rect 10918 35864 11487 35866
rect 10918 35808 11426 35864
rect 11482 35808 11487 35864
rect 10918 35806 11487 35808
rect 11421 35803 11487 35806
rect 12157 35868 12223 35869
rect 12157 35864 12204 35868
rect 12268 35866 12274 35868
rect 16389 35866 16455 35869
rect 18137 35866 18203 35869
rect 12157 35808 12162 35864
rect 12157 35804 12204 35808
rect 12268 35806 12314 35866
rect 16389 35864 18203 35866
rect 16389 35808 16394 35864
rect 16450 35808 18142 35864
rect 18198 35808 18203 35864
rect 16389 35806 18203 35808
rect 12268 35804 12274 35806
rect 12157 35803 12223 35804
rect 16389 35803 16455 35806
rect 18137 35803 18203 35806
rect 21541 35868 21607 35869
rect 21541 35864 21588 35868
rect 21652 35866 21658 35868
rect 21541 35808 21546 35864
rect 21541 35804 21588 35808
rect 21652 35806 21698 35866
rect 21652 35804 21658 35806
rect 21541 35803 21607 35804
rect 2865 35730 2931 35733
rect 3734 35730 3740 35732
rect 2865 35728 3740 35730
rect 2865 35672 2870 35728
rect 2926 35672 3740 35728
rect 2865 35670 3740 35672
rect 2865 35667 2931 35670
rect 3734 35668 3740 35670
rect 3804 35668 3810 35732
rect 9121 35730 9187 35733
rect 9254 35730 9260 35732
rect 9121 35728 9260 35730
rect 9121 35672 9126 35728
rect 9182 35672 9260 35728
rect 9121 35670 9260 35672
rect 9121 35667 9187 35670
rect 9254 35668 9260 35670
rect 9324 35668 9330 35732
rect 15929 35730 15995 35733
rect 18229 35730 18295 35733
rect 15929 35728 18295 35730
rect 15929 35672 15934 35728
rect 15990 35672 18234 35728
rect 18290 35672 18295 35728
rect 15929 35670 18295 35672
rect 15929 35667 15995 35670
rect 18229 35667 18295 35670
rect 19149 35730 19215 35733
rect 20621 35730 20687 35733
rect 19149 35728 20687 35730
rect 19149 35672 19154 35728
rect 19210 35672 20626 35728
rect 20682 35672 20687 35728
rect 19149 35670 20687 35672
rect 19149 35667 19215 35670
rect 20621 35667 20687 35670
rect 21173 35730 21239 35733
rect 27705 35730 27771 35733
rect 21173 35728 27771 35730
rect 21173 35672 21178 35728
rect 21234 35672 27710 35728
rect 27766 35672 27771 35728
rect 21173 35670 27771 35672
rect 21173 35667 21239 35670
rect 27705 35667 27771 35670
rect 6177 35594 6243 35597
rect 12433 35594 12499 35597
rect 15101 35594 15167 35597
rect 15469 35594 15535 35597
rect 6177 35592 15535 35594
rect 6177 35536 6182 35592
rect 6238 35536 12438 35592
rect 12494 35536 15106 35592
rect 15162 35536 15474 35592
rect 15530 35536 15535 35592
rect 6177 35534 15535 35536
rect 6177 35531 6243 35534
rect 12433 35531 12499 35534
rect 15101 35531 15167 35534
rect 15469 35531 15535 35534
rect 16021 35594 16087 35597
rect 19425 35594 19491 35597
rect 16021 35592 19491 35594
rect 16021 35536 16026 35592
rect 16082 35536 19430 35592
rect 19486 35536 19491 35592
rect 16021 35534 19491 35536
rect 16021 35531 16087 35534
rect 19425 35531 19491 35534
rect 22553 35594 22619 35597
rect 22553 35592 25376 35594
rect 22553 35536 22558 35592
rect 22614 35536 25376 35592
rect 22553 35534 25376 35536
rect 22553 35531 22619 35534
rect 0 35458 800 35488
rect 1577 35458 1643 35461
rect 0 35456 1643 35458
rect 0 35400 1582 35456
rect 1638 35400 1643 35456
rect 0 35398 1643 35400
rect 0 35368 800 35398
rect 1577 35395 1643 35398
rect 7741 35458 7807 35461
rect 9489 35458 9555 35461
rect 7741 35456 9555 35458
rect 7741 35400 7746 35456
rect 7802 35400 9494 35456
rect 9550 35400 9555 35456
rect 7741 35398 9555 35400
rect 7741 35395 7807 35398
rect 9489 35395 9555 35398
rect 9949 35458 10015 35461
rect 10726 35458 10732 35460
rect 9949 35456 10732 35458
rect 9949 35400 9954 35456
rect 10010 35400 10732 35456
rect 9949 35398 10732 35400
rect 9949 35395 10015 35398
rect 10726 35396 10732 35398
rect 10796 35396 10802 35460
rect 13813 35458 13879 35461
rect 14038 35458 14044 35460
rect 13813 35456 14044 35458
rect 13813 35400 13818 35456
rect 13874 35400 14044 35456
rect 13813 35398 14044 35400
rect 13813 35395 13879 35398
rect 14038 35396 14044 35398
rect 14108 35396 14114 35460
rect 16614 35396 16620 35460
rect 16684 35458 16690 35460
rect 19333 35458 19399 35461
rect 16684 35456 19399 35458
rect 16684 35400 19338 35456
rect 19394 35400 19399 35456
rect 16684 35398 19399 35400
rect 16684 35396 16690 35398
rect 19333 35395 19399 35398
rect 22829 35458 22895 35461
rect 25129 35458 25195 35461
rect 22829 35456 25195 35458
rect 22829 35400 22834 35456
rect 22890 35400 25134 35456
rect 25190 35400 25195 35456
rect 22829 35398 25195 35400
rect 25316 35458 25376 35534
rect 29200 35458 30000 35488
rect 25316 35398 30000 35458
rect 22829 35395 22895 35398
rect 25129 35395 25195 35398
rect 10944 35392 11264 35393
rect 10944 35328 10952 35392
rect 11016 35328 11032 35392
rect 11096 35328 11112 35392
rect 11176 35328 11192 35392
rect 11256 35328 11264 35392
rect 10944 35327 11264 35328
rect 20944 35392 21264 35393
rect 20944 35328 20952 35392
rect 21016 35328 21032 35392
rect 21096 35328 21112 35392
rect 21176 35328 21192 35392
rect 21256 35328 21264 35392
rect 29200 35368 30000 35398
rect 20944 35327 21264 35328
rect 4613 35322 4679 35325
rect 7414 35322 7420 35324
rect 4613 35320 7420 35322
rect 4613 35264 4618 35320
rect 4674 35264 7420 35320
rect 4613 35262 7420 35264
rect 4613 35259 4679 35262
rect 7414 35260 7420 35262
rect 7484 35322 7490 35324
rect 10317 35322 10383 35325
rect 7484 35320 10383 35322
rect 7484 35264 10322 35320
rect 10378 35264 10383 35320
rect 7484 35262 10383 35264
rect 7484 35260 7490 35262
rect 10317 35259 10383 35262
rect 13721 35322 13787 35325
rect 17585 35322 17651 35325
rect 13721 35320 17651 35322
rect 13721 35264 13726 35320
rect 13782 35264 17590 35320
rect 17646 35264 17651 35320
rect 13721 35262 17651 35264
rect 13721 35259 13787 35262
rect 17585 35259 17651 35262
rect 6637 35186 6703 35189
rect 12525 35186 12591 35189
rect 6637 35184 12591 35186
rect 6637 35128 6642 35184
rect 6698 35128 12530 35184
rect 12586 35128 12591 35184
rect 6637 35126 12591 35128
rect 6637 35123 6703 35126
rect 12525 35123 12591 35126
rect 12985 35186 13051 35189
rect 13302 35186 13308 35188
rect 12985 35184 13308 35186
rect 12985 35128 12990 35184
rect 13046 35128 13308 35184
rect 12985 35126 13308 35128
rect 12985 35123 13051 35126
rect 13302 35124 13308 35126
rect 13372 35124 13378 35188
rect 13629 35186 13695 35189
rect 14549 35186 14615 35189
rect 16849 35186 16915 35189
rect 13629 35184 13738 35186
rect 13629 35128 13634 35184
rect 13690 35128 13738 35184
rect 13629 35123 13738 35128
rect 14549 35184 16915 35186
rect 14549 35128 14554 35184
rect 14610 35128 16854 35184
rect 16910 35128 16915 35184
rect 14549 35126 16915 35128
rect 14549 35123 14615 35126
rect 16849 35123 16915 35126
rect 17769 35186 17835 35189
rect 20897 35186 20963 35189
rect 17769 35184 20963 35186
rect 17769 35128 17774 35184
rect 17830 35128 20902 35184
rect 20958 35128 20963 35184
rect 17769 35126 20963 35128
rect 17769 35123 17835 35126
rect 20897 35123 20963 35126
rect 22001 35186 22067 35189
rect 24301 35186 24367 35189
rect 22001 35184 24367 35186
rect 22001 35128 22006 35184
rect 22062 35128 24306 35184
rect 24362 35128 24367 35184
rect 22001 35126 24367 35128
rect 22001 35123 22067 35126
rect 24301 35123 24367 35126
rect 5993 35050 6059 35053
rect 7833 35050 7899 35053
rect 5993 35048 7899 35050
rect 5993 34992 5998 35048
rect 6054 34992 7838 35048
rect 7894 34992 7899 35048
rect 5993 34990 7899 34992
rect 5993 34987 6059 34990
rect 7833 34987 7899 34990
rect 8937 35050 9003 35053
rect 10593 35050 10659 35053
rect 8937 35048 10659 35050
rect 8937 34992 8942 35048
rect 8998 34992 10598 35048
rect 10654 34992 10659 35048
rect 8937 34990 10659 34992
rect 8937 34987 9003 34990
rect 10593 34987 10659 34990
rect 12801 35050 12867 35053
rect 13678 35050 13738 35123
rect 19425 35050 19491 35053
rect 12801 35048 19491 35050
rect 12801 34992 12806 35048
rect 12862 34992 19430 35048
rect 19486 34992 19491 35048
rect 12801 34990 19491 34992
rect 12801 34987 12867 34990
rect 19425 34987 19491 34990
rect 25446 34988 25452 35052
rect 25516 35050 25522 35052
rect 25516 34990 26434 35050
rect 25516 34988 25522 34990
rect 6913 34914 6979 34917
rect 9121 34916 9187 34917
rect 9070 34914 9076 34916
rect 6913 34912 9076 34914
rect 9140 34914 9187 34916
rect 10685 34914 10751 34917
rect 9140 34912 9268 34914
rect 6913 34856 6918 34912
rect 6974 34856 9076 34912
rect 9182 34856 9268 34912
rect 6913 34854 9076 34856
rect 6913 34851 6979 34854
rect 9070 34852 9076 34854
rect 9140 34854 9268 34856
rect 9492 34912 10751 34914
rect 9492 34856 10690 34912
rect 10746 34856 10751 34912
rect 9492 34854 10751 34856
rect 9140 34852 9187 34854
rect 9121 34851 9187 34852
rect 5944 34848 6264 34849
rect 5944 34784 5952 34848
rect 6016 34784 6032 34848
rect 6096 34784 6112 34848
rect 6176 34784 6192 34848
rect 6256 34784 6264 34848
rect 5944 34783 6264 34784
rect 7925 34778 7991 34781
rect 8477 34778 8543 34781
rect 7925 34776 8543 34778
rect 7925 34720 7930 34776
rect 7986 34720 8482 34776
rect 8538 34720 8543 34776
rect 7925 34718 8543 34720
rect 7925 34715 7991 34718
rect 8477 34715 8543 34718
rect 8937 34778 9003 34781
rect 9492 34778 9552 34854
rect 10685 34851 10751 34854
rect 12065 34914 12131 34917
rect 14549 34914 14615 34917
rect 12065 34912 14615 34914
rect 12065 34856 12070 34912
rect 12126 34856 14554 34912
rect 14610 34856 14615 34912
rect 12065 34854 14615 34856
rect 12065 34851 12131 34854
rect 14549 34851 14615 34854
rect 15944 34848 16264 34849
rect 15944 34784 15952 34848
rect 16016 34784 16032 34848
rect 16096 34784 16112 34848
rect 16176 34784 16192 34848
rect 16256 34784 16264 34848
rect 15944 34783 16264 34784
rect 25944 34848 26264 34849
rect 25944 34784 25952 34848
rect 26016 34784 26032 34848
rect 26096 34784 26112 34848
rect 26176 34784 26192 34848
rect 26256 34784 26264 34848
rect 25944 34783 26264 34784
rect 8937 34776 9552 34778
rect 8937 34720 8942 34776
rect 8998 34720 9552 34776
rect 8937 34718 9552 34720
rect 9673 34778 9739 34781
rect 9806 34778 9812 34780
rect 9673 34776 9812 34778
rect 9673 34720 9678 34776
rect 9734 34720 9812 34776
rect 9673 34718 9812 34720
rect 8937 34715 9003 34718
rect 9673 34715 9739 34718
rect 9806 34716 9812 34718
rect 9876 34716 9882 34780
rect 10542 34716 10548 34780
rect 10612 34778 10618 34780
rect 13813 34778 13879 34781
rect 10612 34776 13879 34778
rect 10612 34720 13818 34776
rect 13874 34720 13879 34776
rect 10612 34718 13879 34720
rect 10612 34716 10618 34718
rect 13813 34715 13879 34718
rect 17953 34778 18019 34781
rect 19057 34778 19123 34781
rect 22461 34778 22527 34781
rect 17953 34776 22527 34778
rect 17953 34720 17958 34776
rect 18014 34720 19062 34776
rect 19118 34720 22466 34776
rect 22522 34720 22527 34776
rect 17953 34718 22527 34720
rect 17953 34715 18019 34718
rect 19057 34715 19123 34718
rect 22188 34645 22248 34718
rect 22461 34715 22527 34718
rect 24301 34778 24367 34781
rect 26374 34778 26434 34990
rect 29200 34778 30000 34808
rect 24301 34776 25376 34778
rect 24301 34720 24306 34776
rect 24362 34720 25376 34776
rect 24301 34718 25376 34720
rect 26374 34718 30000 34778
rect 24301 34715 24367 34718
rect 25316 34645 25376 34718
rect 29200 34688 30000 34718
rect 3877 34642 3943 34645
rect 5901 34642 5967 34645
rect 10501 34642 10567 34645
rect 3877 34640 10567 34642
rect 3877 34584 3882 34640
rect 3938 34584 5906 34640
rect 5962 34584 10506 34640
rect 10562 34584 10567 34640
rect 3877 34582 10567 34584
rect 3877 34579 3943 34582
rect 5901 34579 5967 34582
rect 10501 34579 10567 34582
rect 13261 34642 13327 34645
rect 19057 34642 19123 34645
rect 13261 34640 19123 34642
rect 13261 34584 13266 34640
rect 13322 34584 19062 34640
rect 19118 34584 19123 34640
rect 13261 34582 19123 34584
rect 13261 34579 13327 34582
rect 19057 34579 19123 34582
rect 22185 34640 22251 34645
rect 22185 34584 22190 34640
rect 22246 34584 22251 34640
rect 22185 34579 22251 34584
rect 25313 34640 25379 34645
rect 25313 34584 25318 34640
rect 25374 34584 25379 34640
rect 25313 34579 25379 34584
rect 4337 34506 4403 34509
rect 8661 34506 8727 34509
rect 12893 34506 12959 34509
rect 13629 34506 13695 34509
rect 4337 34504 8727 34506
rect 4337 34448 4342 34504
rect 4398 34448 8666 34504
rect 8722 34448 8727 34504
rect 4337 34446 8727 34448
rect 4337 34443 4403 34446
rect 8661 34443 8727 34446
rect 8894 34504 13695 34506
rect 8894 34448 12898 34504
rect 12954 34448 13634 34504
rect 13690 34448 13695 34504
rect 8894 34446 13695 34448
rect 7097 34370 7163 34373
rect 8894 34370 8954 34446
rect 12893 34443 12959 34446
rect 13629 34443 13695 34446
rect 14590 34444 14596 34508
rect 14660 34506 14666 34508
rect 14733 34506 14799 34509
rect 14660 34504 14799 34506
rect 14660 34448 14738 34504
rect 14794 34448 14799 34504
rect 14660 34446 14799 34448
rect 14660 34444 14666 34446
rect 14733 34443 14799 34446
rect 17217 34506 17283 34509
rect 19885 34506 19951 34509
rect 17217 34504 19951 34506
rect 17217 34448 17222 34504
rect 17278 34448 19890 34504
rect 19946 34448 19951 34504
rect 17217 34446 19951 34448
rect 17217 34443 17283 34446
rect 19885 34443 19951 34446
rect 7097 34368 8954 34370
rect 7097 34312 7102 34368
rect 7158 34312 8954 34368
rect 7097 34310 8954 34312
rect 7097 34307 7163 34310
rect 9438 34308 9444 34372
rect 9508 34370 9514 34372
rect 9581 34370 9647 34373
rect 9508 34368 9647 34370
rect 9508 34312 9586 34368
rect 9642 34312 9647 34368
rect 9508 34310 9647 34312
rect 9508 34308 9514 34310
rect 9581 34307 9647 34310
rect 10133 34370 10199 34373
rect 10358 34370 10364 34372
rect 10133 34368 10364 34370
rect 10133 34312 10138 34368
rect 10194 34312 10364 34368
rect 10133 34310 10364 34312
rect 10133 34307 10199 34310
rect 10358 34308 10364 34310
rect 10428 34308 10434 34372
rect 11973 34370 12039 34373
rect 12566 34370 12572 34372
rect 11973 34368 12572 34370
rect 11973 34312 11978 34368
rect 12034 34312 12572 34368
rect 11973 34310 12572 34312
rect 11973 34307 12039 34310
rect 12566 34308 12572 34310
rect 12636 34370 12642 34372
rect 13077 34370 13143 34373
rect 18781 34370 18847 34373
rect 12636 34368 18847 34370
rect 12636 34312 13082 34368
rect 13138 34312 18786 34368
rect 18842 34312 18847 34368
rect 12636 34310 18847 34312
rect 12636 34308 12642 34310
rect 13077 34307 13143 34310
rect 18781 34307 18847 34310
rect 10944 34304 11264 34305
rect 10944 34240 10952 34304
rect 11016 34240 11032 34304
rect 11096 34240 11112 34304
rect 11176 34240 11192 34304
rect 11256 34240 11264 34304
rect 10944 34239 11264 34240
rect 20944 34304 21264 34305
rect 20944 34240 20952 34304
rect 21016 34240 21032 34304
rect 21096 34240 21112 34304
rect 21176 34240 21192 34304
rect 21256 34240 21264 34304
rect 20944 34239 21264 34240
rect 5349 34234 5415 34237
rect 10501 34234 10567 34237
rect 5349 34232 10567 34234
rect 5349 34176 5354 34232
rect 5410 34176 10506 34232
rect 10562 34176 10567 34232
rect 5349 34174 10567 34176
rect 5349 34171 5415 34174
rect 10501 34171 10567 34174
rect 11697 34234 11763 34237
rect 15009 34234 15075 34237
rect 11697 34232 15075 34234
rect 11697 34176 11702 34232
rect 11758 34176 15014 34232
rect 15070 34176 15075 34232
rect 11697 34174 15075 34176
rect 11697 34171 11763 34174
rect 15009 34171 15075 34174
rect 21633 34234 21699 34237
rect 23565 34234 23631 34237
rect 21633 34232 23631 34234
rect 21633 34176 21638 34232
rect 21694 34176 23570 34232
rect 23626 34176 23631 34232
rect 21633 34174 23631 34176
rect 21633 34171 21699 34174
rect 23565 34171 23631 34174
rect 0 34098 800 34128
rect 2773 34098 2839 34101
rect 0 34096 2839 34098
rect 0 34040 2778 34096
rect 2834 34040 2839 34096
rect 0 34038 2839 34040
rect 0 34008 800 34038
rect 2773 34035 2839 34038
rect 4337 34098 4403 34101
rect 6453 34098 6519 34101
rect 4337 34096 6519 34098
rect 4337 34040 4342 34096
rect 4398 34040 6458 34096
rect 6514 34040 6519 34096
rect 4337 34038 6519 34040
rect 4337 34035 4403 34038
rect 6453 34035 6519 34038
rect 7649 34098 7715 34101
rect 13077 34098 13143 34101
rect 13997 34098 14063 34101
rect 14222 34098 14228 34100
rect 7649 34096 13143 34098
rect 7649 34040 7654 34096
rect 7710 34040 13082 34096
rect 13138 34040 13143 34096
rect 7649 34038 13143 34040
rect 7649 34035 7715 34038
rect 13077 34035 13143 34038
rect 13310 34096 14228 34098
rect 13310 34040 14002 34096
rect 14058 34040 14228 34096
rect 13310 34038 14228 34040
rect 6177 33962 6243 33965
rect 6678 33962 6684 33964
rect 6177 33960 6684 33962
rect 6177 33904 6182 33960
rect 6238 33904 6684 33960
rect 6177 33902 6684 33904
rect 6177 33899 6243 33902
rect 6678 33900 6684 33902
rect 6748 33900 6754 33964
rect 6821 33962 6887 33965
rect 9806 33962 9812 33964
rect 6821 33960 9812 33962
rect 6821 33904 6826 33960
rect 6882 33904 9812 33960
rect 6821 33902 9812 33904
rect 6821 33899 6887 33902
rect 9806 33900 9812 33902
rect 9876 33962 9882 33964
rect 11697 33962 11763 33965
rect 12198 33962 12204 33964
rect 9876 33960 11763 33962
rect 9876 33904 11702 33960
rect 11758 33904 11763 33960
rect 9876 33902 11763 33904
rect 9876 33900 9882 33902
rect 11697 33899 11763 33902
rect 11838 33902 12204 33962
rect 11838 33829 11898 33902
rect 12198 33900 12204 33902
rect 12268 33900 12274 33964
rect 12893 33962 12959 33965
rect 13310 33962 13370 34038
rect 13997 34035 14063 34038
rect 14222 34036 14228 34038
rect 14292 34036 14298 34100
rect 14825 34098 14891 34101
rect 20805 34098 20871 34101
rect 14825 34096 20871 34098
rect 14825 34040 14830 34096
rect 14886 34040 20810 34096
rect 20866 34040 20871 34096
rect 14825 34038 20871 34040
rect 14825 34035 14891 34038
rect 20805 34035 20871 34038
rect 23381 34098 23447 34101
rect 25037 34098 25103 34101
rect 23381 34096 25103 34098
rect 23381 34040 23386 34096
rect 23442 34040 25042 34096
rect 25098 34040 25103 34096
rect 23381 34038 25103 34040
rect 23381 34035 23447 34038
rect 25037 34035 25103 34038
rect 12893 33960 13370 33962
rect 12893 33904 12898 33960
rect 12954 33904 13370 33960
rect 12893 33902 13370 33904
rect 14549 33962 14615 33965
rect 16757 33962 16823 33965
rect 14549 33960 16823 33962
rect 14549 33904 14554 33960
rect 14610 33904 16762 33960
rect 16818 33904 16823 33960
rect 14549 33902 16823 33904
rect 12893 33899 12959 33902
rect 14549 33899 14615 33902
rect 16757 33899 16823 33902
rect 6453 33826 6519 33829
rect 11646 33826 11652 33828
rect 6453 33824 11652 33826
rect 6453 33768 6458 33824
rect 6514 33768 11652 33824
rect 6453 33766 11652 33768
rect 6453 33763 6519 33766
rect 11646 33764 11652 33766
rect 11716 33764 11722 33828
rect 11789 33824 11898 33829
rect 11789 33768 11794 33824
rect 11850 33768 11898 33824
rect 11789 33766 11898 33768
rect 16481 33826 16547 33829
rect 16614 33826 16620 33828
rect 16481 33824 16620 33826
rect 16481 33768 16486 33824
rect 16542 33768 16620 33824
rect 16481 33766 16620 33768
rect 11789 33763 11855 33766
rect 16481 33763 16547 33766
rect 16614 33764 16620 33766
rect 16684 33764 16690 33828
rect 18781 33826 18847 33829
rect 22369 33826 22435 33829
rect 18781 33824 22435 33826
rect 18781 33768 18786 33824
rect 18842 33768 22374 33824
rect 22430 33768 22435 33824
rect 18781 33766 22435 33768
rect 18781 33763 18847 33766
rect 22369 33763 22435 33766
rect 5944 33760 6264 33761
rect 5944 33696 5952 33760
rect 6016 33696 6032 33760
rect 6096 33696 6112 33760
rect 6176 33696 6192 33760
rect 6256 33696 6264 33760
rect 5944 33695 6264 33696
rect 15944 33760 16264 33761
rect 15944 33696 15952 33760
rect 16016 33696 16032 33760
rect 16096 33696 16112 33760
rect 16176 33696 16192 33760
rect 16256 33696 16264 33760
rect 15944 33695 16264 33696
rect 25944 33760 26264 33761
rect 25944 33696 25952 33760
rect 26016 33696 26032 33760
rect 26096 33696 26112 33760
rect 26176 33696 26192 33760
rect 26256 33696 26264 33760
rect 25944 33695 26264 33696
rect 6637 33690 6703 33693
rect 12065 33690 12131 33693
rect 6637 33688 12131 33690
rect 6637 33632 6642 33688
rect 6698 33632 12070 33688
rect 12126 33632 12131 33688
rect 6637 33630 12131 33632
rect 6637 33627 6703 33630
rect 12065 33627 12131 33630
rect 18873 33690 18939 33693
rect 21817 33690 21883 33693
rect 18873 33688 21883 33690
rect 18873 33632 18878 33688
rect 18934 33632 21822 33688
rect 21878 33632 21883 33688
rect 18873 33630 21883 33632
rect 18873 33627 18939 33630
rect 21817 33627 21883 33630
rect 5349 33554 5415 33557
rect 7097 33554 7163 33557
rect 5349 33552 7163 33554
rect 5349 33496 5354 33552
rect 5410 33496 7102 33552
rect 7158 33496 7163 33552
rect 5349 33494 7163 33496
rect 5349 33491 5415 33494
rect 7097 33491 7163 33494
rect 15101 33554 15167 33557
rect 22553 33554 22619 33557
rect 15101 33552 22619 33554
rect 15101 33496 15106 33552
rect 15162 33496 22558 33552
rect 22614 33496 22619 33552
rect 15101 33494 22619 33496
rect 15101 33491 15167 33494
rect 22553 33491 22619 33494
rect 0 33418 800 33448
rect 2865 33418 2931 33421
rect 0 33416 2931 33418
rect 0 33360 2870 33416
rect 2926 33360 2931 33416
rect 0 33358 2931 33360
rect 0 33328 800 33358
rect 2865 33355 2931 33358
rect 3877 33418 3943 33421
rect 8201 33418 8267 33421
rect 3877 33416 8267 33418
rect 3877 33360 3882 33416
rect 3938 33360 8206 33416
rect 8262 33360 8267 33416
rect 3877 33358 8267 33360
rect 3877 33355 3943 33358
rect 8201 33355 8267 33358
rect 11646 33356 11652 33420
rect 11716 33418 11722 33420
rect 14549 33418 14615 33421
rect 11716 33416 14615 33418
rect 11716 33360 14554 33416
rect 14610 33360 14615 33416
rect 11716 33358 14615 33360
rect 11716 33356 11722 33358
rect 14549 33355 14615 33358
rect 15142 33356 15148 33420
rect 15212 33418 15218 33420
rect 15469 33418 15535 33421
rect 15212 33416 15535 33418
rect 15212 33360 15474 33416
rect 15530 33360 15535 33416
rect 15212 33358 15535 33360
rect 15212 33356 15218 33358
rect 15469 33355 15535 33358
rect 16205 33418 16271 33421
rect 21633 33418 21699 33421
rect 16205 33416 21699 33418
rect 16205 33360 16210 33416
rect 16266 33360 21638 33416
rect 21694 33360 21699 33416
rect 16205 33358 21699 33360
rect 16205 33355 16271 33358
rect 21633 33355 21699 33358
rect 25589 33418 25655 33421
rect 29200 33418 30000 33448
rect 25589 33416 30000 33418
rect 25589 33360 25594 33416
rect 25650 33360 30000 33416
rect 25589 33358 30000 33360
rect 25589 33355 25655 33358
rect 29200 33328 30000 33358
rect 6545 33282 6611 33285
rect 10777 33282 10843 33285
rect 6545 33280 10843 33282
rect 6545 33224 6550 33280
rect 6606 33224 10782 33280
rect 10838 33224 10843 33280
rect 6545 33222 10843 33224
rect 6545 33219 6611 33222
rect 10777 33219 10843 33222
rect 12198 33220 12204 33284
rect 12268 33282 12274 33284
rect 12341 33282 12407 33285
rect 12268 33280 12407 33282
rect 12268 33224 12346 33280
rect 12402 33224 12407 33280
rect 12268 33222 12407 33224
rect 12268 33220 12274 33222
rect 12341 33219 12407 33222
rect 12525 33282 12591 33285
rect 13077 33282 13143 33285
rect 12525 33280 13143 33282
rect 12525 33224 12530 33280
rect 12586 33224 13082 33280
rect 13138 33224 13143 33280
rect 12525 33222 13143 33224
rect 12525 33219 12591 33222
rect 13077 33219 13143 33222
rect 14181 33282 14247 33285
rect 14590 33282 14596 33284
rect 14181 33280 14596 33282
rect 14181 33224 14186 33280
rect 14242 33224 14596 33280
rect 14181 33222 14596 33224
rect 14181 33219 14247 33222
rect 14590 33220 14596 33222
rect 14660 33220 14666 33284
rect 15285 33282 15351 33285
rect 16021 33282 16087 33285
rect 19425 33282 19491 33285
rect 15285 33280 19491 33282
rect 15285 33224 15290 33280
rect 15346 33224 16026 33280
rect 16082 33224 19430 33280
rect 19486 33224 19491 33280
rect 15285 33222 19491 33224
rect 10944 33216 11264 33217
rect 10944 33152 10952 33216
rect 11016 33152 11032 33216
rect 11096 33152 11112 33216
rect 11176 33152 11192 33216
rect 11256 33152 11264 33216
rect 10944 33151 11264 33152
rect 4613 33146 4679 33149
rect 6913 33146 6979 33149
rect 4613 33144 6979 33146
rect 4613 33088 4618 33144
rect 4674 33088 6918 33144
rect 6974 33088 6979 33144
rect 4613 33086 6979 33088
rect 4613 33083 4679 33086
rect 6913 33083 6979 33086
rect 7741 33146 7807 33149
rect 12709 33146 12775 33149
rect 12934 33146 12940 33148
rect 7741 33144 10840 33146
rect 7741 33088 7746 33144
rect 7802 33088 10840 33144
rect 7741 33086 10840 33088
rect 7741 33083 7807 33086
rect 5574 32948 5580 33012
rect 5644 33010 5650 33012
rect 5717 33010 5783 33013
rect 5644 33008 5783 33010
rect 5644 32952 5722 33008
rect 5778 32952 5783 33008
rect 5644 32950 5783 32952
rect 5644 32948 5650 32950
rect 5717 32947 5783 32950
rect 5901 33010 5967 33013
rect 9121 33010 9187 33013
rect 5901 33008 9187 33010
rect 5901 32952 5906 33008
rect 5962 32952 9126 33008
rect 9182 32952 9187 33008
rect 5901 32950 9187 32952
rect 5901 32947 5967 32950
rect 9121 32947 9187 32950
rect 9581 33010 9647 33013
rect 10317 33010 10383 33013
rect 9581 33008 10383 33010
rect 9581 32952 9586 33008
rect 9642 32952 10322 33008
rect 10378 32952 10383 33008
rect 9581 32950 10383 32952
rect 10780 33010 10840 33086
rect 12709 33144 12940 33146
rect 12709 33088 12714 33144
rect 12770 33088 12940 33144
rect 12709 33086 12940 33088
rect 12709 33083 12775 33086
rect 12934 33084 12940 33086
rect 13004 33084 13010 33148
rect 14598 33146 14658 33220
rect 15285 33219 15351 33222
rect 16021 33219 16087 33222
rect 19425 33219 19491 33222
rect 19701 33282 19767 33285
rect 20437 33282 20503 33285
rect 19701 33280 20503 33282
rect 19701 33224 19706 33280
rect 19762 33224 20442 33280
rect 20498 33224 20503 33280
rect 19701 33222 20503 33224
rect 19701 33219 19767 33222
rect 20437 33219 20503 33222
rect 21817 33282 21883 33285
rect 23749 33282 23815 33285
rect 27797 33282 27863 33285
rect 21817 33280 27863 33282
rect 21817 33224 21822 33280
rect 21878 33224 23754 33280
rect 23810 33224 27802 33280
rect 27858 33224 27863 33280
rect 21817 33222 27863 33224
rect 21817 33219 21883 33222
rect 23749 33219 23815 33222
rect 27797 33219 27863 33222
rect 20944 33216 21264 33217
rect 20944 33152 20952 33216
rect 21016 33152 21032 33216
rect 21096 33152 21112 33216
rect 21176 33152 21192 33216
rect 21256 33152 21264 33216
rect 20944 33151 21264 33152
rect 20437 33146 20503 33149
rect 14598 33144 20503 33146
rect 14598 33088 20442 33144
rect 20498 33088 20503 33144
rect 14598 33086 20503 33088
rect 20437 33083 20503 33086
rect 11462 33010 11468 33012
rect 10780 32950 11468 33010
rect 9581 32947 9647 32950
rect 10317 32947 10383 32950
rect 11462 32948 11468 32950
rect 11532 33010 11538 33012
rect 12198 33010 12204 33012
rect 11532 32950 12204 33010
rect 11532 32948 11538 32950
rect 12198 32948 12204 32950
rect 12268 32948 12274 33012
rect 14365 33010 14431 33013
rect 15561 33010 15627 33013
rect 14365 33008 15627 33010
rect 14365 32952 14370 33008
rect 14426 32952 15566 33008
rect 15622 32952 15627 33008
rect 14365 32950 15627 32952
rect 14365 32947 14431 32950
rect 15561 32947 15627 32950
rect 15929 33010 15995 33013
rect 22737 33010 22803 33013
rect 15929 33008 22803 33010
rect 15929 32952 15934 33008
rect 15990 32952 22742 33008
rect 22798 32952 22803 33008
rect 15929 32950 22803 32952
rect 15929 32947 15995 32950
rect 22737 32947 22803 32950
rect 4889 32874 4955 32877
rect 13537 32874 13603 32877
rect 4889 32872 13603 32874
rect 4889 32816 4894 32872
rect 4950 32816 13542 32872
rect 13598 32816 13603 32872
rect 4889 32814 13603 32816
rect 4889 32811 4955 32814
rect 13537 32811 13603 32814
rect 13905 32874 13971 32877
rect 14733 32874 14799 32877
rect 22277 32874 22343 32877
rect 13905 32872 14799 32874
rect 13905 32816 13910 32872
rect 13966 32816 14738 32872
rect 14794 32816 14799 32872
rect 13905 32814 14799 32816
rect 13905 32811 13971 32814
rect 14733 32811 14799 32814
rect 14920 32872 22343 32874
rect 14920 32816 22282 32872
rect 22338 32816 22343 32872
rect 14920 32814 22343 32816
rect 9254 32676 9260 32740
rect 9324 32738 9330 32740
rect 13905 32738 13971 32741
rect 14774 32738 14780 32740
rect 9324 32678 13784 32738
rect 9324 32676 9330 32678
rect 5944 32672 6264 32673
rect 5944 32608 5952 32672
rect 6016 32608 6032 32672
rect 6096 32608 6112 32672
rect 6176 32608 6192 32672
rect 6256 32608 6264 32672
rect 5944 32607 6264 32608
rect 7649 32602 7715 32605
rect 10777 32602 10843 32605
rect 7649 32600 10843 32602
rect 7649 32544 7654 32600
rect 7710 32544 10782 32600
rect 10838 32544 10843 32600
rect 7649 32542 10843 32544
rect 13724 32602 13784 32678
rect 13905 32736 14780 32738
rect 13905 32680 13910 32736
rect 13966 32680 14780 32736
rect 13905 32678 14780 32680
rect 13905 32675 13971 32678
rect 14774 32676 14780 32678
rect 14844 32676 14850 32740
rect 14920 32602 14980 32814
rect 22277 32811 22343 32814
rect 17769 32738 17835 32741
rect 19977 32738 20043 32741
rect 17769 32736 20043 32738
rect 17769 32680 17774 32736
rect 17830 32680 19982 32736
rect 20038 32680 20043 32736
rect 17769 32678 20043 32680
rect 17769 32675 17835 32678
rect 19977 32675 20043 32678
rect 20253 32738 20319 32741
rect 21725 32738 21791 32741
rect 20253 32736 21791 32738
rect 20253 32680 20258 32736
rect 20314 32680 21730 32736
rect 21786 32680 21791 32736
rect 20253 32678 21791 32680
rect 20253 32675 20319 32678
rect 21725 32675 21791 32678
rect 15944 32672 16264 32673
rect 15944 32608 15952 32672
rect 16016 32608 16032 32672
rect 16096 32608 16112 32672
rect 16176 32608 16192 32672
rect 16256 32608 16264 32672
rect 15944 32607 16264 32608
rect 25944 32672 26264 32673
rect 25944 32608 25952 32672
rect 26016 32608 26032 32672
rect 26096 32608 26112 32672
rect 26176 32608 26192 32672
rect 26256 32608 26264 32672
rect 25944 32607 26264 32608
rect 13724 32542 14980 32602
rect 7649 32539 7715 32542
rect 10777 32539 10843 32542
rect 3877 32466 3943 32469
rect 6545 32466 6611 32469
rect 3877 32464 6611 32466
rect 3877 32408 3882 32464
rect 3938 32408 6550 32464
rect 6606 32408 6611 32464
rect 3877 32406 6611 32408
rect 3877 32403 3943 32406
rect 6545 32403 6611 32406
rect 8293 32466 8359 32469
rect 11237 32466 11303 32469
rect 8293 32464 11303 32466
rect 8293 32408 8298 32464
rect 8354 32408 11242 32464
rect 11298 32408 11303 32464
rect 8293 32406 11303 32408
rect 8293 32403 8359 32406
rect 11237 32403 11303 32406
rect 11973 32466 12039 32469
rect 15561 32466 15627 32469
rect 20253 32466 20319 32469
rect 11973 32464 20319 32466
rect 11973 32408 11978 32464
rect 12034 32408 15566 32464
rect 15622 32408 20258 32464
rect 20314 32408 20319 32464
rect 11973 32406 20319 32408
rect 11973 32403 12039 32406
rect 15561 32403 15627 32406
rect 20253 32403 20319 32406
rect 21766 32404 21772 32468
rect 21836 32466 21842 32468
rect 22001 32466 22067 32469
rect 21836 32464 22067 32466
rect 21836 32408 22006 32464
rect 22062 32408 22067 32464
rect 21836 32406 22067 32408
rect 21836 32404 21842 32406
rect 22001 32403 22067 32406
rect 5625 32330 5691 32333
rect 13077 32330 13143 32333
rect 16982 32330 16988 32332
rect 5625 32328 13143 32330
rect 5625 32272 5630 32328
rect 5686 32272 13082 32328
rect 13138 32272 13143 32328
rect 5625 32270 13143 32272
rect 5625 32267 5691 32270
rect 13077 32267 13143 32270
rect 14598 32270 16988 32330
rect 5901 32194 5967 32197
rect 9029 32194 9095 32197
rect 10358 32194 10364 32196
rect 5901 32192 10364 32194
rect 5901 32136 5906 32192
rect 5962 32136 9034 32192
rect 9090 32136 10364 32192
rect 5901 32134 10364 32136
rect 5901 32131 5967 32134
rect 9029 32131 9095 32134
rect 10358 32132 10364 32134
rect 10428 32132 10434 32196
rect 14598 32194 14658 32270
rect 16982 32268 16988 32270
rect 17052 32268 17058 32332
rect 12160 32134 14658 32194
rect 14733 32194 14799 32197
rect 16665 32194 16731 32197
rect 14733 32192 16731 32194
rect 14733 32136 14738 32192
rect 14794 32136 16670 32192
rect 16726 32136 16731 32192
rect 14733 32134 16731 32136
rect 10944 32128 11264 32129
rect 0 32058 800 32088
rect 10944 32064 10952 32128
rect 11016 32064 11032 32128
rect 11096 32064 11112 32128
rect 11176 32064 11192 32128
rect 11256 32064 11264 32128
rect 10944 32063 11264 32064
rect 12160 32061 12220 32134
rect 14733 32131 14799 32134
rect 16665 32131 16731 32134
rect 20944 32128 21264 32129
rect 20944 32064 20952 32128
rect 21016 32064 21032 32128
rect 21096 32064 21112 32128
rect 21176 32064 21192 32128
rect 21256 32064 21264 32128
rect 20944 32063 21264 32064
rect 3366 32058 3372 32060
rect 0 31998 3372 32058
rect 0 31968 800 31998
rect 3366 31996 3372 31998
rect 3436 31996 3442 32060
rect 5257 32058 5323 32061
rect 8845 32058 8911 32061
rect 5257 32056 8911 32058
rect 5257 32000 5262 32056
rect 5318 32000 8850 32056
rect 8906 32000 8911 32056
rect 5257 31998 8911 32000
rect 5257 31995 5323 31998
rect 8845 31995 8911 31998
rect 9070 31996 9076 32060
rect 9140 32058 9146 32060
rect 9305 32058 9371 32061
rect 9140 32056 9371 32058
rect 9140 32000 9310 32056
rect 9366 32000 9371 32056
rect 9140 31998 9371 32000
rect 9140 31996 9146 31998
rect 9305 31995 9371 31998
rect 10041 32058 10107 32061
rect 10542 32058 10548 32060
rect 10041 32056 10548 32058
rect 10041 32000 10046 32056
rect 10102 32000 10548 32056
rect 10041 31998 10548 32000
rect 10041 31995 10107 31998
rect 10542 31996 10548 31998
rect 10612 31996 10618 32060
rect 11462 31996 11468 32060
rect 11532 32058 11538 32060
rect 12157 32058 12223 32061
rect 11532 32056 12223 32058
rect 11532 32000 12162 32056
rect 12218 32000 12223 32056
rect 11532 31998 12223 32000
rect 11532 31996 11538 31998
rect 12157 31995 12223 31998
rect 13261 32058 13327 32061
rect 16757 32058 16823 32061
rect 13261 32056 16823 32058
rect 13261 32000 13266 32056
rect 13322 32000 16762 32056
rect 16818 32000 16823 32056
rect 13261 31998 16823 32000
rect 13261 31995 13327 31998
rect 16757 31995 16823 31998
rect 24945 32058 25011 32061
rect 29200 32058 30000 32088
rect 24945 32056 30000 32058
rect 24945 32000 24950 32056
rect 25006 32000 30000 32056
rect 24945 31998 30000 32000
rect 24945 31995 25011 31998
rect 29200 31968 30000 31998
rect 5717 31922 5783 31925
rect 10501 31922 10567 31925
rect 5717 31920 10567 31922
rect 5717 31864 5722 31920
rect 5778 31864 10506 31920
rect 10562 31864 10567 31920
rect 5717 31862 10567 31864
rect 5717 31859 5783 31862
rect 10501 31859 10567 31862
rect 11145 31922 11211 31925
rect 11973 31922 12039 31925
rect 11145 31920 12039 31922
rect 11145 31864 11150 31920
rect 11206 31864 11978 31920
rect 12034 31864 12039 31920
rect 11145 31862 12039 31864
rect 11145 31859 11211 31862
rect 11973 31859 12039 31862
rect 12249 31920 12315 31925
rect 12249 31864 12254 31920
rect 12310 31864 12315 31920
rect 12249 31859 12315 31864
rect 12750 31860 12756 31924
rect 12820 31922 12826 31924
rect 13302 31922 13308 31924
rect 12820 31862 13308 31922
rect 12820 31860 12826 31862
rect 13302 31860 13308 31862
rect 13372 31860 13378 31924
rect 13629 31922 13695 31925
rect 13854 31922 13860 31924
rect 13629 31920 13860 31922
rect 13629 31864 13634 31920
rect 13690 31864 13860 31920
rect 13629 31862 13860 31864
rect 13629 31859 13695 31862
rect 13854 31860 13860 31862
rect 13924 31860 13930 31924
rect 15561 31922 15627 31925
rect 20662 31922 20668 31924
rect 14184 31920 20668 31922
rect 14184 31864 15566 31920
rect 15622 31864 20668 31920
rect 14184 31862 20668 31864
rect 6637 31786 6703 31789
rect 8569 31786 8635 31789
rect 6637 31784 8635 31786
rect 6637 31728 6642 31784
rect 6698 31728 8574 31784
rect 8630 31728 8635 31784
rect 6637 31726 8635 31728
rect 6637 31723 6703 31726
rect 8569 31723 8635 31726
rect 8845 31786 8911 31789
rect 12252 31786 12312 31859
rect 12801 31788 12867 31789
rect 8845 31784 12312 31786
rect 8845 31728 8850 31784
rect 8906 31728 12312 31784
rect 8845 31726 12312 31728
rect 8845 31723 8911 31726
rect 12750 31724 12756 31788
rect 12820 31786 12867 31788
rect 13537 31786 13603 31789
rect 14038 31786 14044 31788
rect 12820 31784 12912 31786
rect 12862 31728 12912 31784
rect 12820 31726 12912 31728
rect 13537 31784 14044 31786
rect 13537 31728 13542 31784
rect 13598 31728 14044 31784
rect 13537 31726 14044 31728
rect 12820 31724 12867 31726
rect 12801 31723 12867 31724
rect 13537 31723 13603 31726
rect 14038 31724 14044 31726
rect 14108 31724 14114 31788
rect 6361 31650 6427 31653
rect 8937 31650 9003 31653
rect 9489 31652 9555 31653
rect 6361 31648 9003 31650
rect 6361 31592 6366 31648
rect 6422 31592 8942 31648
rect 8998 31592 9003 31648
rect 6361 31590 9003 31592
rect 6361 31587 6427 31590
rect 8937 31587 9003 31590
rect 9438 31588 9444 31652
rect 9508 31650 9555 31652
rect 9508 31648 9600 31650
rect 9550 31592 9600 31648
rect 9508 31590 9600 31592
rect 9508 31588 9555 31590
rect 10726 31588 10732 31652
rect 10796 31650 10802 31652
rect 11513 31650 11579 31653
rect 11697 31652 11763 31653
rect 10796 31648 11579 31650
rect 10796 31592 11518 31648
rect 11574 31592 11579 31648
rect 10796 31590 11579 31592
rect 10796 31588 10802 31590
rect 9489 31587 9555 31588
rect 11513 31587 11579 31590
rect 11646 31588 11652 31652
rect 11716 31650 11763 31652
rect 11716 31648 11808 31650
rect 11758 31592 11808 31648
rect 11716 31590 11808 31592
rect 11716 31588 11763 31590
rect 12566 31588 12572 31652
rect 12636 31650 12642 31652
rect 13077 31650 13143 31653
rect 12636 31648 13143 31650
rect 12636 31592 13082 31648
rect 13138 31592 13143 31648
rect 12636 31590 13143 31592
rect 12636 31588 12642 31590
rect 11697 31587 11763 31588
rect 13077 31587 13143 31590
rect 14038 31588 14044 31652
rect 14108 31650 14114 31652
rect 14184 31650 14244 31862
rect 15561 31859 15627 31862
rect 20662 31860 20668 31862
rect 20732 31860 20738 31924
rect 14406 31724 14412 31788
rect 14476 31786 14482 31788
rect 15377 31786 15443 31789
rect 14476 31784 15443 31786
rect 14476 31728 15382 31784
rect 15438 31728 15443 31784
rect 14476 31726 15443 31728
rect 14476 31724 14482 31726
rect 15377 31723 15443 31726
rect 17217 31786 17283 31789
rect 17677 31786 17743 31789
rect 17217 31784 17743 31786
rect 17217 31728 17222 31784
rect 17278 31728 17682 31784
rect 17738 31728 17743 31784
rect 17217 31726 17743 31728
rect 17217 31723 17283 31726
rect 17677 31723 17743 31726
rect 15745 31650 15811 31653
rect 14108 31590 14244 31650
rect 15518 31648 15811 31650
rect 15518 31592 15750 31648
rect 15806 31592 15811 31648
rect 15518 31590 15811 31592
rect 14108 31588 14114 31590
rect 5944 31584 6264 31585
rect 5944 31520 5952 31584
rect 6016 31520 6032 31584
rect 6096 31520 6112 31584
rect 6176 31520 6192 31584
rect 6256 31520 6264 31584
rect 5944 31519 6264 31520
rect 15518 31517 15578 31590
rect 15745 31587 15811 31590
rect 17493 31650 17559 31653
rect 20069 31650 20135 31653
rect 17493 31648 20135 31650
rect 17493 31592 17498 31648
rect 17554 31592 20074 31648
rect 20130 31592 20135 31648
rect 17493 31590 20135 31592
rect 17493 31587 17559 31590
rect 20069 31587 20135 31590
rect 15944 31584 16264 31585
rect 15944 31520 15952 31584
rect 16016 31520 16032 31584
rect 16096 31520 16112 31584
rect 16176 31520 16192 31584
rect 16256 31520 16264 31584
rect 15944 31519 16264 31520
rect 25944 31584 26264 31585
rect 25944 31520 25952 31584
rect 26016 31520 26032 31584
rect 26096 31520 26112 31584
rect 26176 31520 26192 31584
rect 26256 31520 26264 31584
rect 25944 31519 26264 31520
rect 6637 31514 6703 31517
rect 10225 31514 10291 31517
rect 6637 31512 10291 31514
rect 6637 31456 6642 31512
rect 6698 31456 10230 31512
rect 10286 31456 10291 31512
rect 6637 31454 10291 31456
rect 6637 31451 6703 31454
rect 10225 31451 10291 31454
rect 11421 31514 11487 31517
rect 11646 31514 11652 31516
rect 11421 31512 11652 31514
rect 11421 31456 11426 31512
rect 11482 31456 11652 31512
rect 11421 31454 11652 31456
rect 11421 31451 11487 31454
rect 11646 31452 11652 31454
rect 11716 31452 11722 31516
rect 15469 31512 15578 31517
rect 15469 31456 15474 31512
rect 15530 31456 15578 31512
rect 15469 31454 15578 31456
rect 16389 31514 16455 31517
rect 20529 31514 20595 31517
rect 16389 31512 20595 31514
rect 16389 31456 16394 31512
rect 16450 31456 20534 31512
rect 20590 31456 20595 31512
rect 16389 31454 20595 31456
rect 15469 31451 15535 31454
rect 16389 31451 16455 31454
rect 20529 31451 20595 31454
rect 5533 31378 5599 31381
rect 11462 31378 11468 31380
rect 5533 31376 11468 31378
rect 5533 31320 5538 31376
rect 5594 31320 11468 31376
rect 5533 31318 11468 31320
rect 5533 31315 5599 31318
rect 11462 31316 11468 31318
rect 11532 31316 11538 31380
rect 12801 31378 12867 31381
rect 13854 31378 13860 31380
rect 12801 31376 13860 31378
rect 12801 31320 12806 31376
rect 12862 31320 13860 31376
rect 12801 31318 13860 31320
rect 12801 31315 12867 31318
rect 13854 31316 13860 31318
rect 13924 31316 13930 31380
rect 14222 31316 14228 31380
rect 14292 31378 14298 31380
rect 15653 31378 15719 31381
rect 14292 31376 15719 31378
rect 14292 31320 15658 31376
rect 15714 31320 15719 31376
rect 14292 31318 15719 31320
rect 14292 31316 14298 31318
rect 15653 31315 15719 31318
rect 18781 31378 18847 31381
rect 20897 31378 20963 31381
rect 18781 31376 20963 31378
rect 18781 31320 18786 31376
rect 18842 31320 20902 31376
rect 20958 31320 20963 31376
rect 18781 31318 20963 31320
rect 18781 31315 18847 31318
rect 20897 31315 20963 31318
rect 23933 31378 23999 31381
rect 25078 31378 25084 31380
rect 23933 31376 25084 31378
rect 23933 31320 23938 31376
rect 23994 31320 25084 31376
rect 23933 31318 25084 31320
rect 23933 31315 23999 31318
rect 25078 31316 25084 31318
rect 25148 31316 25154 31380
rect 3969 31242 4035 31245
rect 8201 31242 8267 31245
rect 9581 31242 9647 31245
rect 10501 31242 10567 31245
rect 3969 31240 8908 31242
rect 3969 31184 3974 31240
rect 4030 31184 8206 31240
rect 8262 31184 8908 31240
rect 3969 31182 8908 31184
rect 3969 31179 4035 31182
rect 8201 31179 8267 31182
rect 8848 31109 8908 31182
rect 9581 31240 10567 31242
rect 9581 31184 9586 31240
rect 9642 31184 10506 31240
rect 10562 31184 10567 31240
rect 9581 31182 10567 31184
rect 9581 31179 9647 31182
rect 10501 31179 10567 31182
rect 11237 31242 11303 31245
rect 12525 31242 12591 31245
rect 16573 31242 16639 31245
rect 11237 31240 11668 31242
rect 11237 31184 11242 31240
rect 11298 31184 11668 31240
rect 11237 31182 11668 31184
rect 11237 31179 11303 31182
rect 11608 31109 11668 31182
rect 12525 31240 16639 31242
rect 12525 31184 12530 31240
rect 12586 31184 16578 31240
rect 16634 31184 16639 31240
rect 12525 31182 16639 31184
rect 12525 31179 12591 31182
rect 16573 31179 16639 31182
rect 18965 31242 19031 31245
rect 21173 31242 21239 31245
rect 18965 31240 21239 31242
rect 18965 31184 18970 31240
rect 19026 31184 21178 31240
rect 21234 31184 21239 31240
rect 18965 31182 21239 31184
rect 18965 31179 19031 31182
rect 21173 31179 21239 31182
rect 22921 31242 22987 31245
rect 27613 31242 27679 31245
rect 22921 31240 27679 31242
rect 22921 31184 22926 31240
rect 22982 31184 27618 31240
rect 27674 31184 27679 31240
rect 22921 31182 27679 31184
rect 22921 31179 22987 31182
rect 27613 31179 27679 31182
rect 8845 31104 8911 31109
rect 8845 31048 8850 31104
rect 8906 31048 8911 31104
rect 8845 31043 8911 31048
rect 9949 31106 10015 31109
rect 9949 31104 10058 31106
rect 9949 31048 9954 31104
rect 10010 31048 10058 31104
rect 9949 31043 10058 31048
rect 11605 31104 11671 31109
rect 11605 31048 11610 31104
rect 11666 31048 11671 31104
rect 11605 31043 11671 31048
rect 12249 31106 12315 31109
rect 14273 31106 14339 31109
rect 14958 31106 14964 31108
rect 12249 31104 13738 31106
rect 12249 31048 12254 31104
rect 12310 31048 13738 31104
rect 12249 31046 13738 31048
rect 12249 31043 12315 31046
rect 9998 30837 10058 31043
rect 10944 31040 11264 31041
rect 10944 30976 10952 31040
rect 11016 30976 11032 31040
rect 11096 30976 11112 31040
rect 11176 30976 11192 31040
rect 11256 30976 11264 31040
rect 10944 30975 11264 30976
rect 13678 30970 13738 31046
rect 14273 31104 14964 31106
rect 14273 31048 14278 31104
rect 14334 31048 14964 31104
rect 14273 31046 14964 31048
rect 14273 31043 14339 31046
rect 14958 31044 14964 31046
rect 15028 31044 15034 31108
rect 15285 31106 15351 31109
rect 19977 31106 20043 31109
rect 15285 31104 20043 31106
rect 15285 31048 15290 31104
rect 15346 31048 19982 31104
rect 20038 31048 20043 31104
rect 15285 31046 20043 31048
rect 15285 31043 15351 31046
rect 19977 31043 20043 31046
rect 20478 31044 20484 31108
rect 20548 31106 20554 31108
rect 20805 31106 20871 31109
rect 20548 31104 20871 31106
rect 20548 31048 20810 31104
rect 20866 31048 20871 31104
rect 20548 31046 20871 31048
rect 20548 31044 20554 31046
rect 20805 31043 20871 31046
rect 20944 31040 21264 31041
rect 20944 30976 20952 31040
rect 21016 30976 21032 31040
rect 21096 30976 21112 31040
rect 21176 30976 21192 31040
rect 21256 30976 21264 31040
rect 20944 30975 21264 30976
rect 13905 30970 13971 30973
rect 14774 30970 14780 30972
rect 13678 30968 14780 30970
rect 13678 30912 13910 30968
rect 13966 30912 14780 30968
rect 13678 30910 14780 30912
rect 13905 30907 13971 30910
rect 14774 30908 14780 30910
rect 14844 30908 14850 30972
rect 15101 30970 15167 30973
rect 16389 30970 16455 30973
rect 15101 30968 16455 30970
rect 15101 30912 15106 30968
rect 15162 30912 16394 30968
rect 16450 30912 16455 30968
rect 15101 30910 16455 30912
rect 15101 30907 15167 30910
rect 16389 30907 16455 30910
rect 9949 30832 10058 30837
rect 9949 30776 9954 30832
rect 10010 30776 10058 30832
rect 9949 30774 10058 30776
rect 10317 30834 10383 30837
rect 10961 30834 11027 30837
rect 10317 30832 11027 30834
rect 10317 30776 10322 30832
rect 10378 30776 10966 30832
rect 11022 30776 11027 30832
rect 10317 30774 11027 30776
rect 9949 30771 10015 30774
rect 10317 30771 10383 30774
rect 10961 30771 11027 30774
rect 13169 30834 13235 30837
rect 16757 30834 16823 30837
rect 13169 30832 16823 30834
rect 13169 30776 13174 30832
rect 13230 30776 16762 30832
rect 16818 30776 16823 30832
rect 13169 30774 16823 30776
rect 13169 30771 13235 30774
rect 16757 30771 16823 30774
rect 20662 30772 20668 30836
rect 20732 30834 20738 30836
rect 20897 30834 20963 30837
rect 20732 30832 20963 30834
rect 20732 30776 20902 30832
rect 20958 30776 20963 30832
rect 20732 30774 20963 30776
rect 20732 30772 20738 30774
rect 20897 30771 20963 30774
rect 0 30698 800 30728
rect 3601 30698 3667 30701
rect 0 30696 3667 30698
rect 0 30640 3606 30696
rect 3662 30640 3667 30696
rect 0 30638 3667 30640
rect 0 30608 800 30638
rect 3601 30635 3667 30638
rect 5257 30698 5323 30701
rect 11513 30698 11579 30701
rect 13353 30700 13419 30701
rect 13302 30698 13308 30700
rect 5257 30696 11579 30698
rect 5257 30640 5262 30696
rect 5318 30640 11518 30696
rect 11574 30640 11579 30696
rect 5257 30638 11579 30640
rect 13262 30638 13308 30698
rect 13372 30696 13419 30700
rect 13414 30640 13419 30696
rect 5257 30635 5323 30638
rect 11513 30635 11579 30638
rect 13302 30636 13308 30638
rect 13372 30636 13419 30640
rect 13353 30635 13419 30636
rect 13813 30698 13879 30701
rect 16665 30698 16731 30701
rect 21081 30698 21147 30701
rect 13813 30696 16731 30698
rect 13813 30640 13818 30696
rect 13874 30640 16670 30696
rect 16726 30640 16731 30696
rect 13813 30638 16731 30640
rect 13813 30635 13879 30638
rect 16665 30635 16731 30638
rect 16806 30696 21147 30698
rect 16806 30640 21086 30696
rect 21142 30640 21147 30696
rect 16806 30638 21147 30640
rect 3233 30562 3299 30565
rect 5625 30562 5691 30565
rect 3233 30560 5691 30562
rect 3233 30504 3238 30560
rect 3294 30504 5630 30560
rect 5686 30504 5691 30560
rect 3233 30502 5691 30504
rect 3233 30499 3299 30502
rect 5625 30499 5691 30502
rect 8661 30562 8727 30565
rect 12893 30562 12959 30565
rect 8661 30560 12959 30562
rect 8661 30504 8666 30560
rect 8722 30504 12898 30560
rect 12954 30504 12959 30560
rect 8661 30502 12959 30504
rect 8661 30499 8727 30502
rect 12893 30499 12959 30502
rect 13077 30562 13143 30565
rect 15009 30562 15075 30565
rect 16665 30564 16731 30565
rect 16614 30562 16620 30564
rect 13077 30560 15075 30562
rect 13077 30504 13082 30560
rect 13138 30504 15014 30560
rect 15070 30504 15075 30560
rect 13077 30502 15075 30504
rect 16574 30502 16620 30562
rect 16684 30560 16731 30564
rect 16726 30504 16731 30560
rect 13077 30499 13143 30502
rect 15009 30499 15075 30502
rect 16614 30500 16620 30502
rect 16684 30500 16731 30504
rect 16665 30499 16731 30500
rect 5944 30496 6264 30497
rect 5944 30432 5952 30496
rect 6016 30432 6032 30496
rect 6096 30432 6112 30496
rect 6176 30432 6192 30496
rect 6256 30432 6264 30496
rect 5944 30431 6264 30432
rect 15944 30496 16264 30497
rect 15944 30432 15952 30496
rect 16016 30432 16032 30496
rect 16096 30432 16112 30496
rect 16176 30432 16192 30496
rect 16256 30432 16264 30496
rect 15944 30431 16264 30432
rect 6913 30426 6979 30429
rect 12750 30426 12756 30428
rect 6913 30424 12756 30426
rect 6913 30368 6918 30424
rect 6974 30368 12756 30424
rect 6913 30366 12756 30368
rect 6913 30363 6979 30366
rect 12750 30364 12756 30366
rect 12820 30364 12826 30428
rect 12934 30364 12940 30428
rect 13004 30364 13010 30428
rect 16806 30426 16866 30638
rect 21081 30635 21147 30638
rect 25681 30698 25747 30701
rect 29200 30698 30000 30728
rect 25681 30696 30000 30698
rect 25681 30640 25686 30696
rect 25742 30640 30000 30696
rect 25681 30638 30000 30640
rect 25681 30635 25747 30638
rect 29200 30608 30000 30638
rect 18137 30562 18203 30565
rect 16484 30366 16866 30426
rect 18094 30560 18203 30562
rect 18094 30504 18142 30560
rect 18198 30504 18203 30560
rect 18094 30499 18203 30504
rect 12942 30293 13002 30364
rect 16484 30293 16544 30366
rect 12893 30288 13002 30293
rect 12893 30232 12898 30288
rect 12954 30232 13002 30288
rect 12893 30230 13002 30232
rect 14917 30290 14983 30293
rect 16481 30290 16547 30293
rect 14917 30288 16547 30290
rect 14917 30232 14922 30288
rect 14978 30232 16486 30288
rect 16542 30232 16547 30288
rect 14917 30230 16547 30232
rect 12893 30227 12959 30230
rect 14917 30227 14983 30230
rect 16481 30227 16547 30230
rect 16798 30228 16804 30292
rect 16868 30290 16874 30292
rect 17217 30290 17283 30293
rect 16868 30288 17283 30290
rect 16868 30232 17222 30288
rect 17278 30232 17283 30288
rect 16868 30230 17283 30232
rect 16868 30228 16874 30230
rect 17217 30227 17283 30230
rect 17493 30292 17559 30293
rect 17493 30288 17540 30292
rect 17604 30290 17610 30292
rect 17493 30232 17498 30288
rect 17493 30228 17540 30232
rect 17604 30230 17650 30290
rect 17604 30228 17610 30230
rect 17493 30227 17559 30228
rect 11646 30154 11652 30156
rect 8158 30094 11652 30154
rect 0 30018 800 30048
rect 5809 30018 5875 30021
rect 0 30016 5875 30018
rect 0 29960 5814 30016
rect 5870 29960 5875 30016
rect 0 29958 5875 29960
rect 0 29928 800 29958
rect 5809 29955 5875 29958
rect 7097 30018 7163 30021
rect 8158 30018 8218 30094
rect 11646 30092 11652 30094
rect 11716 30154 11722 30156
rect 13854 30154 13860 30156
rect 11716 30094 13860 30154
rect 11716 30092 11722 30094
rect 13854 30092 13860 30094
rect 13924 30092 13930 30156
rect 15929 30154 15995 30157
rect 18094 30154 18154 30499
rect 25944 30496 26264 30497
rect 25944 30432 25952 30496
rect 26016 30432 26032 30496
rect 26096 30432 26112 30496
rect 26176 30432 26192 30496
rect 26256 30432 26264 30496
rect 25944 30431 26264 30432
rect 19241 30290 19307 30293
rect 24945 30290 25011 30293
rect 19241 30288 25011 30290
rect 19241 30232 19246 30288
rect 19302 30232 24950 30288
rect 25006 30232 25011 30288
rect 19241 30230 25011 30232
rect 19241 30227 19307 30230
rect 24945 30227 25011 30230
rect 19425 30154 19491 30157
rect 15929 30152 19491 30154
rect 15929 30096 15934 30152
rect 15990 30096 19430 30152
rect 19486 30096 19491 30152
rect 15929 30094 19491 30096
rect 15929 30091 15995 30094
rect 19425 30091 19491 30094
rect 7097 30016 8218 30018
rect 7097 29960 7102 30016
rect 7158 29960 8218 30016
rect 7097 29958 8218 29960
rect 10133 30018 10199 30021
rect 10358 30018 10364 30020
rect 10133 30016 10364 30018
rect 10133 29960 10138 30016
rect 10194 29960 10364 30016
rect 10133 29958 10364 29960
rect 7097 29955 7163 29958
rect 10133 29955 10199 29958
rect 10358 29956 10364 29958
rect 10428 29956 10434 30020
rect 12341 30018 12407 30021
rect 13302 30018 13308 30020
rect 12341 30016 13308 30018
rect 12341 29960 12346 30016
rect 12402 29960 13308 30016
rect 12341 29958 13308 29960
rect 12341 29955 12407 29958
rect 13302 29956 13308 29958
rect 13372 30018 13378 30020
rect 18689 30018 18755 30021
rect 13372 30016 18755 30018
rect 13372 29960 18694 30016
rect 18750 29960 18755 30016
rect 13372 29958 18755 29960
rect 13372 29956 13378 29958
rect 18689 29955 18755 29958
rect 22645 30018 22711 30021
rect 29200 30018 30000 30048
rect 22645 30016 30000 30018
rect 22645 29960 22650 30016
rect 22706 29960 30000 30016
rect 22645 29958 30000 29960
rect 22645 29955 22711 29958
rect 10944 29952 11264 29953
rect 10944 29888 10952 29952
rect 11016 29888 11032 29952
rect 11096 29888 11112 29952
rect 11176 29888 11192 29952
rect 11256 29888 11264 29952
rect 10944 29887 11264 29888
rect 20944 29952 21264 29953
rect 20944 29888 20952 29952
rect 21016 29888 21032 29952
rect 21096 29888 21112 29952
rect 21176 29888 21192 29952
rect 21256 29888 21264 29952
rect 29200 29928 30000 29958
rect 20944 29887 21264 29888
rect 12934 29820 12940 29884
rect 13004 29882 13010 29884
rect 16849 29882 16915 29885
rect 13004 29880 16915 29882
rect 13004 29824 16854 29880
rect 16910 29824 16915 29880
rect 13004 29822 16915 29824
rect 13004 29820 13010 29822
rect 16849 29819 16915 29822
rect 4981 29746 5047 29749
rect 8753 29746 8819 29749
rect 4981 29744 8819 29746
rect 4981 29688 4986 29744
rect 5042 29688 8758 29744
rect 8814 29688 8819 29744
rect 4981 29686 8819 29688
rect 4981 29683 5047 29686
rect 8753 29683 8819 29686
rect 10133 29746 10199 29749
rect 10542 29746 10548 29748
rect 10133 29744 10548 29746
rect 10133 29688 10138 29744
rect 10194 29688 10548 29744
rect 10133 29686 10548 29688
rect 10133 29683 10199 29686
rect 10542 29684 10548 29686
rect 10612 29684 10618 29748
rect 11513 29746 11579 29749
rect 14089 29748 14155 29749
rect 11646 29746 11652 29748
rect 11513 29744 11652 29746
rect 11513 29688 11518 29744
rect 11574 29688 11652 29744
rect 11513 29686 11652 29688
rect 11513 29683 11579 29686
rect 11646 29684 11652 29686
rect 11716 29684 11722 29748
rect 14038 29684 14044 29748
rect 14108 29746 14155 29748
rect 15101 29746 15167 29749
rect 18045 29746 18111 29749
rect 14108 29744 14200 29746
rect 14150 29688 14200 29744
rect 14108 29686 14200 29688
rect 15101 29744 18111 29746
rect 15101 29688 15106 29744
rect 15162 29688 18050 29744
rect 18106 29688 18111 29744
rect 15101 29686 18111 29688
rect 14108 29684 14155 29686
rect 14089 29683 14155 29684
rect 15101 29683 15167 29686
rect 18045 29683 18111 29686
rect 6637 29610 6703 29613
rect 12893 29610 12959 29613
rect 6637 29608 12959 29610
rect 6637 29552 6642 29608
rect 6698 29552 12898 29608
rect 12954 29552 12959 29608
rect 6637 29550 12959 29552
rect 6637 29547 6703 29550
rect 12893 29547 12959 29550
rect 14222 29548 14228 29612
rect 14292 29610 14298 29612
rect 16205 29610 16271 29613
rect 14292 29608 16271 29610
rect 14292 29552 16210 29608
rect 16266 29552 16271 29608
rect 14292 29550 16271 29552
rect 14292 29548 14298 29550
rect 16205 29547 16271 29550
rect 8201 29474 8267 29477
rect 9254 29474 9260 29476
rect 8201 29472 9260 29474
rect 8201 29416 8206 29472
rect 8262 29416 9260 29472
rect 8201 29414 9260 29416
rect 8201 29411 8267 29414
rect 9254 29412 9260 29414
rect 9324 29412 9330 29476
rect 11513 29474 11579 29477
rect 15745 29474 15811 29477
rect 19057 29474 19123 29477
rect 20989 29474 21055 29477
rect 11513 29472 15811 29474
rect 11513 29416 11518 29472
rect 11574 29416 15750 29472
rect 15806 29416 15811 29472
rect 11513 29414 15811 29416
rect 11513 29411 11579 29414
rect 15745 29411 15811 29414
rect 16438 29472 21055 29474
rect 16438 29416 19062 29472
rect 19118 29416 20994 29472
rect 21050 29416 21055 29472
rect 16438 29414 21055 29416
rect 5944 29408 6264 29409
rect 5944 29344 5952 29408
rect 6016 29344 6032 29408
rect 6096 29344 6112 29408
rect 6176 29344 6192 29408
rect 6256 29344 6264 29408
rect 5944 29343 6264 29344
rect 15944 29408 16264 29409
rect 15944 29344 15952 29408
rect 16016 29344 16032 29408
rect 16096 29344 16112 29408
rect 16176 29344 16192 29408
rect 16256 29344 16264 29408
rect 15944 29343 16264 29344
rect 6821 29338 6887 29341
rect 12750 29338 12756 29340
rect 6821 29336 12756 29338
rect 6821 29280 6826 29336
rect 6882 29280 12756 29336
rect 6821 29278 12756 29280
rect 6821 29275 6887 29278
rect 12750 29276 12756 29278
rect 12820 29338 12826 29340
rect 13118 29338 13124 29340
rect 12820 29278 13124 29338
rect 12820 29276 12826 29278
rect 13118 29276 13124 29278
rect 13188 29276 13194 29340
rect 13721 29338 13787 29341
rect 15745 29338 15811 29341
rect 13721 29336 15811 29338
rect 13721 29280 13726 29336
rect 13782 29280 15750 29336
rect 15806 29280 15811 29336
rect 13721 29278 15811 29280
rect 13721 29275 13787 29278
rect 15745 29275 15811 29278
rect 3141 29202 3207 29205
rect 6177 29202 6243 29205
rect 8293 29202 8359 29205
rect 10869 29202 10935 29205
rect 16438 29202 16498 29414
rect 19057 29411 19123 29414
rect 20989 29411 21055 29414
rect 25944 29408 26264 29409
rect 25944 29344 25952 29408
rect 26016 29344 26032 29408
rect 26096 29344 26112 29408
rect 26176 29344 26192 29408
rect 26256 29344 26264 29408
rect 25944 29343 26264 29344
rect 16573 29338 16639 29341
rect 19885 29338 19951 29341
rect 16573 29336 19951 29338
rect 16573 29280 16578 29336
rect 16634 29280 19890 29336
rect 19946 29280 19951 29336
rect 16573 29278 19951 29280
rect 16573 29275 16639 29278
rect 19885 29275 19951 29278
rect 3141 29200 16498 29202
rect 3141 29144 3146 29200
rect 3202 29144 6182 29200
rect 6238 29144 8298 29200
rect 8354 29144 10874 29200
rect 10930 29144 16498 29200
rect 3141 29142 16498 29144
rect 3141 29139 3207 29142
rect 6177 29139 6243 29142
rect 8293 29139 8359 29142
rect 10869 29139 10935 29142
rect 8109 29066 8175 29069
rect 10133 29066 10199 29069
rect 8109 29064 10199 29066
rect 8109 29008 8114 29064
rect 8170 29008 10138 29064
rect 10194 29008 10199 29064
rect 8109 29006 10199 29008
rect 8109 29003 8175 29006
rect 10133 29003 10199 29006
rect 13169 29066 13235 29069
rect 13721 29066 13787 29069
rect 13169 29064 13787 29066
rect 13169 29008 13174 29064
rect 13230 29008 13726 29064
rect 13782 29008 13787 29064
rect 13169 29006 13787 29008
rect 13169 29003 13235 29006
rect 13721 29003 13787 29006
rect 14273 29066 14339 29069
rect 16849 29066 16915 29069
rect 14273 29064 16915 29066
rect 14273 29008 14278 29064
rect 14334 29008 16854 29064
rect 16910 29008 16915 29064
rect 14273 29006 16915 29008
rect 14273 29003 14339 29006
rect 16849 29003 16915 29006
rect 7414 28868 7420 28932
rect 7484 28930 7490 28932
rect 7925 28930 7991 28933
rect 7484 28928 7991 28930
rect 7484 28872 7930 28928
rect 7986 28872 7991 28928
rect 7484 28870 7991 28872
rect 7484 28868 7490 28870
rect 7925 28867 7991 28870
rect 14733 28930 14799 28933
rect 16757 28930 16823 28933
rect 14733 28928 16823 28930
rect 14733 28872 14738 28928
rect 14794 28872 16762 28928
rect 16818 28872 16823 28928
rect 14733 28870 16823 28872
rect 14733 28867 14799 28870
rect 16757 28867 16823 28870
rect 17033 28930 17099 28933
rect 19333 28930 19399 28933
rect 17033 28928 19399 28930
rect 17033 28872 17038 28928
rect 17094 28872 19338 28928
rect 19394 28872 19399 28928
rect 17033 28870 19399 28872
rect 17033 28867 17099 28870
rect 19333 28867 19399 28870
rect 21633 28930 21699 28933
rect 25865 28930 25931 28933
rect 21633 28928 25931 28930
rect 21633 28872 21638 28928
rect 21694 28872 25870 28928
rect 25926 28872 25931 28928
rect 21633 28870 25931 28872
rect 21633 28867 21699 28870
rect 25865 28867 25931 28870
rect 10944 28864 11264 28865
rect 10944 28800 10952 28864
rect 11016 28800 11032 28864
rect 11096 28800 11112 28864
rect 11176 28800 11192 28864
rect 11256 28800 11264 28864
rect 10944 28799 11264 28800
rect 20944 28864 21264 28865
rect 20944 28800 20952 28864
rect 21016 28800 21032 28864
rect 21096 28800 21112 28864
rect 21176 28800 21192 28864
rect 21256 28800 21264 28864
rect 20944 28799 21264 28800
rect 6545 28794 6611 28797
rect 8385 28794 8451 28797
rect 10685 28794 10751 28797
rect 6545 28792 8451 28794
rect 6545 28736 6550 28792
rect 6606 28736 8390 28792
rect 8446 28736 8451 28792
rect 6545 28734 8451 28736
rect 6545 28731 6611 28734
rect 8385 28731 8451 28734
rect 8526 28792 10751 28794
rect 8526 28736 10690 28792
rect 10746 28736 10751 28792
rect 8526 28734 10751 28736
rect 0 28658 800 28688
rect 4705 28658 4771 28661
rect 0 28656 4771 28658
rect 0 28600 4710 28656
rect 4766 28600 4771 28656
rect 0 28598 4771 28600
rect 0 28568 800 28598
rect 4705 28595 4771 28598
rect 6453 28658 6519 28661
rect 8526 28658 8586 28734
rect 10685 28731 10751 28734
rect 13905 28794 13971 28797
rect 14733 28794 14799 28797
rect 16021 28794 16087 28797
rect 13905 28792 16087 28794
rect 13905 28736 13910 28792
rect 13966 28736 14738 28792
rect 14794 28736 16026 28792
rect 16082 28736 16087 28792
rect 13905 28734 16087 28736
rect 13905 28731 13971 28734
rect 14733 28731 14799 28734
rect 16021 28731 16087 28734
rect 16389 28794 16455 28797
rect 18873 28794 18939 28797
rect 16389 28792 18939 28794
rect 16389 28736 16394 28792
rect 16450 28736 18878 28792
rect 18934 28736 18939 28792
rect 16389 28734 18939 28736
rect 16389 28731 16455 28734
rect 18873 28731 18939 28734
rect 6453 28656 8586 28658
rect 6453 28600 6458 28656
rect 6514 28600 8586 28656
rect 6453 28598 8586 28600
rect 9121 28658 9187 28661
rect 13629 28658 13695 28661
rect 9121 28656 13695 28658
rect 9121 28600 9126 28656
rect 9182 28600 13634 28656
rect 13690 28600 13695 28656
rect 9121 28598 13695 28600
rect 6453 28595 6519 28598
rect 9121 28595 9187 28598
rect 13629 28595 13695 28598
rect 13854 28596 13860 28660
rect 13924 28658 13930 28660
rect 14365 28658 14431 28661
rect 13924 28656 14431 28658
rect 13924 28600 14370 28656
rect 14426 28600 14431 28656
rect 13924 28598 14431 28600
rect 13924 28596 13930 28598
rect 14365 28595 14431 28598
rect 15929 28658 15995 28661
rect 17585 28658 17651 28661
rect 20713 28658 20779 28661
rect 15929 28656 20779 28658
rect 15929 28600 15934 28656
rect 15990 28600 17590 28656
rect 17646 28600 20718 28656
rect 20774 28600 20779 28656
rect 15929 28598 20779 28600
rect 15929 28595 15995 28598
rect 17585 28595 17651 28598
rect 20713 28595 20779 28598
rect 24117 28658 24183 28661
rect 29200 28658 30000 28688
rect 24117 28656 30000 28658
rect 24117 28600 24122 28656
rect 24178 28600 30000 28656
rect 24117 28598 30000 28600
rect 24117 28595 24183 28598
rect 29200 28568 30000 28598
rect 7833 28522 7899 28525
rect 9673 28522 9739 28525
rect 7833 28520 9739 28522
rect 7833 28464 7838 28520
rect 7894 28464 9678 28520
rect 9734 28464 9739 28520
rect 7833 28462 9739 28464
rect 7833 28459 7899 28462
rect 9673 28459 9739 28462
rect 10685 28522 10751 28525
rect 12617 28522 12683 28525
rect 10685 28520 12683 28522
rect 10685 28464 10690 28520
rect 10746 28464 12622 28520
rect 12678 28464 12683 28520
rect 10685 28462 12683 28464
rect 10685 28459 10751 28462
rect 12617 28459 12683 28462
rect 13261 28522 13327 28525
rect 17217 28522 17283 28525
rect 13261 28520 17283 28522
rect 13261 28464 13266 28520
rect 13322 28464 17222 28520
rect 17278 28464 17283 28520
rect 13261 28462 17283 28464
rect 13261 28459 13327 28462
rect 17217 28459 17283 28462
rect 7925 28386 7991 28389
rect 10041 28386 10107 28389
rect 7925 28384 10107 28386
rect 7925 28328 7930 28384
rect 7986 28328 10046 28384
rect 10102 28328 10107 28384
rect 7925 28326 10107 28328
rect 7925 28323 7991 28326
rect 10041 28323 10107 28326
rect 13905 28386 13971 28389
rect 14222 28386 14228 28388
rect 13905 28384 14228 28386
rect 13905 28328 13910 28384
rect 13966 28328 14228 28384
rect 13905 28326 14228 28328
rect 13905 28323 13971 28326
rect 14222 28324 14228 28326
rect 14292 28324 14298 28388
rect 5944 28320 6264 28321
rect 5944 28256 5952 28320
rect 6016 28256 6032 28320
rect 6096 28256 6112 28320
rect 6176 28256 6192 28320
rect 6256 28256 6264 28320
rect 5944 28255 6264 28256
rect 15944 28320 16264 28321
rect 15944 28256 15952 28320
rect 16016 28256 16032 28320
rect 16096 28256 16112 28320
rect 16176 28256 16192 28320
rect 16256 28256 16264 28320
rect 15944 28255 16264 28256
rect 25944 28320 26264 28321
rect 25944 28256 25952 28320
rect 26016 28256 26032 28320
rect 26096 28256 26112 28320
rect 26176 28256 26192 28320
rect 26256 28256 26264 28320
rect 25944 28255 26264 28256
rect 8937 28250 9003 28253
rect 11513 28250 11579 28253
rect 8937 28248 11579 28250
rect 8937 28192 8942 28248
rect 8998 28192 11518 28248
rect 11574 28192 11579 28248
rect 8937 28190 11579 28192
rect 8937 28187 9003 28190
rect 11513 28187 11579 28190
rect 16665 28250 16731 28253
rect 19609 28250 19675 28253
rect 16665 28248 19675 28250
rect 16665 28192 16670 28248
rect 16726 28192 19614 28248
rect 19670 28192 19675 28248
rect 16665 28190 19675 28192
rect 16665 28187 16731 28190
rect 19609 28187 19675 28190
rect 10542 28052 10548 28116
rect 10612 28114 10618 28116
rect 10869 28114 10935 28117
rect 10612 28112 10935 28114
rect 10612 28056 10874 28112
rect 10930 28056 10935 28112
rect 10612 28054 10935 28056
rect 10612 28052 10618 28054
rect 10869 28051 10935 28054
rect 11697 28114 11763 28117
rect 13353 28114 13419 28117
rect 11697 28112 13419 28114
rect 11697 28056 11702 28112
rect 11758 28056 13358 28112
rect 13414 28056 13419 28112
rect 11697 28054 13419 28056
rect 11697 28051 11763 28054
rect 13353 28051 13419 28054
rect 15101 28112 15167 28117
rect 15101 28056 15106 28112
rect 15162 28056 15167 28112
rect 15101 28051 15167 28056
rect 15929 28114 15995 28117
rect 19425 28114 19491 28117
rect 15929 28112 19491 28114
rect 15929 28056 15934 28112
rect 15990 28056 19430 28112
rect 19486 28056 19491 28112
rect 15929 28054 19491 28056
rect 15929 28051 15995 28054
rect 19425 28051 19491 28054
rect 7097 27978 7163 27981
rect 10869 27978 10935 27981
rect 7097 27976 10935 27978
rect 7097 27920 7102 27976
rect 7158 27920 10874 27976
rect 10930 27920 10935 27976
rect 7097 27918 10935 27920
rect 15104 27978 15164 28051
rect 16757 27978 16823 27981
rect 18045 27978 18111 27981
rect 15104 27976 18111 27978
rect 15104 27920 16762 27976
rect 16818 27920 18050 27976
rect 18106 27920 18111 27976
rect 15104 27918 18111 27920
rect 7097 27915 7163 27918
rect 10869 27915 10935 27918
rect 16757 27915 16823 27918
rect 18045 27915 18111 27918
rect 9622 27780 9628 27844
rect 9692 27842 9698 27844
rect 9765 27842 9831 27845
rect 9692 27840 9831 27842
rect 9692 27784 9770 27840
rect 9826 27784 9831 27840
rect 9692 27782 9831 27784
rect 9692 27780 9698 27782
rect 9765 27779 9831 27782
rect 12249 27842 12315 27845
rect 12709 27842 12775 27845
rect 20069 27842 20135 27845
rect 12249 27840 20135 27842
rect 12249 27784 12254 27840
rect 12310 27784 12714 27840
rect 12770 27784 20074 27840
rect 20130 27784 20135 27840
rect 12249 27782 20135 27784
rect 12249 27779 12315 27782
rect 12709 27779 12775 27782
rect 20069 27779 20135 27782
rect 10944 27776 11264 27777
rect 10944 27712 10952 27776
rect 11016 27712 11032 27776
rect 11096 27712 11112 27776
rect 11176 27712 11192 27776
rect 11256 27712 11264 27776
rect 10944 27711 11264 27712
rect 20944 27776 21264 27777
rect 20944 27712 20952 27776
rect 21016 27712 21032 27776
rect 21096 27712 21112 27776
rect 21176 27712 21192 27776
rect 21256 27712 21264 27776
rect 20944 27711 21264 27712
rect 4061 27706 4127 27709
rect 6545 27706 6611 27709
rect 4061 27704 6611 27706
rect 4061 27648 4066 27704
rect 4122 27648 6550 27704
rect 6606 27648 6611 27704
rect 4061 27646 6611 27648
rect 4061 27643 4127 27646
rect 6545 27643 6611 27646
rect 8385 27706 8451 27709
rect 8385 27704 10794 27706
rect 8385 27648 8390 27704
rect 8446 27648 10794 27704
rect 8385 27646 10794 27648
rect 8385 27643 8451 27646
rect 10734 27570 10794 27646
rect 12382 27644 12388 27708
rect 12452 27706 12458 27708
rect 13997 27706 14063 27709
rect 12452 27704 14063 27706
rect 12452 27648 14002 27704
rect 14058 27648 14063 27704
rect 12452 27646 14063 27648
rect 12452 27644 12458 27646
rect 13997 27643 14063 27646
rect 16389 27706 16455 27709
rect 17585 27708 17651 27709
rect 16614 27706 16620 27708
rect 16389 27704 16620 27706
rect 16389 27648 16394 27704
rect 16450 27648 16620 27704
rect 16389 27646 16620 27648
rect 16389 27643 16455 27646
rect 16614 27644 16620 27646
rect 16684 27644 16690 27708
rect 17534 27644 17540 27708
rect 17604 27706 17651 27708
rect 25405 27706 25471 27709
rect 17604 27704 17696 27706
rect 17646 27648 17696 27704
rect 25270 27704 25471 27706
rect 17604 27646 17696 27648
rect 25129 27672 25195 27675
rect 25270 27672 25410 27704
rect 25129 27670 25410 27672
rect 17604 27644 17651 27646
rect 17585 27643 17651 27644
rect 25129 27614 25134 27670
rect 25190 27648 25410 27670
rect 25466 27648 25471 27704
rect 25190 27646 25471 27648
rect 25190 27614 25330 27646
rect 25405 27643 25471 27646
rect 25129 27612 25330 27614
rect 25129 27609 25195 27612
rect 16665 27570 16731 27573
rect 18689 27570 18755 27573
rect 20069 27570 20135 27573
rect 10734 27568 20135 27570
rect 10734 27512 16670 27568
rect 16726 27512 18694 27568
rect 18750 27512 20074 27568
rect 20130 27512 20135 27568
rect 10734 27510 20135 27512
rect 16665 27507 16731 27510
rect 18689 27507 18755 27510
rect 20069 27507 20135 27510
rect 8109 27434 8175 27437
rect 10409 27434 10475 27437
rect 8109 27432 10475 27434
rect 8109 27376 8114 27432
rect 8170 27376 10414 27432
rect 10470 27376 10475 27432
rect 8109 27374 10475 27376
rect 8109 27371 8175 27374
rect 10409 27371 10475 27374
rect 16205 27434 16271 27437
rect 16665 27434 16731 27437
rect 16205 27432 16731 27434
rect 16205 27376 16210 27432
rect 16266 27376 16670 27432
rect 16726 27376 16731 27432
rect 16205 27374 16731 27376
rect 16205 27371 16271 27374
rect 16665 27371 16731 27374
rect 0 27298 800 27328
rect 4153 27298 4219 27301
rect 0 27296 4219 27298
rect 0 27240 4158 27296
rect 4214 27240 4219 27296
rect 0 27238 4219 27240
rect 0 27208 800 27238
rect 4153 27235 4219 27238
rect 8661 27298 8727 27301
rect 12617 27298 12683 27301
rect 8661 27296 12683 27298
rect 8661 27240 8666 27296
rect 8722 27240 12622 27296
rect 12678 27240 12683 27296
rect 8661 27238 12683 27240
rect 8661 27235 8727 27238
rect 12617 27235 12683 27238
rect 15561 27296 15627 27301
rect 29200 27298 30000 27328
rect 15561 27240 15566 27296
rect 15622 27240 15627 27296
rect 15561 27235 15627 27240
rect 26374 27238 30000 27298
rect 5944 27232 6264 27233
rect 5944 27168 5952 27232
rect 6016 27168 6032 27232
rect 6096 27168 6112 27232
rect 6176 27168 6192 27232
rect 6256 27168 6264 27232
rect 5944 27167 6264 27168
rect 6361 27162 6427 27165
rect 12566 27162 12572 27164
rect 6361 27160 12572 27162
rect 6361 27104 6366 27160
rect 6422 27104 12572 27160
rect 6361 27102 12572 27104
rect 6361 27099 6427 27102
rect 12566 27100 12572 27102
rect 12636 27162 12642 27164
rect 13905 27162 13971 27165
rect 12636 27160 13971 27162
rect 12636 27104 13910 27160
rect 13966 27104 13971 27160
rect 12636 27102 13971 27104
rect 12636 27100 12642 27102
rect 13905 27099 13971 27102
rect 12198 26964 12204 27028
rect 12268 27026 12274 27028
rect 12801 27026 12867 27029
rect 12268 27024 12867 27026
rect 12268 26968 12806 27024
rect 12862 26968 12867 27024
rect 12268 26966 12867 26968
rect 15564 27026 15624 27235
rect 15944 27232 16264 27233
rect 15944 27168 15952 27232
rect 16016 27168 16032 27232
rect 16096 27168 16112 27232
rect 16176 27168 16192 27232
rect 16256 27168 16264 27232
rect 15944 27167 16264 27168
rect 25944 27232 26264 27233
rect 25944 27168 25952 27232
rect 26016 27168 26032 27232
rect 26096 27168 26112 27232
rect 26176 27168 26192 27232
rect 26256 27168 26264 27232
rect 25944 27167 26264 27168
rect 16389 27162 16455 27165
rect 18137 27162 18203 27165
rect 16389 27160 18203 27162
rect 16389 27104 16394 27160
rect 16450 27104 18142 27160
rect 18198 27104 18203 27160
rect 16389 27102 18203 27104
rect 16389 27099 16455 27102
rect 18137 27099 18203 27102
rect 18229 27026 18295 27029
rect 15564 27024 18295 27026
rect 15564 26968 18234 27024
rect 18290 26968 18295 27024
rect 15564 26966 18295 26968
rect 12268 26964 12274 26966
rect 12801 26963 12867 26966
rect 18229 26963 18295 26966
rect 18413 27026 18479 27029
rect 26374 27026 26434 27238
rect 29200 27208 30000 27238
rect 18413 27024 26434 27026
rect 18413 26968 18418 27024
rect 18474 26968 26434 27024
rect 18413 26966 26434 26968
rect 18413 26963 18479 26966
rect 9806 26828 9812 26892
rect 9876 26890 9882 26892
rect 13905 26890 13971 26893
rect 9876 26888 13971 26890
rect 9876 26832 13910 26888
rect 13966 26832 13971 26888
rect 9876 26830 13971 26832
rect 9876 26828 9882 26830
rect 13905 26827 13971 26830
rect 13169 26754 13235 26757
rect 17585 26754 17651 26757
rect 13169 26752 17651 26754
rect 13169 26696 13174 26752
rect 13230 26696 17590 26752
rect 17646 26696 17651 26752
rect 13169 26694 17651 26696
rect 13169 26691 13235 26694
rect 17585 26691 17651 26694
rect 10944 26688 11264 26689
rect 0 26618 800 26648
rect 10944 26624 10952 26688
rect 11016 26624 11032 26688
rect 11096 26624 11112 26688
rect 11176 26624 11192 26688
rect 11256 26624 11264 26688
rect 10944 26623 11264 26624
rect 20944 26688 21264 26689
rect 20944 26624 20952 26688
rect 21016 26624 21032 26688
rect 21096 26624 21112 26688
rect 21176 26624 21192 26688
rect 21256 26624 21264 26688
rect 20944 26623 21264 26624
rect 1577 26618 1643 26621
rect 0 26616 1643 26618
rect 0 26560 1582 26616
rect 1638 26560 1643 26616
rect 0 26558 1643 26560
rect 0 26528 800 26558
rect 1577 26555 1643 26558
rect 13537 26618 13603 26621
rect 18137 26618 18203 26621
rect 13537 26616 18203 26618
rect 13537 26560 13542 26616
rect 13598 26560 18142 26616
rect 18198 26560 18203 26616
rect 13537 26558 18203 26560
rect 13537 26555 13603 26558
rect 18137 26555 18203 26558
rect 25497 26618 25563 26621
rect 29200 26618 30000 26648
rect 25497 26616 30000 26618
rect 25497 26560 25502 26616
rect 25558 26560 30000 26616
rect 25497 26558 30000 26560
rect 25497 26555 25563 26558
rect 29200 26528 30000 26558
rect 7465 26346 7531 26349
rect 8753 26346 8819 26349
rect 7465 26344 8819 26346
rect 7465 26288 7470 26344
rect 7526 26288 8758 26344
rect 8814 26288 8819 26344
rect 7465 26286 8819 26288
rect 7465 26283 7531 26286
rect 8753 26283 8819 26286
rect 10726 26284 10732 26348
rect 10796 26346 10802 26348
rect 11237 26346 11303 26349
rect 11462 26346 11468 26348
rect 10796 26344 11468 26346
rect 10796 26288 11242 26344
rect 11298 26288 11468 26344
rect 10796 26286 11468 26288
rect 10796 26284 10802 26286
rect 11237 26283 11303 26286
rect 11462 26284 11468 26286
rect 11532 26284 11538 26348
rect 7189 26210 7255 26213
rect 10317 26210 10383 26213
rect 25681 26210 25747 26213
rect 7189 26208 10383 26210
rect 7189 26152 7194 26208
rect 7250 26152 10322 26208
rect 10378 26152 10383 26208
rect 7189 26150 10383 26152
rect 7189 26147 7255 26150
rect 10317 26147 10383 26150
rect 17220 26208 25747 26210
rect 17220 26152 25686 26208
rect 25742 26152 25747 26208
rect 17220 26150 25747 26152
rect 5944 26144 6264 26145
rect 5944 26080 5952 26144
rect 6016 26080 6032 26144
rect 6096 26080 6112 26144
rect 6176 26080 6192 26144
rect 6256 26080 6264 26144
rect 5944 26079 6264 26080
rect 15944 26144 16264 26145
rect 15944 26080 15952 26144
rect 16016 26080 16032 26144
rect 16096 26080 16112 26144
rect 16176 26080 16192 26144
rect 16256 26080 16264 26144
rect 15944 26079 16264 26080
rect 6545 26074 6611 26077
rect 12157 26074 12223 26077
rect 12525 26074 12591 26077
rect 6545 26072 11346 26074
rect 6545 26016 6550 26072
rect 6606 26016 11346 26072
rect 6545 26014 11346 26016
rect 6545 26011 6611 26014
rect 10174 25876 10180 25940
rect 10244 25938 10250 25940
rect 10317 25938 10383 25941
rect 11145 25938 11211 25941
rect 10244 25936 11211 25938
rect 10244 25880 10322 25936
rect 10378 25880 11150 25936
rect 11206 25880 11211 25936
rect 10244 25878 11211 25880
rect 11286 25938 11346 26014
rect 12157 26072 12591 26074
rect 12157 26016 12162 26072
rect 12218 26016 12530 26072
rect 12586 26016 12591 26072
rect 12157 26014 12591 26016
rect 12157 26011 12223 26014
rect 12525 26011 12591 26014
rect 17220 25938 17280 26150
rect 25681 26147 25747 26150
rect 25944 26144 26264 26145
rect 25944 26080 25952 26144
rect 26016 26080 26032 26144
rect 26096 26080 26112 26144
rect 26176 26080 26192 26144
rect 26256 26080 26264 26144
rect 25944 26079 26264 26080
rect 18413 26074 18479 26077
rect 25037 26074 25103 26077
rect 18413 26072 25103 26074
rect 18413 26016 18418 26072
rect 18474 26016 25042 26072
rect 25098 26016 25103 26072
rect 18413 26014 25103 26016
rect 18413 26011 18479 26014
rect 25037 26011 25103 26014
rect 11286 25878 17280 25938
rect 10244 25876 10250 25878
rect 10317 25875 10383 25878
rect 11145 25875 11211 25878
rect 9121 25802 9187 25805
rect 11237 25802 11303 25805
rect 9121 25800 11303 25802
rect 9121 25744 9126 25800
rect 9182 25744 11242 25800
rect 11298 25744 11303 25800
rect 9121 25742 11303 25744
rect 9121 25739 9187 25742
rect 11237 25739 11303 25742
rect 14733 25802 14799 25805
rect 18413 25802 18479 25805
rect 21633 25802 21699 25805
rect 14733 25800 18479 25802
rect 14733 25744 14738 25800
rect 14794 25744 18418 25800
rect 18474 25744 18479 25800
rect 14733 25742 18479 25744
rect 14733 25739 14799 25742
rect 18413 25739 18479 25742
rect 20670 25800 21699 25802
rect 20670 25744 21638 25800
rect 21694 25744 21699 25800
rect 20670 25742 21699 25744
rect 5809 25666 5875 25669
rect 10685 25668 10751 25669
rect 9622 25666 9628 25668
rect 5809 25664 9628 25666
rect 5809 25608 5814 25664
rect 5870 25608 9628 25664
rect 5809 25606 9628 25608
rect 5809 25603 5875 25606
rect 9622 25604 9628 25606
rect 9692 25666 9698 25668
rect 10542 25666 10548 25668
rect 9692 25606 10548 25666
rect 9692 25604 9698 25606
rect 10542 25604 10548 25606
rect 10612 25604 10618 25668
rect 10685 25664 10732 25668
rect 10796 25666 10802 25668
rect 16205 25666 16271 25669
rect 20670 25666 20730 25742
rect 21633 25739 21699 25742
rect 10685 25608 10690 25664
rect 10685 25604 10732 25608
rect 10796 25606 10842 25666
rect 16205 25664 20730 25666
rect 16205 25608 16210 25664
rect 16266 25608 20730 25664
rect 16205 25606 20730 25608
rect 10796 25604 10802 25606
rect 10685 25603 10751 25604
rect 16205 25603 16271 25606
rect 10944 25600 11264 25601
rect 10944 25536 10952 25600
rect 11016 25536 11032 25600
rect 11096 25536 11112 25600
rect 11176 25536 11192 25600
rect 11256 25536 11264 25600
rect 10944 25535 11264 25536
rect 20944 25600 21264 25601
rect 20944 25536 20952 25600
rect 21016 25536 21032 25600
rect 21096 25536 21112 25600
rect 21176 25536 21192 25600
rect 21256 25536 21264 25600
rect 20944 25535 21264 25536
rect 7373 25394 7439 25397
rect 12382 25394 12388 25396
rect 7373 25392 12388 25394
rect 7373 25336 7378 25392
rect 7434 25336 12388 25392
rect 7373 25334 12388 25336
rect 7373 25331 7439 25334
rect 12382 25332 12388 25334
rect 12452 25394 12458 25396
rect 14406 25394 14412 25396
rect 12452 25334 14412 25394
rect 12452 25332 12458 25334
rect 14406 25332 14412 25334
rect 14476 25332 14482 25396
rect 0 25258 800 25288
rect 2681 25258 2747 25261
rect 0 25256 2747 25258
rect 0 25200 2686 25256
rect 2742 25200 2747 25256
rect 0 25198 2747 25200
rect 0 25168 800 25198
rect 2681 25195 2747 25198
rect 7649 25258 7715 25261
rect 10041 25258 10107 25261
rect 19241 25258 19307 25261
rect 7649 25256 10107 25258
rect 7649 25200 7654 25256
rect 7710 25200 10046 25256
rect 10102 25200 10107 25256
rect 7649 25198 10107 25200
rect 7649 25195 7715 25198
rect 10041 25195 10107 25198
rect 13540 25256 19307 25258
rect 13540 25200 19246 25256
rect 19302 25200 19307 25256
rect 13540 25198 19307 25200
rect 8477 25122 8543 25125
rect 13540 25122 13600 25198
rect 19241 25195 19307 25198
rect 25865 25258 25931 25261
rect 29200 25258 30000 25288
rect 25865 25256 30000 25258
rect 25865 25200 25870 25256
rect 25926 25200 30000 25256
rect 25865 25198 30000 25200
rect 25865 25195 25931 25198
rect 29200 25168 30000 25198
rect 8477 25120 13600 25122
rect 8477 25064 8482 25120
rect 8538 25064 13600 25120
rect 8477 25062 13600 25064
rect 13721 25122 13787 25125
rect 15561 25122 15627 25125
rect 13721 25120 15627 25122
rect 13721 25064 13726 25120
rect 13782 25064 15566 25120
rect 15622 25064 15627 25120
rect 13721 25062 15627 25064
rect 8477 25059 8543 25062
rect 13721 25059 13787 25062
rect 15561 25059 15627 25062
rect 5944 25056 6264 25057
rect 5944 24992 5952 25056
rect 6016 24992 6032 25056
rect 6096 24992 6112 25056
rect 6176 24992 6192 25056
rect 6256 24992 6264 25056
rect 5944 24991 6264 24992
rect 15944 25056 16264 25057
rect 15944 24992 15952 25056
rect 16016 24992 16032 25056
rect 16096 24992 16112 25056
rect 16176 24992 16192 25056
rect 16256 24992 16264 25056
rect 15944 24991 16264 24992
rect 25944 25056 26264 25057
rect 25944 24992 25952 25056
rect 26016 24992 26032 25056
rect 26096 24992 26112 25056
rect 26176 24992 26192 25056
rect 26256 24992 26264 25056
rect 25944 24991 26264 24992
rect 13537 24986 13603 24989
rect 14917 24986 14983 24989
rect 15653 24986 15719 24989
rect 13537 24984 15719 24986
rect 13537 24928 13542 24984
rect 13598 24928 14922 24984
rect 14978 24928 15658 24984
rect 15714 24928 15719 24984
rect 13537 24926 15719 24928
rect 13537 24923 13603 24926
rect 14917 24923 14983 24926
rect 15653 24923 15719 24926
rect 19149 24850 19215 24853
rect 20253 24850 20319 24853
rect 19149 24848 20319 24850
rect 19149 24792 19154 24848
rect 19210 24792 20258 24848
rect 20314 24792 20319 24848
rect 19149 24790 20319 24792
rect 19149 24787 19215 24790
rect 20253 24787 20319 24790
rect 3233 24714 3299 24717
rect 6269 24714 6335 24717
rect 3233 24712 6335 24714
rect 3233 24656 3238 24712
rect 3294 24656 6274 24712
rect 6330 24656 6335 24712
rect 3233 24654 6335 24656
rect 3233 24651 3299 24654
rect 6269 24651 6335 24654
rect 12433 24714 12499 24717
rect 15837 24714 15903 24717
rect 12433 24712 15903 24714
rect 12433 24656 12438 24712
rect 12494 24656 15842 24712
rect 15898 24656 15903 24712
rect 12433 24654 15903 24656
rect 12433 24651 12499 24654
rect 15837 24651 15903 24654
rect 11462 24516 11468 24580
rect 11532 24578 11538 24580
rect 11789 24578 11855 24581
rect 11532 24576 11855 24578
rect 11532 24520 11794 24576
rect 11850 24520 11855 24576
rect 11532 24518 11855 24520
rect 11532 24516 11538 24518
rect 11789 24515 11855 24518
rect 10944 24512 11264 24513
rect 10944 24448 10952 24512
rect 11016 24448 11032 24512
rect 11096 24448 11112 24512
rect 11176 24448 11192 24512
rect 11256 24448 11264 24512
rect 10944 24447 11264 24448
rect 20944 24512 21264 24513
rect 20944 24448 20952 24512
rect 21016 24448 21032 24512
rect 21096 24448 21112 24512
rect 21176 24448 21192 24512
rect 21256 24448 21264 24512
rect 20944 24447 21264 24448
rect 8569 24170 8635 24173
rect 18045 24170 18111 24173
rect 8569 24168 18111 24170
rect 8569 24112 8574 24168
rect 8630 24112 18050 24168
rect 18106 24112 18111 24168
rect 8569 24110 18111 24112
rect 8569 24107 8635 24110
rect 18045 24107 18111 24110
rect 10869 24034 10935 24037
rect 12065 24034 12131 24037
rect 10869 24032 12131 24034
rect 10869 23976 10874 24032
rect 10930 23976 12070 24032
rect 12126 23976 12131 24032
rect 10869 23974 12131 23976
rect 10869 23971 10935 23974
rect 12065 23971 12131 23974
rect 5944 23968 6264 23969
rect 0 23898 800 23928
rect 5944 23904 5952 23968
rect 6016 23904 6032 23968
rect 6096 23904 6112 23968
rect 6176 23904 6192 23968
rect 6256 23904 6264 23968
rect 5944 23903 6264 23904
rect 15944 23968 16264 23969
rect 15944 23904 15952 23968
rect 16016 23904 16032 23968
rect 16096 23904 16112 23968
rect 16176 23904 16192 23968
rect 16256 23904 16264 23968
rect 15944 23903 16264 23904
rect 25944 23968 26264 23969
rect 25944 23904 25952 23968
rect 26016 23904 26032 23968
rect 26096 23904 26112 23968
rect 26176 23904 26192 23968
rect 26256 23904 26264 23968
rect 25944 23903 26264 23904
rect 1945 23898 2011 23901
rect 0 23896 2011 23898
rect 0 23840 1950 23896
rect 2006 23840 2011 23896
rect 0 23838 2011 23840
rect 0 23808 800 23838
rect 1945 23835 2011 23838
rect 26969 23898 27035 23901
rect 29200 23898 30000 23928
rect 26969 23896 30000 23898
rect 26969 23840 26974 23896
rect 27030 23840 30000 23896
rect 26969 23838 30000 23840
rect 26969 23835 27035 23838
rect 29200 23808 30000 23838
rect 6821 23762 6887 23765
rect 16481 23762 16547 23765
rect 6821 23760 16547 23762
rect 6821 23704 6826 23760
rect 6882 23704 16486 23760
rect 16542 23704 16547 23760
rect 6821 23702 16547 23704
rect 6821 23699 6887 23702
rect 16481 23699 16547 23702
rect 16665 23762 16731 23765
rect 21725 23762 21791 23765
rect 16665 23760 21791 23762
rect 16665 23704 16670 23760
rect 16726 23704 21730 23760
rect 21786 23704 21791 23760
rect 16665 23702 21791 23704
rect 16665 23699 16731 23702
rect 21725 23699 21791 23702
rect 11421 23626 11487 23629
rect 12198 23626 12204 23628
rect 11421 23624 12204 23626
rect 11421 23568 11426 23624
rect 11482 23568 12204 23624
rect 11421 23566 12204 23568
rect 11421 23563 11487 23566
rect 12198 23564 12204 23566
rect 12268 23564 12274 23628
rect 16481 23626 16547 23629
rect 16614 23626 16620 23628
rect 16481 23624 16620 23626
rect 16481 23568 16486 23624
rect 16542 23568 16620 23624
rect 16481 23566 16620 23568
rect 16481 23563 16547 23566
rect 16614 23564 16620 23566
rect 16684 23564 16690 23628
rect 18505 23626 18571 23629
rect 25630 23626 25636 23628
rect 18505 23624 25636 23626
rect 18505 23568 18510 23624
rect 18566 23568 25636 23624
rect 18505 23566 25636 23568
rect 18505 23563 18571 23566
rect 25630 23564 25636 23566
rect 25700 23564 25706 23628
rect 10944 23424 11264 23425
rect 10944 23360 10952 23424
rect 11016 23360 11032 23424
rect 11096 23360 11112 23424
rect 11176 23360 11192 23424
rect 11256 23360 11264 23424
rect 10944 23359 11264 23360
rect 20944 23424 21264 23425
rect 20944 23360 20952 23424
rect 21016 23360 21032 23424
rect 21096 23360 21112 23424
rect 21176 23360 21192 23424
rect 21256 23360 21264 23424
rect 20944 23359 21264 23360
rect 9213 23218 9279 23221
rect 11973 23218 12039 23221
rect 9213 23216 12039 23218
rect 9213 23160 9218 23216
rect 9274 23160 11978 23216
rect 12034 23160 12039 23216
rect 9213 23158 12039 23160
rect 9213 23155 9279 23158
rect 11973 23155 12039 23158
rect 13721 23218 13787 23221
rect 15285 23218 15351 23221
rect 13721 23216 15351 23218
rect 13721 23160 13726 23216
rect 13782 23160 15290 23216
rect 15346 23160 15351 23216
rect 13721 23158 15351 23160
rect 13721 23155 13787 23158
rect 15285 23155 15351 23158
rect 23841 23218 23907 23221
rect 29200 23218 30000 23248
rect 23841 23216 30000 23218
rect 23841 23160 23846 23216
rect 23902 23160 30000 23216
rect 23841 23158 30000 23160
rect 23841 23155 23907 23158
rect 29200 23128 30000 23158
rect 9765 22946 9831 22949
rect 12065 22946 12131 22949
rect 9765 22944 12131 22946
rect 9765 22888 9770 22944
rect 9826 22888 12070 22944
rect 12126 22888 12131 22944
rect 9765 22886 12131 22888
rect 9765 22883 9831 22886
rect 12065 22883 12131 22886
rect 14958 22884 14964 22948
rect 15028 22884 15034 22948
rect 5944 22880 6264 22881
rect 5944 22816 5952 22880
rect 6016 22816 6032 22880
rect 6096 22816 6112 22880
rect 6176 22816 6192 22880
rect 6256 22816 6264 22880
rect 5944 22815 6264 22816
rect 14966 22813 15026 22884
rect 15944 22880 16264 22881
rect 15944 22816 15952 22880
rect 16016 22816 16032 22880
rect 16096 22816 16112 22880
rect 16176 22816 16192 22880
rect 16256 22816 16264 22880
rect 15944 22815 16264 22816
rect 25944 22880 26264 22881
rect 25944 22816 25952 22880
rect 26016 22816 26032 22880
rect 26096 22816 26112 22880
rect 26176 22816 26192 22880
rect 26256 22816 26264 22880
rect 25944 22815 26264 22816
rect 7833 22810 7899 22813
rect 7833 22808 12036 22810
rect 7833 22752 7838 22808
rect 7894 22752 12036 22808
rect 7833 22750 12036 22752
rect 7833 22747 7899 22750
rect 11329 22674 11395 22677
rect 11462 22674 11468 22676
rect 11329 22672 11468 22674
rect 11329 22616 11334 22672
rect 11390 22616 11468 22672
rect 11329 22614 11468 22616
rect 11329 22611 11395 22614
rect 11462 22612 11468 22614
rect 11532 22612 11538 22676
rect 11976 22674 12036 22750
rect 14917 22808 15026 22813
rect 14917 22752 14922 22808
rect 14978 22752 15026 22808
rect 14917 22750 15026 22752
rect 14917 22747 14983 22750
rect 12433 22674 12499 22677
rect 11976 22672 12499 22674
rect 11976 22616 12438 22672
rect 12494 22616 12499 22672
rect 11976 22614 12499 22616
rect 12433 22611 12499 22614
rect 15142 22612 15148 22676
rect 15212 22674 15218 22676
rect 15377 22674 15443 22677
rect 15212 22672 15443 22674
rect 15212 22616 15382 22672
rect 15438 22616 15443 22672
rect 15212 22614 15443 22616
rect 15212 22612 15218 22614
rect 15377 22611 15443 22614
rect 0 22538 800 22568
rect 10593 22538 10659 22541
rect 12249 22538 12315 22541
rect 13302 22538 13308 22540
rect 0 22448 858 22538
rect 10593 22536 11714 22538
rect 10593 22480 10598 22536
rect 10654 22480 11714 22536
rect 10593 22478 11714 22480
rect 10593 22475 10659 22478
rect 798 22402 858 22448
rect 11654 22404 11714 22478
rect 12249 22536 13308 22538
rect 12249 22480 12254 22536
rect 12310 22480 13308 22536
rect 12249 22478 13308 22480
rect 12249 22475 12315 22478
rect 13302 22476 13308 22478
rect 13372 22476 13378 22540
rect 798 22342 7666 22402
rect 5533 22130 5599 22133
rect 3190 22128 5599 22130
rect 3190 22072 5538 22128
rect 5594 22072 5599 22128
rect 3190 22070 5599 22072
rect 7606 22130 7666 22342
rect 11646 22340 11652 22404
rect 11716 22402 11722 22404
rect 16573 22402 16639 22405
rect 11716 22400 16639 22402
rect 11716 22344 16578 22400
rect 16634 22344 16639 22400
rect 11716 22342 16639 22344
rect 11716 22340 11722 22342
rect 16573 22339 16639 22342
rect 10944 22336 11264 22337
rect 10944 22272 10952 22336
rect 11016 22272 11032 22336
rect 11096 22272 11112 22336
rect 11176 22272 11192 22336
rect 11256 22272 11264 22336
rect 10944 22271 11264 22272
rect 20944 22336 21264 22337
rect 20944 22272 20952 22336
rect 21016 22272 21032 22336
rect 21096 22272 21112 22336
rect 21176 22272 21192 22336
rect 21256 22272 21264 22336
rect 20944 22271 21264 22272
rect 12198 22204 12204 22268
rect 12268 22266 12274 22268
rect 12341 22266 12407 22269
rect 12268 22264 12407 22266
rect 12268 22208 12346 22264
rect 12402 22208 12407 22264
rect 12268 22206 12407 22208
rect 12268 22204 12274 22206
rect 12341 22203 12407 22206
rect 12934 22204 12940 22268
rect 13004 22266 13010 22268
rect 13353 22266 13419 22269
rect 15101 22266 15167 22269
rect 13004 22264 15167 22266
rect 13004 22208 13358 22264
rect 13414 22208 15106 22264
rect 15162 22208 15167 22264
rect 13004 22206 15167 22208
rect 13004 22204 13010 22206
rect 13353 22203 13419 22206
rect 15101 22203 15167 22206
rect 13486 22130 13492 22132
rect 7606 22070 13492 22130
rect 0 21858 800 21888
rect 3190 21858 3250 22070
rect 5533 22067 5599 22070
rect 13486 22068 13492 22070
rect 13556 22068 13562 22132
rect 9949 21996 10015 21997
rect 9949 21994 9996 21996
rect 9904 21992 9996 21994
rect 9904 21936 9954 21992
rect 9904 21934 9996 21936
rect 9949 21932 9996 21934
rect 10060 21932 10066 21996
rect 14774 21932 14780 21996
rect 14844 21994 14850 21996
rect 15285 21994 15351 21997
rect 14844 21992 15351 21994
rect 14844 21936 15290 21992
rect 15346 21936 15351 21992
rect 14844 21934 15351 21936
rect 14844 21932 14850 21934
rect 9949 21931 10015 21932
rect 15285 21931 15351 21934
rect 0 21798 3250 21858
rect 26325 21858 26391 21861
rect 29200 21858 30000 21888
rect 26325 21856 30000 21858
rect 26325 21800 26330 21856
rect 26386 21800 30000 21856
rect 26325 21798 30000 21800
rect 0 21768 800 21798
rect 26325 21795 26391 21798
rect 5944 21792 6264 21793
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 21727 6264 21728
rect 15944 21792 16264 21793
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 21727 16264 21728
rect 25944 21792 26264 21793
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 29200 21768 30000 21798
rect 25944 21727 26264 21728
rect 6453 21722 6519 21725
rect 7373 21722 7439 21725
rect 10317 21722 10383 21725
rect 10777 21724 10843 21725
rect 6453 21720 10383 21722
rect 6453 21664 6458 21720
rect 6514 21664 7378 21720
rect 7434 21664 10322 21720
rect 10378 21664 10383 21720
rect 6453 21662 10383 21664
rect 6453 21659 6519 21662
rect 7373 21659 7439 21662
rect 10317 21659 10383 21662
rect 10726 21660 10732 21724
rect 10796 21722 10843 21724
rect 18045 21724 18111 21725
rect 10796 21720 10888 21722
rect 10838 21664 10888 21720
rect 10796 21662 10888 21664
rect 18045 21720 18092 21724
rect 18156 21722 18162 21724
rect 18045 21664 18050 21720
rect 10796 21660 10843 21662
rect 10777 21659 10843 21660
rect 18045 21660 18092 21664
rect 18156 21662 18202 21722
rect 18156 21660 18162 21662
rect 18045 21659 18111 21660
rect 1301 21586 1367 21589
rect 2773 21586 2839 21589
rect 1301 21584 2839 21586
rect 1301 21528 1306 21584
rect 1362 21528 2778 21584
rect 2834 21528 2839 21584
rect 1301 21526 2839 21528
rect 1301 21523 1367 21526
rect 2773 21523 2839 21526
rect 3141 21586 3207 21589
rect 6361 21586 6427 21589
rect 8937 21586 9003 21589
rect 15653 21586 15719 21589
rect 17677 21586 17743 21589
rect 3141 21584 15719 21586
rect 3141 21528 3146 21584
rect 3202 21528 6366 21584
rect 6422 21528 8942 21584
rect 8998 21528 15658 21584
rect 15714 21528 15719 21584
rect 3141 21526 15719 21528
rect 3141 21523 3207 21526
rect 6361 21523 6427 21526
rect 8937 21523 9003 21526
rect 15653 21523 15719 21526
rect 16070 21584 17743 21586
rect 16070 21528 17682 21584
rect 17738 21528 17743 21584
rect 16070 21526 17743 21528
rect 8109 21450 8175 21453
rect 9857 21450 9923 21453
rect 16070 21450 16130 21526
rect 17677 21523 17743 21526
rect 8109 21448 16130 21450
rect 8109 21392 8114 21448
rect 8170 21392 9862 21448
rect 9918 21392 16130 21448
rect 8109 21390 16130 21392
rect 16205 21450 16271 21453
rect 18045 21450 18111 21453
rect 19885 21450 19951 21453
rect 16205 21448 19951 21450
rect 16205 21392 16210 21448
rect 16266 21392 18050 21448
rect 18106 21392 19890 21448
rect 19946 21392 19951 21448
rect 16205 21390 19951 21392
rect 8109 21387 8175 21390
rect 9857 21387 9923 21390
rect 16205 21387 16271 21390
rect 18045 21387 18111 21390
rect 19885 21387 19951 21390
rect 14641 21314 14707 21317
rect 19057 21314 19123 21317
rect 14641 21312 19123 21314
rect 14641 21256 14646 21312
rect 14702 21256 19062 21312
rect 19118 21256 19123 21312
rect 14641 21254 19123 21256
rect 14641 21251 14707 21254
rect 19057 21251 19123 21254
rect 10944 21248 11264 21249
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 10944 21183 11264 21184
rect 20944 21248 21264 21249
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 20944 21183 21264 21184
rect 15561 21178 15627 21181
rect 16941 21178 17007 21181
rect 15561 21176 17007 21178
rect 15561 21120 15566 21176
rect 15622 21120 16946 21176
rect 17002 21120 17007 21176
rect 15561 21118 17007 21120
rect 15561 21115 15627 21118
rect 16941 21115 17007 21118
rect 22921 21178 22987 21181
rect 25773 21178 25839 21181
rect 22921 21176 25839 21178
rect 22921 21120 22926 21176
rect 22982 21120 25778 21176
rect 25834 21120 25839 21176
rect 22921 21118 25839 21120
rect 22921 21115 22987 21118
rect 25773 21115 25839 21118
rect 11697 21042 11763 21045
rect 26325 21042 26391 21045
rect 11697 21040 26391 21042
rect 11697 20984 11702 21040
rect 11758 20984 26330 21040
rect 26386 20984 26391 21040
rect 11697 20982 26391 20984
rect 11697 20979 11763 20982
rect 26325 20979 26391 20982
rect 12249 20906 12315 20909
rect 14181 20906 14247 20909
rect 16665 20906 16731 20909
rect 12249 20904 14247 20906
rect 12249 20848 12254 20904
rect 12310 20848 14186 20904
rect 14242 20848 14247 20904
rect 12249 20846 14247 20848
rect 12249 20843 12315 20846
rect 14181 20843 14247 20846
rect 15702 20904 16731 20906
rect 15702 20848 16670 20904
rect 16726 20848 16731 20904
rect 15702 20846 16731 20848
rect 10777 20770 10843 20773
rect 15009 20770 15075 20773
rect 15702 20770 15762 20846
rect 16665 20843 16731 20846
rect 10777 20768 15762 20770
rect 10777 20712 10782 20768
rect 10838 20712 15014 20768
rect 15070 20712 15762 20768
rect 10777 20710 15762 20712
rect 19241 20770 19307 20773
rect 23749 20770 23815 20773
rect 19241 20768 23815 20770
rect 19241 20712 19246 20768
rect 19302 20712 23754 20768
rect 23810 20712 23815 20768
rect 19241 20710 23815 20712
rect 10777 20707 10843 20710
rect 15009 20707 15075 20710
rect 19241 20707 19307 20710
rect 23749 20707 23815 20710
rect 24025 20770 24091 20773
rect 24025 20768 24962 20770
rect 24025 20712 24030 20768
rect 24086 20712 24962 20768
rect 24025 20710 24962 20712
rect 24025 20707 24091 20710
rect 5944 20704 6264 20705
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 20639 6264 20640
rect 15944 20704 16264 20705
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 20639 16264 20640
rect 9489 20634 9555 20637
rect 11053 20634 11119 20637
rect 9489 20632 11119 20634
rect 9489 20576 9494 20632
rect 9550 20576 11058 20632
rect 11114 20576 11119 20632
rect 9489 20574 11119 20576
rect 9489 20571 9555 20574
rect 11053 20571 11119 20574
rect 21725 20634 21791 20637
rect 22277 20634 22343 20637
rect 21725 20632 22343 20634
rect 21725 20576 21730 20632
rect 21786 20576 22282 20632
rect 22338 20576 22343 20632
rect 21725 20574 22343 20576
rect 21725 20571 21791 20574
rect 22277 20571 22343 20574
rect 0 20498 800 20528
rect 1853 20498 1919 20501
rect 0 20496 1919 20498
rect 0 20440 1858 20496
rect 1914 20440 1919 20496
rect 0 20438 1919 20440
rect 0 20408 800 20438
rect 1853 20435 1919 20438
rect 9673 20498 9739 20501
rect 13077 20498 13143 20501
rect 9673 20496 13143 20498
rect 9673 20440 9678 20496
rect 9734 20440 13082 20496
rect 13138 20440 13143 20496
rect 9673 20438 13143 20440
rect 9673 20435 9739 20438
rect 13077 20435 13143 20438
rect 14958 20436 14964 20500
rect 15028 20498 15034 20500
rect 16665 20498 16731 20501
rect 15028 20496 16731 20498
rect 15028 20440 16670 20496
rect 16726 20440 16731 20496
rect 15028 20438 16731 20440
rect 24902 20498 24962 20710
rect 25944 20704 26264 20705
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 20639 26264 20640
rect 29200 20498 30000 20528
rect 24902 20438 30000 20498
rect 15028 20436 15034 20438
rect 16665 20435 16731 20438
rect 29200 20408 30000 20438
rect 8201 20362 8267 20365
rect 9305 20362 9371 20365
rect 12198 20362 12204 20364
rect 8201 20360 12204 20362
rect 8201 20304 8206 20360
rect 8262 20304 9310 20360
rect 9366 20304 12204 20360
rect 8201 20302 12204 20304
rect 8201 20299 8267 20302
rect 9305 20299 9371 20302
rect 12198 20300 12204 20302
rect 12268 20300 12274 20364
rect 13629 20362 13695 20365
rect 19517 20362 19583 20365
rect 27705 20362 27771 20365
rect 13629 20360 19583 20362
rect 13629 20304 13634 20360
rect 13690 20304 19522 20360
rect 19578 20304 19583 20360
rect 13629 20302 19583 20304
rect 13629 20299 13695 20302
rect 19517 20299 19583 20302
rect 19750 20360 27771 20362
rect 19750 20304 27710 20360
rect 27766 20304 27771 20360
rect 19750 20302 27771 20304
rect 9673 20228 9739 20229
rect 9622 20164 9628 20228
rect 9692 20226 9739 20228
rect 15009 20226 15075 20229
rect 19750 20226 19810 20302
rect 27705 20299 27771 20302
rect 9692 20224 9784 20226
rect 9734 20168 9784 20224
rect 9692 20166 9784 20168
rect 15009 20224 19810 20226
rect 15009 20168 15014 20224
rect 15070 20168 19810 20224
rect 15009 20166 19810 20168
rect 21449 20226 21515 20229
rect 25589 20226 25655 20229
rect 21449 20224 25655 20226
rect 21449 20168 21454 20224
rect 21510 20168 25594 20224
rect 25650 20168 25655 20224
rect 21449 20166 25655 20168
rect 9692 20164 9739 20166
rect 9673 20163 9739 20164
rect 15009 20163 15075 20166
rect 21449 20163 21515 20166
rect 25589 20163 25655 20166
rect 10944 20160 11264 20161
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 10944 20095 11264 20096
rect 20944 20160 21264 20161
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 20944 20095 21264 20096
rect 2957 19954 3023 19957
rect 17033 19954 17099 19957
rect 2957 19952 17099 19954
rect 2957 19896 2962 19952
rect 3018 19896 17038 19952
rect 17094 19896 17099 19952
rect 2957 19894 17099 19896
rect 2957 19891 3023 19894
rect 17033 19891 17099 19894
rect 11145 19818 11211 19821
rect 11462 19818 11468 19820
rect 11145 19816 11468 19818
rect 11145 19760 11150 19816
rect 11206 19760 11468 19816
rect 11145 19758 11468 19760
rect 11145 19755 11211 19758
rect 11462 19756 11468 19758
rect 11532 19756 11538 19820
rect 5944 19616 6264 19617
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 19551 6264 19552
rect 15944 19616 16264 19617
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 19551 16264 19552
rect 25944 19616 26264 19617
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 19551 26264 19552
rect 8937 19546 9003 19549
rect 10225 19546 10291 19549
rect 8937 19544 10291 19546
rect 8937 19488 8942 19544
rect 8998 19488 10230 19544
rect 10286 19488 10291 19544
rect 8937 19486 10291 19488
rect 8937 19483 9003 19486
rect 10225 19483 10291 19486
rect 14549 19546 14615 19549
rect 15377 19546 15443 19549
rect 14549 19544 15443 19546
rect 14549 19488 14554 19544
rect 14610 19488 15382 19544
rect 15438 19488 15443 19544
rect 14549 19486 15443 19488
rect 14549 19483 14615 19486
rect 15377 19483 15443 19486
rect 20161 19546 20227 19549
rect 21173 19546 21239 19549
rect 20161 19544 21239 19546
rect 20161 19488 20166 19544
rect 20222 19488 21178 19544
rect 21234 19488 21239 19544
rect 20161 19486 21239 19488
rect 20161 19483 20227 19486
rect 21173 19483 21239 19486
rect 13445 19410 13511 19413
rect 17125 19410 17191 19413
rect 13445 19408 17191 19410
rect 13445 19352 13450 19408
rect 13506 19352 17130 19408
rect 17186 19352 17191 19408
rect 13445 19350 17191 19352
rect 13445 19347 13511 19350
rect 17125 19347 17191 19350
rect 9029 19276 9095 19277
rect 9029 19274 9076 19276
rect 8984 19272 9076 19274
rect 8984 19216 9034 19272
rect 8984 19214 9076 19216
rect 9029 19212 9076 19214
rect 9140 19212 9146 19276
rect 9765 19274 9831 19277
rect 16757 19274 16823 19277
rect 9765 19272 16823 19274
rect 9765 19216 9770 19272
rect 9826 19216 16762 19272
rect 16818 19216 16823 19272
rect 9765 19214 16823 19216
rect 9029 19211 9095 19212
rect 9765 19211 9831 19214
rect 16757 19211 16823 19214
rect 17033 19274 17099 19277
rect 21909 19274 21975 19277
rect 24209 19274 24275 19277
rect 17033 19272 21466 19274
rect 17033 19216 17038 19272
rect 17094 19216 21466 19272
rect 17033 19214 21466 19216
rect 17033 19211 17099 19214
rect 0 19138 800 19168
rect 6729 19138 6795 19141
rect 0 19136 6795 19138
rect 0 19080 6734 19136
rect 6790 19080 6795 19136
rect 0 19078 6795 19080
rect 21406 19138 21466 19214
rect 21909 19272 24275 19274
rect 21909 19216 21914 19272
rect 21970 19216 24214 19272
rect 24270 19216 24275 19272
rect 21909 19214 24275 19216
rect 21909 19211 21975 19214
rect 24209 19211 24275 19214
rect 29200 19138 30000 19168
rect 21406 19078 30000 19138
rect 0 19048 800 19078
rect 6729 19075 6795 19078
rect 10944 19072 11264 19073
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10944 19007 11264 19008
rect 20944 19072 21264 19073
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 29200 19048 30000 19078
rect 20944 19007 21264 19008
rect 10501 18868 10567 18869
rect 10501 18866 10548 18868
rect 10456 18864 10548 18866
rect 10456 18808 10506 18864
rect 10456 18806 10548 18808
rect 10501 18804 10548 18806
rect 10612 18804 10618 18868
rect 10501 18803 10567 18804
rect 25589 18730 25655 18733
rect 25589 18728 26434 18730
rect 25589 18672 25594 18728
rect 25650 18672 26434 18728
rect 25589 18670 26434 18672
rect 25589 18667 25655 18670
rect 5944 18528 6264 18529
rect 0 18458 800 18488
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 18463 6264 18464
rect 15944 18528 16264 18529
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 18463 16264 18464
rect 25944 18528 26264 18529
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25944 18463 26264 18464
rect 3233 18458 3299 18461
rect 0 18456 3299 18458
rect 0 18400 3238 18456
rect 3294 18400 3299 18456
rect 0 18398 3299 18400
rect 26374 18458 26434 18670
rect 29200 18458 30000 18488
rect 26374 18398 30000 18458
rect 0 18368 800 18398
rect 3233 18395 3299 18398
rect 29200 18368 30000 18398
rect 11329 18322 11395 18325
rect 12382 18322 12388 18324
rect 11329 18320 12388 18322
rect 11329 18264 11334 18320
rect 11390 18264 12388 18320
rect 11329 18262 12388 18264
rect 11329 18259 11395 18262
rect 12382 18260 12388 18262
rect 12452 18322 12458 18324
rect 15101 18322 15167 18325
rect 12452 18320 15167 18322
rect 12452 18264 15106 18320
rect 15162 18264 15167 18320
rect 12452 18262 15167 18264
rect 12452 18260 12458 18262
rect 15101 18259 15167 18262
rect 10777 18186 10843 18189
rect 12709 18186 12775 18189
rect 10777 18184 12775 18186
rect 10777 18128 10782 18184
rect 10838 18128 12714 18184
rect 12770 18128 12775 18184
rect 10777 18126 12775 18128
rect 10777 18123 10843 18126
rect 12709 18123 12775 18126
rect 13721 18186 13787 18189
rect 14590 18186 14596 18188
rect 13721 18184 14596 18186
rect 13721 18128 13726 18184
rect 13782 18128 14596 18184
rect 13721 18126 14596 18128
rect 13721 18123 13787 18126
rect 14590 18124 14596 18126
rect 14660 18124 14666 18188
rect 10944 17984 11264 17985
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 17919 11264 17920
rect 20944 17984 21264 17985
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 20944 17919 21264 17920
rect 13261 17914 13327 17917
rect 15561 17914 15627 17917
rect 13261 17912 15627 17914
rect 13261 17856 13266 17912
rect 13322 17856 15566 17912
rect 15622 17856 15627 17912
rect 13261 17854 15627 17856
rect 13261 17851 13327 17854
rect 15561 17851 15627 17854
rect 9581 17778 9647 17781
rect 10501 17778 10567 17781
rect 9581 17776 10567 17778
rect 9581 17720 9586 17776
rect 9642 17720 10506 17776
rect 10562 17720 10567 17776
rect 9581 17718 10567 17720
rect 9581 17715 9647 17718
rect 10501 17715 10567 17718
rect 17166 17716 17172 17780
rect 17236 17778 17242 17780
rect 25497 17778 25563 17781
rect 17236 17776 25563 17778
rect 17236 17720 25502 17776
rect 25558 17720 25563 17776
rect 17236 17718 25563 17720
rect 17236 17716 17242 17718
rect 25497 17715 25563 17718
rect 5944 17440 6264 17441
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 17375 6264 17376
rect 15944 17440 16264 17441
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 17375 16264 17376
rect 25944 17440 26264 17441
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 17375 26264 17376
rect 12985 17370 13051 17373
rect 15561 17370 15627 17373
rect 12985 17368 15627 17370
rect 12985 17312 12990 17368
rect 13046 17312 15566 17368
rect 15622 17312 15627 17368
rect 12985 17310 15627 17312
rect 12985 17307 13051 17310
rect 15561 17307 15627 17310
rect 1669 17234 1735 17237
rect 11421 17234 11487 17237
rect 1669 17232 11487 17234
rect 1669 17176 1674 17232
rect 1730 17176 11426 17232
rect 11482 17176 11487 17232
rect 1669 17174 11487 17176
rect 1669 17171 1735 17174
rect 11421 17171 11487 17174
rect 0 17098 800 17128
rect 1485 17098 1551 17101
rect 0 17096 1551 17098
rect 0 17040 1490 17096
rect 1546 17040 1551 17096
rect 0 17038 1551 17040
rect 0 17008 800 17038
rect 1485 17035 1551 17038
rect 9489 17098 9555 17101
rect 11237 17098 11303 17101
rect 12433 17098 12499 17101
rect 9489 17096 12499 17098
rect 9489 17040 9494 17096
rect 9550 17040 11242 17096
rect 11298 17040 12438 17096
rect 12494 17040 12499 17096
rect 9489 17038 12499 17040
rect 9489 17035 9555 17038
rect 11237 17035 11303 17038
rect 12433 17035 12499 17038
rect 17401 17098 17467 17101
rect 29200 17098 30000 17128
rect 17401 17096 30000 17098
rect 17401 17040 17406 17096
rect 17462 17040 30000 17096
rect 17401 17038 30000 17040
rect 17401 17035 17467 17038
rect 29200 17008 30000 17038
rect 10944 16896 11264 16897
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 16831 11264 16832
rect 20944 16896 21264 16897
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 16831 21264 16832
rect 5944 16352 6264 16353
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 16287 6264 16288
rect 15944 16352 16264 16353
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 16287 16264 16288
rect 25944 16352 26264 16353
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 25944 16287 26264 16288
rect 10593 16146 10659 16149
rect 16205 16146 16271 16149
rect 10593 16144 16271 16146
rect 10593 16088 10598 16144
rect 10654 16088 16210 16144
rect 16266 16088 16271 16144
rect 10593 16086 16271 16088
rect 10593 16083 10659 16086
rect 16205 16083 16271 16086
rect 8661 16010 8727 16013
rect 12525 16010 12591 16013
rect 15377 16010 15443 16013
rect 8661 16008 15443 16010
rect 8661 15952 8666 16008
rect 8722 15952 12530 16008
rect 12586 15952 15382 16008
rect 15438 15952 15443 16008
rect 8661 15950 15443 15952
rect 8661 15947 8727 15950
rect 12525 15947 12591 15950
rect 15377 15947 15443 15950
rect 10944 15808 11264 15809
rect 0 15738 800 15768
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 15743 11264 15744
rect 20944 15808 21264 15809
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 20944 15743 21264 15744
rect 7281 15738 7347 15741
rect 0 15736 7347 15738
rect 0 15680 7286 15736
rect 7342 15680 7347 15736
rect 0 15678 7347 15680
rect 0 15648 800 15678
rect 7281 15675 7347 15678
rect 15009 15738 15075 15741
rect 16849 15738 16915 15741
rect 29200 15738 30000 15768
rect 15009 15736 16915 15738
rect 15009 15680 15014 15736
rect 15070 15680 16854 15736
rect 16910 15680 16915 15736
rect 15009 15678 16915 15680
rect 15009 15675 15075 15678
rect 16849 15675 16915 15678
rect 24350 15678 30000 15738
rect 8109 15602 8175 15605
rect 10041 15602 10107 15605
rect 12249 15602 12315 15605
rect 12433 15602 12499 15605
rect 8109 15600 12499 15602
rect 8109 15544 8114 15600
rect 8170 15544 10046 15600
rect 10102 15544 12254 15600
rect 12310 15544 12438 15600
rect 12494 15544 12499 15600
rect 8109 15542 12499 15544
rect 8109 15539 8175 15542
rect 10041 15539 10107 15542
rect 12249 15539 12315 15542
rect 12433 15539 12499 15542
rect 13353 15602 13419 15605
rect 15469 15602 15535 15605
rect 13353 15600 15535 15602
rect 13353 15544 13358 15600
rect 13414 15544 15474 15600
rect 15530 15544 15535 15600
rect 13353 15542 15535 15544
rect 13353 15539 13419 15542
rect 15469 15539 15535 15542
rect 11421 15466 11487 15469
rect 24350 15466 24410 15678
rect 29200 15648 30000 15678
rect 11421 15464 24410 15466
rect 11421 15408 11426 15464
rect 11482 15408 24410 15464
rect 11421 15406 24410 15408
rect 11421 15403 11487 15406
rect 10317 15330 10383 15333
rect 14181 15330 14247 15333
rect 10317 15328 14247 15330
rect 10317 15272 10322 15328
rect 10378 15272 14186 15328
rect 14242 15272 14247 15328
rect 10317 15270 14247 15272
rect 10317 15267 10383 15270
rect 14181 15267 14247 15270
rect 22461 15330 22527 15333
rect 22461 15328 24962 15330
rect 22461 15272 22466 15328
rect 22522 15272 24962 15328
rect 22461 15270 24962 15272
rect 22461 15267 22527 15270
rect 5944 15264 6264 15265
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 15199 6264 15200
rect 15944 15264 16264 15265
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 15199 16264 15200
rect 0 15058 800 15088
rect 7557 15058 7623 15061
rect 0 15056 7623 15058
rect 0 15000 7562 15056
rect 7618 15000 7623 15056
rect 0 14998 7623 15000
rect 0 14968 800 14998
rect 7557 14995 7623 14998
rect 12617 15058 12683 15061
rect 12750 15058 12756 15060
rect 12617 15056 12756 15058
rect 12617 15000 12622 15056
rect 12678 15000 12756 15056
rect 12617 14998 12756 15000
rect 12617 14995 12683 14998
rect 12750 14996 12756 14998
rect 12820 14996 12826 15060
rect 24902 15058 24962 15270
rect 25944 15264 26264 15265
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 25944 15199 26264 15200
rect 29200 15058 30000 15088
rect 24902 14998 30000 15058
rect 29200 14968 30000 14998
rect 10944 14720 11264 14721
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 10944 14655 11264 14656
rect 20944 14720 21264 14721
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 14655 21264 14656
rect 14641 14650 14707 14653
rect 17401 14650 17467 14653
rect 14641 14648 17467 14650
rect 14641 14592 14646 14648
rect 14702 14592 17406 14648
rect 17462 14592 17467 14648
rect 14641 14590 17467 14592
rect 14641 14587 14707 14590
rect 17401 14587 17467 14590
rect 9949 14378 10015 14381
rect 14917 14378 14983 14381
rect 22553 14378 22619 14381
rect 9949 14376 22619 14378
rect 9949 14320 9954 14376
rect 10010 14320 14922 14376
rect 14978 14320 22558 14376
rect 22614 14320 22619 14376
rect 9949 14318 22619 14320
rect 9949 14315 10015 14318
rect 14917 14315 14983 14318
rect 22553 14315 22619 14318
rect 5944 14176 6264 14177
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 14111 6264 14112
rect 15944 14176 16264 14177
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 14111 16264 14112
rect 25944 14176 26264 14177
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 14111 26264 14112
rect 12985 13970 13051 13973
rect 15561 13970 15627 13973
rect 12985 13968 15627 13970
rect 12985 13912 12990 13968
rect 13046 13912 15566 13968
rect 15622 13912 15627 13968
rect 12985 13910 15627 13912
rect 12985 13907 13051 13910
rect 15561 13907 15627 13910
rect 22001 13970 22067 13973
rect 27613 13970 27679 13973
rect 22001 13968 27679 13970
rect 22001 13912 22006 13968
rect 22062 13912 27618 13968
rect 27674 13912 27679 13968
rect 22001 13910 27679 13912
rect 22001 13907 22067 13910
rect 27613 13907 27679 13910
rect 26233 13834 26299 13837
rect 23246 13832 26299 13834
rect 23246 13776 26238 13832
rect 26294 13776 26299 13832
rect 23246 13774 26299 13776
rect 0 13698 800 13728
rect 2037 13698 2103 13701
rect 0 13696 2103 13698
rect 0 13640 2042 13696
rect 2098 13640 2103 13696
rect 0 13638 2103 13640
rect 0 13608 800 13638
rect 2037 13635 2103 13638
rect 15009 13698 15075 13701
rect 17493 13698 17559 13701
rect 15009 13696 17559 13698
rect 15009 13640 15014 13696
rect 15070 13640 17498 13696
rect 17554 13640 17559 13696
rect 15009 13638 17559 13640
rect 15009 13635 15075 13638
rect 17493 13635 17559 13638
rect 21633 13698 21699 13701
rect 22737 13698 22803 13701
rect 23246 13698 23306 13774
rect 26233 13771 26299 13774
rect 26509 13834 26575 13837
rect 26509 13832 26618 13834
rect 26509 13776 26514 13832
rect 26570 13776 26618 13832
rect 26509 13771 26618 13776
rect 21633 13696 23306 13698
rect 21633 13640 21638 13696
rect 21694 13640 22742 13696
rect 22798 13640 23306 13696
rect 21633 13638 23306 13640
rect 26558 13698 26618 13771
rect 29200 13698 30000 13728
rect 26558 13638 30000 13698
rect 21633 13635 21699 13638
rect 22737 13635 22803 13638
rect 10944 13632 11264 13633
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 10944 13567 11264 13568
rect 20944 13632 21264 13633
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 29200 13608 30000 13638
rect 20944 13567 21264 13568
rect 13537 13562 13603 13565
rect 13670 13562 13676 13564
rect 13537 13560 13676 13562
rect 13537 13504 13542 13560
rect 13598 13504 13676 13560
rect 13537 13502 13676 13504
rect 13537 13499 13603 13502
rect 13670 13500 13676 13502
rect 13740 13500 13746 13564
rect 3049 13426 3115 13429
rect 25405 13426 25471 13429
rect 3049 13424 25471 13426
rect 3049 13368 3054 13424
rect 3110 13368 25410 13424
rect 25466 13368 25471 13424
rect 3049 13366 25471 13368
rect 3049 13363 3115 13366
rect 25405 13363 25471 13366
rect 3325 13290 3391 13293
rect 8385 13290 8451 13293
rect 3325 13288 8451 13290
rect 3325 13232 3330 13288
rect 3386 13232 8390 13288
rect 8446 13232 8451 13288
rect 3325 13230 8451 13232
rect 3325 13227 3391 13230
rect 8385 13227 8451 13230
rect 9765 13290 9831 13293
rect 11973 13290 12039 13293
rect 9765 13288 12039 13290
rect 9765 13232 9770 13288
rect 9826 13232 11978 13288
rect 12034 13232 12039 13288
rect 9765 13230 12039 13232
rect 9765 13227 9831 13230
rect 11973 13227 12039 13230
rect 5944 13088 6264 13089
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 13023 6264 13024
rect 15944 13088 16264 13089
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 13023 16264 13024
rect 25944 13088 26264 13089
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25944 13023 26264 13024
rect 12014 12684 12020 12748
rect 12084 12746 12090 12748
rect 19374 12746 19380 12748
rect 12084 12686 19380 12746
rect 12084 12684 12090 12686
rect 19374 12684 19380 12686
rect 19444 12684 19450 12748
rect 10944 12544 11264 12545
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 12479 11264 12480
rect 20944 12544 21264 12545
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 20944 12479 21264 12480
rect 0 12338 800 12368
rect 1577 12338 1643 12341
rect 0 12336 1643 12338
rect 0 12280 1582 12336
rect 1638 12280 1643 12336
rect 0 12278 1643 12280
rect 0 12248 800 12278
rect 1577 12275 1643 12278
rect 19374 12276 19380 12340
rect 19444 12338 19450 12340
rect 29200 12338 30000 12368
rect 19444 12278 30000 12338
rect 19444 12276 19450 12278
rect 29200 12248 30000 12278
rect 15377 12202 15443 12205
rect 17861 12202 17927 12205
rect 15377 12200 17927 12202
rect 15377 12144 15382 12200
rect 15438 12144 17866 12200
rect 17922 12144 17927 12200
rect 15377 12142 17927 12144
rect 15377 12139 15443 12142
rect 17861 12139 17927 12142
rect 9070 12004 9076 12068
rect 9140 12066 9146 12068
rect 14917 12066 14983 12069
rect 9140 12064 14983 12066
rect 9140 12008 14922 12064
rect 14978 12008 14983 12064
rect 9140 12006 14983 12008
rect 9140 12004 9146 12006
rect 14917 12003 14983 12006
rect 5944 12000 6264 12001
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 11935 6264 11936
rect 15944 12000 16264 12001
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 15944 11935 16264 11936
rect 25944 12000 26264 12001
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25944 11935 26264 11936
rect 17217 11794 17283 11797
rect 22553 11794 22619 11797
rect 17217 11792 22619 11794
rect 17217 11736 17222 11792
rect 17278 11736 22558 11792
rect 22614 11736 22619 11792
rect 17217 11734 22619 11736
rect 17217 11731 17283 11734
rect 22553 11731 22619 11734
rect 18413 11658 18479 11661
rect 25221 11658 25287 11661
rect 29200 11658 30000 11688
rect 18413 11656 24226 11658
rect 18413 11600 18418 11656
rect 18474 11600 24226 11656
rect 18413 11598 24226 11600
rect 18413 11595 18479 11598
rect 24166 11522 24226 11598
rect 25221 11656 30000 11658
rect 25221 11600 25226 11656
rect 25282 11600 30000 11656
rect 25221 11598 30000 11600
rect 25221 11595 25287 11598
rect 29200 11568 30000 11598
rect 26325 11522 26391 11525
rect 24166 11520 26391 11522
rect 24166 11464 26330 11520
rect 26386 11464 26391 11520
rect 24166 11462 26391 11464
rect 26325 11459 26391 11462
rect 10944 11456 11264 11457
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 10944 11391 11264 11392
rect 20944 11456 21264 11457
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 11391 21264 11392
rect 13997 11386 14063 11389
rect 15694 11386 15700 11388
rect 13997 11384 15700 11386
rect 13997 11328 14002 11384
rect 14058 11328 15700 11384
rect 13997 11326 15700 11328
rect 13997 11323 14063 11326
rect 15694 11324 15700 11326
rect 15764 11324 15770 11388
rect 3969 11250 4035 11253
rect 6913 11250 6979 11253
rect 3969 11248 6979 11250
rect 3969 11192 3974 11248
rect 4030 11192 6918 11248
rect 6974 11192 6979 11248
rect 3969 11190 6979 11192
rect 3969 11187 4035 11190
rect 6913 11187 6979 11190
rect 4613 11114 4679 11117
rect 5809 11114 5875 11117
rect 4613 11112 5875 11114
rect 4613 11056 4618 11112
rect 4674 11056 5814 11112
rect 5870 11056 5875 11112
rect 4613 11054 5875 11056
rect 4613 11051 4679 11054
rect 5809 11051 5875 11054
rect 0 10978 800 11008
rect 4061 10978 4127 10981
rect 0 10976 4127 10978
rect 0 10920 4066 10976
rect 4122 10920 4127 10976
rect 0 10918 4127 10920
rect 0 10888 800 10918
rect 4061 10915 4127 10918
rect 5944 10912 6264 10913
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 10847 6264 10848
rect 15944 10912 16264 10913
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 10847 16264 10848
rect 25944 10912 26264 10913
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 10847 26264 10848
rect 10542 10780 10548 10844
rect 10612 10842 10618 10844
rect 11605 10842 11671 10845
rect 10612 10840 11671 10842
rect 10612 10784 11610 10840
rect 11666 10784 11671 10840
rect 10612 10782 11671 10784
rect 10612 10780 10618 10782
rect 11605 10779 11671 10782
rect 2313 10706 2379 10709
rect 22829 10706 22895 10709
rect 2313 10704 22895 10706
rect 2313 10648 2318 10704
rect 2374 10648 22834 10704
rect 22890 10648 22895 10704
rect 2313 10646 22895 10648
rect 2313 10643 2379 10646
rect 22829 10643 22895 10646
rect 3877 10570 3943 10573
rect 19057 10570 19123 10573
rect 3877 10568 19123 10570
rect 3877 10512 3882 10568
rect 3938 10512 19062 10568
rect 19118 10512 19123 10568
rect 3877 10510 19123 10512
rect 3877 10507 3943 10510
rect 19057 10507 19123 10510
rect 10944 10368 11264 10369
rect 0 10298 800 10328
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 10303 11264 10304
rect 20944 10368 21264 10369
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 20944 10303 21264 10304
rect 3509 10298 3575 10301
rect 0 10296 3575 10298
rect 0 10240 3514 10296
rect 3570 10240 3575 10296
rect 0 10238 3575 10240
rect 0 10208 800 10238
rect 3509 10235 3575 10238
rect 21725 10298 21791 10301
rect 29200 10298 30000 10328
rect 21725 10296 30000 10298
rect 21725 10240 21730 10296
rect 21786 10240 30000 10296
rect 21725 10238 30000 10240
rect 21725 10235 21791 10238
rect 29200 10208 30000 10238
rect 4061 10162 4127 10165
rect 13997 10162 14063 10165
rect 4061 10160 14063 10162
rect 4061 10104 4066 10160
rect 4122 10104 14002 10160
rect 14058 10104 14063 10160
rect 4061 10102 14063 10104
rect 4061 10099 4127 10102
rect 13997 10099 14063 10102
rect 5944 9824 6264 9825
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 9759 6264 9760
rect 15944 9824 16264 9825
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 9759 16264 9760
rect 25944 9824 26264 9825
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 25944 9759 26264 9760
rect 10501 9754 10567 9757
rect 10501 9752 13738 9754
rect 10501 9696 10506 9752
rect 10562 9696 13738 9752
rect 10501 9694 13738 9696
rect 10501 9691 10567 9694
rect 13678 9618 13738 9694
rect 14917 9618 14983 9621
rect 13678 9616 14983 9618
rect 13678 9560 14922 9616
rect 14978 9560 14983 9616
rect 13678 9558 14983 9560
rect 14917 9555 14983 9558
rect 14457 9482 14523 9485
rect 16297 9482 16363 9485
rect 14457 9480 16363 9482
rect 14457 9424 14462 9480
rect 14518 9424 16302 9480
rect 16358 9424 16363 9480
rect 14457 9422 16363 9424
rect 14457 9419 14523 9422
rect 16297 9419 16363 9422
rect 10944 9280 11264 9281
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 9215 11264 9216
rect 20944 9280 21264 9281
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 20944 9215 21264 9216
rect 2037 9074 2103 9077
rect 7925 9074 7991 9077
rect 9673 9074 9739 9077
rect 2037 9072 9739 9074
rect 2037 9016 2042 9072
rect 2098 9016 7930 9072
rect 7986 9016 9678 9072
rect 9734 9016 9739 9072
rect 2037 9014 9739 9016
rect 2037 9011 2103 9014
rect 7925 9011 7991 9014
rect 9673 9011 9739 9014
rect 12985 9074 13051 9077
rect 17033 9074 17099 9077
rect 12985 9072 17099 9074
rect 12985 9016 12990 9072
rect 13046 9016 17038 9072
rect 17094 9016 17099 9072
rect 12985 9014 17099 9016
rect 12985 9011 13051 9014
rect 17033 9011 17099 9014
rect 0 8938 800 8968
rect 3325 8938 3391 8941
rect 0 8936 3391 8938
rect 0 8880 3330 8936
rect 3386 8880 3391 8936
rect 0 8878 3391 8880
rect 0 8848 800 8878
rect 3325 8875 3391 8878
rect 16849 8938 16915 8941
rect 29200 8938 30000 8968
rect 16849 8936 30000 8938
rect 16849 8880 16854 8936
rect 16910 8880 30000 8936
rect 16849 8878 30000 8880
rect 16849 8875 16915 8878
rect 29200 8848 30000 8878
rect 5944 8736 6264 8737
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 8671 6264 8672
rect 15944 8736 16264 8737
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 8671 16264 8672
rect 25944 8736 26264 8737
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25944 8671 26264 8672
rect 16481 8530 16547 8533
rect 29453 8530 29519 8533
rect 16481 8528 29519 8530
rect 16481 8472 16486 8528
rect 16542 8472 29458 8528
rect 29514 8472 29519 8528
rect 16481 8470 29519 8472
rect 16481 8467 16547 8470
rect 29453 8467 29519 8470
rect 17033 8394 17099 8397
rect 21817 8394 21883 8397
rect 17033 8392 21883 8394
rect 17033 8336 17038 8392
rect 17094 8336 21822 8392
rect 21878 8336 21883 8392
rect 17033 8334 21883 8336
rect 17033 8331 17099 8334
rect 21817 8331 21883 8334
rect 15193 8258 15259 8261
rect 18137 8258 18203 8261
rect 15193 8256 18203 8258
rect 15193 8200 15198 8256
rect 15254 8200 18142 8256
rect 18198 8200 18203 8256
rect 15193 8198 18203 8200
rect 15193 8195 15259 8198
rect 18137 8195 18203 8198
rect 25262 8196 25268 8260
rect 25332 8258 25338 8260
rect 29200 8258 30000 8288
rect 25332 8198 30000 8258
rect 25332 8196 25338 8198
rect 10944 8192 11264 8193
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 8127 11264 8128
rect 20944 8192 21264 8193
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 29200 8168 30000 8198
rect 20944 8127 21264 8128
rect 14549 8122 14615 8125
rect 15469 8122 15535 8125
rect 14549 8120 15535 8122
rect 14549 8064 14554 8120
rect 14610 8064 15474 8120
rect 15530 8064 15535 8120
rect 14549 8062 15535 8064
rect 14549 8059 14615 8062
rect 15469 8059 15535 8062
rect 13 7986 79 7989
rect 9857 7986 9923 7989
rect 13445 7986 13511 7989
rect 13 7984 7666 7986
rect 13 7928 18 7984
rect 74 7928 7666 7984
rect 13 7926 7666 7928
rect 13 7923 79 7926
rect 7606 7850 7666 7926
rect 9857 7984 13511 7986
rect 9857 7928 9862 7984
rect 9918 7928 13450 7984
rect 13506 7928 13511 7984
rect 9857 7926 13511 7928
rect 9857 7923 9923 7926
rect 13445 7923 13511 7926
rect 15326 7850 15332 7852
rect 7606 7790 15332 7850
rect 15326 7788 15332 7790
rect 15396 7788 15402 7852
rect 5944 7648 6264 7649
rect 0 7578 800 7608
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 7583 6264 7584
rect 15944 7648 16264 7649
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 7583 16264 7584
rect 25944 7648 26264 7649
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 7583 26264 7584
rect 1577 7578 1643 7581
rect 0 7576 1643 7578
rect 0 7520 1582 7576
rect 1638 7520 1643 7576
rect 0 7518 1643 7520
rect 0 7488 800 7518
rect 1577 7515 1643 7518
rect 7649 7578 7715 7581
rect 8293 7578 8359 7581
rect 7649 7576 8359 7578
rect 7649 7520 7654 7576
rect 7710 7520 8298 7576
rect 8354 7520 8359 7576
rect 7649 7518 8359 7520
rect 7649 7515 7715 7518
rect 8293 7515 8359 7518
rect 6269 7442 6335 7445
rect 7741 7442 7807 7445
rect 6269 7440 7807 7442
rect 6269 7384 6274 7440
rect 6330 7384 7746 7440
rect 7802 7384 7807 7440
rect 6269 7382 7807 7384
rect 6269 7379 6335 7382
rect 7741 7379 7807 7382
rect 13721 7442 13787 7445
rect 24945 7442 25011 7445
rect 13721 7440 25011 7442
rect 13721 7384 13726 7440
rect 13782 7384 24950 7440
rect 25006 7384 25011 7440
rect 13721 7382 25011 7384
rect 13721 7379 13787 7382
rect 24945 7379 25011 7382
rect 17769 7306 17835 7309
rect 17769 7304 25698 7306
rect 17769 7248 17774 7304
rect 17830 7248 25698 7304
rect 17769 7246 25698 7248
rect 17769 7243 17835 7246
rect 10944 7104 11264 7105
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 7039 11264 7040
rect 20944 7104 21264 7105
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 7039 21264 7040
rect 4061 7034 4127 7037
rect 9029 7034 9095 7037
rect 4061 7032 9095 7034
rect 4061 6976 4066 7032
rect 4122 6976 9034 7032
rect 9090 6976 9095 7032
rect 4061 6974 9095 6976
rect 4061 6971 4127 6974
rect 9029 6971 9095 6974
rect 0 6898 800 6928
rect 3877 6898 3943 6901
rect 0 6896 3943 6898
rect 0 6840 3882 6896
rect 3938 6840 3943 6896
rect 0 6838 3943 6840
rect 0 6808 800 6838
rect 3877 6835 3943 6838
rect 24393 6898 24459 6901
rect 25313 6898 25379 6901
rect 24393 6896 25379 6898
rect 24393 6840 24398 6896
rect 24454 6840 25318 6896
rect 25374 6840 25379 6896
rect 24393 6838 25379 6840
rect 25638 6898 25698 7246
rect 29200 6898 30000 6928
rect 25638 6838 30000 6898
rect 24393 6835 24459 6838
rect 25313 6835 25379 6838
rect 29200 6808 30000 6838
rect 5944 6560 6264 6561
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 6495 6264 6496
rect 15944 6560 16264 6561
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 6495 16264 6496
rect 25944 6560 26264 6561
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 6495 26264 6496
rect 473 6218 539 6221
rect 22001 6218 22067 6221
rect 473 6216 22067 6218
rect 473 6160 478 6216
rect 534 6160 22006 6216
rect 22062 6160 22067 6216
rect 473 6158 22067 6160
rect 473 6155 539 6158
rect 22001 6155 22067 6158
rect 10944 6016 11264 6017
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 5951 11264 5952
rect 20944 6016 21264 6017
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 5951 21264 5952
rect 0 5538 800 5568
rect 9213 5538 9279 5541
rect 11830 5538 11836 5540
rect 0 5478 5826 5538
rect 0 5448 800 5478
rect 5766 5266 5826 5478
rect 9213 5536 11836 5538
rect 9213 5480 9218 5536
rect 9274 5480 11836 5536
rect 9213 5478 11836 5480
rect 9213 5475 9279 5478
rect 11830 5476 11836 5478
rect 11900 5476 11906 5540
rect 18321 5538 18387 5541
rect 19425 5538 19491 5541
rect 29200 5538 30000 5568
rect 18321 5536 19491 5538
rect 18321 5480 18326 5536
rect 18382 5480 19430 5536
rect 19486 5480 19491 5536
rect 18321 5478 19491 5480
rect 18321 5475 18387 5478
rect 19425 5475 19491 5478
rect 27110 5478 30000 5538
rect 5944 5472 6264 5473
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 5407 6264 5408
rect 15944 5472 16264 5473
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 5407 16264 5408
rect 25944 5472 26264 5473
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 5407 26264 5408
rect 19149 5266 19215 5269
rect 5766 5264 19215 5266
rect 5766 5208 19154 5264
rect 19210 5208 19215 5264
rect 5766 5206 19215 5208
rect 19149 5203 19215 5206
rect 24853 5266 24919 5269
rect 27110 5266 27170 5478
rect 29200 5448 30000 5478
rect 24853 5264 27170 5266
rect 24853 5208 24858 5264
rect 24914 5208 27170 5264
rect 24853 5206 27170 5208
rect 24853 5203 24919 5206
rect 10944 4928 11264 4929
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 4863 11264 4864
rect 20944 4928 21264 4929
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 20944 4863 21264 4864
rect 21449 4858 21515 4861
rect 28533 4858 28599 4861
rect 21449 4856 28599 4858
rect 21449 4800 21454 4856
rect 21510 4800 28538 4856
rect 28594 4800 28599 4856
rect 21449 4798 28599 4800
rect 21449 4795 21515 4798
rect 28533 4795 28599 4798
rect 5944 4384 6264 4385
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 4319 6264 4320
rect 15944 4384 16264 4385
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 4319 16264 4320
rect 25944 4384 26264 4385
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 25944 4319 26264 4320
rect 0 4178 800 4208
rect 3969 4178 4035 4181
rect 0 4176 4035 4178
rect 0 4120 3974 4176
rect 4030 4120 4035 4176
rect 0 4118 4035 4120
rect 0 4088 800 4118
rect 3969 4115 4035 4118
rect 25313 4178 25379 4181
rect 29200 4178 30000 4208
rect 25313 4176 30000 4178
rect 25313 4120 25318 4176
rect 25374 4120 30000 4176
rect 25313 4118 30000 4120
rect 25313 4115 25379 4118
rect 29200 4088 30000 4118
rect 13445 4042 13511 4045
rect 15193 4042 15259 4045
rect 13445 4040 15259 4042
rect 13445 3984 13450 4040
rect 13506 3984 15198 4040
rect 15254 3984 15259 4040
rect 13445 3982 15259 3984
rect 13445 3979 13511 3982
rect 15193 3979 15259 3982
rect 16297 4042 16363 4045
rect 16430 4042 16436 4044
rect 16297 4040 16436 4042
rect 16297 3984 16302 4040
rect 16358 3984 16436 4040
rect 16297 3982 16436 3984
rect 16297 3979 16363 3982
rect 16430 3980 16436 3982
rect 16500 3980 16506 4044
rect 22369 4042 22435 4045
rect 23933 4042 23999 4045
rect 22369 4040 23999 4042
rect 22369 3984 22374 4040
rect 22430 3984 23938 4040
rect 23994 3984 23999 4040
rect 22369 3982 23999 3984
rect 22369 3979 22435 3982
rect 23933 3979 23999 3982
rect 10944 3840 11264 3841
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 3775 11264 3776
rect 20944 3840 21264 3841
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 20944 3775 21264 3776
rect 21398 3708 21404 3772
rect 21468 3770 21474 3772
rect 23013 3770 23079 3773
rect 21468 3768 23079 3770
rect 21468 3712 23018 3768
rect 23074 3712 23079 3768
rect 21468 3710 23079 3712
rect 21468 3708 21474 3710
rect 23013 3707 23079 3710
rect 5073 3634 5139 3637
rect 15142 3634 15148 3636
rect 5073 3632 15148 3634
rect 5073 3576 5078 3632
rect 5134 3576 15148 3632
rect 5073 3574 15148 3576
rect 5073 3571 5139 3574
rect 15142 3572 15148 3574
rect 15212 3572 15218 3636
rect 21633 3634 21699 3637
rect 15334 3632 21699 3634
rect 15334 3576 21638 3632
rect 21694 3576 21699 3632
rect 15334 3574 21699 3576
rect 0 3498 800 3528
rect 4061 3498 4127 3501
rect 0 3496 4127 3498
rect 0 3440 4066 3496
rect 4122 3440 4127 3496
rect 0 3438 4127 3440
rect 0 3408 800 3438
rect 4061 3435 4127 3438
rect 12157 3498 12223 3501
rect 12893 3498 12959 3501
rect 12157 3496 12959 3498
rect 12157 3440 12162 3496
rect 12218 3440 12898 3496
rect 12954 3440 12959 3496
rect 12157 3438 12959 3440
rect 12157 3435 12223 3438
rect 12893 3435 12959 3438
rect 6913 3362 6979 3365
rect 15334 3362 15394 3574
rect 21633 3571 21699 3574
rect 15561 3498 15627 3501
rect 29200 3498 30000 3528
rect 15561 3496 30000 3498
rect 15561 3440 15566 3496
rect 15622 3440 30000 3496
rect 15561 3438 30000 3440
rect 15561 3435 15627 3438
rect 29200 3408 30000 3438
rect 6913 3360 15394 3362
rect 6913 3304 6918 3360
rect 6974 3304 15394 3360
rect 6913 3302 15394 3304
rect 6913 3299 6979 3302
rect 5944 3296 6264 3297
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 3231 6264 3232
rect 15944 3296 16264 3297
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15944 3231 16264 3232
rect 25944 3296 26264 3297
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 25944 3231 26264 3232
rect 7373 3226 7439 3229
rect 15510 3226 15516 3228
rect 7373 3224 15516 3226
rect 7373 3168 7378 3224
rect 7434 3168 15516 3224
rect 7373 3166 15516 3168
rect 7373 3163 7439 3166
rect 15510 3164 15516 3166
rect 15580 3164 15586 3228
rect 10944 2752 11264 2753
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2687 11264 2688
rect 20944 2752 21264 2753
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2687 21264 2688
rect 12801 2682 12867 2685
rect 13997 2682 14063 2685
rect 12801 2680 14063 2682
rect 12801 2624 12806 2680
rect 12862 2624 14002 2680
rect 14058 2624 14063 2680
rect 12801 2622 14063 2624
rect 12801 2619 12867 2622
rect 13997 2619 14063 2622
rect 24894 2620 24900 2684
rect 24964 2682 24970 2684
rect 25313 2682 25379 2685
rect 24964 2680 25379 2682
rect 24964 2624 25318 2680
rect 25374 2624 25379 2680
rect 24964 2622 25379 2624
rect 24964 2620 24970 2622
rect 25313 2619 25379 2622
rect 20897 2410 20963 2413
rect 3374 2408 20963 2410
rect 3374 2352 20902 2408
rect 20958 2352 20963 2408
rect 3374 2350 20963 2352
rect 0 2138 800 2168
rect 3374 2138 3434 2350
rect 20897 2347 20963 2350
rect 5944 2208 6264 2209
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2143 6264 2144
rect 15944 2208 16264 2209
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2143 16264 2144
rect 25944 2208 26264 2209
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2143 26264 2144
rect 0 2078 3434 2138
rect 26509 2138 26575 2141
rect 29200 2138 30000 2168
rect 26509 2136 30000 2138
rect 26509 2080 26514 2136
rect 26570 2080 30000 2136
rect 26509 2078 30000 2080
rect 0 2048 800 2078
rect 26509 2075 26575 2078
rect 29200 2048 30000 2078
rect 3141 2002 3207 2005
rect 17677 2002 17743 2005
rect 3141 2000 17743 2002
rect 3141 1944 3146 2000
rect 3202 1944 17682 2000
rect 17738 1944 17743 2000
rect 3141 1942 17743 1944
rect 3141 1939 3207 1942
rect 17677 1939 17743 1942
rect 18597 2002 18663 2005
rect 28073 2002 28139 2005
rect 18597 2000 28139 2002
rect 18597 1944 18602 2000
rect 18658 1944 28078 2000
rect 28134 1944 28139 2000
rect 18597 1942 28139 1944
rect 18597 1939 18663 1942
rect 28073 1939 28139 1942
rect 2957 914 3023 917
rect 3693 914 3759 917
rect 2957 912 3759 914
rect 2957 856 2962 912
rect 3018 856 3698 912
rect 3754 856 3759 912
rect 2957 854 3759 856
rect 2957 851 3023 854
rect 3693 851 3759 854
rect 20529 914 20595 917
rect 20713 914 20779 917
rect 20529 912 20779 914
rect 20529 856 20534 912
rect 20590 856 20718 912
rect 20774 856 20779 912
rect 20529 854 20779 856
rect 20529 851 20595 854
rect 20713 851 20779 854
rect 0 778 800 808
rect 3141 778 3207 781
rect 0 776 3207 778
rect 0 720 3146 776
rect 3202 720 3207 776
rect 0 718 3207 720
rect 0 688 800 718
rect 3141 715 3207 718
rect 24945 778 25011 781
rect 29200 778 30000 808
rect 24945 776 30000 778
rect 24945 720 24950 776
rect 25006 720 30000 776
rect 24945 718 30000 720
rect 24945 715 25011 718
rect 29200 688 30000 718
rect 25497 98 25563 101
rect 29200 98 30000 128
rect 25497 96 30000 98
rect 25497 40 25502 96
rect 25558 40 30000 96
rect 25497 38 30000 40
rect 25497 35 25563 38
rect 29200 8 30000 38
<< via3 >>
rect 10952 77820 11016 77824
rect 10952 77764 10956 77820
rect 10956 77764 11012 77820
rect 11012 77764 11016 77820
rect 10952 77760 11016 77764
rect 11032 77820 11096 77824
rect 11032 77764 11036 77820
rect 11036 77764 11092 77820
rect 11092 77764 11096 77820
rect 11032 77760 11096 77764
rect 11112 77820 11176 77824
rect 11112 77764 11116 77820
rect 11116 77764 11172 77820
rect 11172 77764 11176 77820
rect 11112 77760 11176 77764
rect 11192 77820 11256 77824
rect 11192 77764 11196 77820
rect 11196 77764 11252 77820
rect 11252 77764 11256 77820
rect 11192 77760 11256 77764
rect 20952 77820 21016 77824
rect 20952 77764 20956 77820
rect 20956 77764 21012 77820
rect 21012 77764 21016 77820
rect 20952 77760 21016 77764
rect 21032 77820 21096 77824
rect 21032 77764 21036 77820
rect 21036 77764 21092 77820
rect 21092 77764 21096 77820
rect 21032 77760 21096 77764
rect 21112 77820 21176 77824
rect 21112 77764 21116 77820
rect 21116 77764 21172 77820
rect 21172 77764 21176 77820
rect 21112 77760 21176 77764
rect 21192 77820 21256 77824
rect 21192 77764 21196 77820
rect 21196 77764 21252 77820
rect 21252 77764 21256 77820
rect 21192 77760 21256 77764
rect 20668 77420 20732 77484
rect 5952 77276 6016 77280
rect 5952 77220 5956 77276
rect 5956 77220 6012 77276
rect 6012 77220 6016 77276
rect 5952 77216 6016 77220
rect 6032 77276 6096 77280
rect 6032 77220 6036 77276
rect 6036 77220 6092 77276
rect 6092 77220 6096 77276
rect 6032 77216 6096 77220
rect 6112 77276 6176 77280
rect 6112 77220 6116 77276
rect 6116 77220 6172 77276
rect 6172 77220 6176 77276
rect 6112 77216 6176 77220
rect 6192 77276 6256 77280
rect 6192 77220 6196 77276
rect 6196 77220 6252 77276
rect 6252 77220 6256 77276
rect 6192 77216 6256 77220
rect 15952 77276 16016 77280
rect 15952 77220 15956 77276
rect 15956 77220 16012 77276
rect 16012 77220 16016 77276
rect 15952 77216 16016 77220
rect 16032 77276 16096 77280
rect 16032 77220 16036 77276
rect 16036 77220 16092 77276
rect 16092 77220 16096 77276
rect 16032 77216 16096 77220
rect 16112 77276 16176 77280
rect 16112 77220 16116 77276
rect 16116 77220 16172 77276
rect 16172 77220 16176 77276
rect 16112 77216 16176 77220
rect 16192 77276 16256 77280
rect 16192 77220 16196 77276
rect 16196 77220 16252 77276
rect 16252 77220 16256 77276
rect 16192 77216 16256 77220
rect 25952 77276 26016 77280
rect 25952 77220 25956 77276
rect 25956 77220 26012 77276
rect 26012 77220 26016 77276
rect 25952 77216 26016 77220
rect 26032 77276 26096 77280
rect 26032 77220 26036 77276
rect 26036 77220 26092 77276
rect 26092 77220 26096 77276
rect 26032 77216 26096 77220
rect 26112 77276 26176 77280
rect 26112 77220 26116 77276
rect 26116 77220 26172 77276
rect 26172 77220 26176 77276
rect 26112 77216 26176 77220
rect 26192 77276 26256 77280
rect 26192 77220 26196 77276
rect 26196 77220 26252 77276
rect 26252 77220 26256 77276
rect 26192 77216 26256 77220
rect 10952 76732 11016 76736
rect 10952 76676 10956 76732
rect 10956 76676 11012 76732
rect 11012 76676 11016 76732
rect 10952 76672 11016 76676
rect 11032 76732 11096 76736
rect 11032 76676 11036 76732
rect 11036 76676 11092 76732
rect 11092 76676 11096 76732
rect 11032 76672 11096 76676
rect 11112 76732 11176 76736
rect 11112 76676 11116 76732
rect 11116 76676 11172 76732
rect 11172 76676 11176 76732
rect 11112 76672 11176 76676
rect 11192 76732 11256 76736
rect 11192 76676 11196 76732
rect 11196 76676 11252 76732
rect 11252 76676 11256 76732
rect 11192 76672 11256 76676
rect 20952 76732 21016 76736
rect 20952 76676 20956 76732
rect 20956 76676 21012 76732
rect 21012 76676 21016 76732
rect 20952 76672 21016 76676
rect 21032 76732 21096 76736
rect 21032 76676 21036 76732
rect 21036 76676 21092 76732
rect 21092 76676 21096 76732
rect 21032 76672 21096 76676
rect 21112 76732 21176 76736
rect 21112 76676 21116 76732
rect 21116 76676 21172 76732
rect 21172 76676 21176 76732
rect 21112 76672 21176 76676
rect 21192 76732 21256 76736
rect 21192 76676 21196 76732
rect 21196 76676 21252 76732
rect 21252 76676 21256 76732
rect 21192 76672 21256 76676
rect 5952 76188 6016 76192
rect 5952 76132 5956 76188
rect 5956 76132 6012 76188
rect 6012 76132 6016 76188
rect 5952 76128 6016 76132
rect 6032 76188 6096 76192
rect 6032 76132 6036 76188
rect 6036 76132 6092 76188
rect 6092 76132 6096 76188
rect 6032 76128 6096 76132
rect 6112 76188 6176 76192
rect 6112 76132 6116 76188
rect 6116 76132 6172 76188
rect 6172 76132 6176 76188
rect 6112 76128 6176 76132
rect 6192 76188 6256 76192
rect 6192 76132 6196 76188
rect 6196 76132 6252 76188
rect 6252 76132 6256 76188
rect 6192 76128 6256 76132
rect 15952 76188 16016 76192
rect 15952 76132 15956 76188
rect 15956 76132 16012 76188
rect 16012 76132 16016 76188
rect 15952 76128 16016 76132
rect 16032 76188 16096 76192
rect 16032 76132 16036 76188
rect 16036 76132 16092 76188
rect 16092 76132 16096 76188
rect 16032 76128 16096 76132
rect 16112 76188 16176 76192
rect 16112 76132 16116 76188
rect 16116 76132 16172 76188
rect 16172 76132 16176 76188
rect 16112 76128 16176 76132
rect 16192 76188 16256 76192
rect 16192 76132 16196 76188
rect 16196 76132 16252 76188
rect 16252 76132 16256 76188
rect 16192 76128 16256 76132
rect 25952 76188 26016 76192
rect 25952 76132 25956 76188
rect 25956 76132 26012 76188
rect 26012 76132 26016 76188
rect 25952 76128 26016 76132
rect 26032 76188 26096 76192
rect 26032 76132 26036 76188
rect 26036 76132 26092 76188
rect 26092 76132 26096 76188
rect 26032 76128 26096 76132
rect 26112 76188 26176 76192
rect 26112 76132 26116 76188
rect 26116 76132 26172 76188
rect 26172 76132 26176 76188
rect 26112 76128 26176 76132
rect 26192 76188 26256 76192
rect 26192 76132 26196 76188
rect 26196 76132 26252 76188
rect 26252 76132 26256 76188
rect 26192 76128 26256 76132
rect 11836 75652 11900 75716
rect 10952 75644 11016 75648
rect 10952 75588 10956 75644
rect 10956 75588 11012 75644
rect 11012 75588 11016 75644
rect 10952 75584 11016 75588
rect 11032 75644 11096 75648
rect 11032 75588 11036 75644
rect 11036 75588 11092 75644
rect 11092 75588 11096 75644
rect 11032 75584 11096 75588
rect 11112 75644 11176 75648
rect 11112 75588 11116 75644
rect 11116 75588 11172 75644
rect 11172 75588 11176 75644
rect 11112 75584 11176 75588
rect 11192 75644 11256 75648
rect 11192 75588 11196 75644
rect 11196 75588 11252 75644
rect 11252 75588 11256 75644
rect 11192 75584 11256 75588
rect 20952 75644 21016 75648
rect 20952 75588 20956 75644
rect 20956 75588 21012 75644
rect 21012 75588 21016 75644
rect 20952 75584 21016 75588
rect 21032 75644 21096 75648
rect 21032 75588 21036 75644
rect 21036 75588 21092 75644
rect 21092 75588 21096 75644
rect 21032 75584 21096 75588
rect 21112 75644 21176 75648
rect 21112 75588 21116 75644
rect 21116 75588 21172 75644
rect 21172 75588 21176 75644
rect 21112 75584 21176 75588
rect 21192 75644 21256 75648
rect 21192 75588 21196 75644
rect 21196 75588 21252 75644
rect 21252 75588 21256 75644
rect 21192 75584 21256 75588
rect 5952 75100 6016 75104
rect 5952 75044 5956 75100
rect 5956 75044 6012 75100
rect 6012 75044 6016 75100
rect 5952 75040 6016 75044
rect 6032 75100 6096 75104
rect 6032 75044 6036 75100
rect 6036 75044 6092 75100
rect 6092 75044 6096 75100
rect 6032 75040 6096 75044
rect 6112 75100 6176 75104
rect 6112 75044 6116 75100
rect 6116 75044 6172 75100
rect 6172 75044 6176 75100
rect 6112 75040 6176 75044
rect 6192 75100 6256 75104
rect 6192 75044 6196 75100
rect 6196 75044 6252 75100
rect 6252 75044 6256 75100
rect 6192 75040 6256 75044
rect 15952 75100 16016 75104
rect 15952 75044 15956 75100
rect 15956 75044 16012 75100
rect 16012 75044 16016 75100
rect 15952 75040 16016 75044
rect 16032 75100 16096 75104
rect 16032 75044 16036 75100
rect 16036 75044 16092 75100
rect 16092 75044 16096 75100
rect 16032 75040 16096 75044
rect 16112 75100 16176 75104
rect 16112 75044 16116 75100
rect 16116 75044 16172 75100
rect 16172 75044 16176 75100
rect 16112 75040 16176 75044
rect 16192 75100 16256 75104
rect 16192 75044 16196 75100
rect 16196 75044 16252 75100
rect 16252 75044 16256 75100
rect 16192 75040 16256 75044
rect 25952 75100 26016 75104
rect 25952 75044 25956 75100
rect 25956 75044 26012 75100
rect 26012 75044 26016 75100
rect 25952 75040 26016 75044
rect 26032 75100 26096 75104
rect 26032 75044 26036 75100
rect 26036 75044 26092 75100
rect 26092 75044 26096 75100
rect 26032 75040 26096 75044
rect 26112 75100 26176 75104
rect 26112 75044 26116 75100
rect 26116 75044 26172 75100
rect 26172 75044 26176 75100
rect 26112 75040 26176 75044
rect 26192 75100 26256 75104
rect 26192 75044 26196 75100
rect 26196 75044 26252 75100
rect 26252 75044 26256 75100
rect 26192 75040 26256 75044
rect 9996 74700 10060 74764
rect 25084 74564 25148 74628
rect 10952 74556 11016 74560
rect 10952 74500 10956 74556
rect 10956 74500 11012 74556
rect 11012 74500 11016 74556
rect 10952 74496 11016 74500
rect 11032 74556 11096 74560
rect 11032 74500 11036 74556
rect 11036 74500 11092 74556
rect 11092 74500 11096 74556
rect 11032 74496 11096 74500
rect 11112 74556 11176 74560
rect 11112 74500 11116 74556
rect 11116 74500 11172 74556
rect 11172 74500 11176 74556
rect 11112 74496 11176 74500
rect 11192 74556 11256 74560
rect 11192 74500 11196 74556
rect 11196 74500 11252 74556
rect 11252 74500 11256 74556
rect 11192 74496 11256 74500
rect 20952 74556 21016 74560
rect 20952 74500 20956 74556
rect 20956 74500 21012 74556
rect 21012 74500 21016 74556
rect 20952 74496 21016 74500
rect 21032 74556 21096 74560
rect 21032 74500 21036 74556
rect 21036 74500 21092 74556
rect 21092 74500 21096 74556
rect 21032 74496 21096 74500
rect 21112 74556 21176 74560
rect 21112 74500 21116 74556
rect 21116 74500 21172 74556
rect 21172 74500 21176 74556
rect 21112 74496 21176 74500
rect 21192 74556 21256 74560
rect 21192 74500 21196 74556
rect 21196 74500 21252 74556
rect 21252 74500 21256 74556
rect 21192 74496 21256 74500
rect 24900 74428 24964 74492
rect 5952 74012 6016 74016
rect 5952 73956 5956 74012
rect 5956 73956 6012 74012
rect 6012 73956 6016 74012
rect 5952 73952 6016 73956
rect 6032 74012 6096 74016
rect 6032 73956 6036 74012
rect 6036 73956 6092 74012
rect 6092 73956 6096 74012
rect 6032 73952 6096 73956
rect 6112 74012 6176 74016
rect 6112 73956 6116 74012
rect 6116 73956 6172 74012
rect 6172 73956 6176 74012
rect 6112 73952 6176 73956
rect 6192 74012 6256 74016
rect 6192 73956 6196 74012
rect 6196 73956 6252 74012
rect 6252 73956 6256 74012
rect 6192 73952 6256 73956
rect 15952 74012 16016 74016
rect 15952 73956 15956 74012
rect 15956 73956 16012 74012
rect 16012 73956 16016 74012
rect 15952 73952 16016 73956
rect 16032 74012 16096 74016
rect 16032 73956 16036 74012
rect 16036 73956 16092 74012
rect 16092 73956 16096 74012
rect 16032 73952 16096 73956
rect 16112 74012 16176 74016
rect 16112 73956 16116 74012
rect 16116 73956 16172 74012
rect 16172 73956 16176 74012
rect 16112 73952 16176 73956
rect 16192 74012 16256 74016
rect 16192 73956 16196 74012
rect 16196 73956 16252 74012
rect 16252 73956 16256 74012
rect 16192 73952 16256 73956
rect 25952 74012 26016 74016
rect 25952 73956 25956 74012
rect 25956 73956 26012 74012
rect 26012 73956 26016 74012
rect 25952 73952 26016 73956
rect 26032 74012 26096 74016
rect 26032 73956 26036 74012
rect 26036 73956 26092 74012
rect 26092 73956 26096 74012
rect 26032 73952 26096 73956
rect 26112 74012 26176 74016
rect 26112 73956 26116 74012
rect 26116 73956 26172 74012
rect 26172 73956 26176 74012
rect 26112 73952 26176 73956
rect 26192 74012 26256 74016
rect 26192 73956 26196 74012
rect 26196 73956 26252 74012
rect 26252 73956 26256 74012
rect 26192 73952 26256 73956
rect 10952 73468 11016 73472
rect 10952 73412 10956 73468
rect 10956 73412 11012 73468
rect 11012 73412 11016 73468
rect 10952 73408 11016 73412
rect 11032 73468 11096 73472
rect 11032 73412 11036 73468
rect 11036 73412 11092 73468
rect 11092 73412 11096 73468
rect 11032 73408 11096 73412
rect 11112 73468 11176 73472
rect 11112 73412 11116 73468
rect 11116 73412 11172 73468
rect 11172 73412 11176 73468
rect 11112 73408 11176 73412
rect 11192 73468 11256 73472
rect 11192 73412 11196 73468
rect 11196 73412 11252 73468
rect 11252 73412 11256 73468
rect 11192 73408 11256 73412
rect 20952 73468 21016 73472
rect 20952 73412 20956 73468
rect 20956 73412 21012 73468
rect 21012 73412 21016 73468
rect 20952 73408 21016 73412
rect 21032 73468 21096 73472
rect 21032 73412 21036 73468
rect 21036 73412 21092 73468
rect 21092 73412 21096 73468
rect 21032 73408 21096 73412
rect 21112 73468 21176 73472
rect 21112 73412 21116 73468
rect 21116 73412 21172 73468
rect 21172 73412 21176 73468
rect 21112 73408 21176 73412
rect 21192 73468 21256 73472
rect 21192 73412 21196 73468
rect 21196 73412 21252 73468
rect 21252 73412 21256 73468
rect 21192 73408 21256 73412
rect 5952 72924 6016 72928
rect 5952 72868 5956 72924
rect 5956 72868 6012 72924
rect 6012 72868 6016 72924
rect 5952 72864 6016 72868
rect 6032 72924 6096 72928
rect 6032 72868 6036 72924
rect 6036 72868 6092 72924
rect 6092 72868 6096 72924
rect 6032 72864 6096 72868
rect 6112 72924 6176 72928
rect 6112 72868 6116 72924
rect 6116 72868 6172 72924
rect 6172 72868 6176 72924
rect 6112 72864 6176 72868
rect 6192 72924 6256 72928
rect 6192 72868 6196 72924
rect 6196 72868 6252 72924
rect 6252 72868 6256 72924
rect 6192 72864 6256 72868
rect 15952 72924 16016 72928
rect 15952 72868 15956 72924
rect 15956 72868 16012 72924
rect 16012 72868 16016 72924
rect 15952 72864 16016 72868
rect 16032 72924 16096 72928
rect 16032 72868 16036 72924
rect 16036 72868 16092 72924
rect 16092 72868 16096 72924
rect 16032 72864 16096 72868
rect 16112 72924 16176 72928
rect 16112 72868 16116 72924
rect 16116 72868 16172 72924
rect 16172 72868 16176 72924
rect 16112 72864 16176 72868
rect 16192 72924 16256 72928
rect 16192 72868 16196 72924
rect 16196 72868 16252 72924
rect 16252 72868 16256 72924
rect 16192 72864 16256 72868
rect 25952 72924 26016 72928
rect 25952 72868 25956 72924
rect 25956 72868 26012 72924
rect 26012 72868 26016 72924
rect 25952 72864 26016 72868
rect 26032 72924 26096 72928
rect 26032 72868 26036 72924
rect 26036 72868 26092 72924
rect 26092 72868 26096 72924
rect 26032 72864 26096 72868
rect 26112 72924 26176 72928
rect 26112 72868 26116 72924
rect 26116 72868 26172 72924
rect 26172 72868 26176 72924
rect 26112 72864 26176 72868
rect 26192 72924 26256 72928
rect 26192 72868 26196 72924
rect 26196 72868 26252 72924
rect 26252 72868 26256 72924
rect 26192 72864 26256 72868
rect 10952 72380 11016 72384
rect 10952 72324 10956 72380
rect 10956 72324 11012 72380
rect 11012 72324 11016 72380
rect 10952 72320 11016 72324
rect 11032 72380 11096 72384
rect 11032 72324 11036 72380
rect 11036 72324 11092 72380
rect 11092 72324 11096 72380
rect 11032 72320 11096 72324
rect 11112 72380 11176 72384
rect 11112 72324 11116 72380
rect 11116 72324 11172 72380
rect 11172 72324 11176 72380
rect 11112 72320 11176 72324
rect 11192 72380 11256 72384
rect 11192 72324 11196 72380
rect 11196 72324 11252 72380
rect 11252 72324 11256 72380
rect 11192 72320 11256 72324
rect 20952 72380 21016 72384
rect 20952 72324 20956 72380
rect 20956 72324 21012 72380
rect 21012 72324 21016 72380
rect 20952 72320 21016 72324
rect 21032 72380 21096 72384
rect 21032 72324 21036 72380
rect 21036 72324 21092 72380
rect 21092 72324 21096 72380
rect 21032 72320 21096 72324
rect 21112 72380 21176 72384
rect 21112 72324 21116 72380
rect 21116 72324 21172 72380
rect 21172 72324 21176 72380
rect 21112 72320 21176 72324
rect 21192 72380 21256 72384
rect 21192 72324 21196 72380
rect 21196 72324 21252 72380
rect 21252 72324 21256 72380
rect 21192 72320 21256 72324
rect 5952 71836 6016 71840
rect 5952 71780 5956 71836
rect 5956 71780 6012 71836
rect 6012 71780 6016 71836
rect 5952 71776 6016 71780
rect 6032 71836 6096 71840
rect 6032 71780 6036 71836
rect 6036 71780 6092 71836
rect 6092 71780 6096 71836
rect 6032 71776 6096 71780
rect 6112 71836 6176 71840
rect 6112 71780 6116 71836
rect 6116 71780 6172 71836
rect 6172 71780 6176 71836
rect 6112 71776 6176 71780
rect 6192 71836 6256 71840
rect 6192 71780 6196 71836
rect 6196 71780 6252 71836
rect 6252 71780 6256 71836
rect 6192 71776 6256 71780
rect 15952 71836 16016 71840
rect 15952 71780 15956 71836
rect 15956 71780 16012 71836
rect 16012 71780 16016 71836
rect 15952 71776 16016 71780
rect 16032 71836 16096 71840
rect 16032 71780 16036 71836
rect 16036 71780 16092 71836
rect 16092 71780 16096 71836
rect 16032 71776 16096 71780
rect 16112 71836 16176 71840
rect 16112 71780 16116 71836
rect 16116 71780 16172 71836
rect 16172 71780 16176 71836
rect 16112 71776 16176 71780
rect 16192 71836 16256 71840
rect 16192 71780 16196 71836
rect 16196 71780 16252 71836
rect 16252 71780 16256 71836
rect 16192 71776 16256 71780
rect 25952 71836 26016 71840
rect 25952 71780 25956 71836
rect 25956 71780 26012 71836
rect 26012 71780 26016 71836
rect 25952 71776 26016 71780
rect 26032 71836 26096 71840
rect 26032 71780 26036 71836
rect 26036 71780 26092 71836
rect 26092 71780 26096 71836
rect 26032 71776 26096 71780
rect 26112 71836 26176 71840
rect 26112 71780 26116 71836
rect 26116 71780 26172 71836
rect 26172 71780 26176 71836
rect 26112 71776 26176 71780
rect 26192 71836 26256 71840
rect 26192 71780 26196 71836
rect 26196 71780 26252 71836
rect 26252 71780 26256 71836
rect 26192 71776 26256 71780
rect 10952 71292 11016 71296
rect 10952 71236 10956 71292
rect 10956 71236 11012 71292
rect 11012 71236 11016 71292
rect 10952 71232 11016 71236
rect 11032 71292 11096 71296
rect 11032 71236 11036 71292
rect 11036 71236 11092 71292
rect 11092 71236 11096 71292
rect 11032 71232 11096 71236
rect 11112 71292 11176 71296
rect 11112 71236 11116 71292
rect 11116 71236 11172 71292
rect 11172 71236 11176 71292
rect 11112 71232 11176 71236
rect 11192 71292 11256 71296
rect 11192 71236 11196 71292
rect 11196 71236 11252 71292
rect 11252 71236 11256 71292
rect 11192 71232 11256 71236
rect 20952 71292 21016 71296
rect 20952 71236 20956 71292
rect 20956 71236 21012 71292
rect 21012 71236 21016 71292
rect 20952 71232 21016 71236
rect 21032 71292 21096 71296
rect 21032 71236 21036 71292
rect 21036 71236 21092 71292
rect 21092 71236 21096 71292
rect 21032 71232 21096 71236
rect 21112 71292 21176 71296
rect 21112 71236 21116 71292
rect 21116 71236 21172 71292
rect 21172 71236 21176 71292
rect 21112 71232 21176 71236
rect 21192 71292 21256 71296
rect 21192 71236 21196 71292
rect 21196 71236 21252 71292
rect 21252 71236 21256 71292
rect 21192 71232 21256 71236
rect 5952 70748 6016 70752
rect 5952 70692 5956 70748
rect 5956 70692 6012 70748
rect 6012 70692 6016 70748
rect 5952 70688 6016 70692
rect 6032 70748 6096 70752
rect 6032 70692 6036 70748
rect 6036 70692 6092 70748
rect 6092 70692 6096 70748
rect 6032 70688 6096 70692
rect 6112 70748 6176 70752
rect 6112 70692 6116 70748
rect 6116 70692 6172 70748
rect 6172 70692 6176 70748
rect 6112 70688 6176 70692
rect 6192 70748 6256 70752
rect 6192 70692 6196 70748
rect 6196 70692 6252 70748
rect 6252 70692 6256 70748
rect 6192 70688 6256 70692
rect 15952 70748 16016 70752
rect 15952 70692 15956 70748
rect 15956 70692 16012 70748
rect 16012 70692 16016 70748
rect 15952 70688 16016 70692
rect 16032 70748 16096 70752
rect 16032 70692 16036 70748
rect 16036 70692 16092 70748
rect 16092 70692 16096 70748
rect 16032 70688 16096 70692
rect 16112 70748 16176 70752
rect 16112 70692 16116 70748
rect 16116 70692 16172 70748
rect 16172 70692 16176 70748
rect 16112 70688 16176 70692
rect 16192 70748 16256 70752
rect 16192 70692 16196 70748
rect 16196 70692 16252 70748
rect 16252 70692 16256 70748
rect 16192 70688 16256 70692
rect 25952 70748 26016 70752
rect 25952 70692 25956 70748
rect 25956 70692 26012 70748
rect 26012 70692 26016 70748
rect 25952 70688 26016 70692
rect 26032 70748 26096 70752
rect 26032 70692 26036 70748
rect 26036 70692 26092 70748
rect 26092 70692 26096 70748
rect 26032 70688 26096 70692
rect 26112 70748 26176 70752
rect 26112 70692 26116 70748
rect 26116 70692 26172 70748
rect 26172 70692 26176 70748
rect 26112 70688 26176 70692
rect 26192 70748 26256 70752
rect 26192 70692 26196 70748
rect 26196 70692 26252 70748
rect 26252 70692 26256 70748
rect 26192 70688 26256 70692
rect 10952 70204 11016 70208
rect 10952 70148 10956 70204
rect 10956 70148 11012 70204
rect 11012 70148 11016 70204
rect 10952 70144 11016 70148
rect 11032 70204 11096 70208
rect 11032 70148 11036 70204
rect 11036 70148 11092 70204
rect 11092 70148 11096 70204
rect 11032 70144 11096 70148
rect 11112 70204 11176 70208
rect 11112 70148 11116 70204
rect 11116 70148 11172 70204
rect 11172 70148 11176 70204
rect 11112 70144 11176 70148
rect 11192 70204 11256 70208
rect 11192 70148 11196 70204
rect 11196 70148 11252 70204
rect 11252 70148 11256 70204
rect 11192 70144 11256 70148
rect 20952 70204 21016 70208
rect 20952 70148 20956 70204
rect 20956 70148 21012 70204
rect 21012 70148 21016 70204
rect 20952 70144 21016 70148
rect 21032 70204 21096 70208
rect 21032 70148 21036 70204
rect 21036 70148 21092 70204
rect 21092 70148 21096 70204
rect 21032 70144 21096 70148
rect 21112 70204 21176 70208
rect 21112 70148 21116 70204
rect 21116 70148 21172 70204
rect 21172 70148 21176 70204
rect 21112 70144 21176 70148
rect 21192 70204 21256 70208
rect 21192 70148 21196 70204
rect 21196 70148 21252 70204
rect 21252 70148 21256 70204
rect 21192 70144 21256 70148
rect 5952 69660 6016 69664
rect 5952 69604 5956 69660
rect 5956 69604 6012 69660
rect 6012 69604 6016 69660
rect 5952 69600 6016 69604
rect 6032 69660 6096 69664
rect 6032 69604 6036 69660
rect 6036 69604 6092 69660
rect 6092 69604 6096 69660
rect 6032 69600 6096 69604
rect 6112 69660 6176 69664
rect 6112 69604 6116 69660
rect 6116 69604 6172 69660
rect 6172 69604 6176 69660
rect 6112 69600 6176 69604
rect 6192 69660 6256 69664
rect 6192 69604 6196 69660
rect 6196 69604 6252 69660
rect 6252 69604 6256 69660
rect 6192 69600 6256 69604
rect 15952 69660 16016 69664
rect 15952 69604 15956 69660
rect 15956 69604 16012 69660
rect 16012 69604 16016 69660
rect 15952 69600 16016 69604
rect 16032 69660 16096 69664
rect 16032 69604 16036 69660
rect 16036 69604 16092 69660
rect 16092 69604 16096 69660
rect 16032 69600 16096 69604
rect 16112 69660 16176 69664
rect 16112 69604 16116 69660
rect 16116 69604 16172 69660
rect 16172 69604 16176 69660
rect 16112 69600 16176 69604
rect 16192 69660 16256 69664
rect 16192 69604 16196 69660
rect 16196 69604 16252 69660
rect 16252 69604 16256 69660
rect 16192 69600 16256 69604
rect 25952 69660 26016 69664
rect 25952 69604 25956 69660
rect 25956 69604 26012 69660
rect 26012 69604 26016 69660
rect 25952 69600 26016 69604
rect 26032 69660 26096 69664
rect 26032 69604 26036 69660
rect 26036 69604 26092 69660
rect 26092 69604 26096 69660
rect 26032 69600 26096 69604
rect 26112 69660 26176 69664
rect 26112 69604 26116 69660
rect 26116 69604 26172 69660
rect 26172 69604 26176 69660
rect 26112 69600 26176 69604
rect 26192 69660 26256 69664
rect 26192 69604 26196 69660
rect 26196 69604 26252 69660
rect 26252 69604 26256 69660
rect 26192 69600 26256 69604
rect 17172 69260 17236 69324
rect 10952 69116 11016 69120
rect 10952 69060 10956 69116
rect 10956 69060 11012 69116
rect 11012 69060 11016 69116
rect 10952 69056 11016 69060
rect 11032 69116 11096 69120
rect 11032 69060 11036 69116
rect 11036 69060 11092 69116
rect 11092 69060 11096 69116
rect 11032 69056 11096 69060
rect 11112 69116 11176 69120
rect 11112 69060 11116 69116
rect 11116 69060 11172 69116
rect 11172 69060 11176 69116
rect 11112 69056 11176 69060
rect 11192 69116 11256 69120
rect 11192 69060 11196 69116
rect 11196 69060 11252 69116
rect 11252 69060 11256 69116
rect 11192 69056 11256 69060
rect 20952 69116 21016 69120
rect 20952 69060 20956 69116
rect 20956 69060 21012 69116
rect 21012 69060 21016 69116
rect 20952 69056 21016 69060
rect 21032 69116 21096 69120
rect 21032 69060 21036 69116
rect 21036 69060 21092 69116
rect 21092 69060 21096 69116
rect 21032 69056 21096 69060
rect 21112 69116 21176 69120
rect 21112 69060 21116 69116
rect 21116 69060 21172 69116
rect 21172 69060 21176 69116
rect 21112 69056 21176 69060
rect 21192 69116 21256 69120
rect 21192 69060 21196 69116
rect 21196 69060 21252 69116
rect 21252 69060 21256 69116
rect 21192 69056 21256 69060
rect 25636 68716 25700 68780
rect 5952 68572 6016 68576
rect 5952 68516 5956 68572
rect 5956 68516 6012 68572
rect 6012 68516 6016 68572
rect 5952 68512 6016 68516
rect 6032 68572 6096 68576
rect 6032 68516 6036 68572
rect 6036 68516 6092 68572
rect 6092 68516 6096 68572
rect 6032 68512 6096 68516
rect 6112 68572 6176 68576
rect 6112 68516 6116 68572
rect 6116 68516 6172 68572
rect 6172 68516 6176 68572
rect 6112 68512 6176 68516
rect 6192 68572 6256 68576
rect 6192 68516 6196 68572
rect 6196 68516 6252 68572
rect 6252 68516 6256 68572
rect 6192 68512 6256 68516
rect 15952 68572 16016 68576
rect 15952 68516 15956 68572
rect 15956 68516 16012 68572
rect 16012 68516 16016 68572
rect 15952 68512 16016 68516
rect 16032 68572 16096 68576
rect 16032 68516 16036 68572
rect 16036 68516 16092 68572
rect 16092 68516 16096 68572
rect 16032 68512 16096 68516
rect 16112 68572 16176 68576
rect 16112 68516 16116 68572
rect 16116 68516 16172 68572
rect 16172 68516 16176 68572
rect 16112 68512 16176 68516
rect 16192 68572 16256 68576
rect 16192 68516 16196 68572
rect 16196 68516 16252 68572
rect 16252 68516 16256 68572
rect 16192 68512 16256 68516
rect 25952 68572 26016 68576
rect 25952 68516 25956 68572
rect 25956 68516 26012 68572
rect 26012 68516 26016 68572
rect 25952 68512 26016 68516
rect 26032 68572 26096 68576
rect 26032 68516 26036 68572
rect 26036 68516 26092 68572
rect 26092 68516 26096 68572
rect 26032 68512 26096 68516
rect 26112 68572 26176 68576
rect 26112 68516 26116 68572
rect 26116 68516 26172 68572
rect 26172 68516 26176 68572
rect 26112 68512 26176 68516
rect 26192 68572 26256 68576
rect 26192 68516 26196 68572
rect 26196 68516 26252 68572
rect 26252 68516 26256 68572
rect 26192 68512 26256 68516
rect 10952 68028 11016 68032
rect 10952 67972 10956 68028
rect 10956 67972 11012 68028
rect 11012 67972 11016 68028
rect 10952 67968 11016 67972
rect 11032 68028 11096 68032
rect 11032 67972 11036 68028
rect 11036 67972 11092 68028
rect 11092 67972 11096 68028
rect 11032 67968 11096 67972
rect 11112 68028 11176 68032
rect 11112 67972 11116 68028
rect 11116 67972 11172 68028
rect 11172 67972 11176 68028
rect 11112 67968 11176 67972
rect 11192 68028 11256 68032
rect 11192 67972 11196 68028
rect 11196 67972 11252 68028
rect 11252 67972 11256 68028
rect 11192 67968 11256 67972
rect 20952 68028 21016 68032
rect 20952 67972 20956 68028
rect 20956 67972 21012 68028
rect 21012 67972 21016 68028
rect 20952 67968 21016 67972
rect 21032 68028 21096 68032
rect 21032 67972 21036 68028
rect 21036 67972 21092 68028
rect 21092 67972 21096 68028
rect 21032 67968 21096 67972
rect 21112 68028 21176 68032
rect 21112 67972 21116 68028
rect 21116 67972 21172 68028
rect 21172 67972 21176 68028
rect 21112 67968 21176 67972
rect 21192 68028 21256 68032
rect 21192 67972 21196 68028
rect 21196 67972 21252 68028
rect 21252 67972 21256 68028
rect 21192 67968 21256 67972
rect 5952 67484 6016 67488
rect 5952 67428 5956 67484
rect 5956 67428 6012 67484
rect 6012 67428 6016 67484
rect 5952 67424 6016 67428
rect 6032 67484 6096 67488
rect 6032 67428 6036 67484
rect 6036 67428 6092 67484
rect 6092 67428 6096 67484
rect 6032 67424 6096 67428
rect 6112 67484 6176 67488
rect 6112 67428 6116 67484
rect 6116 67428 6172 67484
rect 6172 67428 6176 67484
rect 6112 67424 6176 67428
rect 6192 67484 6256 67488
rect 6192 67428 6196 67484
rect 6196 67428 6252 67484
rect 6252 67428 6256 67484
rect 6192 67424 6256 67428
rect 15952 67484 16016 67488
rect 15952 67428 15956 67484
rect 15956 67428 16012 67484
rect 16012 67428 16016 67484
rect 15952 67424 16016 67428
rect 16032 67484 16096 67488
rect 16032 67428 16036 67484
rect 16036 67428 16092 67484
rect 16092 67428 16096 67484
rect 16032 67424 16096 67428
rect 16112 67484 16176 67488
rect 16112 67428 16116 67484
rect 16116 67428 16172 67484
rect 16172 67428 16176 67484
rect 16112 67424 16176 67428
rect 16192 67484 16256 67488
rect 16192 67428 16196 67484
rect 16196 67428 16252 67484
rect 16252 67428 16256 67484
rect 16192 67424 16256 67428
rect 25952 67484 26016 67488
rect 25952 67428 25956 67484
rect 25956 67428 26012 67484
rect 26012 67428 26016 67484
rect 25952 67424 26016 67428
rect 26032 67484 26096 67488
rect 26032 67428 26036 67484
rect 26036 67428 26092 67484
rect 26092 67428 26096 67484
rect 26032 67424 26096 67428
rect 26112 67484 26176 67488
rect 26112 67428 26116 67484
rect 26116 67428 26172 67484
rect 26172 67428 26176 67484
rect 26112 67424 26176 67428
rect 26192 67484 26256 67488
rect 26192 67428 26196 67484
rect 26196 67428 26252 67484
rect 26252 67428 26256 67484
rect 26192 67424 26256 67428
rect 10952 66940 11016 66944
rect 10952 66884 10956 66940
rect 10956 66884 11012 66940
rect 11012 66884 11016 66940
rect 10952 66880 11016 66884
rect 11032 66940 11096 66944
rect 11032 66884 11036 66940
rect 11036 66884 11092 66940
rect 11092 66884 11096 66940
rect 11032 66880 11096 66884
rect 11112 66940 11176 66944
rect 11112 66884 11116 66940
rect 11116 66884 11172 66940
rect 11172 66884 11176 66940
rect 11112 66880 11176 66884
rect 11192 66940 11256 66944
rect 11192 66884 11196 66940
rect 11196 66884 11252 66940
rect 11252 66884 11256 66940
rect 11192 66880 11256 66884
rect 20952 66940 21016 66944
rect 20952 66884 20956 66940
rect 20956 66884 21012 66940
rect 21012 66884 21016 66940
rect 20952 66880 21016 66884
rect 21032 66940 21096 66944
rect 21032 66884 21036 66940
rect 21036 66884 21092 66940
rect 21092 66884 21096 66940
rect 21032 66880 21096 66884
rect 21112 66940 21176 66944
rect 21112 66884 21116 66940
rect 21116 66884 21172 66940
rect 21172 66884 21176 66940
rect 21112 66880 21176 66884
rect 21192 66940 21256 66944
rect 21192 66884 21196 66940
rect 21196 66884 21252 66940
rect 21252 66884 21256 66940
rect 21192 66880 21256 66884
rect 5952 66396 6016 66400
rect 5952 66340 5956 66396
rect 5956 66340 6012 66396
rect 6012 66340 6016 66396
rect 5952 66336 6016 66340
rect 6032 66396 6096 66400
rect 6032 66340 6036 66396
rect 6036 66340 6092 66396
rect 6092 66340 6096 66396
rect 6032 66336 6096 66340
rect 6112 66396 6176 66400
rect 6112 66340 6116 66396
rect 6116 66340 6172 66396
rect 6172 66340 6176 66396
rect 6112 66336 6176 66340
rect 6192 66396 6256 66400
rect 6192 66340 6196 66396
rect 6196 66340 6252 66396
rect 6252 66340 6256 66396
rect 6192 66336 6256 66340
rect 15952 66396 16016 66400
rect 15952 66340 15956 66396
rect 15956 66340 16012 66396
rect 16012 66340 16016 66396
rect 15952 66336 16016 66340
rect 16032 66396 16096 66400
rect 16032 66340 16036 66396
rect 16036 66340 16092 66396
rect 16092 66340 16096 66396
rect 16032 66336 16096 66340
rect 16112 66396 16176 66400
rect 16112 66340 16116 66396
rect 16116 66340 16172 66396
rect 16172 66340 16176 66396
rect 16112 66336 16176 66340
rect 16192 66396 16256 66400
rect 16192 66340 16196 66396
rect 16196 66340 16252 66396
rect 16252 66340 16256 66396
rect 16192 66336 16256 66340
rect 25952 66396 26016 66400
rect 25952 66340 25956 66396
rect 25956 66340 26012 66396
rect 26012 66340 26016 66396
rect 25952 66336 26016 66340
rect 26032 66396 26096 66400
rect 26032 66340 26036 66396
rect 26036 66340 26092 66396
rect 26092 66340 26096 66396
rect 26032 66336 26096 66340
rect 26112 66396 26176 66400
rect 26112 66340 26116 66396
rect 26116 66340 26172 66396
rect 26172 66340 26176 66396
rect 26112 66336 26176 66340
rect 26192 66396 26256 66400
rect 26192 66340 26196 66396
rect 26196 66340 26252 66396
rect 26252 66340 26256 66396
rect 26192 66336 26256 66340
rect 27844 66132 27908 66196
rect 10952 65852 11016 65856
rect 10952 65796 10956 65852
rect 10956 65796 11012 65852
rect 11012 65796 11016 65852
rect 10952 65792 11016 65796
rect 11032 65852 11096 65856
rect 11032 65796 11036 65852
rect 11036 65796 11092 65852
rect 11092 65796 11096 65852
rect 11032 65792 11096 65796
rect 11112 65852 11176 65856
rect 11112 65796 11116 65852
rect 11116 65796 11172 65852
rect 11172 65796 11176 65852
rect 11112 65792 11176 65796
rect 11192 65852 11256 65856
rect 11192 65796 11196 65852
rect 11196 65796 11252 65852
rect 11252 65796 11256 65852
rect 11192 65792 11256 65796
rect 20952 65852 21016 65856
rect 20952 65796 20956 65852
rect 20956 65796 21012 65852
rect 21012 65796 21016 65852
rect 20952 65792 21016 65796
rect 21032 65852 21096 65856
rect 21032 65796 21036 65852
rect 21036 65796 21092 65852
rect 21092 65796 21096 65852
rect 21032 65792 21096 65796
rect 21112 65852 21176 65856
rect 21112 65796 21116 65852
rect 21116 65796 21172 65852
rect 21172 65796 21176 65852
rect 21112 65792 21176 65796
rect 21192 65852 21256 65856
rect 21192 65796 21196 65852
rect 21196 65796 21252 65852
rect 21252 65796 21256 65852
rect 21192 65792 21256 65796
rect 21956 65452 22020 65516
rect 5952 65308 6016 65312
rect 5952 65252 5956 65308
rect 5956 65252 6012 65308
rect 6012 65252 6016 65308
rect 5952 65248 6016 65252
rect 6032 65308 6096 65312
rect 6032 65252 6036 65308
rect 6036 65252 6092 65308
rect 6092 65252 6096 65308
rect 6032 65248 6096 65252
rect 6112 65308 6176 65312
rect 6112 65252 6116 65308
rect 6116 65252 6172 65308
rect 6172 65252 6176 65308
rect 6112 65248 6176 65252
rect 6192 65308 6256 65312
rect 6192 65252 6196 65308
rect 6196 65252 6252 65308
rect 6252 65252 6256 65308
rect 6192 65248 6256 65252
rect 15952 65308 16016 65312
rect 15952 65252 15956 65308
rect 15956 65252 16012 65308
rect 16012 65252 16016 65308
rect 15952 65248 16016 65252
rect 16032 65308 16096 65312
rect 16032 65252 16036 65308
rect 16036 65252 16092 65308
rect 16092 65252 16096 65308
rect 16032 65248 16096 65252
rect 16112 65308 16176 65312
rect 16112 65252 16116 65308
rect 16116 65252 16172 65308
rect 16172 65252 16176 65308
rect 16112 65248 16176 65252
rect 16192 65308 16256 65312
rect 16192 65252 16196 65308
rect 16196 65252 16252 65308
rect 16252 65252 16256 65308
rect 16192 65248 16256 65252
rect 25952 65308 26016 65312
rect 25952 65252 25956 65308
rect 25956 65252 26012 65308
rect 26012 65252 26016 65308
rect 25952 65248 26016 65252
rect 26032 65308 26096 65312
rect 26032 65252 26036 65308
rect 26036 65252 26092 65308
rect 26092 65252 26096 65308
rect 26032 65248 26096 65252
rect 26112 65308 26176 65312
rect 26112 65252 26116 65308
rect 26116 65252 26172 65308
rect 26172 65252 26176 65308
rect 26112 65248 26176 65252
rect 26192 65308 26256 65312
rect 26192 65252 26196 65308
rect 26196 65252 26252 65308
rect 26252 65252 26256 65308
rect 26192 65248 26256 65252
rect 10952 64764 11016 64768
rect 10952 64708 10956 64764
rect 10956 64708 11012 64764
rect 11012 64708 11016 64764
rect 10952 64704 11016 64708
rect 11032 64764 11096 64768
rect 11032 64708 11036 64764
rect 11036 64708 11092 64764
rect 11092 64708 11096 64764
rect 11032 64704 11096 64708
rect 11112 64764 11176 64768
rect 11112 64708 11116 64764
rect 11116 64708 11172 64764
rect 11172 64708 11176 64764
rect 11112 64704 11176 64708
rect 11192 64764 11256 64768
rect 11192 64708 11196 64764
rect 11196 64708 11252 64764
rect 11252 64708 11256 64764
rect 11192 64704 11256 64708
rect 20952 64764 21016 64768
rect 20952 64708 20956 64764
rect 20956 64708 21012 64764
rect 21012 64708 21016 64764
rect 20952 64704 21016 64708
rect 21032 64764 21096 64768
rect 21032 64708 21036 64764
rect 21036 64708 21092 64764
rect 21092 64708 21096 64764
rect 21032 64704 21096 64708
rect 21112 64764 21176 64768
rect 21112 64708 21116 64764
rect 21116 64708 21172 64764
rect 21172 64708 21176 64764
rect 21112 64704 21176 64708
rect 21192 64764 21256 64768
rect 21192 64708 21196 64764
rect 21196 64708 21252 64764
rect 21252 64708 21256 64764
rect 21192 64704 21256 64708
rect 21588 64500 21652 64564
rect 5952 64220 6016 64224
rect 5952 64164 5956 64220
rect 5956 64164 6012 64220
rect 6012 64164 6016 64220
rect 5952 64160 6016 64164
rect 6032 64220 6096 64224
rect 6032 64164 6036 64220
rect 6036 64164 6092 64220
rect 6092 64164 6096 64220
rect 6032 64160 6096 64164
rect 6112 64220 6176 64224
rect 6112 64164 6116 64220
rect 6116 64164 6172 64220
rect 6172 64164 6176 64220
rect 6112 64160 6176 64164
rect 6192 64220 6256 64224
rect 6192 64164 6196 64220
rect 6196 64164 6252 64220
rect 6252 64164 6256 64220
rect 6192 64160 6256 64164
rect 15952 64220 16016 64224
rect 15952 64164 15956 64220
rect 15956 64164 16012 64220
rect 16012 64164 16016 64220
rect 15952 64160 16016 64164
rect 16032 64220 16096 64224
rect 16032 64164 16036 64220
rect 16036 64164 16092 64220
rect 16092 64164 16096 64220
rect 16032 64160 16096 64164
rect 16112 64220 16176 64224
rect 16112 64164 16116 64220
rect 16116 64164 16172 64220
rect 16172 64164 16176 64220
rect 16112 64160 16176 64164
rect 16192 64220 16256 64224
rect 16192 64164 16196 64220
rect 16196 64164 16252 64220
rect 16252 64164 16256 64220
rect 16192 64160 16256 64164
rect 25952 64220 26016 64224
rect 25952 64164 25956 64220
rect 25956 64164 26012 64220
rect 26012 64164 26016 64220
rect 25952 64160 26016 64164
rect 26032 64220 26096 64224
rect 26032 64164 26036 64220
rect 26036 64164 26092 64220
rect 26092 64164 26096 64220
rect 26032 64160 26096 64164
rect 26112 64220 26176 64224
rect 26112 64164 26116 64220
rect 26116 64164 26172 64220
rect 26172 64164 26176 64220
rect 26112 64160 26176 64164
rect 26192 64220 26256 64224
rect 26192 64164 26196 64220
rect 26196 64164 26252 64220
rect 26252 64164 26256 64220
rect 26192 64160 26256 64164
rect 10952 63676 11016 63680
rect 10952 63620 10956 63676
rect 10956 63620 11012 63676
rect 11012 63620 11016 63676
rect 10952 63616 11016 63620
rect 11032 63676 11096 63680
rect 11032 63620 11036 63676
rect 11036 63620 11092 63676
rect 11092 63620 11096 63676
rect 11032 63616 11096 63620
rect 11112 63676 11176 63680
rect 11112 63620 11116 63676
rect 11116 63620 11172 63676
rect 11172 63620 11176 63676
rect 11112 63616 11176 63620
rect 11192 63676 11256 63680
rect 11192 63620 11196 63676
rect 11196 63620 11252 63676
rect 11252 63620 11256 63676
rect 11192 63616 11256 63620
rect 20952 63676 21016 63680
rect 20952 63620 20956 63676
rect 20956 63620 21012 63676
rect 21012 63620 21016 63676
rect 20952 63616 21016 63620
rect 21032 63676 21096 63680
rect 21032 63620 21036 63676
rect 21036 63620 21092 63676
rect 21092 63620 21096 63676
rect 21032 63616 21096 63620
rect 21112 63676 21176 63680
rect 21112 63620 21116 63676
rect 21116 63620 21172 63676
rect 21172 63620 21176 63676
rect 21112 63616 21176 63620
rect 21192 63676 21256 63680
rect 21192 63620 21196 63676
rect 21196 63620 21252 63676
rect 21252 63620 21256 63676
rect 21192 63616 21256 63620
rect 5952 63132 6016 63136
rect 5952 63076 5956 63132
rect 5956 63076 6012 63132
rect 6012 63076 6016 63132
rect 5952 63072 6016 63076
rect 6032 63132 6096 63136
rect 6032 63076 6036 63132
rect 6036 63076 6092 63132
rect 6092 63076 6096 63132
rect 6032 63072 6096 63076
rect 6112 63132 6176 63136
rect 6112 63076 6116 63132
rect 6116 63076 6172 63132
rect 6172 63076 6176 63132
rect 6112 63072 6176 63076
rect 6192 63132 6256 63136
rect 6192 63076 6196 63132
rect 6196 63076 6252 63132
rect 6252 63076 6256 63132
rect 6192 63072 6256 63076
rect 15952 63132 16016 63136
rect 15952 63076 15956 63132
rect 15956 63076 16012 63132
rect 16012 63076 16016 63132
rect 15952 63072 16016 63076
rect 16032 63132 16096 63136
rect 16032 63076 16036 63132
rect 16036 63076 16092 63132
rect 16092 63076 16096 63132
rect 16032 63072 16096 63076
rect 16112 63132 16176 63136
rect 16112 63076 16116 63132
rect 16116 63076 16172 63132
rect 16172 63076 16176 63132
rect 16112 63072 16176 63076
rect 16192 63132 16256 63136
rect 16192 63076 16196 63132
rect 16196 63076 16252 63132
rect 16252 63076 16256 63132
rect 16192 63072 16256 63076
rect 25952 63132 26016 63136
rect 25952 63076 25956 63132
rect 25956 63076 26012 63132
rect 26012 63076 26016 63132
rect 25952 63072 26016 63076
rect 26032 63132 26096 63136
rect 26032 63076 26036 63132
rect 26036 63076 26092 63132
rect 26092 63076 26096 63132
rect 26032 63072 26096 63076
rect 26112 63132 26176 63136
rect 26112 63076 26116 63132
rect 26116 63076 26172 63132
rect 26172 63076 26176 63132
rect 26112 63072 26176 63076
rect 26192 63132 26256 63136
rect 26192 63076 26196 63132
rect 26196 63076 26252 63132
rect 26252 63076 26256 63132
rect 26192 63072 26256 63076
rect 18092 62868 18156 62932
rect 10952 62588 11016 62592
rect 10952 62532 10956 62588
rect 10956 62532 11012 62588
rect 11012 62532 11016 62588
rect 10952 62528 11016 62532
rect 11032 62588 11096 62592
rect 11032 62532 11036 62588
rect 11036 62532 11092 62588
rect 11092 62532 11096 62588
rect 11032 62528 11096 62532
rect 11112 62588 11176 62592
rect 11112 62532 11116 62588
rect 11116 62532 11172 62588
rect 11172 62532 11176 62588
rect 11112 62528 11176 62532
rect 11192 62588 11256 62592
rect 11192 62532 11196 62588
rect 11196 62532 11252 62588
rect 11252 62532 11256 62588
rect 11192 62528 11256 62532
rect 20952 62588 21016 62592
rect 20952 62532 20956 62588
rect 20956 62532 21012 62588
rect 21012 62532 21016 62588
rect 20952 62528 21016 62532
rect 21032 62588 21096 62592
rect 21032 62532 21036 62588
rect 21036 62532 21092 62588
rect 21092 62532 21096 62588
rect 21032 62528 21096 62532
rect 21112 62588 21176 62592
rect 21112 62532 21116 62588
rect 21116 62532 21172 62588
rect 21172 62532 21176 62588
rect 21112 62528 21176 62532
rect 21192 62588 21256 62592
rect 21192 62532 21196 62588
rect 21196 62532 21252 62588
rect 21252 62532 21256 62588
rect 21192 62528 21256 62532
rect 5952 62044 6016 62048
rect 5952 61988 5956 62044
rect 5956 61988 6012 62044
rect 6012 61988 6016 62044
rect 5952 61984 6016 61988
rect 6032 62044 6096 62048
rect 6032 61988 6036 62044
rect 6036 61988 6092 62044
rect 6092 61988 6096 62044
rect 6032 61984 6096 61988
rect 6112 62044 6176 62048
rect 6112 61988 6116 62044
rect 6116 61988 6172 62044
rect 6172 61988 6176 62044
rect 6112 61984 6176 61988
rect 6192 62044 6256 62048
rect 6192 61988 6196 62044
rect 6196 61988 6252 62044
rect 6252 61988 6256 62044
rect 6192 61984 6256 61988
rect 15952 62044 16016 62048
rect 15952 61988 15956 62044
rect 15956 61988 16012 62044
rect 16012 61988 16016 62044
rect 15952 61984 16016 61988
rect 16032 62044 16096 62048
rect 16032 61988 16036 62044
rect 16036 61988 16092 62044
rect 16092 61988 16096 62044
rect 16032 61984 16096 61988
rect 16112 62044 16176 62048
rect 16112 61988 16116 62044
rect 16116 61988 16172 62044
rect 16172 61988 16176 62044
rect 16112 61984 16176 61988
rect 16192 62044 16256 62048
rect 16192 61988 16196 62044
rect 16196 61988 16252 62044
rect 16252 61988 16256 62044
rect 16192 61984 16256 61988
rect 25952 62044 26016 62048
rect 25952 61988 25956 62044
rect 25956 61988 26012 62044
rect 26012 61988 26016 62044
rect 25952 61984 26016 61988
rect 26032 62044 26096 62048
rect 26032 61988 26036 62044
rect 26036 61988 26092 62044
rect 26092 61988 26096 62044
rect 26032 61984 26096 61988
rect 26112 62044 26176 62048
rect 26112 61988 26116 62044
rect 26116 61988 26172 62044
rect 26172 61988 26176 62044
rect 26112 61984 26176 61988
rect 26192 62044 26256 62048
rect 26192 61988 26196 62044
rect 26196 61988 26252 62044
rect 26252 61988 26256 62044
rect 26192 61984 26256 61988
rect 10952 61500 11016 61504
rect 10952 61444 10956 61500
rect 10956 61444 11012 61500
rect 11012 61444 11016 61500
rect 10952 61440 11016 61444
rect 11032 61500 11096 61504
rect 11032 61444 11036 61500
rect 11036 61444 11092 61500
rect 11092 61444 11096 61500
rect 11032 61440 11096 61444
rect 11112 61500 11176 61504
rect 11112 61444 11116 61500
rect 11116 61444 11172 61500
rect 11172 61444 11176 61500
rect 11112 61440 11176 61444
rect 11192 61500 11256 61504
rect 11192 61444 11196 61500
rect 11196 61444 11252 61500
rect 11252 61444 11256 61500
rect 11192 61440 11256 61444
rect 20952 61500 21016 61504
rect 20952 61444 20956 61500
rect 20956 61444 21012 61500
rect 21012 61444 21016 61500
rect 20952 61440 21016 61444
rect 21032 61500 21096 61504
rect 21032 61444 21036 61500
rect 21036 61444 21092 61500
rect 21092 61444 21096 61500
rect 21032 61440 21096 61444
rect 21112 61500 21176 61504
rect 21112 61444 21116 61500
rect 21116 61444 21172 61500
rect 21172 61444 21176 61500
rect 21112 61440 21176 61444
rect 21192 61500 21256 61504
rect 21192 61444 21196 61500
rect 21196 61444 21252 61500
rect 21252 61444 21256 61500
rect 21192 61440 21256 61444
rect 5952 60956 6016 60960
rect 5952 60900 5956 60956
rect 5956 60900 6012 60956
rect 6012 60900 6016 60956
rect 5952 60896 6016 60900
rect 6032 60956 6096 60960
rect 6032 60900 6036 60956
rect 6036 60900 6092 60956
rect 6092 60900 6096 60956
rect 6032 60896 6096 60900
rect 6112 60956 6176 60960
rect 6112 60900 6116 60956
rect 6116 60900 6172 60956
rect 6172 60900 6176 60956
rect 6112 60896 6176 60900
rect 6192 60956 6256 60960
rect 6192 60900 6196 60956
rect 6196 60900 6252 60956
rect 6252 60900 6256 60956
rect 6192 60896 6256 60900
rect 15952 60956 16016 60960
rect 15952 60900 15956 60956
rect 15956 60900 16012 60956
rect 16012 60900 16016 60956
rect 15952 60896 16016 60900
rect 16032 60956 16096 60960
rect 16032 60900 16036 60956
rect 16036 60900 16092 60956
rect 16092 60900 16096 60956
rect 16032 60896 16096 60900
rect 16112 60956 16176 60960
rect 16112 60900 16116 60956
rect 16116 60900 16172 60956
rect 16172 60900 16176 60956
rect 16112 60896 16176 60900
rect 16192 60956 16256 60960
rect 16192 60900 16196 60956
rect 16196 60900 16252 60956
rect 16252 60900 16256 60956
rect 16192 60896 16256 60900
rect 25952 60956 26016 60960
rect 25952 60900 25956 60956
rect 25956 60900 26012 60956
rect 26012 60900 26016 60956
rect 25952 60896 26016 60900
rect 26032 60956 26096 60960
rect 26032 60900 26036 60956
rect 26036 60900 26092 60956
rect 26092 60900 26096 60956
rect 26032 60896 26096 60900
rect 26112 60956 26176 60960
rect 26112 60900 26116 60956
rect 26116 60900 26172 60956
rect 26172 60900 26176 60956
rect 26112 60896 26176 60900
rect 26192 60956 26256 60960
rect 26192 60900 26196 60956
rect 26196 60900 26252 60956
rect 26252 60900 26256 60956
rect 26192 60896 26256 60900
rect 10952 60412 11016 60416
rect 10952 60356 10956 60412
rect 10956 60356 11012 60412
rect 11012 60356 11016 60412
rect 10952 60352 11016 60356
rect 11032 60412 11096 60416
rect 11032 60356 11036 60412
rect 11036 60356 11092 60412
rect 11092 60356 11096 60412
rect 11032 60352 11096 60356
rect 11112 60412 11176 60416
rect 11112 60356 11116 60412
rect 11116 60356 11172 60412
rect 11172 60356 11176 60412
rect 11112 60352 11176 60356
rect 11192 60412 11256 60416
rect 11192 60356 11196 60412
rect 11196 60356 11252 60412
rect 11252 60356 11256 60412
rect 11192 60352 11256 60356
rect 20952 60412 21016 60416
rect 20952 60356 20956 60412
rect 20956 60356 21012 60412
rect 21012 60356 21016 60412
rect 20952 60352 21016 60356
rect 21032 60412 21096 60416
rect 21032 60356 21036 60412
rect 21036 60356 21092 60412
rect 21092 60356 21096 60412
rect 21032 60352 21096 60356
rect 21112 60412 21176 60416
rect 21112 60356 21116 60412
rect 21116 60356 21172 60412
rect 21172 60356 21176 60412
rect 21112 60352 21176 60356
rect 21192 60412 21256 60416
rect 21192 60356 21196 60412
rect 21196 60356 21252 60412
rect 21252 60356 21256 60412
rect 21192 60352 21256 60356
rect 5952 59868 6016 59872
rect 5952 59812 5956 59868
rect 5956 59812 6012 59868
rect 6012 59812 6016 59868
rect 5952 59808 6016 59812
rect 6032 59868 6096 59872
rect 6032 59812 6036 59868
rect 6036 59812 6092 59868
rect 6092 59812 6096 59868
rect 6032 59808 6096 59812
rect 6112 59868 6176 59872
rect 6112 59812 6116 59868
rect 6116 59812 6172 59868
rect 6172 59812 6176 59868
rect 6112 59808 6176 59812
rect 6192 59868 6256 59872
rect 6192 59812 6196 59868
rect 6196 59812 6252 59868
rect 6252 59812 6256 59868
rect 6192 59808 6256 59812
rect 15952 59868 16016 59872
rect 15952 59812 15956 59868
rect 15956 59812 16012 59868
rect 16012 59812 16016 59868
rect 15952 59808 16016 59812
rect 16032 59868 16096 59872
rect 16032 59812 16036 59868
rect 16036 59812 16092 59868
rect 16092 59812 16096 59868
rect 16032 59808 16096 59812
rect 16112 59868 16176 59872
rect 16112 59812 16116 59868
rect 16116 59812 16172 59868
rect 16172 59812 16176 59868
rect 16112 59808 16176 59812
rect 16192 59868 16256 59872
rect 16192 59812 16196 59868
rect 16196 59812 16252 59868
rect 16252 59812 16256 59868
rect 16192 59808 16256 59812
rect 25952 59868 26016 59872
rect 25952 59812 25956 59868
rect 25956 59812 26012 59868
rect 26012 59812 26016 59868
rect 25952 59808 26016 59812
rect 26032 59868 26096 59872
rect 26032 59812 26036 59868
rect 26036 59812 26092 59868
rect 26092 59812 26096 59868
rect 26032 59808 26096 59812
rect 26112 59868 26176 59872
rect 26112 59812 26116 59868
rect 26116 59812 26172 59868
rect 26172 59812 26176 59868
rect 26112 59808 26176 59812
rect 26192 59868 26256 59872
rect 26192 59812 26196 59868
rect 26196 59812 26252 59868
rect 26252 59812 26256 59868
rect 26192 59808 26256 59812
rect 10952 59324 11016 59328
rect 10952 59268 10956 59324
rect 10956 59268 11012 59324
rect 11012 59268 11016 59324
rect 10952 59264 11016 59268
rect 11032 59324 11096 59328
rect 11032 59268 11036 59324
rect 11036 59268 11092 59324
rect 11092 59268 11096 59324
rect 11032 59264 11096 59268
rect 11112 59324 11176 59328
rect 11112 59268 11116 59324
rect 11116 59268 11172 59324
rect 11172 59268 11176 59324
rect 11112 59264 11176 59268
rect 11192 59324 11256 59328
rect 11192 59268 11196 59324
rect 11196 59268 11252 59324
rect 11252 59268 11256 59324
rect 11192 59264 11256 59268
rect 20952 59324 21016 59328
rect 20952 59268 20956 59324
rect 20956 59268 21012 59324
rect 21012 59268 21016 59324
rect 20952 59264 21016 59268
rect 21032 59324 21096 59328
rect 21032 59268 21036 59324
rect 21036 59268 21092 59324
rect 21092 59268 21096 59324
rect 21032 59264 21096 59268
rect 21112 59324 21176 59328
rect 21112 59268 21116 59324
rect 21116 59268 21172 59324
rect 21172 59268 21176 59324
rect 21112 59264 21176 59268
rect 21192 59324 21256 59328
rect 21192 59268 21196 59324
rect 21196 59268 21252 59324
rect 21252 59268 21256 59324
rect 21192 59264 21256 59268
rect 5952 58780 6016 58784
rect 5952 58724 5956 58780
rect 5956 58724 6012 58780
rect 6012 58724 6016 58780
rect 5952 58720 6016 58724
rect 6032 58780 6096 58784
rect 6032 58724 6036 58780
rect 6036 58724 6092 58780
rect 6092 58724 6096 58780
rect 6032 58720 6096 58724
rect 6112 58780 6176 58784
rect 6112 58724 6116 58780
rect 6116 58724 6172 58780
rect 6172 58724 6176 58780
rect 6112 58720 6176 58724
rect 6192 58780 6256 58784
rect 6192 58724 6196 58780
rect 6196 58724 6252 58780
rect 6252 58724 6256 58780
rect 6192 58720 6256 58724
rect 15952 58780 16016 58784
rect 15952 58724 15956 58780
rect 15956 58724 16012 58780
rect 16012 58724 16016 58780
rect 15952 58720 16016 58724
rect 16032 58780 16096 58784
rect 16032 58724 16036 58780
rect 16036 58724 16092 58780
rect 16092 58724 16096 58780
rect 16032 58720 16096 58724
rect 16112 58780 16176 58784
rect 16112 58724 16116 58780
rect 16116 58724 16172 58780
rect 16172 58724 16176 58780
rect 16112 58720 16176 58724
rect 16192 58780 16256 58784
rect 16192 58724 16196 58780
rect 16196 58724 16252 58780
rect 16252 58724 16256 58780
rect 16192 58720 16256 58724
rect 25952 58780 26016 58784
rect 25952 58724 25956 58780
rect 25956 58724 26012 58780
rect 26012 58724 26016 58780
rect 25952 58720 26016 58724
rect 26032 58780 26096 58784
rect 26032 58724 26036 58780
rect 26036 58724 26092 58780
rect 26092 58724 26096 58780
rect 26032 58720 26096 58724
rect 26112 58780 26176 58784
rect 26112 58724 26116 58780
rect 26116 58724 26172 58780
rect 26172 58724 26176 58780
rect 26112 58720 26176 58724
rect 26192 58780 26256 58784
rect 26192 58724 26196 58780
rect 26196 58724 26252 58780
rect 26252 58724 26256 58780
rect 26192 58720 26256 58724
rect 10952 58236 11016 58240
rect 10952 58180 10956 58236
rect 10956 58180 11012 58236
rect 11012 58180 11016 58236
rect 10952 58176 11016 58180
rect 11032 58236 11096 58240
rect 11032 58180 11036 58236
rect 11036 58180 11092 58236
rect 11092 58180 11096 58236
rect 11032 58176 11096 58180
rect 11112 58236 11176 58240
rect 11112 58180 11116 58236
rect 11116 58180 11172 58236
rect 11172 58180 11176 58236
rect 11112 58176 11176 58180
rect 11192 58236 11256 58240
rect 11192 58180 11196 58236
rect 11196 58180 11252 58236
rect 11252 58180 11256 58236
rect 11192 58176 11256 58180
rect 20952 58236 21016 58240
rect 20952 58180 20956 58236
rect 20956 58180 21012 58236
rect 21012 58180 21016 58236
rect 20952 58176 21016 58180
rect 21032 58236 21096 58240
rect 21032 58180 21036 58236
rect 21036 58180 21092 58236
rect 21092 58180 21096 58236
rect 21032 58176 21096 58180
rect 21112 58236 21176 58240
rect 21112 58180 21116 58236
rect 21116 58180 21172 58236
rect 21172 58180 21176 58236
rect 21112 58176 21176 58180
rect 21192 58236 21256 58240
rect 21192 58180 21196 58236
rect 21196 58180 21252 58236
rect 21252 58180 21256 58236
rect 21192 58176 21256 58180
rect 11468 58032 11532 58036
rect 11468 57976 11518 58032
rect 11518 57976 11532 58032
rect 11468 57972 11532 57976
rect 5952 57692 6016 57696
rect 5952 57636 5956 57692
rect 5956 57636 6012 57692
rect 6012 57636 6016 57692
rect 5952 57632 6016 57636
rect 6032 57692 6096 57696
rect 6032 57636 6036 57692
rect 6036 57636 6092 57692
rect 6092 57636 6096 57692
rect 6032 57632 6096 57636
rect 6112 57692 6176 57696
rect 6112 57636 6116 57692
rect 6116 57636 6172 57692
rect 6172 57636 6176 57692
rect 6112 57632 6176 57636
rect 6192 57692 6256 57696
rect 6192 57636 6196 57692
rect 6196 57636 6252 57692
rect 6252 57636 6256 57692
rect 6192 57632 6256 57636
rect 15952 57692 16016 57696
rect 15952 57636 15956 57692
rect 15956 57636 16012 57692
rect 16012 57636 16016 57692
rect 15952 57632 16016 57636
rect 16032 57692 16096 57696
rect 16032 57636 16036 57692
rect 16036 57636 16092 57692
rect 16092 57636 16096 57692
rect 16032 57632 16096 57636
rect 16112 57692 16176 57696
rect 16112 57636 16116 57692
rect 16116 57636 16172 57692
rect 16172 57636 16176 57692
rect 16112 57632 16176 57636
rect 16192 57692 16256 57696
rect 16192 57636 16196 57692
rect 16196 57636 16252 57692
rect 16252 57636 16256 57692
rect 16192 57632 16256 57636
rect 25952 57692 26016 57696
rect 25952 57636 25956 57692
rect 25956 57636 26012 57692
rect 26012 57636 26016 57692
rect 25952 57632 26016 57636
rect 26032 57692 26096 57696
rect 26032 57636 26036 57692
rect 26036 57636 26092 57692
rect 26092 57636 26096 57692
rect 26032 57632 26096 57636
rect 26112 57692 26176 57696
rect 26112 57636 26116 57692
rect 26116 57636 26172 57692
rect 26172 57636 26176 57692
rect 26112 57632 26176 57636
rect 26192 57692 26256 57696
rect 26192 57636 26196 57692
rect 26196 57636 26252 57692
rect 26252 57636 26256 57692
rect 26192 57632 26256 57636
rect 20484 57292 20548 57356
rect 10952 57148 11016 57152
rect 10952 57092 10956 57148
rect 10956 57092 11012 57148
rect 11012 57092 11016 57148
rect 10952 57088 11016 57092
rect 11032 57148 11096 57152
rect 11032 57092 11036 57148
rect 11036 57092 11092 57148
rect 11092 57092 11096 57148
rect 11032 57088 11096 57092
rect 11112 57148 11176 57152
rect 11112 57092 11116 57148
rect 11116 57092 11172 57148
rect 11172 57092 11176 57148
rect 11112 57088 11176 57092
rect 11192 57148 11256 57152
rect 11192 57092 11196 57148
rect 11196 57092 11252 57148
rect 11252 57092 11256 57148
rect 11192 57088 11256 57092
rect 20952 57148 21016 57152
rect 20952 57092 20956 57148
rect 20956 57092 21012 57148
rect 21012 57092 21016 57148
rect 20952 57088 21016 57092
rect 21032 57148 21096 57152
rect 21032 57092 21036 57148
rect 21036 57092 21092 57148
rect 21092 57092 21096 57148
rect 21032 57088 21096 57092
rect 21112 57148 21176 57152
rect 21112 57092 21116 57148
rect 21116 57092 21172 57148
rect 21172 57092 21176 57148
rect 21112 57088 21176 57092
rect 21192 57148 21256 57152
rect 21192 57092 21196 57148
rect 21196 57092 21252 57148
rect 21252 57092 21256 57148
rect 21192 57088 21256 57092
rect 15700 56672 15764 56676
rect 15700 56616 15750 56672
rect 15750 56616 15764 56672
rect 15700 56612 15764 56616
rect 5952 56604 6016 56608
rect 5952 56548 5956 56604
rect 5956 56548 6012 56604
rect 6012 56548 6016 56604
rect 5952 56544 6016 56548
rect 6032 56604 6096 56608
rect 6032 56548 6036 56604
rect 6036 56548 6092 56604
rect 6092 56548 6096 56604
rect 6032 56544 6096 56548
rect 6112 56604 6176 56608
rect 6112 56548 6116 56604
rect 6116 56548 6172 56604
rect 6172 56548 6176 56604
rect 6112 56544 6176 56548
rect 6192 56604 6256 56608
rect 6192 56548 6196 56604
rect 6196 56548 6252 56604
rect 6252 56548 6256 56604
rect 6192 56544 6256 56548
rect 15952 56604 16016 56608
rect 15952 56548 15956 56604
rect 15956 56548 16012 56604
rect 16012 56548 16016 56604
rect 15952 56544 16016 56548
rect 16032 56604 16096 56608
rect 16032 56548 16036 56604
rect 16036 56548 16092 56604
rect 16092 56548 16096 56604
rect 16032 56544 16096 56548
rect 16112 56604 16176 56608
rect 16112 56548 16116 56604
rect 16116 56548 16172 56604
rect 16172 56548 16176 56604
rect 16112 56544 16176 56548
rect 16192 56604 16256 56608
rect 16192 56548 16196 56604
rect 16196 56548 16252 56604
rect 16252 56548 16256 56604
rect 16192 56544 16256 56548
rect 27844 56612 27908 56676
rect 25952 56604 26016 56608
rect 25952 56548 25956 56604
rect 25956 56548 26012 56604
rect 26012 56548 26016 56604
rect 25952 56544 26016 56548
rect 26032 56604 26096 56608
rect 26032 56548 26036 56604
rect 26036 56548 26092 56604
rect 26092 56548 26096 56604
rect 26032 56544 26096 56548
rect 26112 56604 26176 56608
rect 26112 56548 26116 56604
rect 26116 56548 26172 56604
rect 26172 56548 26176 56604
rect 26112 56544 26176 56548
rect 26192 56604 26256 56608
rect 26192 56548 26196 56604
rect 26196 56548 26252 56604
rect 26252 56548 26256 56604
rect 26192 56544 26256 56548
rect 17724 56476 17788 56540
rect 10952 56060 11016 56064
rect 10952 56004 10956 56060
rect 10956 56004 11012 56060
rect 11012 56004 11016 56060
rect 10952 56000 11016 56004
rect 11032 56060 11096 56064
rect 11032 56004 11036 56060
rect 11036 56004 11092 56060
rect 11092 56004 11096 56060
rect 11032 56000 11096 56004
rect 11112 56060 11176 56064
rect 11112 56004 11116 56060
rect 11116 56004 11172 56060
rect 11172 56004 11176 56060
rect 11112 56000 11176 56004
rect 11192 56060 11256 56064
rect 11192 56004 11196 56060
rect 11196 56004 11252 56060
rect 11252 56004 11256 56060
rect 11192 56000 11256 56004
rect 20952 56060 21016 56064
rect 20952 56004 20956 56060
rect 20956 56004 21012 56060
rect 21012 56004 21016 56060
rect 20952 56000 21016 56004
rect 21032 56060 21096 56064
rect 21032 56004 21036 56060
rect 21036 56004 21092 56060
rect 21092 56004 21096 56060
rect 21032 56000 21096 56004
rect 21112 56060 21176 56064
rect 21112 56004 21116 56060
rect 21116 56004 21172 56060
rect 21172 56004 21176 56060
rect 21112 56000 21176 56004
rect 21192 56060 21256 56064
rect 21192 56004 21196 56060
rect 21196 56004 21252 56060
rect 21252 56004 21256 56060
rect 21192 56000 21256 56004
rect 5952 55516 6016 55520
rect 5952 55460 5956 55516
rect 5956 55460 6012 55516
rect 6012 55460 6016 55516
rect 5952 55456 6016 55460
rect 6032 55516 6096 55520
rect 6032 55460 6036 55516
rect 6036 55460 6092 55516
rect 6092 55460 6096 55516
rect 6032 55456 6096 55460
rect 6112 55516 6176 55520
rect 6112 55460 6116 55516
rect 6116 55460 6172 55516
rect 6172 55460 6176 55516
rect 6112 55456 6176 55460
rect 6192 55516 6256 55520
rect 6192 55460 6196 55516
rect 6196 55460 6252 55516
rect 6252 55460 6256 55516
rect 6192 55456 6256 55460
rect 15952 55516 16016 55520
rect 15952 55460 15956 55516
rect 15956 55460 16012 55516
rect 16012 55460 16016 55516
rect 15952 55456 16016 55460
rect 16032 55516 16096 55520
rect 16032 55460 16036 55516
rect 16036 55460 16092 55516
rect 16092 55460 16096 55516
rect 16032 55456 16096 55460
rect 16112 55516 16176 55520
rect 16112 55460 16116 55516
rect 16116 55460 16172 55516
rect 16172 55460 16176 55516
rect 16112 55456 16176 55460
rect 16192 55516 16256 55520
rect 16192 55460 16196 55516
rect 16196 55460 16252 55516
rect 16252 55460 16256 55516
rect 16192 55456 16256 55460
rect 25952 55516 26016 55520
rect 25952 55460 25956 55516
rect 25956 55460 26012 55516
rect 26012 55460 26016 55516
rect 25952 55456 26016 55460
rect 26032 55516 26096 55520
rect 26032 55460 26036 55516
rect 26036 55460 26092 55516
rect 26092 55460 26096 55516
rect 26032 55456 26096 55460
rect 26112 55516 26176 55520
rect 26112 55460 26116 55516
rect 26116 55460 26172 55516
rect 26172 55460 26176 55516
rect 26112 55456 26176 55460
rect 26192 55516 26256 55520
rect 26192 55460 26196 55516
rect 26196 55460 26252 55516
rect 26252 55460 26256 55516
rect 26192 55456 26256 55460
rect 21404 55252 21468 55316
rect 10952 54972 11016 54976
rect 10952 54916 10956 54972
rect 10956 54916 11012 54972
rect 11012 54916 11016 54972
rect 10952 54912 11016 54916
rect 11032 54972 11096 54976
rect 11032 54916 11036 54972
rect 11036 54916 11092 54972
rect 11092 54916 11096 54972
rect 11032 54912 11096 54916
rect 11112 54972 11176 54976
rect 11112 54916 11116 54972
rect 11116 54916 11172 54972
rect 11172 54916 11176 54972
rect 11112 54912 11176 54916
rect 11192 54972 11256 54976
rect 11192 54916 11196 54972
rect 11196 54916 11252 54972
rect 11252 54916 11256 54972
rect 11192 54912 11256 54916
rect 20952 54972 21016 54976
rect 20952 54916 20956 54972
rect 20956 54916 21012 54972
rect 21012 54916 21016 54972
rect 20952 54912 21016 54916
rect 21032 54972 21096 54976
rect 21032 54916 21036 54972
rect 21036 54916 21092 54972
rect 21092 54916 21096 54972
rect 21032 54912 21096 54916
rect 21112 54972 21176 54976
rect 21112 54916 21116 54972
rect 21116 54916 21172 54972
rect 21172 54916 21176 54972
rect 21112 54912 21176 54916
rect 21192 54972 21256 54976
rect 21192 54916 21196 54972
rect 21196 54916 21252 54972
rect 21252 54916 21256 54972
rect 21192 54912 21256 54916
rect 5952 54428 6016 54432
rect 5952 54372 5956 54428
rect 5956 54372 6012 54428
rect 6012 54372 6016 54428
rect 5952 54368 6016 54372
rect 6032 54428 6096 54432
rect 6032 54372 6036 54428
rect 6036 54372 6092 54428
rect 6092 54372 6096 54428
rect 6032 54368 6096 54372
rect 6112 54428 6176 54432
rect 6112 54372 6116 54428
rect 6116 54372 6172 54428
rect 6172 54372 6176 54428
rect 6112 54368 6176 54372
rect 6192 54428 6256 54432
rect 6192 54372 6196 54428
rect 6196 54372 6252 54428
rect 6252 54372 6256 54428
rect 6192 54368 6256 54372
rect 15952 54428 16016 54432
rect 15952 54372 15956 54428
rect 15956 54372 16012 54428
rect 16012 54372 16016 54428
rect 15952 54368 16016 54372
rect 16032 54428 16096 54432
rect 16032 54372 16036 54428
rect 16036 54372 16092 54428
rect 16092 54372 16096 54428
rect 16032 54368 16096 54372
rect 16112 54428 16176 54432
rect 16112 54372 16116 54428
rect 16116 54372 16172 54428
rect 16172 54372 16176 54428
rect 16112 54368 16176 54372
rect 16192 54428 16256 54432
rect 16192 54372 16196 54428
rect 16196 54372 16252 54428
rect 16252 54372 16256 54428
rect 16192 54368 16256 54372
rect 25952 54428 26016 54432
rect 25952 54372 25956 54428
rect 25956 54372 26012 54428
rect 26012 54372 26016 54428
rect 25952 54368 26016 54372
rect 26032 54428 26096 54432
rect 26032 54372 26036 54428
rect 26036 54372 26092 54428
rect 26092 54372 26096 54428
rect 26032 54368 26096 54372
rect 26112 54428 26176 54432
rect 26112 54372 26116 54428
rect 26116 54372 26172 54428
rect 26172 54372 26176 54428
rect 26112 54368 26176 54372
rect 26192 54428 26256 54432
rect 26192 54372 26196 54428
rect 26196 54372 26252 54428
rect 26252 54372 26256 54428
rect 26192 54368 26256 54372
rect 10952 53884 11016 53888
rect 10952 53828 10956 53884
rect 10956 53828 11012 53884
rect 11012 53828 11016 53884
rect 10952 53824 11016 53828
rect 11032 53884 11096 53888
rect 11032 53828 11036 53884
rect 11036 53828 11092 53884
rect 11092 53828 11096 53884
rect 11032 53824 11096 53828
rect 11112 53884 11176 53888
rect 11112 53828 11116 53884
rect 11116 53828 11172 53884
rect 11172 53828 11176 53884
rect 11112 53824 11176 53828
rect 11192 53884 11256 53888
rect 11192 53828 11196 53884
rect 11196 53828 11252 53884
rect 11252 53828 11256 53884
rect 11192 53824 11256 53828
rect 20952 53884 21016 53888
rect 20952 53828 20956 53884
rect 20956 53828 21012 53884
rect 21012 53828 21016 53884
rect 20952 53824 21016 53828
rect 21032 53884 21096 53888
rect 21032 53828 21036 53884
rect 21036 53828 21092 53884
rect 21092 53828 21096 53884
rect 21032 53824 21096 53828
rect 21112 53884 21176 53888
rect 21112 53828 21116 53884
rect 21116 53828 21172 53884
rect 21172 53828 21176 53884
rect 21112 53824 21176 53828
rect 21192 53884 21256 53888
rect 21192 53828 21196 53884
rect 21196 53828 21252 53884
rect 21252 53828 21256 53884
rect 21192 53824 21256 53828
rect 5952 53340 6016 53344
rect 5952 53284 5956 53340
rect 5956 53284 6012 53340
rect 6012 53284 6016 53340
rect 5952 53280 6016 53284
rect 6032 53340 6096 53344
rect 6032 53284 6036 53340
rect 6036 53284 6092 53340
rect 6092 53284 6096 53340
rect 6032 53280 6096 53284
rect 6112 53340 6176 53344
rect 6112 53284 6116 53340
rect 6116 53284 6172 53340
rect 6172 53284 6176 53340
rect 6112 53280 6176 53284
rect 6192 53340 6256 53344
rect 6192 53284 6196 53340
rect 6196 53284 6252 53340
rect 6252 53284 6256 53340
rect 6192 53280 6256 53284
rect 15952 53340 16016 53344
rect 15952 53284 15956 53340
rect 15956 53284 16012 53340
rect 16012 53284 16016 53340
rect 15952 53280 16016 53284
rect 16032 53340 16096 53344
rect 16032 53284 16036 53340
rect 16036 53284 16092 53340
rect 16092 53284 16096 53340
rect 16032 53280 16096 53284
rect 16112 53340 16176 53344
rect 16112 53284 16116 53340
rect 16116 53284 16172 53340
rect 16172 53284 16176 53340
rect 16112 53280 16176 53284
rect 16192 53340 16256 53344
rect 16192 53284 16196 53340
rect 16196 53284 16252 53340
rect 16252 53284 16256 53340
rect 16192 53280 16256 53284
rect 25952 53340 26016 53344
rect 25952 53284 25956 53340
rect 25956 53284 26012 53340
rect 26012 53284 26016 53340
rect 25952 53280 26016 53284
rect 26032 53340 26096 53344
rect 26032 53284 26036 53340
rect 26036 53284 26092 53340
rect 26092 53284 26096 53340
rect 26032 53280 26096 53284
rect 26112 53340 26176 53344
rect 26112 53284 26116 53340
rect 26116 53284 26172 53340
rect 26172 53284 26176 53340
rect 26112 53280 26176 53284
rect 26192 53340 26256 53344
rect 26192 53284 26196 53340
rect 26196 53284 26252 53340
rect 26252 53284 26256 53340
rect 26192 53280 26256 53284
rect 21772 53076 21836 53140
rect 25452 52940 25516 53004
rect 10952 52796 11016 52800
rect 10952 52740 10956 52796
rect 10956 52740 11012 52796
rect 11012 52740 11016 52796
rect 10952 52736 11016 52740
rect 11032 52796 11096 52800
rect 11032 52740 11036 52796
rect 11036 52740 11092 52796
rect 11092 52740 11096 52796
rect 11032 52736 11096 52740
rect 11112 52796 11176 52800
rect 11112 52740 11116 52796
rect 11116 52740 11172 52796
rect 11172 52740 11176 52796
rect 11112 52736 11176 52740
rect 11192 52796 11256 52800
rect 11192 52740 11196 52796
rect 11196 52740 11252 52796
rect 11252 52740 11256 52796
rect 11192 52736 11256 52740
rect 20952 52796 21016 52800
rect 20952 52740 20956 52796
rect 20956 52740 21012 52796
rect 21012 52740 21016 52796
rect 20952 52736 21016 52740
rect 21032 52796 21096 52800
rect 21032 52740 21036 52796
rect 21036 52740 21092 52796
rect 21092 52740 21096 52796
rect 21032 52736 21096 52740
rect 21112 52796 21176 52800
rect 21112 52740 21116 52796
rect 21116 52740 21172 52796
rect 21172 52740 21176 52796
rect 21112 52736 21176 52740
rect 21192 52796 21256 52800
rect 21192 52740 21196 52796
rect 21196 52740 21252 52796
rect 21252 52740 21256 52796
rect 21192 52736 21256 52740
rect 12020 52532 12084 52596
rect 16436 52592 16500 52596
rect 16436 52536 16486 52592
rect 16486 52536 16500 52592
rect 16436 52532 16500 52536
rect 5952 52252 6016 52256
rect 5952 52196 5956 52252
rect 5956 52196 6012 52252
rect 6012 52196 6016 52252
rect 5952 52192 6016 52196
rect 6032 52252 6096 52256
rect 6032 52196 6036 52252
rect 6036 52196 6092 52252
rect 6092 52196 6096 52252
rect 6032 52192 6096 52196
rect 6112 52252 6176 52256
rect 6112 52196 6116 52252
rect 6116 52196 6172 52252
rect 6172 52196 6176 52252
rect 6112 52192 6176 52196
rect 6192 52252 6256 52256
rect 6192 52196 6196 52252
rect 6196 52196 6252 52252
rect 6252 52196 6256 52252
rect 6192 52192 6256 52196
rect 15952 52252 16016 52256
rect 15952 52196 15956 52252
rect 15956 52196 16012 52252
rect 16012 52196 16016 52252
rect 15952 52192 16016 52196
rect 16032 52252 16096 52256
rect 16032 52196 16036 52252
rect 16036 52196 16092 52252
rect 16092 52196 16096 52252
rect 16032 52192 16096 52196
rect 16112 52252 16176 52256
rect 16112 52196 16116 52252
rect 16116 52196 16172 52252
rect 16172 52196 16176 52252
rect 16112 52192 16176 52196
rect 16192 52252 16256 52256
rect 16192 52196 16196 52252
rect 16196 52196 16252 52252
rect 16252 52196 16256 52252
rect 16192 52192 16256 52196
rect 25952 52252 26016 52256
rect 25952 52196 25956 52252
rect 25956 52196 26012 52252
rect 26012 52196 26016 52252
rect 25952 52192 26016 52196
rect 26032 52252 26096 52256
rect 26032 52196 26036 52252
rect 26036 52196 26092 52252
rect 26092 52196 26096 52252
rect 26032 52192 26096 52196
rect 26112 52252 26176 52256
rect 26112 52196 26116 52252
rect 26116 52196 26172 52252
rect 26172 52196 26176 52252
rect 26112 52192 26176 52196
rect 26192 52252 26256 52256
rect 26192 52196 26196 52252
rect 26196 52196 26252 52252
rect 26252 52196 26256 52252
rect 26192 52192 26256 52196
rect 17724 52124 17788 52188
rect 10952 51708 11016 51712
rect 10952 51652 10956 51708
rect 10956 51652 11012 51708
rect 11012 51652 11016 51708
rect 10952 51648 11016 51652
rect 11032 51708 11096 51712
rect 11032 51652 11036 51708
rect 11036 51652 11092 51708
rect 11092 51652 11096 51708
rect 11032 51648 11096 51652
rect 11112 51708 11176 51712
rect 11112 51652 11116 51708
rect 11116 51652 11172 51708
rect 11172 51652 11176 51708
rect 11112 51648 11176 51652
rect 11192 51708 11256 51712
rect 11192 51652 11196 51708
rect 11196 51652 11252 51708
rect 11252 51652 11256 51708
rect 11192 51648 11256 51652
rect 15516 51308 15580 51372
rect 20952 51708 21016 51712
rect 20952 51652 20956 51708
rect 20956 51652 21012 51708
rect 21012 51652 21016 51708
rect 20952 51648 21016 51652
rect 21032 51708 21096 51712
rect 21032 51652 21036 51708
rect 21036 51652 21092 51708
rect 21092 51652 21096 51708
rect 21032 51648 21096 51652
rect 21112 51708 21176 51712
rect 21112 51652 21116 51708
rect 21116 51652 21172 51708
rect 21172 51652 21176 51708
rect 21112 51648 21176 51652
rect 21192 51708 21256 51712
rect 21192 51652 21196 51708
rect 21196 51652 21252 51708
rect 21252 51652 21256 51708
rect 21192 51648 21256 51652
rect 5952 51164 6016 51168
rect 5952 51108 5956 51164
rect 5956 51108 6012 51164
rect 6012 51108 6016 51164
rect 5952 51104 6016 51108
rect 6032 51164 6096 51168
rect 6032 51108 6036 51164
rect 6036 51108 6092 51164
rect 6092 51108 6096 51164
rect 6032 51104 6096 51108
rect 6112 51164 6176 51168
rect 6112 51108 6116 51164
rect 6116 51108 6172 51164
rect 6172 51108 6176 51164
rect 6112 51104 6176 51108
rect 6192 51164 6256 51168
rect 6192 51108 6196 51164
rect 6196 51108 6252 51164
rect 6252 51108 6256 51164
rect 6192 51104 6256 51108
rect 15952 51164 16016 51168
rect 15952 51108 15956 51164
rect 15956 51108 16012 51164
rect 16012 51108 16016 51164
rect 15952 51104 16016 51108
rect 16032 51164 16096 51168
rect 16032 51108 16036 51164
rect 16036 51108 16092 51164
rect 16092 51108 16096 51164
rect 16032 51104 16096 51108
rect 16112 51164 16176 51168
rect 16112 51108 16116 51164
rect 16116 51108 16172 51164
rect 16172 51108 16176 51164
rect 16112 51104 16176 51108
rect 16192 51164 16256 51168
rect 16192 51108 16196 51164
rect 16196 51108 16252 51164
rect 16252 51108 16256 51164
rect 16192 51104 16256 51108
rect 25952 51164 26016 51168
rect 25952 51108 25956 51164
rect 25956 51108 26012 51164
rect 26012 51108 26016 51164
rect 25952 51104 26016 51108
rect 26032 51164 26096 51168
rect 26032 51108 26036 51164
rect 26036 51108 26092 51164
rect 26092 51108 26096 51164
rect 26032 51104 26096 51108
rect 26112 51164 26176 51168
rect 26112 51108 26116 51164
rect 26116 51108 26172 51164
rect 26172 51108 26176 51164
rect 26112 51104 26176 51108
rect 26192 51164 26256 51168
rect 26192 51108 26196 51164
rect 26196 51108 26252 51164
rect 26252 51108 26256 51164
rect 26192 51104 26256 51108
rect 15516 50764 15580 50828
rect 10952 50620 11016 50624
rect 10952 50564 10956 50620
rect 10956 50564 11012 50620
rect 11012 50564 11016 50620
rect 10952 50560 11016 50564
rect 11032 50620 11096 50624
rect 11032 50564 11036 50620
rect 11036 50564 11092 50620
rect 11092 50564 11096 50620
rect 11032 50560 11096 50564
rect 11112 50620 11176 50624
rect 11112 50564 11116 50620
rect 11116 50564 11172 50620
rect 11172 50564 11176 50620
rect 11112 50560 11176 50564
rect 11192 50620 11256 50624
rect 11192 50564 11196 50620
rect 11196 50564 11252 50620
rect 11252 50564 11256 50620
rect 11192 50560 11256 50564
rect 20952 50620 21016 50624
rect 20952 50564 20956 50620
rect 20956 50564 21012 50620
rect 21012 50564 21016 50620
rect 20952 50560 21016 50564
rect 21032 50620 21096 50624
rect 21032 50564 21036 50620
rect 21036 50564 21092 50620
rect 21092 50564 21096 50620
rect 21032 50560 21096 50564
rect 21112 50620 21176 50624
rect 21112 50564 21116 50620
rect 21116 50564 21172 50620
rect 21172 50564 21176 50620
rect 21112 50560 21176 50564
rect 21192 50620 21256 50624
rect 21192 50564 21196 50620
rect 21196 50564 21252 50620
rect 21252 50564 21256 50620
rect 21192 50560 21256 50564
rect 5952 50076 6016 50080
rect 5952 50020 5956 50076
rect 5956 50020 6012 50076
rect 6012 50020 6016 50076
rect 5952 50016 6016 50020
rect 6032 50076 6096 50080
rect 6032 50020 6036 50076
rect 6036 50020 6092 50076
rect 6092 50020 6096 50076
rect 6032 50016 6096 50020
rect 6112 50076 6176 50080
rect 6112 50020 6116 50076
rect 6116 50020 6172 50076
rect 6172 50020 6176 50076
rect 6112 50016 6176 50020
rect 6192 50076 6256 50080
rect 6192 50020 6196 50076
rect 6196 50020 6252 50076
rect 6252 50020 6256 50076
rect 6192 50016 6256 50020
rect 15952 50076 16016 50080
rect 15952 50020 15956 50076
rect 15956 50020 16012 50076
rect 16012 50020 16016 50076
rect 15952 50016 16016 50020
rect 16032 50076 16096 50080
rect 16032 50020 16036 50076
rect 16036 50020 16092 50076
rect 16092 50020 16096 50076
rect 16032 50016 16096 50020
rect 16112 50076 16176 50080
rect 16112 50020 16116 50076
rect 16116 50020 16172 50076
rect 16172 50020 16176 50076
rect 16112 50016 16176 50020
rect 16192 50076 16256 50080
rect 16192 50020 16196 50076
rect 16196 50020 16252 50076
rect 16252 50020 16256 50076
rect 16192 50016 16256 50020
rect 25952 50076 26016 50080
rect 25952 50020 25956 50076
rect 25956 50020 26012 50076
rect 26012 50020 26016 50076
rect 25952 50016 26016 50020
rect 26032 50076 26096 50080
rect 26032 50020 26036 50076
rect 26036 50020 26092 50076
rect 26092 50020 26096 50076
rect 26032 50016 26096 50020
rect 26112 50076 26176 50080
rect 26112 50020 26116 50076
rect 26116 50020 26172 50076
rect 26172 50020 26176 50076
rect 26112 50016 26176 50020
rect 26192 50076 26256 50080
rect 26192 50020 26196 50076
rect 26196 50020 26252 50076
rect 26252 50020 26256 50076
rect 26192 50016 26256 50020
rect 20300 49948 20364 50012
rect 16436 49540 16500 49604
rect 10952 49532 11016 49536
rect 10952 49476 10956 49532
rect 10956 49476 11012 49532
rect 11012 49476 11016 49532
rect 10952 49472 11016 49476
rect 11032 49532 11096 49536
rect 11032 49476 11036 49532
rect 11036 49476 11092 49532
rect 11092 49476 11096 49532
rect 11032 49472 11096 49476
rect 11112 49532 11176 49536
rect 11112 49476 11116 49532
rect 11116 49476 11172 49532
rect 11172 49476 11176 49532
rect 11112 49472 11176 49476
rect 11192 49532 11256 49536
rect 11192 49476 11196 49532
rect 11196 49476 11252 49532
rect 11252 49476 11256 49532
rect 11192 49472 11256 49476
rect 20952 49532 21016 49536
rect 20952 49476 20956 49532
rect 20956 49476 21012 49532
rect 21012 49476 21016 49532
rect 20952 49472 21016 49476
rect 21032 49532 21096 49536
rect 21032 49476 21036 49532
rect 21036 49476 21092 49532
rect 21092 49476 21096 49532
rect 21032 49472 21096 49476
rect 21112 49532 21176 49536
rect 21112 49476 21116 49532
rect 21116 49476 21172 49532
rect 21172 49476 21176 49532
rect 21112 49472 21176 49476
rect 21192 49532 21256 49536
rect 21192 49476 21196 49532
rect 21196 49476 21252 49532
rect 21252 49476 21256 49532
rect 21192 49472 21256 49476
rect 20484 49404 20548 49468
rect 20300 49132 20364 49196
rect 5952 48988 6016 48992
rect 5952 48932 5956 48988
rect 5956 48932 6012 48988
rect 6012 48932 6016 48988
rect 5952 48928 6016 48932
rect 6032 48988 6096 48992
rect 6032 48932 6036 48988
rect 6036 48932 6092 48988
rect 6092 48932 6096 48988
rect 6032 48928 6096 48932
rect 6112 48988 6176 48992
rect 6112 48932 6116 48988
rect 6116 48932 6172 48988
rect 6172 48932 6176 48988
rect 6112 48928 6176 48932
rect 6192 48988 6256 48992
rect 6192 48932 6196 48988
rect 6196 48932 6252 48988
rect 6252 48932 6256 48988
rect 6192 48928 6256 48932
rect 15952 48988 16016 48992
rect 15952 48932 15956 48988
rect 15956 48932 16012 48988
rect 16012 48932 16016 48988
rect 15952 48928 16016 48932
rect 16032 48988 16096 48992
rect 16032 48932 16036 48988
rect 16036 48932 16092 48988
rect 16092 48932 16096 48988
rect 16032 48928 16096 48932
rect 16112 48988 16176 48992
rect 16112 48932 16116 48988
rect 16116 48932 16172 48988
rect 16172 48932 16176 48988
rect 16112 48928 16176 48932
rect 16192 48988 16256 48992
rect 16192 48932 16196 48988
rect 16196 48932 16252 48988
rect 16252 48932 16256 48988
rect 16192 48928 16256 48932
rect 25952 48988 26016 48992
rect 25952 48932 25956 48988
rect 25956 48932 26012 48988
rect 26012 48932 26016 48988
rect 25952 48928 26016 48932
rect 26032 48988 26096 48992
rect 26032 48932 26036 48988
rect 26036 48932 26092 48988
rect 26092 48932 26096 48988
rect 26032 48928 26096 48932
rect 26112 48988 26176 48992
rect 26112 48932 26116 48988
rect 26116 48932 26172 48988
rect 26172 48932 26176 48988
rect 26112 48928 26176 48932
rect 26192 48988 26256 48992
rect 26192 48932 26196 48988
rect 26196 48932 26252 48988
rect 26252 48932 26256 48988
rect 26192 48928 26256 48932
rect 10952 48444 11016 48448
rect 10952 48388 10956 48444
rect 10956 48388 11012 48444
rect 11012 48388 11016 48444
rect 10952 48384 11016 48388
rect 11032 48444 11096 48448
rect 11032 48388 11036 48444
rect 11036 48388 11092 48444
rect 11092 48388 11096 48444
rect 11032 48384 11096 48388
rect 11112 48444 11176 48448
rect 11112 48388 11116 48444
rect 11116 48388 11172 48444
rect 11172 48388 11176 48444
rect 11112 48384 11176 48388
rect 11192 48444 11256 48448
rect 11192 48388 11196 48444
rect 11196 48388 11252 48444
rect 11252 48388 11256 48444
rect 11192 48384 11256 48388
rect 20952 48444 21016 48448
rect 20952 48388 20956 48444
rect 20956 48388 21012 48444
rect 21012 48388 21016 48444
rect 20952 48384 21016 48388
rect 21032 48444 21096 48448
rect 21032 48388 21036 48444
rect 21036 48388 21092 48444
rect 21092 48388 21096 48444
rect 21032 48384 21096 48388
rect 21112 48444 21176 48448
rect 21112 48388 21116 48444
rect 21116 48388 21172 48444
rect 21172 48388 21176 48444
rect 21112 48384 21176 48388
rect 21192 48444 21256 48448
rect 21192 48388 21196 48444
rect 21196 48388 21252 48444
rect 21252 48388 21256 48444
rect 21192 48384 21256 48388
rect 15332 48316 15396 48380
rect 21772 48512 21836 48516
rect 21772 48456 21822 48512
rect 21822 48456 21836 48512
rect 21772 48452 21836 48456
rect 19932 47908 19996 47972
rect 5952 47900 6016 47904
rect 5952 47844 5956 47900
rect 5956 47844 6012 47900
rect 6012 47844 6016 47900
rect 5952 47840 6016 47844
rect 6032 47900 6096 47904
rect 6032 47844 6036 47900
rect 6036 47844 6092 47900
rect 6092 47844 6096 47900
rect 6032 47840 6096 47844
rect 6112 47900 6176 47904
rect 6112 47844 6116 47900
rect 6116 47844 6172 47900
rect 6172 47844 6176 47900
rect 6112 47840 6176 47844
rect 6192 47900 6256 47904
rect 6192 47844 6196 47900
rect 6196 47844 6252 47900
rect 6252 47844 6256 47900
rect 6192 47840 6256 47844
rect 15952 47900 16016 47904
rect 15952 47844 15956 47900
rect 15956 47844 16012 47900
rect 16012 47844 16016 47900
rect 15952 47840 16016 47844
rect 16032 47900 16096 47904
rect 16032 47844 16036 47900
rect 16036 47844 16092 47900
rect 16092 47844 16096 47900
rect 16032 47840 16096 47844
rect 16112 47900 16176 47904
rect 16112 47844 16116 47900
rect 16116 47844 16172 47900
rect 16172 47844 16176 47900
rect 16112 47840 16176 47844
rect 16192 47900 16256 47904
rect 16192 47844 16196 47900
rect 16196 47844 16252 47900
rect 16252 47844 16256 47900
rect 16192 47840 16256 47844
rect 25952 47900 26016 47904
rect 25952 47844 25956 47900
rect 25956 47844 26012 47900
rect 26012 47844 26016 47900
rect 25952 47840 26016 47844
rect 26032 47900 26096 47904
rect 26032 47844 26036 47900
rect 26036 47844 26092 47900
rect 26092 47844 26096 47900
rect 26032 47840 26096 47844
rect 26112 47900 26176 47904
rect 26112 47844 26116 47900
rect 26116 47844 26172 47900
rect 26172 47844 26176 47900
rect 26112 47840 26176 47844
rect 26192 47900 26256 47904
rect 26192 47844 26196 47900
rect 26196 47844 26252 47900
rect 26252 47844 26256 47900
rect 26192 47840 26256 47844
rect 23980 47636 24044 47700
rect 10952 47356 11016 47360
rect 10952 47300 10956 47356
rect 10956 47300 11012 47356
rect 11012 47300 11016 47356
rect 10952 47296 11016 47300
rect 11032 47356 11096 47360
rect 11032 47300 11036 47356
rect 11036 47300 11092 47356
rect 11092 47300 11096 47356
rect 11032 47296 11096 47300
rect 11112 47356 11176 47360
rect 11112 47300 11116 47356
rect 11116 47300 11172 47356
rect 11172 47300 11176 47356
rect 11112 47296 11176 47300
rect 11192 47356 11256 47360
rect 11192 47300 11196 47356
rect 11196 47300 11252 47356
rect 11252 47300 11256 47356
rect 11192 47296 11256 47300
rect 20952 47356 21016 47360
rect 20952 47300 20956 47356
rect 20956 47300 21012 47356
rect 21012 47300 21016 47356
rect 20952 47296 21016 47300
rect 21032 47356 21096 47360
rect 21032 47300 21036 47356
rect 21036 47300 21092 47356
rect 21092 47300 21096 47356
rect 21032 47296 21096 47300
rect 21112 47356 21176 47360
rect 21112 47300 21116 47356
rect 21116 47300 21172 47356
rect 21172 47300 21176 47356
rect 21112 47296 21176 47300
rect 21192 47356 21256 47360
rect 21192 47300 21196 47356
rect 21196 47300 21252 47356
rect 21252 47300 21256 47356
rect 21192 47296 21256 47300
rect 9628 46956 9692 47020
rect 15516 46956 15580 47020
rect 16436 47016 16500 47020
rect 16436 46960 16486 47016
rect 16486 46960 16500 47016
rect 16436 46956 16500 46960
rect 5952 46812 6016 46816
rect 5952 46756 5956 46812
rect 5956 46756 6012 46812
rect 6012 46756 6016 46812
rect 5952 46752 6016 46756
rect 6032 46812 6096 46816
rect 6032 46756 6036 46812
rect 6036 46756 6092 46812
rect 6092 46756 6096 46812
rect 6032 46752 6096 46756
rect 6112 46812 6176 46816
rect 6112 46756 6116 46812
rect 6116 46756 6172 46812
rect 6172 46756 6176 46812
rect 6112 46752 6176 46756
rect 6192 46812 6256 46816
rect 6192 46756 6196 46812
rect 6196 46756 6252 46812
rect 6252 46756 6256 46812
rect 6192 46752 6256 46756
rect 15952 46812 16016 46816
rect 15952 46756 15956 46812
rect 15956 46756 16012 46812
rect 16012 46756 16016 46812
rect 15952 46752 16016 46756
rect 16032 46812 16096 46816
rect 16032 46756 16036 46812
rect 16036 46756 16092 46812
rect 16092 46756 16096 46812
rect 16032 46752 16096 46756
rect 16112 46812 16176 46816
rect 16112 46756 16116 46812
rect 16116 46756 16172 46812
rect 16172 46756 16176 46812
rect 16112 46752 16176 46756
rect 16192 46812 16256 46816
rect 16192 46756 16196 46812
rect 16196 46756 16252 46812
rect 16252 46756 16256 46812
rect 16192 46752 16256 46756
rect 25952 46812 26016 46816
rect 25952 46756 25956 46812
rect 25956 46756 26012 46812
rect 26012 46756 26016 46812
rect 25952 46752 26016 46756
rect 26032 46812 26096 46816
rect 26032 46756 26036 46812
rect 26036 46756 26092 46812
rect 26092 46756 26096 46812
rect 26032 46752 26096 46756
rect 26112 46812 26176 46816
rect 26112 46756 26116 46812
rect 26116 46756 26172 46812
rect 26172 46756 26176 46812
rect 26112 46752 26176 46756
rect 26192 46812 26256 46816
rect 26192 46756 26196 46812
rect 26196 46756 26252 46812
rect 26252 46756 26256 46812
rect 26192 46752 26256 46756
rect 20116 46684 20180 46748
rect 10952 46268 11016 46272
rect 10952 46212 10956 46268
rect 10956 46212 11012 46268
rect 11012 46212 11016 46268
rect 10952 46208 11016 46212
rect 11032 46268 11096 46272
rect 11032 46212 11036 46268
rect 11036 46212 11092 46268
rect 11092 46212 11096 46268
rect 11032 46208 11096 46212
rect 11112 46268 11176 46272
rect 11112 46212 11116 46268
rect 11116 46212 11172 46268
rect 11172 46212 11176 46268
rect 11112 46208 11176 46212
rect 11192 46268 11256 46272
rect 11192 46212 11196 46268
rect 11196 46212 11252 46268
rect 11252 46212 11256 46268
rect 11192 46208 11256 46212
rect 20952 46268 21016 46272
rect 20952 46212 20956 46268
rect 20956 46212 21012 46268
rect 21012 46212 21016 46268
rect 20952 46208 21016 46212
rect 21032 46268 21096 46272
rect 21032 46212 21036 46268
rect 21036 46212 21092 46268
rect 21092 46212 21096 46268
rect 21032 46208 21096 46212
rect 21112 46268 21176 46272
rect 21112 46212 21116 46268
rect 21116 46212 21172 46268
rect 21172 46212 21176 46268
rect 21112 46208 21176 46212
rect 21192 46268 21256 46272
rect 21192 46212 21196 46268
rect 21196 46212 21252 46268
rect 21252 46212 21256 46268
rect 21192 46208 21256 46212
rect 5952 45724 6016 45728
rect 5952 45668 5956 45724
rect 5956 45668 6012 45724
rect 6012 45668 6016 45724
rect 5952 45664 6016 45668
rect 6032 45724 6096 45728
rect 6032 45668 6036 45724
rect 6036 45668 6092 45724
rect 6092 45668 6096 45724
rect 6032 45664 6096 45668
rect 6112 45724 6176 45728
rect 6112 45668 6116 45724
rect 6116 45668 6172 45724
rect 6172 45668 6176 45724
rect 6112 45664 6176 45668
rect 6192 45724 6256 45728
rect 6192 45668 6196 45724
rect 6196 45668 6252 45724
rect 6252 45668 6256 45724
rect 6192 45664 6256 45668
rect 15952 45724 16016 45728
rect 15952 45668 15956 45724
rect 15956 45668 16012 45724
rect 16012 45668 16016 45724
rect 15952 45664 16016 45668
rect 16032 45724 16096 45728
rect 16032 45668 16036 45724
rect 16036 45668 16092 45724
rect 16092 45668 16096 45724
rect 16032 45664 16096 45668
rect 16112 45724 16176 45728
rect 16112 45668 16116 45724
rect 16116 45668 16172 45724
rect 16172 45668 16176 45724
rect 16112 45664 16176 45668
rect 16192 45724 16256 45728
rect 16192 45668 16196 45724
rect 16196 45668 16252 45724
rect 16252 45668 16256 45724
rect 16192 45664 16256 45668
rect 25952 45724 26016 45728
rect 25952 45668 25956 45724
rect 25956 45668 26012 45724
rect 26012 45668 26016 45724
rect 25952 45664 26016 45668
rect 26032 45724 26096 45728
rect 26032 45668 26036 45724
rect 26036 45668 26092 45724
rect 26092 45668 26096 45724
rect 26032 45664 26096 45668
rect 26112 45724 26176 45728
rect 26112 45668 26116 45724
rect 26116 45668 26172 45724
rect 26172 45668 26176 45724
rect 26112 45664 26176 45668
rect 26192 45724 26256 45728
rect 26192 45668 26196 45724
rect 26196 45668 26252 45724
rect 26252 45668 26256 45724
rect 26192 45664 26256 45668
rect 20116 45596 20180 45660
rect 25268 45596 25332 45660
rect 10952 45180 11016 45184
rect 10952 45124 10956 45180
rect 10956 45124 11012 45180
rect 11012 45124 11016 45180
rect 10952 45120 11016 45124
rect 11032 45180 11096 45184
rect 11032 45124 11036 45180
rect 11036 45124 11092 45180
rect 11092 45124 11096 45180
rect 11032 45120 11096 45124
rect 11112 45180 11176 45184
rect 11112 45124 11116 45180
rect 11116 45124 11172 45180
rect 11172 45124 11176 45180
rect 11112 45120 11176 45124
rect 11192 45180 11256 45184
rect 11192 45124 11196 45180
rect 11196 45124 11252 45180
rect 11252 45124 11256 45180
rect 11192 45120 11256 45124
rect 20952 45180 21016 45184
rect 20952 45124 20956 45180
rect 20956 45124 21012 45180
rect 21012 45124 21016 45180
rect 20952 45120 21016 45124
rect 21032 45180 21096 45184
rect 21032 45124 21036 45180
rect 21036 45124 21092 45180
rect 21092 45124 21096 45180
rect 21032 45120 21096 45124
rect 21112 45180 21176 45184
rect 21112 45124 21116 45180
rect 21116 45124 21172 45180
rect 21172 45124 21176 45180
rect 21112 45120 21176 45124
rect 21192 45180 21256 45184
rect 21192 45124 21196 45180
rect 21196 45124 21252 45180
rect 21252 45124 21256 45180
rect 21192 45120 21256 45124
rect 20300 44840 20364 44844
rect 20300 44784 20350 44840
rect 20350 44784 20364 44840
rect 20300 44780 20364 44784
rect 23060 44644 23124 44708
rect 5952 44636 6016 44640
rect 5952 44580 5956 44636
rect 5956 44580 6012 44636
rect 6012 44580 6016 44636
rect 5952 44576 6016 44580
rect 6032 44636 6096 44640
rect 6032 44580 6036 44636
rect 6036 44580 6092 44636
rect 6092 44580 6096 44636
rect 6032 44576 6096 44580
rect 6112 44636 6176 44640
rect 6112 44580 6116 44636
rect 6116 44580 6172 44636
rect 6172 44580 6176 44636
rect 6112 44576 6176 44580
rect 6192 44636 6256 44640
rect 6192 44580 6196 44636
rect 6196 44580 6252 44636
rect 6252 44580 6256 44636
rect 6192 44576 6256 44580
rect 15952 44636 16016 44640
rect 15952 44580 15956 44636
rect 15956 44580 16012 44636
rect 16012 44580 16016 44636
rect 15952 44576 16016 44580
rect 16032 44636 16096 44640
rect 16032 44580 16036 44636
rect 16036 44580 16092 44636
rect 16092 44580 16096 44636
rect 16032 44576 16096 44580
rect 16112 44636 16176 44640
rect 16112 44580 16116 44636
rect 16116 44580 16172 44636
rect 16172 44580 16176 44636
rect 16112 44576 16176 44580
rect 16192 44636 16256 44640
rect 16192 44580 16196 44636
rect 16196 44580 16252 44636
rect 16252 44580 16256 44636
rect 16192 44576 16256 44580
rect 25952 44636 26016 44640
rect 25952 44580 25956 44636
rect 25956 44580 26012 44636
rect 26012 44580 26016 44636
rect 25952 44576 26016 44580
rect 26032 44636 26096 44640
rect 26032 44580 26036 44636
rect 26036 44580 26092 44636
rect 26092 44580 26096 44636
rect 26032 44576 26096 44580
rect 26112 44636 26176 44640
rect 26112 44580 26116 44636
rect 26116 44580 26172 44636
rect 26172 44580 26176 44636
rect 26112 44576 26176 44580
rect 26192 44636 26256 44640
rect 26192 44580 26196 44636
rect 26196 44580 26252 44636
rect 26252 44580 26256 44636
rect 26192 44576 26256 44580
rect 3188 44508 3252 44572
rect 10952 44092 11016 44096
rect 10952 44036 10956 44092
rect 10956 44036 11012 44092
rect 11012 44036 11016 44092
rect 10952 44032 11016 44036
rect 11032 44092 11096 44096
rect 11032 44036 11036 44092
rect 11036 44036 11092 44092
rect 11092 44036 11096 44092
rect 11032 44032 11096 44036
rect 11112 44092 11176 44096
rect 11112 44036 11116 44092
rect 11116 44036 11172 44092
rect 11172 44036 11176 44092
rect 11112 44032 11176 44036
rect 11192 44092 11256 44096
rect 11192 44036 11196 44092
rect 11196 44036 11252 44092
rect 11252 44036 11256 44092
rect 11192 44032 11256 44036
rect 20952 44092 21016 44096
rect 20952 44036 20956 44092
rect 20956 44036 21012 44092
rect 21012 44036 21016 44092
rect 20952 44032 21016 44036
rect 21032 44092 21096 44096
rect 21032 44036 21036 44092
rect 21036 44036 21092 44092
rect 21092 44036 21096 44092
rect 21032 44032 21096 44036
rect 21112 44092 21176 44096
rect 21112 44036 21116 44092
rect 21116 44036 21172 44092
rect 21172 44036 21176 44092
rect 21112 44032 21176 44036
rect 21192 44092 21256 44096
rect 21192 44036 21196 44092
rect 21196 44036 21252 44092
rect 21252 44036 21256 44092
rect 21192 44032 21256 44036
rect 5952 43548 6016 43552
rect 5952 43492 5956 43548
rect 5956 43492 6012 43548
rect 6012 43492 6016 43548
rect 5952 43488 6016 43492
rect 6032 43548 6096 43552
rect 6032 43492 6036 43548
rect 6036 43492 6092 43548
rect 6092 43492 6096 43548
rect 6032 43488 6096 43492
rect 6112 43548 6176 43552
rect 6112 43492 6116 43548
rect 6116 43492 6172 43548
rect 6172 43492 6176 43548
rect 6112 43488 6176 43492
rect 6192 43548 6256 43552
rect 6192 43492 6196 43548
rect 6196 43492 6252 43548
rect 6252 43492 6256 43548
rect 6192 43488 6256 43492
rect 15952 43548 16016 43552
rect 15952 43492 15956 43548
rect 15956 43492 16012 43548
rect 16012 43492 16016 43548
rect 15952 43488 16016 43492
rect 16032 43548 16096 43552
rect 16032 43492 16036 43548
rect 16036 43492 16092 43548
rect 16092 43492 16096 43548
rect 16032 43488 16096 43492
rect 16112 43548 16176 43552
rect 16112 43492 16116 43548
rect 16116 43492 16172 43548
rect 16172 43492 16176 43548
rect 16112 43488 16176 43492
rect 16192 43548 16256 43552
rect 16192 43492 16196 43548
rect 16196 43492 16252 43548
rect 16252 43492 16256 43548
rect 16192 43488 16256 43492
rect 25952 43548 26016 43552
rect 25952 43492 25956 43548
rect 25956 43492 26012 43548
rect 26012 43492 26016 43548
rect 25952 43488 26016 43492
rect 26032 43548 26096 43552
rect 26032 43492 26036 43548
rect 26036 43492 26092 43548
rect 26092 43492 26096 43548
rect 26032 43488 26096 43492
rect 26112 43548 26176 43552
rect 26112 43492 26116 43548
rect 26116 43492 26172 43548
rect 26172 43492 26176 43548
rect 26112 43488 26176 43492
rect 26192 43548 26256 43552
rect 26192 43492 26196 43548
rect 26196 43492 26252 43548
rect 26252 43492 26256 43548
rect 26192 43488 26256 43492
rect 10952 43004 11016 43008
rect 10952 42948 10956 43004
rect 10956 42948 11012 43004
rect 11012 42948 11016 43004
rect 10952 42944 11016 42948
rect 11032 43004 11096 43008
rect 11032 42948 11036 43004
rect 11036 42948 11092 43004
rect 11092 42948 11096 43004
rect 11032 42944 11096 42948
rect 11112 43004 11176 43008
rect 11112 42948 11116 43004
rect 11116 42948 11172 43004
rect 11172 42948 11176 43004
rect 11112 42944 11176 42948
rect 11192 43004 11256 43008
rect 11192 42948 11196 43004
rect 11196 42948 11252 43004
rect 11252 42948 11256 43004
rect 11192 42944 11256 42948
rect 20952 43004 21016 43008
rect 20952 42948 20956 43004
rect 20956 42948 21012 43004
rect 21012 42948 21016 43004
rect 20952 42944 21016 42948
rect 21032 43004 21096 43008
rect 21032 42948 21036 43004
rect 21036 42948 21092 43004
rect 21092 42948 21096 43004
rect 21032 42944 21096 42948
rect 21112 43004 21176 43008
rect 21112 42948 21116 43004
rect 21116 42948 21172 43004
rect 21172 42948 21176 43004
rect 21112 42944 21176 42948
rect 21192 43004 21256 43008
rect 21192 42948 21196 43004
rect 21196 42948 21252 43004
rect 21252 42948 21256 43004
rect 21192 42944 21256 42948
rect 13676 42876 13740 42940
rect 5952 42460 6016 42464
rect 5952 42404 5956 42460
rect 5956 42404 6012 42460
rect 6012 42404 6016 42460
rect 5952 42400 6016 42404
rect 6032 42460 6096 42464
rect 6032 42404 6036 42460
rect 6036 42404 6092 42460
rect 6092 42404 6096 42460
rect 6032 42400 6096 42404
rect 6112 42460 6176 42464
rect 6112 42404 6116 42460
rect 6116 42404 6172 42460
rect 6172 42404 6176 42460
rect 6112 42400 6176 42404
rect 6192 42460 6256 42464
rect 6192 42404 6196 42460
rect 6196 42404 6252 42460
rect 6252 42404 6256 42460
rect 6192 42400 6256 42404
rect 15952 42460 16016 42464
rect 15952 42404 15956 42460
rect 15956 42404 16012 42460
rect 16012 42404 16016 42460
rect 15952 42400 16016 42404
rect 16032 42460 16096 42464
rect 16032 42404 16036 42460
rect 16036 42404 16092 42460
rect 16092 42404 16096 42460
rect 16032 42400 16096 42404
rect 16112 42460 16176 42464
rect 16112 42404 16116 42460
rect 16116 42404 16172 42460
rect 16172 42404 16176 42460
rect 16112 42400 16176 42404
rect 16192 42460 16256 42464
rect 16192 42404 16196 42460
rect 16196 42404 16252 42460
rect 16252 42404 16256 42460
rect 16192 42400 16256 42404
rect 25952 42460 26016 42464
rect 25952 42404 25956 42460
rect 25956 42404 26012 42460
rect 26012 42404 26016 42460
rect 25952 42400 26016 42404
rect 26032 42460 26096 42464
rect 26032 42404 26036 42460
rect 26036 42404 26092 42460
rect 26092 42404 26096 42460
rect 26032 42400 26096 42404
rect 26112 42460 26176 42464
rect 26112 42404 26116 42460
rect 26116 42404 26172 42460
rect 26172 42404 26176 42460
rect 26112 42400 26176 42404
rect 26192 42460 26256 42464
rect 26192 42404 26196 42460
rect 26196 42404 26252 42460
rect 26252 42404 26256 42460
rect 26192 42400 26256 42404
rect 19932 42392 19996 42396
rect 19932 42336 19946 42392
rect 19946 42336 19996 42392
rect 19932 42332 19996 42336
rect 12388 42060 12452 42124
rect 20116 41984 20180 41988
rect 20116 41928 20130 41984
rect 20130 41928 20180 41984
rect 20116 41924 20180 41928
rect 10952 41916 11016 41920
rect 10952 41860 10956 41916
rect 10956 41860 11012 41916
rect 11012 41860 11016 41916
rect 10952 41856 11016 41860
rect 11032 41916 11096 41920
rect 11032 41860 11036 41916
rect 11036 41860 11092 41916
rect 11092 41860 11096 41916
rect 11032 41856 11096 41860
rect 11112 41916 11176 41920
rect 11112 41860 11116 41916
rect 11116 41860 11172 41916
rect 11172 41860 11176 41916
rect 11112 41856 11176 41860
rect 11192 41916 11256 41920
rect 11192 41860 11196 41916
rect 11196 41860 11252 41916
rect 11252 41860 11256 41916
rect 11192 41856 11256 41860
rect 20952 41916 21016 41920
rect 20952 41860 20956 41916
rect 20956 41860 21012 41916
rect 21012 41860 21016 41916
rect 20952 41856 21016 41860
rect 21032 41916 21096 41920
rect 21032 41860 21036 41916
rect 21036 41860 21092 41916
rect 21092 41860 21096 41916
rect 21032 41856 21096 41860
rect 21112 41916 21176 41920
rect 21112 41860 21116 41916
rect 21116 41860 21172 41916
rect 21172 41860 21176 41916
rect 21112 41856 21176 41860
rect 21192 41916 21256 41920
rect 21192 41860 21196 41916
rect 21196 41860 21252 41916
rect 21252 41860 21256 41916
rect 21192 41856 21256 41860
rect 12940 41788 13004 41852
rect 20484 41516 20548 41580
rect 24716 41516 24780 41580
rect 20484 41380 20548 41444
rect 23060 41380 23124 41444
rect 5952 41372 6016 41376
rect 5952 41316 5956 41372
rect 5956 41316 6012 41372
rect 6012 41316 6016 41372
rect 5952 41312 6016 41316
rect 6032 41372 6096 41376
rect 6032 41316 6036 41372
rect 6036 41316 6092 41372
rect 6092 41316 6096 41372
rect 6032 41312 6096 41316
rect 6112 41372 6176 41376
rect 6112 41316 6116 41372
rect 6116 41316 6172 41372
rect 6172 41316 6176 41372
rect 6112 41312 6176 41316
rect 6192 41372 6256 41376
rect 6192 41316 6196 41372
rect 6196 41316 6252 41372
rect 6252 41316 6256 41372
rect 6192 41312 6256 41316
rect 15952 41372 16016 41376
rect 15952 41316 15956 41372
rect 15956 41316 16012 41372
rect 16012 41316 16016 41372
rect 15952 41312 16016 41316
rect 16032 41372 16096 41376
rect 16032 41316 16036 41372
rect 16036 41316 16092 41372
rect 16092 41316 16096 41372
rect 16032 41312 16096 41316
rect 16112 41372 16176 41376
rect 16112 41316 16116 41372
rect 16116 41316 16172 41372
rect 16172 41316 16176 41372
rect 16112 41312 16176 41316
rect 16192 41372 16256 41376
rect 16192 41316 16196 41372
rect 16196 41316 16252 41372
rect 16252 41316 16256 41372
rect 16192 41312 16256 41316
rect 25952 41372 26016 41376
rect 25952 41316 25956 41372
rect 25956 41316 26012 41372
rect 26012 41316 26016 41372
rect 25952 41312 26016 41316
rect 26032 41372 26096 41376
rect 26032 41316 26036 41372
rect 26036 41316 26092 41372
rect 26092 41316 26096 41372
rect 26032 41312 26096 41316
rect 26112 41372 26176 41376
rect 26112 41316 26116 41372
rect 26116 41316 26172 41372
rect 26172 41316 26176 41372
rect 26112 41312 26176 41316
rect 26192 41372 26256 41376
rect 26192 41316 26196 41372
rect 26196 41316 26252 41372
rect 26252 41316 26256 41372
rect 26192 41312 26256 41316
rect 20484 41168 20548 41172
rect 20484 41112 20534 41168
rect 20534 41112 20548 41168
rect 20484 41108 20548 41112
rect 20668 41108 20732 41172
rect 20484 40836 20548 40900
rect 10952 40828 11016 40832
rect 10952 40772 10956 40828
rect 10956 40772 11012 40828
rect 11012 40772 11016 40828
rect 10952 40768 11016 40772
rect 11032 40828 11096 40832
rect 11032 40772 11036 40828
rect 11036 40772 11092 40828
rect 11092 40772 11096 40828
rect 11032 40768 11096 40772
rect 11112 40828 11176 40832
rect 11112 40772 11116 40828
rect 11116 40772 11172 40828
rect 11172 40772 11176 40828
rect 11112 40768 11176 40772
rect 11192 40828 11256 40832
rect 11192 40772 11196 40828
rect 11196 40772 11252 40828
rect 11252 40772 11256 40828
rect 11192 40768 11256 40772
rect 20952 40828 21016 40832
rect 20952 40772 20956 40828
rect 20956 40772 21012 40828
rect 21012 40772 21016 40828
rect 20952 40768 21016 40772
rect 21032 40828 21096 40832
rect 21032 40772 21036 40828
rect 21036 40772 21092 40828
rect 21092 40772 21096 40828
rect 21032 40768 21096 40772
rect 21112 40828 21176 40832
rect 21112 40772 21116 40828
rect 21116 40772 21172 40828
rect 21172 40772 21176 40828
rect 21112 40768 21176 40772
rect 21192 40828 21256 40832
rect 21192 40772 21196 40828
rect 21196 40772 21252 40828
rect 21252 40772 21256 40828
rect 21192 40768 21256 40772
rect 23980 40836 24044 40900
rect 5952 40284 6016 40288
rect 5952 40228 5956 40284
rect 5956 40228 6012 40284
rect 6012 40228 6016 40284
rect 5952 40224 6016 40228
rect 6032 40284 6096 40288
rect 6032 40228 6036 40284
rect 6036 40228 6092 40284
rect 6092 40228 6096 40284
rect 6032 40224 6096 40228
rect 6112 40284 6176 40288
rect 6112 40228 6116 40284
rect 6116 40228 6172 40284
rect 6172 40228 6176 40284
rect 6112 40224 6176 40228
rect 6192 40284 6256 40288
rect 6192 40228 6196 40284
rect 6196 40228 6252 40284
rect 6252 40228 6256 40284
rect 6192 40224 6256 40228
rect 15952 40284 16016 40288
rect 15952 40228 15956 40284
rect 15956 40228 16012 40284
rect 16012 40228 16016 40284
rect 15952 40224 16016 40228
rect 16032 40284 16096 40288
rect 16032 40228 16036 40284
rect 16036 40228 16092 40284
rect 16092 40228 16096 40284
rect 16032 40224 16096 40228
rect 16112 40284 16176 40288
rect 16112 40228 16116 40284
rect 16116 40228 16172 40284
rect 16172 40228 16176 40284
rect 16112 40224 16176 40228
rect 16192 40284 16256 40288
rect 16192 40228 16196 40284
rect 16196 40228 16252 40284
rect 16252 40228 16256 40284
rect 16192 40224 16256 40228
rect 25952 40284 26016 40288
rect 25952 40228 25956 40284
rect 25956 40228 26012 40284
rect 26012 40228 26016 40284
rect 25952 40224 26016 40228
rect 26032 40284 26096 40288
rect 26032 40228 26036 40284
rect 26036 40228 26092 40284
rect 26092 40228 26096 40284
rect 26032 40224 26096 40228
rect 26112 40284 26176 40288
rect 26112 40228 26116 40284
rect 26116 40228 26172 40284
rect 26172 40228 26176 40284
rect 26112 40224 26176 40228
rect 26192 40284 26256 40288
rect 26192 40228 26196 40284
rect 26196 40228 26252 40284
rect 26252 40228 26256 40284
rect 26192 40224 26256 40228
rect 13492 39748 13556 39812
rect 10952 39740 11016 39744
rect 10952 39684 10956 39740
rect 10956 39684 11012 39740
rect 11012 39684 11016 39740
rect 10952 39680 11016 39684
rect 11032 39740 11096 39744
rect 11032 39684 11036 39740
rect 11036 39684 11092 39740
rect 11092 39684 11096 39740
rect 11032 39680 11096 39684
rect 11112 39740 11176 39744
rect 11112 39684 11116 39740
rect 11116 39684 11172 39740
rect 11172 39684 11176 39740
rect 11112 39680 11176 39684
rect 11192 39740 11256 39744
rect 11192 39684 11196 39740
rect 11196 39684 11252 39740
rect 11252 39684 11256 39740
rect 11192 39680 11256 39684
rect 20952 39740 21016 39744
rect 20952 39684 20956 39740
rect 20956 39684 21012 39740
rect 21012 39684 21016 39740
rect 20952 39680 21016 39684
rect 21032 39740 21096 39744
rect 21032 39684 21036 39740
rect 21036 39684 21092 39740
rect 21092 39684 21096 39740
rect 21032 39680 21096 39684
rect 21112 39740 21176 39744
rect 21112 39684 21116 39740
rect 21116 39684 21172 39740
rect 21172 39684 21176 39740
rect 21112 39680 21176 39684
rect 21192 39740 21256 39744
rect 21192 39684 21196 39740
rect 21196 39684 21252 39740
rect 21252 39684 21256 39740
rect 21192 39680 21256 39684
rect 12756 39612 12820 39676
rect 13308 39612 13372 39676
rect 13308 39340 13372 39404
rect 5952 39196 6016 39200
rect 5952 39140 5956 39196
rect 5956 39140 6012 39196
rect 6012 39140 6016 39196
rect 5952 39136 6016 39140
rect 6032 39196 6096 39200
rect 6032 39140 6036 39196
rect 6036 39140 6092 39196
rect 6092 39140 6096 39196
rect 6032 39136 6096 39140
rect 6112 39196 6176 39200
rect 6112 39140 6116 39196
rect 6116 39140 6172 39196
rect 6172 39140 6176 39196
rect 6112 39136 6176 39140
rect 6192 39196 6256 39200
rect 6192 39140 6196 39196
rect 6196 39140 6252 39196
rect 6252 39140 6256 39196
rect 6192 39136 6256 39140
rect 15952 39196 16016 39200
rect 15952 39140 15956 39196
rect 15956 39140 16012 39196
rect 16012 39140 16016 39196
rect 15952 39136 16016 39140
rect 16032 39196 16096 39200
rect 16032 39140 16036 39196
rect 16036 39140 16092 39196
rect 16092 39140 16096 39196
rect 16032 39136 16096 39140
rect 16112 39196 16176 39200
rect 16112 39140 16116 39196
rect 16116 39140 16172 39196
rect 16172 39140 16176 39196
rect 16112 39136 16176 39140
rect 16192 39196 16256 39200
rect 16192 39140 16196 39196
rect 16196 39140 16252 39196
rect 16252 39140 16256 39196
rect 16192 39136 16256 39140
rect 24716 39204 24780 39268
rect 25952 39196 26016 39200
rect 25952 39140 25956 39196
rect 25956 39140 26012 39196
rect 26012 39140 26016 39196
rect 25952 39136 26016 39140
rect 26032 39196 26096 39200
rect 26032 39140 26036 39196
rect 26036 39140 26092 39196
rect 26092 39140 26096 39196
rect 26032 39136 26096 39140
rect 26112 39196 26176 39200
rect 26112 39140 26116 39196
rect 26116 39140 26172 39196
rect 26172 39140 26176 39196
rect 26112 39136 26176 39140
rect 26192 39196 26256 39200
rect 26192 39140 26196 39196
rect 26196 39140 26252 39196
rect 26252 39140 26256 39196
rect 26192 39136 26256 39140
rect 10952 38652 11016 38656
rect 10952 38596 10956 38652
rect 10956 38596 11012 38652
rect 11012 38596 11016 38652
rect 10952 38592 11016 38596
rect 11032 38652 11096 38656
rect 11032 38596 11036 38652
rect 11036 38596 11092 38652
rect 11092 38596 11096 38652
rect 11032 38592 11096 38596
rect 11112 38652 11176 38656
rect 11112 38596 11116 38652
rect 11116 38596 11172 38652
rect 11172 38596 11176 38652
rect 11112 38592 11176 38596
rect 11192 38652 11256 38656
rect 11192 38596 11196 38652
rect 11196 38596 11252 38652
rect 11252 38596 11256 38652
rect 11192 38592 11256 38596
rect 13124 38388 13188 38452
rect 21772 38660 21836 38724
rect 20952 38652 21016 38656
rect 20952 38596 20956 38652
rect 20956 38596 21012 38652
rect 21012 38596 21016 38652
rect 20952 38592 21016 38596
rect 21032 38652 21096 38656
rect 21032 38596 21036 38652
rect 21036 38596 21092 38652
rect 21092 38596 21096 38652
rect 21032 38592 21096 38596
rect 21112 38652 21176 38656
rect 21112 38596 21116 38652
rect 21116 38596 21172 38652
rect 21172 38596 21176 38652
rect 21112 38592 21176 38596
rect 21192 38652 21256 38656
rect 21192 38596 21196 38652
rect 21196 38596 21252 38652
rect 21252 38596 21256 38652
rect 21192 38592 21256 38596
rect 25452 38584 25516 38588
rect 25452 38528 25502 38584
rect 25502 38528 25516 38584
rect 25452 38524 25516 38528
rect 24348 38388 24412 38452
rect 25452 38388 25516 38452
rect 5952 38108 6016 38112
rect 5952 38052 5956 38108
rect 5956 38052 6012 38108
rect 6012 38052 6016 38108
rect 5952 38048 6016 38052
rect 6032 38108 6096 38112
rect 6032 38052 6036 38108
rect 6036 38052 6092 38108
rect 6092 38052 6096 38108
rect 6032 38048 6096 38052
rect 6112 38108 6176 38112
rect 6112 38052 6116 38108
rect 6116 38052 6172 38108
rect 6172 38052 6176 38108
rect 6112 38048 6176 38052
rect 6192 38108 6256 38112
rect 6192 38052 6196 38108
rect 6196 38052 6252 38108
rect 6252 38052 6256 38108
rect 6192 38048 6256 38052
rect 15952 38108 16016 38112
rect 15952 38052 15956 38108
rect 15956 38052 16012 38108
rect 16012 38052 16016 38108
rect 15952 38048 16016 38052
rect 16032 38108 16096 38112
rect 16032 38052 16036 38108
rect 16036 38052 16092 38108
rect 16092 38052 16096 38108
rect 16032 38048 16096 38052
rect 16112 38108 16176 38112
rect 16112 38052 16116 38108
rect 16116 38052 16172 38108
rect 16172 38052 16176 38108
rect 16112 38048 16176 38052
rect 16192 38108 16256 38112
rect 16192 38052 16196 38108
rect 16196 38052 16252 38108
rect 16252 38052 16256 38108
rect 16192 38048 16256 38052
rect 25952 38108 26016 38112
rect 25952 38052 25956 38108
rect 25956 38052 26012 38108
rect 26012 38052 26016 38108
rect 25952 38048 26016 38052
rect 26032 38108 26096 38112
rect 26032 38052 26036 38108
rect 26036 38052 26092 38108
rect 26092 38052 26096 38108
rect 26032 38048 26096 38052
rect 26112 38108 26176 38112
rect 26112 38052 26116 38108
rect 26116 38052 26172 38108
rect 26172 38052 26176 38108
rect 26112 38048 26176 38052
rect 26192 38108 26256 38112
rect 26192 38052 26196 38108
rect 26196 38052 26252 38108
rect 26252 38052 26256 38108
rect 26192 38048 26256 38052
rect 10364 37708 10428 37772
rect 9812 37632 9876 37636
rect 19380 37708 19444 37772
rect 9812 37576 9862 37632
rect 9862 37576 9876 37632
rect 9812 37572 9876 37576
rect 14596 37572 14660 37636
rect 10952 37564 11016 37568
rect 10952 37508 10956 37564
rect 10956 37508 11012 37564
rect 11012 37508 11016 37564
rect 10952 37504 11016 37508
rect 11032 37564 11096 37568
rect 11032 37508 11036 37564
rect 11036 37508 11092 37564
rect 11092 37508 11096 37564
rect 11032 37504 11096 37508
rect 11112 37564 11176 37568
rect 11112 37508 11116 37564
rect 11116 37508 11172 37564
rect 11172 37508 11176 37564
rect 11112 37504 11176 37508
rect 11192 37564 11256 37568
rect 11192 37508 11196 37564
rect 11196 37508 11252 37564
rect 11252 37508 11256 37564
rect 11192 37504 11256 37508
rect 20952 37564 21016 37568
rect 20952 37508 20956 37564
rect 20956 37508 21012 37564
rect 21012 37508 21016 37564
rect 20952 37504 21016 37508
rect 21032 37564 21096 37568
rect 21032 37508 21036 37564
rect 21036 37508 21092 37564
rect 21092 37508 21096 37564
rect 21032 37504 21096 37508
rect 21112 37564 21176 37568
rect 21112 37508 21116 37564
rect 21116 37508 21172 37564
rect 21172 37508 21176 37564
rect 21112 37504 21176 37508
rect 21192 37564 21256 37568
rect 21192 37508 21196 37564
rect 21196 37508 21252 37564
rect 21252 37508 21256 37564
rect 21192 37504 21256 37508
rect 16804 37436 16868 37500
rect 9628 37300 9692 37364
rect 10180 37300 10244 37364
rect 16620 37164 16684 37228
rect 10548 37028 10612 37092
rect 23796 37028 23860 37092
rect 5952 37020 6016 37024
rect 5952 36964 5956 37020
rect 5956 36964 6012 37020
rect 6012 36964 6016 37020
rect 5952 36960 6016 36964
rect 6032 37020 6096 37024
rect 6032 36964 6036 37020
rect 6036 36964 6092 37020
rect 6092 36964 6096 37020
rect 6032 36960 6096 36964
rect 6112 37020 6176 37024
rect 6112 36964 6116 37020
rect 6116 36964 6172 37020
rect 6172 36964 6176 37020
rect 6112 36960 6176 36964
rect 6192 37020 6256 37024
rect 6192 36964 6196 37020
rect 6196 36964 6252 37020
rect 6252 36964 6256 37020
rect 6192 36960 6256 36964
rect 15952 37020 16016 37024
rect 15952 36964 15956 37020
rect 15956 36964 16012 37020
rect 16012 36964 16016 37020
rect 15952 36960 16016 36964
rect 16032 37020 16096 37024
rect 16032 36964 16036 37020
rect 16036 36964 16092 37020
rect 16092 36964 16096 37020
rect 16032 36960 16096 36964
rect 16112 37020 16176 37024
rect 16112 36964 16116 37020
rect 16116 36964 16172 37020
rect 16172 36964 16176 37020
rect 16112 36960 16176 36964
rect 16192 37020 16256 37024
rect 16192 36964 16196 37020
rect 16196 36964 16252 37020
rect 16252 36964 16256 37020
rect 16192 36960 16256 36964
rect 25952 37020 26016 37024
rect 25952 36964 25956 37020
rect 25956 36964 26012 37020
rect 26012 36964 26016 37020
rect 25952 36960 26016 36964
rect 26032 37020 26096 37024
rect 26032 36964 26036 37020
rect 26036 36964 26092 37020
rect 26092 36964 26096 37020
rect 26032 36960 26096 36964
rect 26112 37020 26176 37024
rect 26112 36964 26116 37020
rect 26116 36964 26172 37020
rect 26172 36964 26176 37020
rect 26112 36960 26176 36964
rect 26192 37020 26256 37024
rect 26192 36964 26196 37020
rect 26196 36964 26252 37020
rect 26252 36964 26256 37020
rect 26192 36960 26256 36964
rect 10952 36476 11016 36480
rect 10952 36420 10956 36476
rect 10956 36420 11012 36476
rect 11012 36420 11016 36476
rect 10952 36416 11016 36420
rect 11032 36476 11096 36480
rect 11032 36420 11036 36476
rect 11036 36420 11092 36476
rect 11092 36420 11096 36476
rect 11032 36416 11096 36420
rect 11112 36476 11176 36480
rect 11112 36420 11116 36476
rect 11116 36420 11172 36476
rect 11172 36420 11176 36476
rect 11112 36416 11176 36420
rect 11192 36476 11256 36480
rect 11192 36420 11196 36476
rect 11196 36420 11252 36476
rect 11252 36420 11256 36476
rect 11192 36416 11256 36420
rect 20952 36476 21016 36480
rect 20952 36420 20956 36476
rect 20956 36420 21012 36476
rect 21012 36420 21016 36476
rect 20952 36416 21016 36420
rect 21032 36476 21096 36480
rect 21032 36420 21036 36476
rect 21036 36420 21092 36476
rect 21092 36420 21096 36476
rect 21032 36416 21096 36420
rect 21112 36476 21176 36480
rect 21112 36420 21116 36476
rect 21116 36420 21172 36476
rect 21172 36420 21176 36476
rect 21112 36416 21176 36420
rect 21192 36476 21256 36480
rect 21192 36420 21196 36476
rect 21196 36420 21252 36476
rect 21252 36420 21256 36476
rect 21192 36416 21256 36420
rect 16620 36348 16684 36412
rect 21956 36348 22020 36412
rect 9628 36000 9692 36004
rect 9628 35944 9678 36000
rect 9678 35944 9692 36000
rect 9628 35940 9692 35944
rect 5952 35932 6016 35936
rect 5952 35876 5956 35932
rect 5956 35876 6012 35932
rect 6012 35876 6016 35932
rect 5952 35872 6016 35876
rect 6032 35932 6096 35936
rect 6032 35876 6036 35932
rect 6036 35876 6092 35932
rect 6092 35876 6096 35932
rect 6032 35872 6096 35876
rect 6112 35932 6176 35936
rect 6112 35876 6116 35932
rect 6116 35876 6172 35932
rect 6172 35876 6176 35932
rect 6112 35872 6176 35876
rect 6192 35932 6256 35936
rect 6192 35876 6196 35932
rect 6196 35876 6252 35932
rect 6252 35876 6256 35932
rect 6192 35872 6256 35876
rect 11652 35940 11716 36004
rect 16988 35940 17052 36004
rect 15952 35932 16016 35936
rect 15952 35876 15956 35932
rect 15956 35876 16012 35932
rect 16012 35876 16016 35932
rect 15952 35872 16016 35876
rect 16032 35932 16096 35936
rect 16032 35876 16036 35932
rect 16036 35876 16092 35932
rect 16092 35876 16096 35932
rect 16032 35872 16096 35876
rect 16112 35932 16176 35936
rect 16112 35876 16116 35932
rect 16116 35876 16172 35932
rect 16172 35876 16176 35932
rect 16112 35872 16176 35876
rect 16192 35932 16256 35936
rect 16192 35876 16196 35932
rect 16196 35876 16252 35932
rect 16252 35876 16256 35932
rect 16192 35872 16256 35876
rect 25952 35932 26016 35936
rect 25952 35876 25956 35932
rect 25956 35876 26012 35932
rect 26012 35876 26016 35932
rect 25952 35872 26016 35876
rect 26032 35932 26096 35936
rect 26032 35876 26036 35932
rect 26036 35876 26092 35932
rect 26092 35876 26096 35932
rect 26032 35872 26096 35876
rect 26112 35932 26176 35936
rect 26112 35876 26116 35932
rect 26116 35876 26172 35932
rect 26172 35876 26176 35932
rect 26112 35872 26176 35876
rect 26192 35932 26256 35936
rect 26192 35876 26196 35932
rect 26196 35876 26252 35932
rect 26252 35876 26256 35932
rect 26192 35872 26256 35876
rect 12204 35864 12268 35868
rect 12204 35808 12218 35864
rect 12218 35808 12268 35864
rect 12204 35804 12268 35808
rect 21588 35864 21652 35868
rect 21588 35808 21602 35864
rect 21602 35808 21652 35864
rect 21588 35804 21652 35808
rect 3740 35668 3804 35732
rect 9260 35668 9324 35732
rect 10732 35396 10796 35460
rect 14044 35396 14108 35460
rect 16620 35396 16684 35460
rect 10952 35388 11016 35392
rect 10952 35332 10956 35388
rect 10956 35332 11012 35388
rect 11012 35332 11016 35388
rect 10952 35328 11016 35332
rect 11032 35388 11096 35392
rect 11032 35332 11036 35388
rect 11036 35332 11092 35388
rect 11092 35332 11096 35388
rect 11032 35328 11096 35332
rect 11112 35388 11176 35392
rect 11112 35332 11116 35388
rect 11116 35332 11172 35388
rect 11172 35332 11176 35388
rect 11112 35328 11176 35332
rect 11192 35388 11256 35392
rect 11192 35332 11196 35388
rect 11196 35332 11252 35388
rect 11252 35332 11256 35388
rect 11192 35328 11256 35332
rect 20952 35388 21016 35392
rect 20952 35332 20956 35388
rect 20956 35332 21012 35388
rect 21012 35332 21016 35388
rect 20952 35328 21016 35332
rect 21032 35388 21096 35392
rect 21032 35332 21036 35388
rect 21036 35332 21092 35388
rect 21092 35332 21096 35388
rect 21032 35328 21096 35332
rect 21112 35388 21176 35392
rect 21112 35332 21116 35388
rect 21116 35332 21172 35388
rect 21172 35332 21176 35388
rect 21112 35328 21176 35332
rect 21192 35388 21256 35392
rect 21192 35332 21196 35388
rect 21196 35332 21252 35388
rect 21252 35332 21256 35388
rect 21192 35328 21256 35332
rect 7420 35260 7484 35324
rect 13308 35124 13372 35188
rect 25452 34988 25516 35052
rect 9076 34912 9140 34916
rect 9076 34856 9126 34912
rect 9126 34856 9140 34912
rect 9076 34852 9140 34856
rect 5952 34844 6016 34848
rect 5952 34788 5956 34844
rect 5956 34788 6012 34844
rect 6012 34788 6016 34844
rect 5952 34784 6016 34788
rect 6032 34844 6096 34848
rect 6032 34788 6036 34844
rect 6036 34788 6092 34844
rect 6092 34788 6096 34844
rect 6032 34784 6096 34788
rect 6112 34844 6176 34848
rect 6112 34788 6116 34844
rect 6116 34788 6172 34844
rect 6172 34788 6176 34844
rect 6112 34784 6176 34788
rect 6192 34844 6256 34848
rect 6192 34788 6196 34844
rect 6196 34788 6252 34844
rect 6252 34788 6256 34844
rect 6192 34784 6256 34788
rect 15952 34844 16016 34848
rect 15952 34788 15956 34844
rect 15956 34788 16012 34844
rect 16012 34788 16016 34844
rect 15952 34784 16016 34788
rect 16032 34844 16096 34848
rect 16032 34788 16036 34844
rect 16036 34788 16092 34844
rect 16092 34788 16096 34844
rect 16032 34784 16096 34788
rect 16112 34844 16176 34848
rect 16112 34788 16116 34844
rect 16116 34788 16172 34844
rect 16172 34788 16176 34844
rect 16112 34784 16176 34788
rect 16192 34844 16256 34848
rect 16192 34788 16196 34844
rect 16196 34788 16252 34844
rect 16252 34788 16256 34844
rect 16192 34784 16256 34788
rect 25952 34844 26016 34848
rect 25952 34788 25956 34844
rect 25956 34788 26012 34844
rect 26012 34788 26016 34844
rect 25952 34784 26016 34788
rect 26032 34844 26096 34848
rect 26032 34788 26036 34844
rect 26036 34788 26092 34844
rect 26092 34788 26096 34844
rect 26032 34784 26096 34788
rect 26112 34844 26176 34848
rect 26112 34788 26116 34844
rect 26116 34788 26172 34844
rect 26172 34788 26176 34844
rect 26112 34784 26176 34788
rect 26192 34844 26256 34848
rect 26192 34788 26196 34844
rect 26196 34788 26252 34844
rect 26252 34788 26256 34844
rect 26192 34784 26256 34788
rect 9812 34716 9876 34780
rect 10548 34716 10612 34780
rect 14596 34444 14660 34508
rect 9444 34308 9508 34372
rect 10364 34308 10428 34372
rect 12572 34308 12636 34372
rect 10952 34300 11016 34304
rect 10952 34244 10956 34300
rect 10956 34244 11012 34300
rect 11012 34244 11016 34300
rect 10952 34240 11016 34244
rect 11032 34300 11096 34304
rect 11032 34244 11036 34300
rect 11036 34244 11092 34300
rect 11092 34244 11096 34300
rect 11032 34240 11096 34244
rect 11112 34300 11176 34304
rect 11112 34244 11116 34300
rect 11116 34244 11172 34300
rect 11172 34244 11176 34300
rect 11112 34240 11176 34244
rect 11192 34300 11256 34304
rect 11192 34244 11196 34300
rect 11196 34244 11252 34300
rect 11252 34244 11256 34300
rect 11192 34240 11256 34244
rect 20952 34300 21016 34304
rect 20952 34244 20956 34300
rect 20956 34244 21012 34300
rect 21012 34244 21016 34300
rect 20952 34240 21016 34244
rect 21032 34300 21096 34304
rect 21032 34244 21036 34300
rect 21036 34244 21092 34300
rect 21092 34244 21096 34300
rect 21032 34240 21096 34244
rect 21112 34300 21176 34304
rect 21112 34244 21116 34300
rect 21116 34244 21172 34300
rect 21172 34244 21176 34300
rect 21112 34240 21176 34244
rect 21192 34300 21256 34304
rect 21192 34244 21196 34300
rect 21196 34244 21252 34300
rect 21252 34244 21256 34300
rect 21192 34240 21256 34244
rect 6684 33900 6748 33964
rect 9812 33900 9876 33964
rect 12204 33900 12268 33964
rect 14228 34036 14292 34100
rect 11652 33764 11716 33828
rect 16620 33764 16684 33828
rect 5952 33756 6016 33760
rect 5952 33700 5956 33756
rect 5956 33700 6012 33756
rect 6012 33700 6016 33756
rect 5952 33696 6016 33700
rect 6032 33756 6096 33760
rect 6032 33700 6036 33756
rect 6036 33700 6092 33756
rect 6092 33700 6096 33756
rect 6032 33696 6096 33700
rect 6112 33756 6176 33760
rect 6112 33700 6116 33756
rect 6116 33700 6172 33756
rect 6172 33700 6176 33756
rect 6112 33696 6176 33700
rect 6192 33756 6256 33760
rect 6192 33700 6196 33756
rect 6196 33700 6252 33756
rect 6252 33700 6256 33756
rect 6192 33696 6256 33700
rect 15952 33756 16016 33760
rect 15952 33700 15956 33756
rect 15956 33700 16012 33756
rect 16012 33700 16016 33756
rect 15952 33696 16016 33700
rect 16032 33756 16096 33760
rect 16032 33700 16036 33756
rect 16036 33700 16092 33756
rect 16092 33700 16096 33756
rect 16032 33696 16096 33700
rect 16112 33756 16176 33760
rect 16112 33700 16116 33756
rect 16116 33700 16172 33756
rect 16172 33700 16176 33756
rect 16112 33696 16176 33700
rect 16192 33756 16256 33760
rect 16192 33700 16196 33756
rect 16196 33700 16252 33756
rect 16252 33700 16256 33756
rect 16192 33696 16256 33700
rect 25952 33756 26016 33760
rect 25952 33700 25956 33756
rect 25956 33700 26012 33756
rect 26012 33700 26016 33756
rect 25952 33696 26016 33700
rect 26032 33756 26096 33760
rect 26032 33700 26036 33756
rect 26036 33700 26092 33756
rect 26092 33700 26096 33756
rect 26032 33696 26096 33700
rect 26112 33756 26176 33760
rect 26112 33700 26116 33756
rect 26116 33700 26172 33756
rect 26172 33700 26176 33756
rect 26112 33696 26176 33700
rect 26192 33756 26256 33760
rect 26192 33700 26196 33756
rect 26196 33700 26252 33756
rect 26252 33700 26256 33756
rect 26192 33696 26256 33700
rect 11652 33356 11716 33420
rect 15148 33356 15212 33420
rect 12204 33220 12268 33284
rect 14596 33220 14660 33284
rect 10952 33212 11016 33216
rect 10952 33156 10956 33212
rect 10956 33156 11012 33212
rect 11012 33156 11016 33212
rect 10952 33152 11016 33156
rect 11032 33212 11096 33216
rect 11032 33156 11036 33212
rect 11036 33156 11092 33212
rect 11092 33156 11096 33212
rect 11032 33152 11096 33156
rect 11112 33212 11176 33216
rect 11112 33156 11116 33212
rect 11116 33156 11172 33212
rect 11172 33156 11176 33212
rect 11112 33152 11176 33156
rect 11192 33212 11256 33216
rect 11192 33156 11196 33212
rect 11196 33156 11252 33212
rect 11252 33156 11256 33212
rect 11192 33152 11256 33156
rect 5580 32948 5644 33012
rect 12940 33084 13004 33148
rect 20952 33212 21016 33216
rect 20952 33156 20956 33212
rect 20956 33156 21012 33212
rect 21012 33156 21016 33212
rect 20952 33152 21016 33156
rect 21032 33212 21096 33216
rect 21032 33156 21036 33212
rect 21036 33156 21092 33212
rect 21092 33156 21096 33212
rect 21032 33152 21096 33156
rect 21112 33212 21176 33216
rect 21112 33156 21116 33212
rect 21116 33156 21172 33212
rect 21172 33156 21176 33212
rect 21112 33152 21176 33156
rect 21192 33212 21256 33216
rect 21192 33156 21196 33212
rect 21196 33156 21252 33212
rect 21252 33156 21256 33212
rect 21192 33152 21256 33156
rect 11468 32948 11532 33012
rect 12204 32948 12268 33012
rect 9260 32676 9324 32740
rect 5952 32668 6016 32672
rect 5952 32612 5956 32668
rect 5956 32612 6012 32668
rect 6012 32612 6016 32668
rect 5952 32608 6016 32612
rect 6032 32668 6096 32672
rect 6032 32612 6036 32668
rect 6036 32612 6092 32668
rect 6092 32612 6096 32668
rect 6032 32608 6096 32612
rect 6112 32668 6176 32672
rect 6112 32612 6116 32668
rect 6116 32612 6172 32668
rect 6172 32612 6176 32668
rect 6112 32608 6176 32612
rect 6192 32668 6256 32672
rect 6192 32612 6196 32668
rect 6196 32612 6252 32668
rect 6252 32612 6256 32668
rect 6192 32608 6256 32612
rect 14780 32676 14844 32740
rect 15952 32668 16016 32672
rect 15952 32612 15956 32668
rect 15956 32612 16012 32668
rect 16012 32612 16016 32668
rect 15952 32608 16016 32612
rect 16032 32668 16096 32672
rect 16032 32612 16036 32668
rect 16036 32612 16092 32668
rect 16092 32612 16096 32668
rect 16032 32608 16096 32612
rect 16112 32668 16176 32672
rect 16112 32612 16116 32668
rect 16116 32612 16172 32668
rect 16172 32612 16176 32668
rect 16112 32608 16176 32612
rect 16192 32668 16256 32672
rect 16192 32612 16196 32668
rect 16196 32612 16252 32668
rect 16252 32612 16256 32668
rect 16192 32608 16256 32612
rect 25952 32668 26016 32672
rect 25952 32612 25956 32668
rect 25956 32612 26012 32668
rect 26012 32612 26016 32668
rect 25952 32608 26016 32612
rect 26032 32668 26096 32672
rect 26032 32612 26036 32668
rect 26036 32612 26092 32668
rect 26092 32612 26096 32668
rect 26032 32608 26096 32612
rect 26112 32668 26176 32672
rect 26112 32612 26116 32668
rect 26116 32612 26172 32668
rect 26172 32612 26176 32668
rect 26112 32608 26176 32612
rect 26192 32668 26256 32672
rect 26192 32612 26196 32668
rect 26196 32612 26252 32668
rect 26252 32612 26256 32668
rect 26192 32608 26256 32612
rect 21772 32404 21836 32468
rect 10364 32132 10428 32196
rect 16988 32268 17052 32332
rect 10952 32124 11016 32128
rect 10952 32068 10956 32124
rect 10956 32068 11012 32124
rect 11012 32068 11016 32124
rect 10952 32064 11016 32068
rect 11032 32124 11096 32128
rect 11032 32068 11036 32124
rect 11036 32068 11092 32124
rect 11092 32068 11096 32124
rect 11032 32064 11096 32068
rect 11112 32124 11176 32128
rect 11112 32068 11116 32124
rect 11116 32068 11172 32124
rect 11172 32068 11176 32124
rect 11112 32064 11176 32068
rect 11192 32124 11256 32128
rect 11192 32068 11196 32124
rect 11196 32068 11252 32124
rect 11252 32068 11256 32124
rect 11192 32064 11256 32068
rect 20952 32124 21016 32128
rect 20952 32068 20956 32124
rect 20956 32068 21012 32124
rect 21012 32068 21016 32124
rect 20952 32064 21016 32068
rect 21032 32124 21096 32128
rect 21032 32068 21036 32124
rect 21036 32068 21092 32124
rect 21092 32068 21096 32124
rect 21032 32064 21096 32068
rect 21112 32124 21176 32128
rect 21112 32068 21116 32124
rect 21116 32068 21172 32124
rect 21172 32068 21176 32124
rect 21112 32064 21176 32068
rect 21192 32124 21256 32128
rect 21192 32068 21196 32124
rect 21196 32068 21252 32124
rect 21252 32068 21256 32124
rect 21192 32064 21256 32068
rect 3372 31996 3436 32060
rect 9076 31996 9140 32060
rect 10548 31996 10612 32060
rect 11468 31996 11532 32060
rect 12756 31860 12820 31924
rect 13308 31860 13372 31924
rect 13860 31860 13924 31924
rect 12756 31784 12820 31788
rect 12756 31728 12806 31784
rect 12806 31728 12820 31784
rect 12756 31724 12820 31728
rect 14044 31724 14108 31788
rect 9444 31648 9508 31652
rect 9444 31592 9494 31648
rect 9494 31592 9508 31648
rect 9444 31588 9508 31592
rect 10732 31588 10796 31652
rect 11652 31648 11716 31652
rect 11652 31592 11702 31648
rect 11702 31592 11716 31648
rect 11652 31588 11716 31592
rect 12572 31588 12636 31652
rect 14044 31588 14108 31652
rect 20668 31860 20732 31924
rect 14412 31724 14476 31788
rect 5952 31580 6016 31584
rect 5952 31524 5956 31580
rect 5956 31524 6012 31580
rect 6012 31524 6016 31580
rect 5952 31520 6016 31524
rect 6032 31580 6096 31584
rect 6032 31524 6036 31580
rect 6036 31524 6092 31580
rect 6092 31524 6096 31580
rect 6032 31520 6096 31524
rect 6112 31580 6176 31584
rect 6112 31524 6116 31580
rect 6116 31524 6172 31580
rect 6172 31524 6176 31580
rect 6112 31520 6176 31524
rect 6192 31580 6256 31584
rect 6192 31524 6196 31580
rect 6196 31524 6252 31580
rect 6252 31524 6256 31580
rect 6192 31520 6256 31524
rect 15952 31580 16016 31584
rect 15952 31524 15956 31580
rect 15956 31524 16012 31580
rect 16012 31524 16016 31580
rect 15952 31520 16016 31524
rect 16032 31580 16096 31584
rect 16032 31524 16036 31580
rect 16036 31524 16092 31580
rect 16092 31524 16096 31580
rect 16032 31520 16096 31524
rect 16112 31580 16176 31584
rect 16112 31524 16116 31580
rect 16116 31524 16172 31580
rect 16172 31524 16176 31580
rect 16112 31520 16176 31524
rect 16192 31580 16256 31584
rect 16192 31524 16196 31580
rect 16196 31524 16252 31580
rect 16252 31524 16256 31580
rect 16192 31520 16256 31524
rect 25952 31580 26016 31584
rect 25952 31524 25956 31580
rect 25956 31524 26012 31580
rect 26012 31524 26016 31580
rect 25952 31520 26016 31524
rect 26032 31580 26096 31584
rect 26032 31524 26036 31580
rect 26036 31524 26092 31580
rect 26092 31524 26096 31580
rect 26032 31520 26096 31524
rect 26112 31580 26176 31584
rect 26112 31524 26116 31580
rect 26116 31524 26172 31580
rect 26172 31524 26176 31580
rect 26112 31520 26176 31524
rect 26192 31580 26256 31584
rect 26192 31524 26196 31580
rect 26196 31524 26252 31580
rect 26252 31524 26256 31580
rect 26192 31520 26256 31524
rect 11652 31452 11716 31516
rect 11468 31316 11532 31380
rect 13860 31316 13924 31380
rect 14228 31316 14292 31380
rect 25084 31316 25148 31380
rect 10952 31036 11016 31040
rect 10952 30980 10956 31036
rect 10956 30980 11012 31036
rect 11012 30980 11016 31036
rect 10952 30976 11016 30980
rect 11032 31036 11096 31040
rect 11032 30980 11036 31036
rect 11036 30980 11092 31036
rect 11092 30980 11096 31036
rect 11032 30976 11096 30980
rect 11112 31036 11176 31040
rect 11112 30980 11116 31036
rect 11116 30980 11172 31036
rect 11172 30980 11176 31036
rect 11112 30976 11176 30980
rect 11192 31036 11256 31040
rect 11192 30980 11196 31036
rect 11196 30980 11252 31036
rect 11252 30980 11256 31036
rect 11192 30976 11256 30980
rect 14964 31044 15028 31108
rect 20484 31044 20548 31108
rect 20952 31036 21016 31040
rect 20952 30980 20956 31036
rect 20956 30980 21012 31036
rect 21012 30980 21016 31036
rect 20952 30976 21016 30980
rect 21032 31036 21096 31040
rect 21032 30980 21036 31036
rect 21036 30980 21092 31036
rect 21092 30980 21096 31036
rect 21032 30976 21096 30980
rect 21112 31036 21176 31040
rect 21112 30980 21116 31036
rect 21116 30980 21172 31036
rect 21172 30980 21176 31036
rect 21112 30976 21176 30980
rect 21192 31036 21256 31040
rect 21192 30980 21196 31036
rect 21196 30980 21252 31036
rect 21252 30980 21256 31036
rect 21192 30976 21256 30980
rect 14780 30908 14844 30972
rect 20668 30772 20732 30836
rect 13308 30696 13372 30700
rect 13308 30640 13358 30696
rect 13358 30640 13372 30696
rect 13308 30636 13372 30640
rect 16620 30560 16684 30564
rect 16620 30504 16670 30560
rect 16670 30504 16684 30560
rect 16620 30500 16684 30504
rect 5952 30492 6016 30496
rect 5952 30436 5956 30492
rect 5956 30436 6012 30492
rect 6012 30436 6016 30492
rect 5952 30432 6016 30436
rect 6032 30492 6096 30496
rect 6032 30436 6036 30492
rect 6036 30436 6092 30492
rect 6092 30436 6096 30492
rect 6032 30432 6096 30436
rect 6112 30492 6176 30496
rect 6112 30436 6116 30492
rect 6116 30436 6172 30492
rect 6172 30436 6176 30492
rect 6112 30432 6176 30436
rect 6192 30492 6256 30496
rect 6192 30436 6196 30492
rect 6196 30436 6252 30492
rect 6252 30436 6256 30492
rect 6192 30432 6256 30436
rect 15952 30492 16016 30496
rect 15952 30436 15956 30492
rect 15956 30436 16012 30492
rect 16012 30436 16016 30492
rect 15952 30432 16016 30436
rect 16032 30492 16096 30496
rect 16032 30436 16036 30492
rect 16036 30436 16092 30492
rect 16092 30436 16096 30492
rect 16032 30432 16096 30436
rect 16112 30492 16176 30496
rect 16112 30436 16116 30492
rect 16116 30436 16172 30492
rect 16172 30436 16176 30492
rect 16112 30432 16176 30436
rect 16192 30492 16256 30496
rect 16192 30436 16196 30492
rect 16196 30436 16252 30492
rect 16252 30436 16256 30492
rect 16192 30432 16256 30436
rect 12756 30364 12820 30428
rect 12940 30364 13004 30428
rect 16804 30228 16868 30292
rect 17540 30288 17604 30292
rect 17540 30232 17554 30288
rect 17554 30232 17604 30288
rect 17540 30228 17604 30232
rect 11652 30092 11716 30156
rect 13860 30092 13924 30156
rect 25952 30492 26016 30496
rect 25952 30436 25956 30492
rect 25956 30436 26012 30492
rect 26012 30436 26016 30492
rect 25952 30432 26016 30436
rect 26032 30492 26096 30496
rect 26032 30436 26036 30492
rect 26036 30436 26092 30492
rect 26092 30436 26096 30492
rect 26032 30432 26096 30436
rect 26112 30492 26176 30496
rect 26112 30436 26116 30492
rect 26116 30436 26172 30492
rect 26172 30436 26176 30492
rect 26112 30432 26176 30436
rect 26192 30492 26256 30496
rect 26192 30436 26196 30492
rect 26196 30436 26252 30492
rect 26252 30436 26256 30492
rect 26192 30432 26256 30436
rect 10364 29956 10428 30020
rect 13308 29956 13372 30020
rect 10952 29948 11016 29952
rect 10952 29892 10956 29948
rect 10956 29892 11012 29948
rect 11012 29892 11016 29948
rect 10952 29888 11016 29892
rect 11032 29948 11096 29952
rect 11032 29892 11036 29948
rect 11036 29892 11092 29948
rect 11092 29892 11096 29948
rect 11032 29888 11096 29892
rect 11112 29948 11176 29952
rect 11112 29892 11116 29948
rect 11116 29892 11172 29948
rect 11172 29892 11176 29948
rect 11112 29888 11176 29892
rect 11192 29948 11256 29952
rect 11192 29892 11196 29948
rect 11196 29892 11252 29948
rect 11252 29892 11256 29948
rect 11192 29888 11256 29892
rect 20952 29948 21016 29952
rect 20952 29892 20956 29948
rect 20956 29892 21012 29948
rect 21012 29892 21016 29948
rect 20952 29888 21016 29892
rect 21032 29948 21096 29952
rect 21032 29892 21036 29948
rect 21036 29892 21092 29948
rect 21092 29892 21096 29948
rect 21032 29888 21096 29892
rect 21112 29948 21176 29952
rect 21112 29892 21116 29948
rect 21116 29892 21172 29948
rect 21172 29892 21176 29948
rect 21112 29888 21176 29892
rect 21192 29948 21256 29952
rect 21192 29892 21196 29948
rect 21196 29892 21252 29948
rect 21252 29892 21256 29948
rect 21192 29888 21256 29892
rect 12940 29820 13004 29884
rect 10548 29684 10612 29748
rect 11652 29684 11716 29748
rect 14044 29744 14108 29748
rect 14044 29688 14094 29744
rect 14094 29688 14108 29744
rect 14044 29684 14108 29688
rect 14228 29548 14292 29612
rect 9260 29412 9324 29476
rect 5952 29404 6016 29408
rect 5952 29348 5956 29404
rect 5956 29348 6012 29404
rect 6012 29348 6016 29404
rect 5952 29344 6016 29348
rect 6032 29404 6096 29408
rect 6032 29348 6036 29404
rect 6036 29348 6092 29404
rect 6092 29348 6096 29404
rect 6032 29344 6096 29348
rect 6112 29404 6176 29408
rect 6112 29348 6116 29404
rect 6116 29348 6172 29404
rect 6172 29348 6176 29404
rect 6112 29344 6176 29348
rect 6192 29404 6256 29408
rect 6192 29348 6196 29404
rect 6196 29348 6252 29404
rect 6252 29348 6256 29404
rect 6192 29344 6256 29348
rect 15952 29404 16016 29408
rect 15952 29348 15956 29404
rect 15956 29348 16012 29404
rect 16012 29348 16016 29404
rect 15952 29344 16016 29348
rect 16032 29404 16096 29408
rect 16032 29348 16036 29404
rect 16036 29348 16092 29404
rect 16092 29348 16096 29404
rect 16032 29344 16096 29348
rect 16112 29404 16176 29408
rect 16112 29348 16116 29404
rect 16116 29348 16172 29404
rect 16172 29348 16176 29404
rect 16112 29344 16176 29348
rect 16192 29404 16256 29408
rect 16192 29348 16196 29404
rect 16196 29348 16252 29404
rect 16252 29348 16256 29404
rect 16192 29344 16256 29348
rect 12756 29276 12820 29340
rect 13124 29276 13188 29340
rect 25952 29404 26016 29408
rect 25952 29348 25956 29404
rect 25956 29348 26012 29404
rect 26012 29348 26016 29404
rect 25952 29344 26016 29348
rect 26032 29404 26096 29408
rect 26032 29348 26036 29404
rect 26036 29348 26092 29404
rect 26092 29348 26096 29404
rect 26032 29344 26096 29348
rect 26112 29404 26176 29408
rect 26112 29348 26116 29404
rect 26116 29348 26172 29404
rect 26172 29348 26176 29404
rect 26112 29344 26176 29348
rect 26192 29404 26256 29408
rect 26192 29348 26196 29404
rect 26196 29348 26252 29404
rect 26252 29348 26256 29404
rect 26192 29344 26256 29348
rect 7420 28868 7484 28932
rect 10952 28860 11016 28864
rect 10952 28804 10956 28860
rect 10956 28804 11012 28860
rect 11012 28804 11016 28860
rect 10952 28800 11016 28804
rect 11032 28860 11096 28864
rect 11032 28804 11036 28860
rect 11036 28804 11092 28860
rect 11092 28804 11096 28860
rect 11032 28800 11096 28804
rect 11112 28860 11176 28864
rect 11112 28804 11116 28860
rect 11116 28804 11172 28860
rect 11172 28804 11176 28860
rect 11112 28800 11176 28804
rect 11192 28860 11256 28864
rect 11192 28804 11196 28860
rect 11196 28804 11252 28860
rect 11252 28804 11256 28860
rect 11192 28800 11256 28804
rect 20952 28860 21016 28864
rect 20952 28804 20956 28860
rect 20956 28804 21012 28860
rect 21012 28804 21016 28860
rect 20952 28800 21016 28804
rect 21032 28860 21096 28864
rect 21032 28804 21036 28860
rect 21036 28804 21092 28860
rect 21092 28804 21096 28860
rect 21032 28800 21096 28804
rect 21112 28860 21176 28864
rect 21112 28804 21116 28860
rect 21116 28804 21172 28860
rect 21172 28804 21176 28860
rect 21112 28800 21176 28804
rect 21192 28860 21256 28864
rect 21192 28804 21196 28860
rect 21196 28804 21252 28860
rect 21252 28804 21256 28860
rect 21192 28800 21256 28804
rect 13860 28596 13924 28660
rect 14228 28324 14292 28388
rect 5952 28316 6016 28320
rect 5952 28260 5956 28316
rect 5956 28260 6012 28316
rect 6012 28260 6016 28316
rect 5952 28256 6016 28260
rect 6032 28316 6096 28320
rect 6032 28260 6036 28316
rect 6036 28260 6092 28316
rect 6092 28260 6096 28316
rect 6032 28256 6096 28260
rect 6112 28316 6176 28320
rect 6112 28260 6116 28316
rect 6116 28260 6172 28316
rect 6172 28260 6176 28316
rect 6112 28256 6176 28260
rect 6192 28316 6256 28320
rect 6192 28260 6196 28316
rect 6196 28260 6252 28316
rect 6252 28260 6256 28316
rect 6192 28256 6256 28260
rect 15952 28316 16016 28320
rect 15952 28260 15956 28316
rect 15956 28260 16012 28316
rect 16012 28260 16016 28316
rect 15952 28256 16016 28260
rect 16032 28316 16096 28320
rect 16032 28260 16036 28316
rect 16036 28260 16092 28316
rect 16092 28260 16096 28316
rect 16032 28256 16096 28260
rect 16112 28316 16176 28320
rect 16112 28260 16116 28316
rect 16116 28260 16172 28316
rect 16172 28260 16176 28316
rect 16112 28256 16176 28260
rect 16192 28316 16256 28320
rect 16192 28260 16196 28316
rect 16196 28260 16252 28316
rect 16252 28260 16256 28316
rect 16192 28256 16256 28260
rect 25952 28316 26016 28320
rect 25952 28260 25956 28316
rect 25956 28260 26012 28316
rect 26012 28260 26016 28316
rect 25952 28256 26016 28260
rect 26032 28316 26096 28320
rect 26032 28260 26036 28316
rect 26036 28260 26092 28316
rect 26092 28260 26096 28316
rect 26032 28256 26096 28260
rect 26112 28316 26176 28320
rect 26112 28260 26116 28316
rect 26116 28260 26172 28316
rect 26172 28260 26176 28316
rect 26112 28256 26176 28260
rect 26192 28316 26256 28320
rect 26192 28260 26196 28316
rect 26196 28260 26252 28316
rect 26252 28260 26256 28316
rect 26192 28256 26256 28260
rect 10548 28052 10612 28116
rect 9628 27780 9692 27844
rect 10952 27772 11016 27776
rect 10952 27716 10956 27772
rect 10956 27716 11012 27772
rect 11012 27716 11016 27772
rect 10952 27712 11016 27716
rect 11032 27772 11096 27776
rect 11032 27716 11036 27772
rect 11036 27716 11092 27772
rect 11092 27716 11096 27772
rect 11032 27712 11096 27716
rect 11112 27772 11176 27776
rect 11112 27716 11116 27772
rect 11116 27716 11172 27772
rect 11172 27716 11176 27772
rect 11112 27712 11176 27716
rect 11192 27772 11256 27776
rect 11192 27716 11196 27772
rect 11196 27716 11252 27772
rect 11252 27716 11256 27772
rect 11192 27712 11256 27716
rect 20952 27772 21016 27776
rect 20952 27716 20956 27772
rect 20956 27716 21012 27772
rect 21012 27716 21016 27772
rect 20952 27712 21016 27716
rect 21032 27772 21096 27776
rect 21032 27716 21036 27772
rect 21036 27716 21092 27772
rect 21092 27716 21096 27772
rect 21032 27712 21096 27716
rect 21112 27772 21176 27776
rect 21112 27716 21116 27772
rect 21116 27716 21172 27772
rect 21172 27716 21176 27772
rect 21112 27712 21176 27716
rect 21192 27772 21256 27776
rect 21192 27716 21196 27772
rect 21196 27716 21252 27772
rect 21252 27716 21256 27772
rect 21192 27712 21256 27716
rect 12388 27644 12452 27708
rect 16620 27644 16684 27708
rect 17540 27704 17604 27708
rect 17540 27648 17590 27704
rect 17590 27648 17604 27704
rect 17540 27644 17604 27648
rect 5952 27228 6016 27232
rect 5952 27172 5956 27228
rect 5956 27172 6012 27228
rect 6012 27172 6016 27228
rect 5952 27168 6016 27172
rect 6032 27228 6096 27232
rect 6032 27172 6036 27228
rect 6036 27172 6092 27228
rect 6092 27172 6096 27228
rect 6032 27168 6096 27172
rect 6112 27228 6176 27232
rect 6112 27172 6116 27228
rect 6116 27172 6172 27228
rect 6172 27172 6176 27228
rect 6112 27168 6176 27172
rect 6192 27228 6256 27232
rect 6192 27172 6196 27228
rect 6196 27172 6252 27228
rect 6252 27172 6256 27228
rect 6192 27168 6256 27172
rect 12572 27100 12636 27164
rect 12204 26964 12268 27028
rect 15952 27228 16016 27232
rect 15952 27172 15956 27228
rect 15956 27172 16012 27228
rect 16012 27172 16016 27228
rect 15952 27168 16016 27172
rect 16032 27228 16096 27232
rect 16032 27172 16036 27228
rect 16036 27172 16092 27228
rect 16092 27172 16096 27228
rect 16032 27168 16096 27172
rect 16112 27228 16176 27232
rect 16112 27172 16116 27228
rect 16116 27172 16172 27228
rect 16172 27172 16176 27228
rect 16112 27168 16176 27172
rect 16192 27228 16256 27232
rect 16192 27172 16196 27228
rect 16196 27172 16252 27228
rect 16252 27172 16256 27228
rect 16192 27168 16256 27172
rect 25952 27228 26016 27232
rect 25952 27172 25956 27228
rect 25956 27172 26012 27228
rect 26012 27172 26016 27228
rect 25952 27168 26016 27172
rect 26032 27228 26096 27232
rect 26032 27172 26036 27228
rect 26036 27172 26092 27228
rect 26092 27172 26096 27228
rect 26032 27168 26096 27172
rect 26112 27228 26176 27232
rect 26112 27172 26116 27228
rect 26116 27172 26172 27228
rect 26172 27172 26176 27228
rect 26112 27168 26176 27172
rect 26192 27228 26256 27232
rect 26192 27172 26196 27228
rect 26196 27172 26252 27228
rect 26252 27172 26256 27228
rect 26192 27168 26256 27172
rect 9812 26828 9876 26892
rect 10952 26684 11016 26688
rect 10952 26628 10956 26684
rect 10956 26628 11012 26684
rect 11012 26628 11016 26684
rect 10952 26624 11016 26628
rect 11032 26684 11096 26688
rect 11032 26628 11036 26684
rect 11036 26628 11092 26684
rect 11092 26628 11096 26684
rect 11032 26624 11096 26628
rect 11112 26684 11176 26688
rect 11112 26628 11116 26684
rect 11116 26628 11172 26684
rect 11172 26628 11176 26684
rect 11112 26624 11176 26628
rect 11192 26684 11256 26688
rect 11192 26628 11196 26684
rect 11196 26628 11252 26684
rect 11252 26628 11256 26684
rect 11192 26624 11256 26628
rect 20952 26684 21016 26688
rect 20952 26628 20956 26684
rect 20956 26628 21012 26684
rect 21012 26628 21016 26684
rect 20952 26624 21016 26628
rect 21032 26684 21096 26688
rect 21032 26628 21036 26684
rect 21036 26628 21092 26684
rect 21092 26628 21096 26684
rect 21032 26624 21096 26628
rect 21112 26684 21176 26688
rect 21112 26628 21116 26684
rect 21116 26628 21172 26684
rect 21172 26628 21176 26684
rect 21112 26624 21176 26628
rect 21192 26684 21256 26688
rect 21192 26628 21196 26684
rect 21196 26628 21252 26684
rect 21252 26628 21256 26684
rect 21192 26624 21256 26628
rect 10732 26284 10796 26348
rect 11468 26284 11532 26348
rect 5952 26140 6016 26144
rect 5952 26084 5956 26140
rect 5956 26084 6012 26140
rect 6012 26084 6016 26140
rect 5952 26080 6016 26084
rect 6032 26140 6096 26144
rect 6032 26084 6036 26140
rect 6036 26084 6092 26140
rect 6092 26084 6096 26140
rect 6032 26080 6096 26084
rect 6112 26140 6176 26144
rect 6112 26084 6116 26140
rect 6116 26084 6172 26140
rect 6172 26084 6176 26140
rect 6112 26080 6176 26084
rect 6192 26140 6256 26144
rect 6192 26084 6196 26140
rect 6196 26084 6252 26140
rect 6252 26084 6256 26140
rect 6192 26080 6256 26084
rect 15952 26140 16016 26144
rect 15952 26084 15956 26140
rect 15956 26084 16012 26140
rect 16012 26084 16016 26140
rect 15952 26080 16016 26084
rect 16032 26140 16096 26144
rect 16032 26084 16036 26140
rect 16036 26084 16092 26140
rect 16092 26084 16096 26140
rect 16032 26080 16096 26084
rect 16112 26140 16176 26144
rect 16112 26084 16116 26140
rect 16116 26084 16172 26140
rect 16172 26084 16176 26140
rect 16112 26080 16176 26084
rect 16192 26140 16256 26144
rect 16192 26084 16196 26140
rect 16196 26084 16252 26140
rect 16252 26084 16256 26140
rect 16192 26080 16256 26084
rect 10180 25876 10244 25940
rect 25952 26140 26016 26144
rect 25952 26084 25956 26140
rect 25956 26084 26012 26140
rect 26012 26084 26016 26140
rect 25952 26080 26016 26084
rect 26032 26140 26096 26144
rect 26032 26084 26036 26140
rect 26036 26084 26092 26140
rect 26092 26084 26096 26140
rect 26032 26080 26096 26084
rect 26112 26140 26176 26144
rect 26112 26084 26116 26140
rect 26116 26084 26172 26140
rect 26172 26084 26176 26140
rect 26112 26080 26176 26084
rect 26192 26140 26256 26144
rect 26192 26084 26196 26140
rect 26196 26084 26252 26140
rect 26252 26084 26256 26140
rect 26192 26080 26256 26084
rect 9628 25604 9692 25668
rect 10548 25604 10612 25668
rect 10732 25664 10796 25668
rect 10732 25608 10746 25664
rect 10746 25608 10796 25664
rect 10732 25604 10796 25608
rect 10952 25596 11016 25600
rect 10952 25540 10956 25596
rect 10956 25540 11012 25596
rect 11012 25540 11016 25596
rect 10952 25536 11016 25540
rect 11032 25596 11096 25600
rect 11032 25540 11036 25596
rect 11036 25540 11092 25596
rect 11092 25540 11096 25596
rect 11032 25536 11096 25540
rect 11112 25596 11176 25600
rect 11112 25540 11116 25596
rect 11116 25540 11172 25596
rect 11172 25540 11176 25596
rect 11112 25536 11176 25540
rect 11192 25596 11256 25600
rect 11192 25540 11196 25596
rect 11196 25540 11252 25596
rect 11252 25540 11256 25596
rect 11192 25536 11256 25540
rect 20952 25596 21016 25600
rect 20952 25540 20956 25596
rect 20956 25540 21012 25596
rect 21012 25540 21016 25596
rect 20952 25536 21016 25540
rect 21032 25596 21096 25600
rect 21032 25540 21036 25596
rect 21036 25540 21092 25596
rect 21092 25540 21096 25596
rect 21032 25536 21096 25540
rect 21112 25596 21176 25600
rect 21112 25540 21116 25596
rect 21116 25540 21172 25596
rect 21172 25540 21176 25596
rect 21112 25536 21176 25540
rect 21192 25596 21256 25600
rect 21192 25540 21196 25596
rect 21196 25540 21252 25596
rect 21252 25540 21256 25596
rect 21192 25536 21256 25540
rect 12388 25332 12452 25396
rect 14412 25332 14476 25396
rect 5952 25052 6016 25056
rect 5952 24996 5956 25052
rect 5956 24996 6012 25052
rect 6012 24996 6016 25052
rect 5952 24992 6016 24996
rect 6032 25052 6096 25056
rect 6032 24996 6036 25052
rect 6036 24996 6092 25052
rect 6092 24996 6096 25052
rect 6032 24992 6096 24996
rect 6112 25052 6176 25056
rect 6112 24996 6116 25052
rect 6116 24996 6172 25052
rect 6172 24996 6176 25052
rect 6112 24992 6176 24996
rect 6192 25052 6256 25056
rect 6192 24996 6196 25052
rect 6196 24996 6252 25052
rect 6252 24996 6256 25052
rect 6192 24992 6256 24996
rect 15952 25052 16016 25056
rect 15952 24996 15956 25052
rect 15956 24996 16012 25052
rect 16012 24996 16016 25052
rect 15952 24992 16016 24996
rect 16032 25052 16096 25056
rect 16032 24996 16036 25052
rect 16036 24996 16092 25052
rect 16092 24996 16096 25052
rect 16032 24992 16096 24996
rect 16112 25052 16176 25056
rect 16112 24996 16116 25052
rect 16116 24996 16172 25052
rect 16172 24996 16176 25052
rect 16112 24992 16176 24996
rect 16192 25052 16256 25056
rect 16192 24996 16196 25052
rect 16196 24996 16252 25052
rect 16252 24996 16256 25052
rect 16192 24992 16256 24996
rect 25952 25052 26016 25056
rect 25952 24996 25956 25052
rect 25956 24996 26012 25052
rect 26012 24996 26016 25052
rect 25952 24992 26016 24996
rect 26032 25052 26096 25056
rect 26032 24996 26036 25052
rect 26036 24996 26092 25052
rect 26092 24996 26096 25052
rect 26032 24992 26096 24996
rect 26112 25052 26176 25056
rect 26112 24996 26116 25052
rect 26116 24996 26172 25052
rect 26172 24996 26176 25052
rect 26112 24992 26176 24996
rect 26192 25052 26256 25056
rect 26192 24996 26196 25052
rect 26196 24996 26252 25052
rect 26252 24996 26256 25052
rect 26192 24992 26256 24996
rect 11468 24516 11532 24580
rect 10952 24508 11016 24512
rect 10952 24452 10956 24508
rect 10956 24452 11012 24508
rect 11012 24452 11016 24508
rect 10952 24448 11016 24452
rect 11032 24508 11096 24512
rect 11032 24452 11036 24508
rect 11036 24452 11092 24508
rect 11092 24452 11096 24508
rect 11032 24448 11096 24452
rect 11112 24508 11176 24512
rect 11112 24452 11116 24508
rect 11116 24452 11172 24508
rect 11172 24452 11176 24508
rect 11112 24448 11176 24452
rect 11192 24508 11256 24512
rect 11192 24452 11196 24508
rect 11196 24452 11252 24508
rect 11252 24452 11256 24508
rect 11192 24448 11256 24452
rect 20952 24508 21016 24512
rect 20952 24452 20956 24508
rect 20956 24452 21012 24508
rect 21012 24452 21016 24508
rect 20952 24448 21016 24452
rect 21032 24508 21096 24512
rect 21032 24452 21036 24508
rect 21036 24452 21092 24508
rect 21092 24452 21096 24508
rect 21032 24448 21096 24452
rect 21112 24508 21176 24512
rect 21112 24452 21116 24508
rect 21116 24452 21172 24508
rect 21172 24452 21176 24508
rect 21112 24448 21176 24452
rect 21192 24508 21256 24512
rect 21192 24452 21196 24508
rect 21196 24452 21252 24508
rect 21252 24452 21256 24508
rect 21192 24448 21256 24452
rect 5952 23964 6016 23968
rect 5952 23908 5956 23964
rect 5956 23908 6012 23964
rect 6012 23908 6016 23964
rect 5952 23904 6016 23908
rect 6032 23964 6096 23968
rect 6032 23908 6036 23964
rect 6036 23908 6092 23964
rect 6092 23908 6096 23964
rect 6032 23904 6096 23908
rect 6112 23964 6176 23968
rect 6112 23908 6116 23964
rect 6116 23908 6172 23964
rect 6172 23908 6176 23964
rect 6112 23904 6176 23908
rect 6192 23964 6256 23968
rect 6192 23908 6196 23964
rect 6196 23908 6252 23964
rect 6252 23908 6256 23964
rect 6192 23904 6256 23908
rect 15952 23964 16016 23968
rect 15952 23908 15956 23964
rect 15956 23908 16012 23964
rect 16012 23908 16016 23964
rect 15952 23904 16016 23908
rect 16032 23964 16096 23968
rect 16032 23908 16036 23964
rect 16036 23908 16092 23964
rect 16092 23908 16096 23964
rect 16032 23904 16096 23908
rect 16112 23964 16176 23968
rect 16112 23908 16116 23964
rect 16116 23908 16172 23964
rect 16172 23908 16176 23964
rect 16112 23904 16176 23908
rect 16192 23964 16256 23968
rect 16192 23908 16196 23964
rect 16196 23908 16252 23964
rect 16252 23908 16256 23964
rect 16192 23904 16256 23908
rect 25952 23964 26016 23968
rect 25952 23908 25956 23964
rect 25956 23908 26012 23964
rect 26012 23908 26016 23964
rect 25952 23904 26016 23908
rect 26032 23964 26096 23968
rect 26032 23908 26036 23964
rect 26036 23908 26092 23964
rect 26092 23908 26096 23964
rect 26032 23904 26096 23908
rect 26112 23964 26176 23968
rect 26112 23908 26116 23964
rect 26116 23908 26172 23964
rect 26172 23908 26176 23964
rect 26112 23904 26176 23908
rect 26192 23964 26256 23968
rect 26192 23908 26196 23964
rect 26196 23908 26252 23964
rect 26252 23908 26256 23964
rect 26192 23904 26256 23908
rect 12204 23564 12268 23628
rect 16620 23564 16684 23628
rect 25636 23564 25700 23628
rect 10952 23420 11016 23424
rect 10952 23364 10956 23420
rect 10956 23364 11012 23420
rect 11012 23364 11016 23420
rect 10952 23360 11016 23364
rect 11032 23420 11096 23424
rect 11032 23364 11036 23420
rect 11036 23364 11092 23420
rect 11092 23364 11096 23420
rect 11032 23360 11096 23364
rect 11112 23420 11176 23424
rect 11112 23364 11116 23420
rect 11116 23364 11172 23420
rect 11172 23364 11176 23420
rect 11112 23360 11176 23364
rect 11192 23420 11256 23424
rect 11192 23364 11196 23420
rect 11196 23364 11252 23420
rect 11252 23364 11256 23420
rect 11192 23360 11256 23364
rect 20952 23420 21016 23424
rect 20952 23364 20956 23420
rect 20956 23364 21012 23420
rect 21012 23364 21016 23420
rect 20952 23360 21016 23364
rect 21032 23420 21096 23424
rect 21032 23364 21036 23420
rect 21036 23364 21092 23420
rect 21092 23364 21096 23420
rect 21032 23360 21096 23364
rect 21112 23420 21176 23424
rect 21112 23364 21116 23420
rect 21116 23364 21172 23420
rect 21172 23364 21176 23420
rect 21112 23360 21176 23364
rect 21192 23420 21256 23424
rect 21192 23364 21196 23420
rect 21196 23364 21252 23420
rect 21252 23364 21256 23420
rect 21192 23360 21256 23364
rect 14964 22884 15028 22948
rect 5952 22876 6016 22880
rect 5952 22820 5956 22876
rect 5956 22820 6012 22876
rect 6012 22820 6016 22876
rect 5952 22816 6016 22820
rect 6032 22876 6096 22880
rect 6032 22820 6036 22876
rect 6036 22820 6092 22876
rect 6092 22820 6096 22876
rect 6032 22816 6096 22820
rect 6112 22876 6176 22880
rect 6112 22820 6116 22876
rect 6116 22820 6172 22876
rect 6172 22820 6176 22876
rect 6112 22816 6176 22820
rect 6192 22876 6256 22880
rect 6192 22820 6196 22876
rect 6196 22820 6252 22876
rect 6252 22820 6256 22876
rect 6192 22816 6256 22820
rect 15952 22876 16016 22880
rect 15952 22820 15956 22876
rect 15956 22820 16012 22876
rect 16012 22820 16016 22876
rect 15952 22816 16016 22820
rect 16032 22876 16096 22880
rect 16032 22820 16036 22876
rect 16036 22820 16092 22876
rect 16092 22820 16096 22876
rect 16032 22816 16096 22820
rect 16112 22876 16176 22880
rect 16112 22820 16116 22876
rect 16116 22820 16172 22876
rect 16172 22820 16176 22876
rect 16112 22816 16176 22820
rect 16192 22876 16256 22880
rect 16192 22820 16196 22876
rect 16196 22820 16252 22876
rect 16252 22820 16256 22876
rect 16192 22816 16256 22820
rect 25952 22876 26016 22880
rect 25952 22820 25956 22876
rect 25956 22820 26012 22876
rect 26012 22820 26016 22876
rect 25952 22816 26016 22820
rect 26032 22876 26096 22880
rect 26032 22820 26036 22876
rect 26036 22820 26092 22876
rect 26092 22820 26096 22876
rect 26032 22816 26096 22820
rect 26112 22876 26176 22880
rect 26112 22820 26116 22876
rect 26116 22820 26172 22876
rect 26172 22820 26176 22876
rect 26112 22816 26176 22820
rect 26192 22876 26256 22880
rect 26192 22820 26196 22876
rect 26196 22820 26252 22876
rect 26252 22820 26256 22876
rect 26192 22816 26256 22820
rect 11468 22612 11532 22676
rect 15148 22612 15212 22676
rect 13308 22476 13372 22540
rect 11652 22340 11716 22404
rect 10952 22332 11016 22336
rect 10952 22276 10956 22332
rect 10956 22276 11012 22332
rect 11012 22276 11016 22332
rect 10952 22272 11016 22276
rect 11032 22332 11096 22336
rect 11032 22276 11036 22332
rect 11036 22276 11092 22332
rect 11092 22276 11096 22332
rect 11032 22272 11096 22276
rect 11112 22332 11176 22336
rect 11112 22276 11116 22332
rect 11116 22276 11172 22332
rect 11172 22276 11176 22332
rect 11112 22272 11176 22276
rect 11192 22332 11256 22336
rect 11192 22276 11196 22332
rect 11196 22276 11252 22332
rect 11252 22276 11256 22332
rect 11192 22272 11256 22276
rect 20952 22332 21016 22336
rect 20952 22276 20956 22332
rect 20956 22276 21012 22332
rect 21012 22276 21016 22332
rect 20952 22272 21016 22276
rect 21032 22332 21096 22336
rect 21032 22276 21036 22332
rect 21036 22276 21092 22332
rect 21092 22276 21096 22332
rect 21032 22272 21096 22276
rect 21112 22332 21176 22336
rect 21112 22276 21116 22332
rect 21116 22276 21172 22332
rect 21172 22276 21176 22332
rect 21112 22272 21176 22276
rect 21192 22332 21256 22336
rect 21192 22276 21196 22332
rect 21196 22276 21252 22332
rect 21252 22276 21256 22332
rect 21192 22272 21256 22276
rect 12204 22204 12268 22268
rect 12940 22204 13004 22268
rect 13492 22068 13556 22132
rect 9996 21992 10060 21996
rect 9996 21936 10010 21992
rect 10010 21936 10060 21992
rect 9996 21932 10060 21936
rect 14780 21932 14844 21996
rect 5952 21788 6016 21792
rect 5952 21732 5956 21788
rect 5956 21732 6012 21788
rect 6012 21732 6016 21788
rect 5952 21728 6016 21732
rect 6032 21788 6096 21792
rect 6032 21732 6036 21788
rect 6036 21732 6092 21788
rect 6092 21732 6096 21788
rect 6032 21728 6096 21732
rect 6112 21788 6176 21792
rect 6112 21732 6116 21788
rect 6116 21732 6172 21788
rect 6172 21732 6176 21788
rect 6112 21728 6176 21732
rect 6192 21788 6256 21792
rect 6192 21732 6196 21788
rect 6196 21732 6252 21788
rect 6252 21732 6256 21788
rect 6192 21728 6256 21732
rect 15952 21788 16016 21792
rect 15952 21732 15956 21788
rect 15956 21732 16012 21788
rect 16012 21732 16016 21788
rect 15952 21728 16016 21732
rect 16032 21788 16096 21792
rect 16032 21732 16036 21788
rect 16036 21732 16092 21788
rect 16092 21732 16096 21788
rect 16032 21728 16096 21732
rect 16112 21788 16176 21792
rect 16112 21732 16116 21788
rect 16116 21732 16172 21788
rect 16172 21732 16176 21788
rect 16112 21728 16176 21732
rect 16192 21788 16256 21792
rect 16192 21732 16196 21788
rect 16196 21732 16252 21788
rect 16252 21732 16256 21788
rect 16192 21728 16256 21732
rect 25952 21788 26016 21792
rect 25952 21732 25956 21788
rect 25956 21732 26012 21788
rect 26012 21732 26016 21788
rect 25952 21728 26016 21732
rect 26032 21788 26096 21792
rect 26032 21732 26036 21788
rect 26036 21732 26092 21788
rect 26092 21732 26096 21788
rect 26032 21728 26096 21732
rect 26112 21788 26176 21792
rect 26112 21732 26116 21788
rect 26116 21732 26172 21788
rect 26172 21732 26176 21788
rect 26112 21728 26176 21732
rect 26192 21788 26256 21792
rect 26192 21732 26196 21788
rect 26196 21732 26252 21788
rect 26252 21732 26256 21788
rect 26192 21728 26256 21732
rect 10732 21720 10796 21724
rect 10732 21664 10782 21720
rect 10782 21664 10796 21720
rect 10732 21660 10796 21664
rect 18092 21720 18156 21724
rect 18092 21664 18106 21720
rect 18106 21664 18156 21720
rect 18092 21660 18156 21664
rect 10952 21244 11016 21248
rect 10952 21188 10956 21244
rect 10956 21188 11012 21244
rect 11012 21188 11016 21244
rect 10952 21184 11016 21188
rect 11032 21244 11096 21248
rect 11032 21188 11036 21244
rect 11036 21188 11092 21244
rect 11092 21188 11096 21244
rect 11032 21184 11096 21188
rect 11112 21244 11176 21248
rect 11112 21188 11116 21244
rect 11116 21188 11172 21244
rect 11172 21188 11176 21244
rect 11112 21184 11176 21188
rect 11192 21244 11256 21248
rect 11192 21188 11196 21244
rect 11196 21188 11252 21244
rect 11252 21188 11256 21244
rect 11192 21184 11256 21188
rect 20952 21244 21016 21248
rect 20952 21188 20956 21244
rect 20956 21188 21012 21244
rect 21012 21188 21016 21244
rect 20952 21184 21016 21188
rect 21032 21244 21096 21248
rect 21032 21188 21036 21244
rect 21036 21188 21092 21244
rect 21092 21188 21096 21244
rect 21032 21184 21096 21188
rect 21112 21244 21176 21248
rect 21112 21188 21116 21244
rect 21116 21188 21172 21244
rect 21172 21188 21176 21244
rect 21112 21184 21176 21188
rect 21192 21244 21256 21248
rect 21192 21188 21196 21244
rect 21196 21188 21252 21244
rect 21252 21188 21256 21244
rect 21192 21184 21256 21188
rect 5952 20700 6016 20704
rect 5952 20644 5956 20700
rect 5956 20644 6012 20700
rect 6012 20644 6016 20700
rect 5952 20640 6016 20644
rect 6032 20700 6096 20704
rect 6032 20644 6036 20700
rect 6036 20644 6092 20700
rect 6092 20644 6096 20700
rect 6032 20640 6096 20644
rect 6112 20700 6176 20704
rect 6112 20644 6116 20700
rect 6116 20644 6172 20700
rect 6172 20644 6176 20700
rect 6112 20640 6176 20644
rect 6192 20700 6256 20704
rect 6192 20644 6196 20700
rect 6196 20644 6252 20700
rect 6252 20644 6256 20700
rect 6192 20640 6256 20644
rect 15952 20700 16016 20704
rect 15952 20644 15956 20700
rect 15956 20644 16012 20700
rect 16012 20644 16016 20700
rect 15952 20640 16016 20644
rect 16032 20700 16096 20704
rect 16032 20644 16036 20700
rect 16036 20644 16092 20700
rect 16092 20644 16096 20700
rect 16032 20640 16096 20644
rect 16112 20700 16176 20704
rect 16112 20644 16116 20700
rect 16116 20644 16172 20700
rect 16172 20644 16176 20700
rect 16112 20640 16176 20644
rect 16192 20700 16256 20704
rect 16192 20644 16196 20700
rect 16196 20644 16252 20700
rect 16252 20644 16256 20700
rect 16192 20640 16256 20644
rect 14964 20436 15028 20500
rect 25952 20700 26016 20704
rect 25952 20644 25956 20700
rect 25956 20644 26012 20700
rect 26012 20644 26016 20700
rect 25952 20640 26016 20644
rect 26032 20700 26096 20704
rect 26032 20644 26036 20700
rect 26036 20644 26092 20700
rect 26092 20644 26096 20700
rect 26032 20640 26096 20644
rect 26112 20700 26176 20704
rect 26112 20644 26116 20700
rect 26116 20644 26172 20700
rect 26172 20644 26176 20700
rect 26112 20640 26176 20644
rect 26192 20700 26256 20704
rect 26192 20644 26196 20700
rect 26196 20644 26252 20700
rect 26252 20644 26256 20700
rect 26192 20640 26256 20644
rect 12204 20300 12268 20364
rect 9628 20224 9692 20228
rect 9628 20168 9678 20224
rect 9678 20168 9692 20224
rect 9628 20164 9692 20168
rect 10952 20156 11016 20160
rect 10952 20100 10956 20156
rect 10956 20100 11012 20156
rect 11012 20100 11016 20156
rect 10952 20096 11016 20100
rect 11032 20156 11096 20160
rect 11032 20100 11036 20156
rect 11036 20100 11092 20156
rect 11092 20100 11096 20156
rect 11032 20096 11096 20100
rect 11112 20156 11176 20160
rect 11112 20100 11116 20156
rect 11116 20100 11172 20156
rect 11172 20100 11176 20156
rect 11112 20096 11176 20100
rect 11192 20156 11256 20160
rect 11192 20100 11196 20156
rect 11196 20100 11252 20156
rect 11252 20100 11256 20156
rect 11192 20096 11256 20100
rect 20952 20156 21016 20160
rect 20952 20100 20956 20156
rect 20956 20100 21012 20156
rect 21012 20100 21016 20156
rect 20952 20096 21016 20100
rect 21032 20156 21096 20160
rect 21032 20100 21036 20156
rect 21036 20100 21092 20156
rect 21092 20100 21096 20156
rect 21032 20096 21096 20100
rect 21112 20156 21176 20160
rect 21112 20100 21116 20156
rect 21116 20100 21172 20156
rect 21172 20100 21176 20156
rect 21112 20096 21176 20100
rect 21192 20156 21256 20160
rect 21192 20100 21196 20156
rect 21196 20100 21252 20156
rect 21252 20100 21256 20156
rect 21192 20096 21256 20100
rect 11468 19756 11532 19820
rect 5952 19612 6016 19616
rect 5952 19556 5956 19612
rect 5956 19556 6012 19612
rect 6012 19556 6016 19612
rect 5952 19552 6016 19556
rect 6032 19612 6096 19616
rect 6032 19556 6036 19612
rect 6036 19556 6092 19612
rect 6092 19556 6096 19612
rect 6032 19552 6096 19556
rect 6112 19612 6176 19616
rect 6112 19556 6116 19612
rect 6116 19556 6172 19612
rect 6172 19556 6176 19612
rect 6112 19552 6176 19556
rect 6192 19612 6256 19616
rect 6192 19556 6196 19612
rect 6196 19556 6252 19612
rect 6252 19556 6256 19612
rect 6192 19552 6256 19556
rect 15952 19612 16016 19616
rect 15952 19556 15956 19612
rect 15956 19556 16012 19612
rect 16012 19556 16016 19612
rect 15952 19552 16016 19556
rect 16032 19612 16096 19616
rect 16032 19556 16036 19612
rect 16036 19556 16092 19612
rect 16092 19556 16096 19612
rect 16032 19552 16096 19556
rect 16112 19612 16176 19616
rect 16112 19556 16116 19612
rect 16116 19556 16172 19612
rect 16172 19556 16176 19612
rect 16112 19552 16176 19556
rect 16192 19612 16256 19616
rect 16192 19556 16196 19612
rect 16196 19556 16252 19612
rect 16252 19556 16256 19612
rect 16192 19552 16256 19556
rect 25952 19612 26016 19616
rect 25952 19556 25956 19612
rect 25956 19556 26012 19612
rect 26012 19556 26016 19612
rect 25952 19552 26016 19556
rect 26032 19612 26096 19616
rect 26032 19556 26036 19612
rect 26036 19556 26092 19612
rect 26092 19556 26096 19612
rect 26032 19552 26096 19556
rect 26112 19612 26176 19616
rect 26112 19556 26116 19612
rect 26116 19556 26172 19612
rect 26172 19556 26176 19612
rect 26112 19552 26176 19556
rect 26192 19612 26256 19616
rect 26192 19556 26196 19612
rect 26196 19556 26252 19612
rect 26252 19556 26256 19612
rect 26192 19552 26256 19556
rect 9076 19272 9140 19276
rect 9076 19216 9090 19272
rect 9090 19216 9140 19272
rect 9076 19212 9140 19216
rect 10952 19068 11016 19072
rect 10952 19012 10956 19068
rect 10956 19012 11012 19068
rect 11012 19012 11016 19068
rect 10952 19008 11016 19012
rect 11032 19068 11096 19072
rect 11032 19012 11036 19068
rect 11036 19012 11092 19068
rect 11092 19012 11096 19068
rect 11032 19008 11096 19012
rect 11112 19068 11176 19072
rect 11112 19012 11116 19068
rect 11116 19012 11172 19068
rect 11172 19012 11176 19068
rect 11112 19008 11176 19012
rect 11192 19068 11256 19072
rect 11192 19012 11196 19068
rect 11196 19012 11252 19068
rect 11252 19012 11256 19068
rect 11192 19008 11256 19012
rect 20952 19068 21016 19072
rect 20952 19012 20956 19068
rect 20956 19012 21012 19068
rect 21012 19012 21016 19068
rect 20952 19008 21016 19012
rect 21032 19068 21096 19072
rect 21032 19012 21036 19068
rect 21036 19012 21092 19068
rect 21092 19012 21096 19068
rect 21032 19008 21096 19012
rect 21112 19068 21176 19072
rect 21112 19012 21116 19068
rect 21116 19012 21172 19068
rect 21172 19012 21176 19068
rect 21112 19008 21176 19012
rect 21192 19068 21256 19072
rect 21192 19012 21196 19068
rect 21196 19012 21252 19068
rect 21252 19012 21256 19068
rect 21192 19008 21256 19012
rect 10548 18864 10612 18868
rect 10548 18808 10562 18864
rect 10562 18808 10612 18864
rect 10548 18804 10612 18808
rect 5952 18524 6016 18528
rect 5952 18468 5956 18524
rect 5956 18468 6012 18524
rect 6012 18468 6016 18524
rect 5952 18464 6016 18468
rect 6032 18524 6096 18528
rect 6032 18468 6036 18524
rect 6036 18468 6092 18524
rect 6092 18468 6096 18524
rect 6032 18464 6096 18468
rect 6112 18524 6176 18528
rect 6112 18468 6116 18524
rect 6116 18468 6172 18524
rect 6172 18468 6176 18524
rect 6112 18464 6176 18468
rect 6192 18524 6256 18528
rect 6192 18468 6196 18524
rect 6196 18468 6252 18524
rect 6252 18468 6256 18524
rect 6192 18464 6256 18468
rect 15952 18524 16016 18528
rect 15952 18468 15956 18524
rect 15956 18468 16012 18524
rect 16012 18468 16016 18524
rect 15952 18464 16016 18468
rect 16032 18524 16096 18528
rect 16032 18468 16036 18524
rect 16036 18468 16092 18524
rect 16092 18468 16096 18524
rect 16032 18464 16096 18468
rect 16112 18524 16176 18528
rect 16112 18468 16116 18524
rect 16116 18468 16172 18524
rect 16172 18468 16176 18524
rect 16112 18464 16176 18468
rect 16192 18524 16256 18528
rect 16192 18468 16196 18524
rect 16196 18468 16252 18524
rect 16252 18468 16256 18524
rect 16192 18464 16256 18468
rect 25952 18524 26016 18528
rect 25952 18468 25956 18524
rect 25956 18468 26012 18524
rect 26012 18468 26016 18524
rect 25952 18464 26016 18468
rect 26032 18524 26096 18528
rect 26032 18468 26036 18524
rect 26036 18468 26092 18524
rect 26092 18468 26096 18524
rect 26032 18464 26096 18468
rect 26112 18524 26176 18528
rect 26112 18468 26116 18524
rect 26116 18468 26172 18524
rect 26172 18468 26176 18524
rect 26112 18464 26176 18468
rect 26192 18524 26256 18528
rect 26192 18468 26196 18524
rect 26196 18468 26252 18524
rect 26252 18468 26256 18524
rect 26192 18464 26256 18468
rect 12388 18260 12452 18324
rect 14596 18124 14660 18188
rect 10952 17980 11016 17984
rect 10952 17924 10956 17980
rect 10956 17924 11012 17980
rect 11012 17924 11016 17980
rect 10952 17920 11016 17924
rect 11032 17980 11096 17984
rect 11032 17924 11036 17980
rect 11036 17924 11092 17980
rect 11092 17924 11096 17980
rect 11032 17920 11096 17924
rect 11112 17980 11176 17984
rect 11112 17924 11116 17980
rect 11116 17924 11172 17980
rect 11172 17924 11176 17980
rect 11112 17920 11176 17924
rect 11192 17980 11256 17984
rect 11192 17924 11196 17980
rect 11196 17924 11252 17980
rect 11252 17924 11256 17980
rect 11192 17920 11256 17924
rect 20952 17980 21016 17984
rect 20952 17924 20956 17980
rect 20956 17924 21012 17980
rect 21012 17924 21016 17980
rect 20952 17920 21016 17924
rect 21032 17980 21096 17984
rect 21032 17924 21036 17980
rect 21036 17924 21092 17980
rect 21092 17924 21096 17980
rect 21032 17920 21096 17924
rect 21112 17980 21176 17984
rect 21112 17924 21116 17980
rect 21116 17924 21172 17980
rect 21172 17924 21176 17980
rect 21112 17920 21176 17924
rect 21192 17980 21256 17984
rect 21192 17924 21196 17980
rect 21196 17924 21252 17980
rect 21252 17924 21256 17980
rect 21192 17920 21256 17924
rect 17172 17716 17236 17780
rect 5952 17436 6016 17440
rect 5952 17380 5956 17436
rect 5956 17380 6012 17436
rect 6012 17380 6016 17436
rect 5952 17376 6016 17380
rect 6032 17436 6096 17440
rect 6032 17380 6036 17436
rect 6036 17380 6092 17436
rect 6092 17380 6096 17436
rect 6032 17376 6096 17380
rect 6112 17436 6176 17440
rect 6112 17380 6116 17436
rect 6116 17380 6172 17436
rect 6172 17380 6176 17436
rect 6112 17376 6176 17380
rect 6192 17436 6256 17440
rect 6192 17380 6196 17436
rect 6196 17380 6252 17436
rect 6252 17380 6256 17436
rect 6192 17376 6256 17380
rect 15952 17436 16016 17440
rect 15952 17380 15956 17436
rect 15956 17380 16012 17436
rect 16012 17380 16016 17436
rect 15952 17376 16016 17380
rect 16032 17436 16096 17440
rect 16032 17380 16036 17436
rect 16036 17380 16092 17436
rect 16092 17380 16096 17436
rect 16032 17376 16096 17380
rect 16112 17436 16176 17440
rect 16112 17380 16116 17436
rect 16116 17380 16172 17436
rect 16172 17380 16176 17436
rect 16112 17376 16176 17380
rect 16192 17436 16256 17440
rect 16192 17380 16196 17436
rect 16196 17380 16252 17436
rect 16252 17380 16256 17436
rect 16192 17376 16256 17380
rect 25952 17436 26016 17440
rect 25952 17380 25956 17436
rect 25956 17380 26012 17436
rect 26012 17380 26016 17436
rect 25952 17376 26016 17380
rect 26032 17436 26096 17440
rect 26032 17380 26036 17436
rect 26036 17380 26092 17436
rect 26092 17380 26096 17436
rect 26032 17376 26096 17380
rect 26112 17436 26176 17440
rect 26112 17380 26116 17436
rect 26116 17380 26172 17436
rect 26172 17380 26176 17436
rect 26112 17376 26176 17380
rect 26192 17436 26256 17440
rect 26192 17380 26196 17436
rect 26196 17380 26252 17436
rect 26252 17380 26256 17436
rect 26192 17376 26256 17380
rect 10952 16892 11016 16896
rect 10952 16836 10956 16892
rect 10956 16836 11012 16892
rect 11012 16836 11016 16892
rect 10952 16832 11016 16836
rect 11032 16892 11096 16896
rect 11032 16836 11036 16892
rect 11036 16836 11092 16892
rect 11092 16836 11096 16892
rect 11032 16832 11096 16836
rect 11112 16892 11176 16896
rect 11112 16836 11116 16892
rect 11116 16836 11172 16892
rect 11172 16836 11176 16892
rect 11112 16832 11176 16836
rect 11192 16892 11256 16896
rect 11192 16836 11196 16892
rect 11196 16836 11252 16892
rect 11252 16836 11256 16892
rect 11192 16832 11256 16836
rect 20952 16892 21016 16896
rect 20952 16836 20956 16892
rect 20956 16836 21012 16892
rect 21012 16836 21016 16892
rect 20952 16832 21016 16836
rect 21032 16892 21096 16896
rect 21032 16836 21036 16892
rect 21036 16836 21092 16892
rect 21092 16836 21096 16892
rect 21032 16832 21096 16836
rect 21112 16892 21176 16896
rect 21112 16836 21116 16892
rect 21116 16836 21172 16892
rect 21172 16836 21176 16892
rect 21112 16832 21176 16836
rect 21192 16892 21256 16896
rect 21192 16836 21196 16892
rect 21196 16836 21252 16892
rect 21252 16836 21256 16892
rect 21192 16832 21256 16836
rect 5952 16348 6016 16352
rect 5952 16292 5956 16348
rect 5956 16292 6012 16348
rect 6012 16292 6016 16348
rect 5952 16288 6016 16292
rect 6032 16348 6096 16352
rect 6032 16292 6036 16348
rect 6036 16292 6092 16348
rect 6092 16292 6096 16348
rect 6032 16288 6096 16292
rect 6112 16348 6176 16352
rect 6112 16292 6116 16348
rect 6116 16292 6172 16348
rect 6172 16292 6176 16348
rect 6112 16288 6176 16292
rect 6192 16348 6256 16352
rect 6192 16292 6196 16348
rect 6196 16292 6252 16348
rect 6252 16292 6256 16348
rect 6192 16288 6256 16292
rect 15952 16348 16016 16352
rect 15952 16292 15956 16348
rect 15956 16292 16012 16348
rect 16012 16292 16016 16348
rect 15952 16288 16016 16292
rect 16032 16348 16096 16352
rect 16032 16292 16036 16348
rect 16036 16292 16092 16348
rect 16092 16292 16096 16348
rect 16032 16288 16096 16292
rect 16112 16348 16176 16352
rect 16112 16292 16116 16348
rect 16116 16292 16172 16348
rect 16172 16292 16176 16348
rect 16112 16288 16176 16292
rect 16192 16348 16256 16352
rect 16192 16292 16196 16348
rect 16196 16292 16252 16348
rect 16252 16292 16256 16348
rect 16192 16288 16256 16292
rect 25952 16348 26016 16352
rect 25952 16292 25956 16348
rect 25956 16292 26012 16348
rect 26012 16292 26016 16348
rect 25952 16288 26016 16292
rect 26032 16348 26096 16352
rect 26032 16292 26036 16348
rect 26036 16292 26092 16348
rect 26092 16292 26096 16348
rect 26032 16288 26096 16292
rect 26112 16348 26176 16352
rect 26112 16292 26116 16348
rect 26116 16292 26172 16348
rect 26172 16292 26176 16348
rect 26112 16288 26176 16292
rect 26192 16348 26256 16352
rect 26192 16292 26196 16348
rect 26196 16292 26252 16348
rect 26252 16292 26256 16348
rect 26192 16288 26256 16292
rect 10952 15804 11016 15808
rect 10952 15748 10956 15804
rect 10956 15748 11012 15804
rect 11012 15748 11016 15804
rect 10952 15744 11016 15748
rect 11032 15804 11096 15808
rect 11032 15748 11036 15804
rect 11036 15748 11092 15804
rect 11092 15748 11096 15804
rect 11032 15744 11096 15748
rect 11112 15804 11176 15808
rect 11112 15748 11116 15804
rect 11116 15748 11172 15804
rect 11172 15748 11176 15804
rect 11112 15744 11176 15748
rect 11192 15804 11256 15808
rect 11192 15748 11196 15804
rect 11196 15748 11252 15804
rect 11252 15748 11256 15804
rect 11192 15744 11256 15748
rect 20952 15804 21016 15808
rect 20952 15748 20956 15804
rect 20956 15748 21012 15804
rect 21012 15748 21016 15804
rect 20952 15744 21016 15748
rect 21032 15804 21096 15808
rect 21032 15748 21036 15804
rect 21036 15748 21092 15804
rect 21092 15748 21096 15804
rect 21032 15744 21096 15748
rect 21112 15804 21176 15808
rect 21112 15748 21116 15804
rect 21116 15748 21172 15804
rect 21172 15748 21176 15804
rect 21112 15744 21176 15748
rect 21192 15804 21256 15808
rect 21192 15748 21196 15804
rect 21196 15748 21252 15804
rect 21252 15748 21256 15804
rect 21192 15744 21256 15748
rect 5952 15260 6016 15264
rect 5952 15204 5956 15260
rect 5956 15204 6012 15260
rect 6012 15204 6016 15260
rect 5952 15200 6016 15204
rect 6032 15260 6096 15264
rect 6032 15204 6036 15260
rect 6036 15204 6092 15260
rect 6092 15204 6096 15260
rect 6032 15200 6096 15204
rect 6112 15260 6176 15264
rect 6112 15204 6116 15260
rect 6116 15204 6172 15260
rect 6172 15204 6176 15260
rect 6112 15200 6176 15204
rect 6192 15260 6256 15264
rect 6192 15204 6196 15260
rect 6196 15204 6252 15260
rect 6252 15204 6256 15260
rect 6192 15200 6256 15204
rect 15952 15260 16016 15264
rect 15952 15204 15956 15260
rect 15956 15204 16012 15260
rect 16012 15204 16016 15260
rect 15952 15200 16016 15204
rect 16032 15260 16096 15264
rect 16032 15204 16036 15260
rect 16036 15204 16092 15260
rect 16092 15204 16096 15260
rect 16032 15200 16096 15204
rect 16112 15260 16176 15264
rect 16112 15204 16116 15260
rect 16116 15204 16172 15260
rect 16172 15204 16176 15260
rect 16112 15200 16176 15204
rect 16192 15260 16256 15264
rect 16192 15204 16196 15260
rect 16196 15204 16252 15260
rect 16252 15204 16256 15260
rect 16192 15200 16256 15204
rect 12756 14996 12820 15060
rect 25952 15260 26016 15264
rect 25952 15204 25956 15260
rect 25956 15204 26012 15260
rect 26012 15204 26016 15260
rect 25952 15200 26016 15204
rect 26032 15260 26096 15264
rect 26032 15204 26036 15260
rect 26036 15204 26092 15260
rect 26092 15204 26096 15260
rect 26032 15200 26096 15204
rect 26112 15260 26176 15264
rect 26112 15204 26116 15260
rect 26116 15204 26172 15260
rect 26172 15204 26176 15260
rect 26112 15200 26176 15204
rect 26192 15260 26256 15264
rect 26192 15204 26196 15260
rect 26196 15204 26252 15260
rect 26252 15204 26256 15260
rect 26192 15200 26256 15204
rect 10952 14716 11016 14720
rect 10952 14660 10956 14716
rect 10956 14660 11012 14716
rect 11012 14660 11016 14716
rect 10952 14656 11016 14660
rect 11032 14716 11096 14720
rect 11032 14660 11036 14716
rect 11036 14660 11092 14716
rect 11092 14660 11096 14716
rect 11032 14656 11096 14660
rect 11112 14716 11176 14720
rect 11112 14660 11116 14716
rect 11116 14660 11172 14716
rect 11172 14660 11176 14716
rect 11112 14656 11176 14660
rect 11192 14716 11256 14720
rect 11192 14660 11196 14716
rect 11196 14660 11252 14716
rect 11252 14660 11256 14716
rect 11192 14656 11256 14660
rect 20952 14716 21016 14720
rect 20952 14660 20956 14716
rect 20956 14660 21012 14716
rect 21012 14660 21016 14716
rect 20952 14656 21016 14660
rect 21032 14716 21096 14720
rect 21032 14660 21036 14716
rect 21036 14660 21092 14716
rect 21092 14660 21096 14716
rect 21032 14656 21096 14660
rect 21112 14716 21176 14720
rect 21112 14660 21116 14716
rect 21116 14660 21172 14716
rect 21172 14660 21176 14716
rect 21112 14656 21176 14660
rect 21192 14716 21256 14720
rect 21192 14660 21196 14716
rect 21196 14660 21252 14716
rect 21252 14660 21256 14716
rect 21192 14656 21256 14660
rect 5952 14172 6016 14176
rect 5952 14116 5956 14172
rect 5956 14116 6012 14172
rect 6012 14116 6016 14172
rect 5952 14112 6016 14116
rect 6032 14172 6096 14176
rect 6032 14116 6036 14172
rect 6036 14116 6092 14172
rect 6092 14116 6096 14172
rect 6032 14112 6096 14116
rect 6112 14172 6176 14176
rect 6112 14116 6116 14172
rect 6116 14116 6172 14172
rect 6172 14116 6176 14172
rect 6112 14112 6176 14116
rect 6192 14172 6256 14176
rect 6192 14116 6196 14172
rect 6196 14116 6252 14172
rect 6252 14116 6256 14172
rect 6192 14112 6256 14116
rect 15952 14172 16016 14176
rect 15952 14116 15956 14172
rect 15956 14116 16012 14172
rect 16012 14116 16016 14172
rect 15952 14112 16016 14116
rect 16032 14172 16096 14176
rect 16032 14116 16036 14172
rect 16036 14116 16092 14172
rect 16092 14116 16096 14172
rect 16032 14112 16096 14116
rect 16112 14172 16176 14176
rect 16112 14116 16116 14172
rect 16116 14116 16172 14172
rect 16172 14116 16176 14172
rect 16112 14112 16176 14116
rect 16192 14172 16256 14176
rect 16192 14116 16196 14172
rect 16196 14116 16252 14172
rect 16252 14116 16256 14172
rect 16192 14112 16256 14116
rect 25952 14172 26016 14176
rect 25952 14116 25956 14172
rect 25956 14116 26012 14172
rect 26012 14116 26016 14172
rect 25952 14112 26016 14116
rect 26032 14172 26096 14176
rect 26032 14116 26036 14172
rect 26036 14116 26092 14172
rect 26092 14116 26096 14172
rect 26032 14112 26096 14116
rect 26112 14172 26176 14176
rect 26112 14116 26116 14172
rect 26116 14116 26172 14172
rect 26172 14116 26176 14172
rect 26112 14112 26176 14116
rect 26192 14172 26256 14176
rect 26192 14116 26196 14172
rect 26196 14116 26252 14172
rect 26252 14116 26256 14172
rect 26192 14112 26256 14116
rect 10952 13628 11016 13632
rect 10952 13572 10956 13628
rect 10956 13572 11012 13628
rect 11012 13572 11016 13628
rect 10952 13568 11016 13572
rect 11032 13628 11096 13632
rect 11032 13572 11036 13628
rect 11036 13572 11092 13628
rect 11092 13572 11096 13628
rect 11032 13568 11096 13572
rect 11112 13628 11176 13632
rect 11112 13572 11116 13628
rect 11116 13572 11172 13628
rect 11172 13572 11176 13628
rect 11112 13568 11176 13572
rect 11192 13628 11256 13632
rect 11192 13572 11196 13628
rect 11196 13572 11252 13628
rect 11252 13572 11256 13628
rect 11192 13568 11256 13572
rect 20952 13628 21016 13632
rect 20952 13572 20956 13628
rect 20956 13572 21012 13628
rect 21012 13572 21016 13628
rect 20952 13568 21016 13572
rect 21032 13628 21096 13632
rect 21032 13572 21036 13628
rect 21036 13572 21092 13628
rect 21092 13572 21096 13628
rect 21032 13568 21096 13572
rect 21112 13628 21176 13632
rect 21112 13572 21116 13628
rect 21116 13572 21172 13628
rect 21172 13572 21176 13628
rect 21112 13568 21176 13572
rect 21192 13628 21256 13632
rect 21192 13572 21196 13628
rect 21196 13572 21252 13628
rect 21252 13572 21256 13628
rect 21192 13568 21256 13572
rect 13676 13500 13740 13564
rect 5952 13084 6016 13088
rect 5952 13028 5956 13084
rect 5956 13028 6012 13084
rect 6012 13028 6016 13084
rect 5952 13024 6016 13028
rect 6032 13084 6096 13088
rect 6032 13028 6036 13084
rect 6036 13028 6092 13084
rect 6092 13028 6096 13084
rect 6032 13024 6096 13028
rect 6112 13084 6176 13088
rect 6112 13028 6116 13084
rect 6116 13028 6172 13084
rect 6172 13028 6176 13084
rect 6112 13024 6176 13028
rect 6192 13084 6256 13088
rect 6192 13028 6196 13084
rect 6196 13028 6252 13084
rect 6252 13028 6256 13084
rect 6192 13024 6256 13028
rect 15952 13084 16016 13088
rect 15952 13028 15956 13084
rect 15956 13028 16012 13084
rect 16012 13028 16016 13084
rect 15952 13024 16016 13028
rect 16032 13084 16096 13088
rect 16032 13028 16036 13084
rect 16036 13028 16092 13084
rect 16092 13028 16096 13084
rect 16032 13024 16096 13028
rect 16112 13084 16176 13088
rect 16112 13028 16116 13084
rect 16116 13028 16172 13084
rect 16172 13028 16176 13084
rect 16112 13024 16176 13028
rect 16192 13084 16256 13088
rect 16192 13028 16196 13084
rect 16196 13028 16252 13084
rect 16252 13028 16256 13084
rect 16192 13024 16256 13028
rect 25952 13084 26016 13088
rect 25952 13028 25956 13084
rect 25956 13028 26012 13084
rect 26012 13028 26016 13084
rect 25952 13024 26016 13028
rect 26032 13084 26096 13088
rect 26032 13028 26036 13084
rect 26036 13028 26092 13084
rect 26092 13028 26096 13084
rect 26032 13024 26096 13028
rect 26112 13084 26176 13088
rect 26112 13028 26116 13084
rect 26116 13028 26172 13084
rect 26172 13028 26176 13084
rect 26112 13024 26176 13028
rect 26192 13084 26256 13088
rect 26192 13028 26196 13084
rect 26196 13028 26252 13084
rect 26252 13028 26256 13084
rect 26192 13024 26256 13028
rect 12020 12684 12084 12748
rect 19380 12684 19444 12748
rect 10952 12540 11016 12544
rect 10952 12484 10956 12540
rect 10956 12484 11012 12540
rect 11012 12484 11016 12540
rect 10952 12480 11016 12484
rect 11032 12540 11096 12544
rect 11032 12484 11036 12540
rect 11036 12484 11092 12540
rect 11092 12484 11096 12540
rect 11032 12480 11096 12484
rect 11112 12540 11176 12544
rect 11112 12484 11116 12540
rect 11116 12484 11172 12540
rect 11172 12484 11176 12540
rect 11112 12480 11176 12484
rect 11192 12540 11256 12544
rect 11192 12484 11196 12540
rect 11196 12484 11252 12540
rect 11252 12484 11256 12540
rect 11192 12480 11256 12484
rect 20952 12540 21016 12544
rect 20952 12484 20956 12540
rect 20956 12484 21012 12540
rect 21012 12484 21016 12540
rect 20952 12480 21016 12484
rect 21032 12540 21096 12544
rect 21032 12484 21036 12540
rect 21036 12484 21092 12540
rect 21092 12484 21096 12540
rect 21032 12480 21096 12484
rect 21112 12540 21176 12544
rect 21112 12484 21116 12540
rect 21116 12484 21172 12540
rect 21172 12484 21176 12540
rect 21112 12480 21176 12484
rect 21192 12540 21256 12544
rect 21192 12484 21196 12540
rect 21196 12484 21252 12540
rect 21252 12484 21256 12540
rect 21192 12480 21256 12484
rect 19380 12276 19444 12340
rect 9076 12004 9140 12068
rect 5952 11996 6016 12000
rect 5952 11940 5956 11996
rect 5956 11940 6012 11996
rect 6012 11940 6016 11996
rect 5952 11936 6016 11940
rect 6032 11996 6096 12000
rect 6032 11940 6036 11996
rect 6036 11940 6092 11996
rect 6092 11940 6096 11996
rect 6032 11936 6096 11940
rect 6112 11996 6176 12000
rect 6112 11940 6116 11996
rect 6116 11940 6172 11996
rect 6172 11940 6176 11996
rect 6112 11936 6176 11940
rect 6192 11996 6256 12000
rect 6192 11940 6196 11996
rect 6196 11940 6252 11996
rect 6252 11940 6256 11996
rect 6192 11936 6256 11940
rect 15952 11996 16016 12000
rect 15952 11940 15956 11996
rect 15956 11940 16012 11996
rect 16012 11940 16016 11996
rect 15952 11936 16016 11940
rect 16032 11996 16096 12000
rect 16032 11940 16036 11996
rect 16036 11940 16092 11996
rect 16092 11940 16096 11996
rect 16032 11936 16096 11940
rect 16112 11996 16176 12000
rect 16112 11940 16116 11996
rect 16116 11940 16172 11996
rect 16172 11940 16176 11996
rect 16112 11936 16176 11940
rect 16192 11996 16256 12000
rect 16192 11940 16196 11996
rect 16196 11940 16252 11996
rect 16252 11940 16256 11996
rect 16192 11936 16256 11940
rect 25952 11996 26016 12000
rect 25952 11940 25956 11996
rect 25956 11940 26012 11996
rect 26012 11940 26016 11996
rect 25952 11936 26016 11940
rect 26032 11996 26096 12000
rect 26032 11940 26036 11996
rect 26036 11940 26092 11996
rect 26092 11940 26096 11996
rect 26032 11936 26096 11940
rect 26112 11996 26176 12000
rect 26112 11940 26116 11996
rect 26116 11940 26172 11996
rect 26172 11940 26176 11996
rect 26112 11936 26176 11940
rect 26192 11996 26256 12000
rect 26192 11940 26196 11996
rect 26196 11940 26252 11996
rect 26252 11940 26256 11996
rect 26192 11936 26256 11940
rect 10952 11452 11016 11456
rect 10952 11396 10956 11452
rect 10956 11396 11012 11452
rect 11012 11396 11016 11452
rect 10952 11392 11016 11396
rect 11032 11452 11096 11456
rect 11032 11396 11036 11452
rect 11036 11396 11092 11452
rect 11092 11396 11096 11452
rect 11032 11392 11096 11396
rect 11112 11452 11176 11456
rect 11112 11396 11116 11452
rect 11116 11396 11172 11452
rect 11172 11396 11176 11452
rect 11112 11392 11176 11396
rect 11192 11452 11256 11456
rect 11192 11396 11196 11452
rect 11196 11396 11252 11452
rect 11252 11396 11256 11452
rect 11192 11392 11256 11396
rect 20952 11452 21016 11456
rect 20952 11396 20956 11452
rect 20956 11396 21012 11452
rect 21012 11396 21016 11452
rect 20952 11392 21016 11396
rect 21032 11452 21096 11456
rect 21032 11396 21036 11452
rect 21036 11396 21092 11452
rect 21092 11396 21096 11452
rect 21032 11392 21096 11396
rect 21112 11452 21176 11456
rect 21112 11396 21116 11452
rect 21116 11396 21172 11452
rect 21172 11396 21176 11452
rect 21112 11392 21176 11396
rect 21192 11452 21256 11456
rect 21192 11396 21196 11452
rect 21196 11396 21252 11452
rect 21252 11396 21256 11452
rect 21192 11392 21256 11396
rect 15700 11324 15764 11388
rect 5952 10908 6016 10912
rect 5952 10852 5956 10908
rect 5956 10852 6012 10908
rect 6012 10852 6016 10908
rect 5952 10848 6016 10852
rect 6032 10908 6096 10912
rect 6032 10852 6036 10908
rect 6036 10852 6092 10908
rect 6092 10852 6096 10908
rect 6032 10848 6096 10852
rect 6112 10908 6176 10912
rect 6112 10852 6116 10908
rect 6116 10852 6172 10908
rect 6172 10852 6176 10908
rect 6112 10848 6176 10852
rect 6192 10908 6256 10912
rect 6192 10852 6196 10908
rect 6196 10852 6252 10908
rect 6252 10852 6256 10908
rect 6192 10848 6256 10852
rect 15952 10908 16016 10912
rect 15952 10852 15956 10908
rect 15956 10852 16012 10908
rect 16012 10852 16016 10908
rect 15952 10848 16016 10852
rect 16032 10908 16096 10912
rect 16032 10852 16036 10908
rect 16036 10852 16092 10908
rect 16092 10852 16096 10908
rect 16032 10848 16096 10852
rect 16112 10908 16176 10912
rect 16112 10852 16116 10908
rect 16116 10852 16172 10908
rect 16172 10852 16176 10908
rect 16112 10848 16176 10852
rect 16192 10908 16256 10912
rect 16192 10852 16196 10908
rect 16196 10852 16252 10908
rect 16252 10852 16256 10908
rect 16192 10848 16256 10852
rect 25952 10908 26016 10912
rect 25952 10852 25956 10908
rect 25956 10852 26012 10908
rect 26012 10852 26016 10908
rect 25952 10848 26016 10852
rect 26032 10908 26096 10912
rect 26032 10852 26036 10908
rect 26036 10852 26092 10908
rect 26092 10852 26096 10908
rect 26032 10848 26096 10852
rect 26112 10908 26176 10912
rect 26112 10852 26116 10908
rect 26116 10852 26172 10908
rect 26172 10852 26176 10908
rect 26112 10848 26176 10852
rect 26192 10908 26256 10912
rect 26192 10852 26196 10908
rect 26196 10852 26252 10908
rect 26252 10852 26256 10908
rect 26192 10848 26256 10852
rect 10548 10780 10612 10844
rect 10952 10364 11016 10368
rect 10952 10308 10956 10364
rect 10956 10308 11012 10364
rect 11012 10308 11016 10364
rect 10952 10304 11016 10308
rect 11032 10364 11096 10368
rect 11032 10308 11036 10364
rect 11036 10308 11092 10364
rect 11092 10308 11096 10364
rect 11032 10304 11096 10308
rect 11112 10364 11176 10368
rect 11112 10308 11116 10364
rect 11116 10308 11172 10364
rect 11172 10308 11176 10364
rect 11112 10304 11176 10308
rect 11192 10364 11256 10368
rect 11192 10308 11196 10364
rect 11196 10308 11252 10364
rect 11252 10308 11256 10364
rect 11192 10304 11256 10308
rect 20952 10364 21016 10368
rect 20952 10308 20956 10364
rect 20956 10308 21012 10364
rect 21012 10308 21016 10364
rect 20952 10304 21016 10308
rect 21032 10364 21096 10368
rect 21032 10308 21036 10364
rect 21036 10308 21092 10364
rect 21092 10308 21096 10364
rect 21032 10304 21096 10308
rect 21112 10364 21176 10368
rect 21112 10308 21116 10364
rect 21116 10308 21172 10364
rect 21172 10308 21176 10364
rect 21112 10304 21176 10308
rect 21192 10364 21256 10368
rect 21192 10308 21196 10364
rect 21196 10308 21252 10364
rect 21252 10308 21256 10364
rect 21192 10304 21256 10308
rect 5952 9820 6016 9824
rect 5952 9764 5956 9820
rect 5956 9764 6012 9820
rect 6012 9764 6016 9820
rect 5952 9760 6016 9764
rect 6032 9820 6096 9824
rect 6032 9764 6036 9820
rect 6036 9764 6092 9820
rect 6092 9764 6096 9820
rect 6032 9760 6096 9764
rect 6112 9820 6176 9824
rect 6112 9764 6116 9820
rect 6116 9764 6172 9820
rect 6172 9764 6176 9820
rect 6112 9760 6176 9764
rect 6192 9820 6256 9824
rect 6192 9764 6196 9820
rect 6196 9764 6252 9820
rect 6252 9764 6256 9820
rect 6192 9760 6256 9764
rect 15952 9820 16016 9824
rect 15952 9764 15956 9820
rect 15956 9764 16012 9820
rect 16012 9764 16016 9820
rect 15952 9760 16016 9764
rect 16032 9820 16096 9824
rect 16032 9764 16036 9820
rect 16036 9764 16092 9820
rect 16092 9764 16096 9820
rect 16032 9760 16096 9764
rect 16112 9820 16176 9824
rect 16112 9764 16116 9820
rect 16116 9764 16172 9820
rect 16172 9764 16176 9820
rect 16112 9760 16176 9764
rect 16192 9820 16256 9824
rect 16192 9764 16196 9820
rect 16196 9764 16252 9820
rect 16252 9764 16256 9820
rect 16192 9760 16256 9764
rect 25952 9820 26016 9824
rect 25952 9764 25956 9820
rect 25956 9764 26012 9820
rect 26012 9764 26016 9820
rect 25952 9760 26016 9764
rect 26032 9820 26096 9824
rect 26032 9764 26036 9820
rect 26036 9764 26092 9820
rect 26092 9764 26096 9820
rect 26032 9760 26096 9764
rect 26112 9820 26176 9824
rect 26112 9764 26116 9820
rect 26116 9764 26172 9820
rect 26172 9764 26176 9820
rect 26112 9760 26176 9764
rect 26192 9820 26256 9824
rect 26192 9764 26196 9820
rect 26196 9764 26252 9820
rect 26252 9764 26256 9820
rect 26192 9760 26256 9764
rect 10952 9276 11016 9280
rect 10952 9220 10956 9276
rect 10956 9220 11012 9276
rect 11012 9220 11016 9276
rect 10952 9216 11016 9220
rect 11032 9276 11096 9280
rect 11032 9220 11036 9276
rect 11036 9220 11092 9276
rect 11092 9220 11096 9276
rect 11032 9216 11096 9220
rect 11112 9276 11176 9280
rect 11112 9220 11116 9276
rect 11116 9220 11172 9276
rect 11172 9220 11176 9276
rect 11112 9216 11176 9220
rect 11192 9276 11256 9280
rect 11192 9220 11196 9276
rect 11196 9220 11252 9276
rect 11252 9220 11256 9276
rect 11192 9216 11256 9220
rect 20952 9276 21016 9280
rect 20952 9220 20956 9276
rect 20956 9220 21012 9276
rect 21012 9220 21016 9276
rect 20952 9216 21016 9220
rect 21032 9276 21096 9280
rect 21032 9220 21036 9276
rect 21036 9220 21092 9276
rect 21092 9220 21096 9276
rect 21032 9216 21096 9220
rect 21112 9276 21176 9280
rect 21112 9220 21116 9276
rect 21116 9220 21172 9276
rect 21172 9220 21176 9276
rect 21112 9216 21176 9220
rect 21192 9276 21256 9280
rect 21192 9220 21196 9276
rect 21196 9220 21252 9276
rect 21252 9220 21256 9276
rect 21192 9216 21256 9220
rect 5952 8732 6016 8736
rect 5952 8676 5956 8732
rect 5956 8676 6012 8732
rect 6012 8676 6016 8732
rect 5952 8672 6016 8676
rect 6032 8732 6096 8736
rect 6032 8676 6036 8732
rect 6036 8676 6092 8732
rect 6092 8676 6096 8732
rect 6032 8672 6096 8676
rect 6112 8732 6176 8736
rect 6112 8676 6116 8732
rect 6116 8676 6172 8732
rect 6172 8676 6176 8732
rect 6112 8672 6176 8676
rect 6192 8732 6256 8736
rect 6192 8676 6196 8732
rect 6196 8676 6252 8732
rect 6252 8676 6256 8732
rect 6192 8672 6256 8676
rect 15952 8732 16016 8736
rect 15952 8676 15956 8732
rect 15956 8676 16012 8732
rect 16012 8676 16016 8732
rect 15952 8672 16016 8676
rect 16032 8732 16096 8736
rect 16032 8676 16036 8732
rect 16036 8676 16092 8732
rect 16092 8676 16096 8732
rect 16032 8672 16096 8676
rect 16112 8732 16176 8736
rect 16112 8676 16116 8732
rect 16116 8676 16172 8732
rect 16172 8676 16176 8732
rect 16112 8672 16176 8676
rect 16192 8732 16256 8736
rect 16192 8676 16196 8732
rect 16196 8676 16252 8732
rect 16252 8676 16256 8732
rect 16192 8672 16256 8676
rect 25952 8732 26016 8736
rect 25952 8676 25956 8732
rect 25956 8676 26012 8732
rect 26012 8676 26016 8732
rect 25952 8672 26016 8676
rect 26032 8732 26096 8736
rect 26032 8676 26036 8732
rect 26036 8676 26092 8732
rect 26092 8676 26096 8732
rect 26032 8672 26096 8676
rect 26112 8732 26176 8736
rect 26112 8676 26116 8732
rect 26116 8676 26172 8732
rect 26172 8676 26176 8732
rect 26112 8672 26176 8676
rect 26192 8732 26256 8736
rect 26192 8676 26196 8732
rect 26196 8676 26252 8732
rect 26252 8676 26256 8732
rect 26192 8672 26256 8676
rect 25268 8196 25332 8260
rect 10952 8188 11016 8192
rect 10952 8132 10956 8188
rect 10956 8132 11012 8188
rect 11012 8132 11016 8188
rect 10952 8128 11016 8132
rect 11032 8188 11096 8192
rect 11032 8132 11036 8188
rect 11036 8132 11092 8188
rect 11092 8132 11096 8188
rect 11032 8128 11096 8132
rect 11112 8188 11176 8192
rect 11112 8132 11116 8188
rect 11116 8132 11172 8188
rect 11172 8132 11176 8188
rect 11112 8128 11176 8132
rect 11192 8188 11256 8192
rect 11192 8132 11196 8188
rect 11196 8132 11252 8188
rect 11252 8132 11256 8188
rect 11192 8128 11256 8132
rect 20952 8188 21016 8192
rect 20952 8132 20956 8188
rect 20956 8132 21012 8188
rect 21012 8132 21016 8188
rect 20952 8128 21016 8132
rect 21032 8188 21096 8192
rect 21032 8132 21036 8188
rect 21036 8132 21092 8188
rect 21092 8132 21096 8188
rect 21032 8128 21096 8132
rect 21112 8188 21176 8192
rect 21112 8132 21116 8188
rect 21116 8132 21172 8188
rect 21172 8132 21176 8188
rect 21112 8128 21176 8132
rect 21192 8188 21256 8192
rect 21192 8132 21196 8188
rect 21196 8132 21252 8188
rect 21252 8132 21256 8188
rect 21192 8128 21256 8132
rect 15332 7788 15396 7852
rect 5952 7644 6016 7648
rect 5952 7588 5956 7644
rect 5956 7588 6012 7644
rect 6012 7588 6016 7644
rect 5952 7584 6016 7588
rect 6032 7644 6096 7648
rect 6032 7588 6036 7644
rect 6036 7588 6092 7644
rect 6092 7588 6096 7644
rect 6032 7584 6096 7588
rect 6112 7644 6176 7648
rect 6112 7588 6116 7644
rect 6116 7588 6172 7644
rect 6172 7588 6176 7644
rect 6112 7584 6176 7588
rect 6192 7644 6256 7648
rect 6192 7588 6196 7644
rect 6196 7588 6252 7644
rect 6252 7588 6256 7644
rect 6192 7584 6256 7588
rect 15952 7644 16016 7648
rect 15952 7588 15956 7644
rect 15956 7588 16012 7644
rect 16012 7588 16016 7644
rect 15952 7584 16016 7588
rect 16032 7644 16096 7648
rect 16032 7588 16036 7644
rect 16036 7588 16092 7644
rect 16092 7588 16096 7644
rect 16032 7584 16096 7588
rect 16112 7644 16176 7648
rect 16112 7588 16116 7644
rect 16116 7588 16172 7644
rect 16172 7588 16176 7644
rect 16112 7584 16176 7588
rect 16192 7644 16256 7648
rect 16192 7588 16196 7644
rect 16196 7588 16252 7644
rect 16252 7588 16256 7644
rect 16192 7584 16256 7588
rect 25952 7644 26016 7648
rect 25952 7588 25956 7644
rect 25956 7588 26012 7644
rect 26012 7588 26016 7644
rect 25952 7584 26016 7588
rect 26032 7644 26096 7648
rect 26032 7588 26036 7644
rect 26036 7588 26092 7644
rect 26092 7588 26096 7644
rect 26032 7584 26096 7588
rect 26112 7644 26176 7648
rect 26112 7588 26116 7644
rect 26116 7588 26172 7644
rect 26172 7588 26176 7644
rect 26112 7584 26176 7588
rect 26192 7644 26256 7648
rect 26192 7588 26196 7644
rect 26196 7588 26252 7644
rect 26252 7588 26256 7644
rect 26192 7584 26256 7588
rect 10952 7100 11016 7104
rect 10952 7044 10956 7100
rect 10956 7044 11012 7100
rect 11012 7044 11016 7100
rect 10952 7040 11016 7044
rect 11032 7100 11096 7104
rect 11032 7044 11036 7100
rect 11036 7044 11092 7100
rect 11092 7044 11096 7100
rect 11032 7040 11096 7044
rect 11112 7100 11176 7104
rect 11112 7044 11116 7100
rect 11116 7044 11172 7100
rect 11172 7044 11176 7100
rect 11112 7040 11176 7044
rect 11192 7100 11256 7104
rect 11192 7044 11196 7100
rect 11196 7044 11252 7100
rect 11252 7044 11256 7100
rect 11192 7040 11256 7044
rect 20952 7100 21016 7104
rect 20952 7044 20956 7100
rect 20956 7044 21012 7100
rect 21012 7044 21016 7100
rect 20952 7040 21016 7044
rect 21032 7100 21096 7104
rect 21032 7044 21036 7100
rect 21036 7044 21092 7100
rect 21092 7044 21096 7100
rect 21032 7040 21096 7044
rect 21112 7100 21176 7104
rect 21112 7044 21116 7100
rect 21116 7044 21172 7100
rect 21172 7044 21176 7100
rect 21112 7040 21176 7044
rect 21192 7100 21256 7104
rect 21192 7044 21196 7100
rect 21196 7044 21252 7100
rect 21252 7044 21256 7100
rect 21192 7040 21256 7044
rect 5952 6556 6016 6560
rect 5952 6500 5956 6556
rect 5956 6500 6012 6556
rect 6012 6500 6016 6556
rect 5952 6496 6016 6500
rect 6032 6556 6096 6560
rect 6032 6500 6036 6556
rect 6036 6500 6092 6556
rect 6092 6500 6096 6556
rect 6032 6496 6096 6500
rect 6112 6556 6176 6560
rect 6112 6500 6116 6556
rect 6116 6500 6172 6556
rect 6172 6500 6176 6556
rect 6112 6496 6176 6500
rect 6192 6556 6256 6560
rect 6192 6500 6196 6556
rect 6196 6500 6252 6556
rect 6252 6500 6256 6556
rect 6192 6496 6256 6500
rect 15952 6556 16016 6560
rect 15952 6500 15956 6556
rect 15956 6500 16012 6556
rect 16012 6500 16016 6556
rect 15952 6496 16016 6500
rect 16032 6556 16096 6560
rect 16032 6500 16036 6556
rect 16036 6500 16092 6556
rect 16092 6500 16096 6556
rect 16032 6496 16096 6500
rect 16112 6556 16176 6560
rect 16112 6500 16116 6556
rect 16116 6500 16172 6556
rect 16172 6500 16176 6556
rect 16112 6496 16176 6500
rect 16192 6556 16256 6560
rect 16192 6500 16196 6556
rect 16196 6500 16252 6556
rect 16252 6500 16256 6556
rect 16192 6496 16256 6500
rect 25952 6556 26016 6560
rect 25952 6500 25956 6556
rect 25956 6500 26012 6556
rect 26012 6500 26016 6556
rect 25952 6496 26016 6500
rect 26032 6556 26096 6560
rect 26032 6500 26036 6556
rect 26036 6500 26092 6556
rect 26092 6500 26096 6556
rect 26032 6496 26096 6500
rect 26112 6556 26176 6560
rect 26112 6500 26116 6556
rect 26116 6500 26172 6556
rect 26172 6500 26176 6556
rect 26112 6496 26176 6500
rect 26192 6556 26256 6560
rect 26192 6500 26196 6556
rect 26196 6500 26252 6556
rect 26252 6500 26256 6556
rect 26192 6496 26256 6500
rect 10952 6012 11016 6016
rect 10952 5956 10956 6012
rect 10956 5956 11012 6012
rect 11012 5956 11016 6012
rect 10952 5952 11016 5956
rect 11032 6012 11096 6016
rect 11032 5956 11036 6012
rect 11036 5956 11092 6012
rect 11092 5956 11096 6012
rect 11032 5952 11096 5956
rect 11112 6012 11176 6016
rect 11112 5956 11116 6012
rect 11116 5956 11172 6012
rect 11172 5956 11176 6012
rect 11112 5952 11176 5956
rect 11192 6012 11256 6016
rect 11192 5956 11196 6012
rect 11196 5956 11252 6012
rect 11252 5956 11256 6012
rect 11192 5952 11256 5956
rect 20952 6012 21016 6016
rect 20952 5956 20956 6012
rect 20956 5956 21012 6012
rect 21012 5956 21016 6012
rect 20952 5952 21016 5956
rect 21032 6012 21096 6016
rect 21032 5956 21036 6012
rect 21036 5956 21092 6012
rect 21092 5956 21096 6012
rect 21032 5952 21096 5956
rect 21112 6012 21176 6016
rect 21112 5956 21116 6012
rect 21116 5956 21172 6012
rect 21172 5956 21176 6012
rect 21112 5952 21176 5956
rect 21192 6012 21256 6016
rect 21192 5956 21196 6012
rect 21196 5956 21252 6012
rect 21252 5956 21256 6012
rect 21192 5952 21256 5956
rect 11836 5476 11900 5540
rect 5952 5468 6016 5472
rect 5952 5412 5956 5468
rect 5956 5412 6012 5468
rect 6012 5412 6016 5468
rect 5952 5408 6016 5412
rect 6032 5468 6096 5472
rect 6032 5412 6036 5468
rect 6036 5412 6092 5468
rect 6092 5412 6096 5468
rect 6032 5408 6096 5412
rect 6112 5468 6176 5472
rect 6112 5412 6116 5468
rect 6116 5412 6172 5468
rect 6172 5412 6176 5468
rect 6112 5408 6176 5412
rect 6192 5468 6256 5472
rect 6192 5412 6196 5468
rect 6196 5412 6252 5468
rect 6252 5412 6256 5468
rect 6192 5408 6256 5412
rect 15952 5468 16016 5472
rect 15952 5412 15956 5468
rect 15956 5412 16012 5468
rect 16012 5412 16016 5468
rect 15952 5408 16016 5412
rect 16032 5468 16096 5472
rect 16032 5412 16036 5468
rect 16036 5412 16092 5468
rect 16092 5412 16096 5468
rect 16032 5408 16096 5412
rect 16112 5468 16176 5472
rect 16112 5412 16116 5468
rect 16116 5412 16172 5468
rect 16172 5412 16176 5468
rect 16112 5408 16176 5412
rect 16192 5468 16256 5472
rect 16192 5412 16196 5468
rect 16196 5412 16252 5468
rect 16252 5412 16256 5468
rect 16192 5408 16256 5412
rect 25952 5468 26016 5472
rect 25952 5412 25956 5468
rect 25956 5412 26012 5468
rect 26012 5412 26016 5468
rect 25952 5408 26016 5412
rect 26032 5468 26096 5472
rect 26032 5412 26036 5468
rect 26036 5412 26092 5468
rect 26092 5412 26096 5468
rect 26032 5408 26096 5412
rect 26112 5468 26176 5472
rect 26112 5412 26116 5468
rect 26116 5412 26172 5468
rect 26172 5412 26176 5468
rect 26112 5408 26176 5412
rect 26192 5468 26256 5472
rect 26192 5412 26196 5468
rect 26196 5412 26252 5468
rect 26252 5412 26256 5468
rect 26192 5408 26256 5412
rect 10952 4924 11016 4928
rect 10952 4868 10956 4924
rect 10956 4868 11012 4924
rect 11012 4868 11016 4924
rect 10952 4864 11016 4868
rect 11032 4924 11096 4928
rect 11032 4868 11036 4924
rect 11036 4868 11092 4924
rect 11092 4868 11096 4924
rect 11032 4864 11096 4868
rect 11112 4924 11176 4928
rect 11112 4868 11116 4924
rect 11116 4868 11172 4924
rect 11172 4868 11176 4924
rect 11112 4864 11176 4868
rect 11192 4924 11256 4928
rect 11192 4868 11196 4924
rect 11196 4868 11252 4924
rect 11252 4868 11256 4924
rect 11192 4864 11256 4868
rect 20952 4924 21016 4928
rect 20952 4868 20956 4924
rect 20956 4868 21012 4924
rect 21012 4868 21016 4924
rect 20952 4864 21016 4868
rect 21032 4924 21096 4928
rect 21032 4868 21036 4924
rect 21036 4868 21092 4924
rect 21092 4868 21096 4924
rect 21032 4864 21096 4868
rect 21112 4924 21176 4928
rect 21112 4868 21116 4924
rect 21116 4868 21172 4924
rect 21172 4868 21176 4924
rect 21112 4864 21176 4868
rect 21192 4924 21256 4928
rect 21192 4868 21196 4924
rect 21196 4868 21252 4924
rect 21252 4868 21256 4924
rect 21192 4864 21256 4868
rect 5952 4380 6016 4384
rect 5952 4324 5956 4380
rect 5956 4324 6012 4380
rect 6012 4324 6016 4380
rect 5952 4320 6016 4324
rect 6032 4380 6096 4384
rect 6032 4324 6036 4380
rect 6036 4324 6092 4380
rect 6092 4324 6096 4380
rect 6032 4320 6096 4324
rect 6112 4380 6176 4384
rect 6112 4324 6116 4380
rect 6116 4324 6172 4380
rect 6172 4324 6176 4380
rect 6112 4320 6176 4324
rect 6192 4380 6256 4384
rect 6192 4324 6196 4380
rect 6196 4324 6252 4380
rect 6252 4324 6256 4380
rect 6192 4320 6256 4324
rect 15952 4380 16016 4384
rect 15952 4324 15956 4380
rect 15956 4324 16012 4380
rect 16012 4324 16016 4380
rect 15952 4320 16016 4324
rect 16032 4380 16096 4384
rect 16032 4324 16036 4380
rect 16036 4324 16092 4380
rect 16092 4324 16096 4380
rect 16032 4320 16096 4324
rect 16112 4380 16176 4384
rect 16112 4324 16116 4380
rect 16116 4324 16172 4380
rect 16172 4324 16176 4380
rect 16112 4320 16176 4324
rect 16192 4380 16256 4384
rect 16192 4324 16196 4380
rect 16196 4324 16252 4380
rect 16252 4324 16256 4380
rect 16192 4320 16256 4324
rect 25952 4380 26016 4384
rect 25952 4324 25956 4380
rect 25956 4324 26012 4380
rect 26012 4324 26016 4380
rect 25952 4320 26016 4324
rect 26032 4380 26096 4384
rect 26032 4324 26036 4380
rect 26036 4324 26092 4380
rect 26092 4324 26096 4380
rect 26032 4320 26096 4324
rect 26112 4380 26176 4384
rect 26112 4324 26116 4380
rect 26116 4324 26172 4380
rect 26172 4324 26176 4380
rect 26112 4320 26176 4324
rect 26192 4380 26256 4384
rect 26192 4324 26196 4380
rect 26196 4324 26252 4380
rect 26252 4324 26256 4380
rect 26192 4320 26256 4324
rect 16436 3980 16500 4044
rect 10952 3836 11016 3840
rect 10952 3780 10956 3836
rect 10956 3780 11012 3836
rect 11012 3780 11016 3836
rect 10952 3776 11016 3780
rect 11032 3836 11096 3840
rect 11032 3780 11036 3836
rect 11036 3780 11092 3836
rect 11092 3780 11096 3836
rect 11032 3776 11096 3780
rect 11112 3836 11176 3840
rect 11112 3780 11116 3836
rect 11116 3780 11172 3836
rect 11172 3780 11176 3836
rect 11112 3776 11176 3780
rect 11192 3836 11256 3840
rect 11192 3780 11196 3836
rect 11196 3780 11252 3836
rect 11252 3780 11256 3836
rect 11192 3776 11256 3780
rect 20952 3836 21016 3840
rect 20952 3780 20956 3836
rect 20956 3780 21012 3836
rect 21012 3780 21016 3836
rect 20952 3776 21016 3780
rect 21032 3836 21096 3840
rect 21032 3780 21036 3836
rect 21036 3780 21092 3836
rect 21092 3780 21096 3836
rect 21032 3776 21096 3780
rect 21112 3836 21176 3840
rect 21112 3780 21116 3836
rect 21116 3780 21172 3836
rect 21172 3780 21176 3836
rect 21112 3776 21176 3780
rect 21192 3836 21256 3840
rect 21192 3780 21196 3836
rect 21196 3780 21252 3836
rect 21252 3780 21256 3836
rect 21192 3776 21256 3780
rect 21404 3708 21468 3772
rect 15148 3572 15212 3636
rect 5952 3292 6016 3296
rect 5952 3236 5956 3292
rect 5956 3236 6012 3292
rect 6012 3236 6016 3292
rect 5952 3232 6016 3236
rect 6032 3292 6096 3296
rect 6032 3236 6036 3292
rect 6036 3236 6092 3292
rect 6092 3236 6096 3292
rect 6032 3232 6096 3236
rect 6112 3292 6176 3296
rect 6112 3236 6116 3292
rect 6116 3236 6172 3292
rect 6172 3236 6176 3292
rect 6112 3232 6176 3236
rect 6192 3292 6256 3296
rect 6192 3236 6196 3292
rect 6196 3236 6252 3292
rect 6252 3236 6256 3292
rect 6192 3232 6256 3236
rect 15952 3292 16016 3296
rect 15952 3236 15956 3292
rect 15956 3236 16012 3292
rect 16012 3236 16016 3292
rect 15952 3232 16016 3236
rect 16032 3292 16096 3296
rect 16032 3236 16036 3292
rect 16036 3236 16092 3292
rect 16092 3236 16096 3292
rect 16032 3232 16096 3236
rect 16112 3292 16176 3296
rect 16112 3236 16116 3292
rect 16116 3236 16172 3292
rect 16172 3236 16176 3292
rect 16112 3232 16176 3236
rect 16192 3292 16256 3296
rect 16192 3236 16196 3292
rect 16196 3236 16252 3292
rect 16252 3236 16256 3292
rect 16192 3232 16256 3236
rect 25952 3292 26016 3296
rect 25952 3236 25956 3292
rect 25956 3236 26012 3292
rect 26012 3236 26016 3292
rect 25952 3232 26016 3236
rect 26032 3292 26096 3296
rect 26032 3236 26036 3292
rect 26036 3236 26092 3292
rect 26092 3236 26096 3292
rect 26032 3232 26096 3236
rect 26112 3292 26176 3296
rect 26112 3236 26116 3292
rect 26116 3236 26172 3292
rect 26172 3236 26176 3292
rect 26112 3232 26176 3236
rect 26192 3292 26256 3296
rect 26192 3236 26196 3292
rect 26196 3236 26252 3292
rect 26252 3236 26256 3292
rect 26192 3232 26256 3236
rect 15516 3164 15580 3228
rect 10952 2748 11016 2752
rect 10952 2692 10956 2748
rect 10956 2692 11012 2748
rect 11012 2692 11016 2748
rect 10952 2688 11016 2692
rect 11032 2748 11096 2752
rect 11032 2692 11036 2748
rect 11036 2692 11092 2748
rect 11092 2692 11096 2748
rect 11032 2688 11096 2692
rect 11112 2748 11176 2752
rect 11112 2692 11116 2748
rect 11116 2692 11172 2748
rect 11172 2692 11176 2748
rect 11112 2688 11176 2692
rect 11192 2748 11256 2752
rect 11192 2692 11196 2748
rect 11196 2692 11252 2748
rect 11252 2692 11256 2748
rect 11192 2688 11256 2692
rect 20952 2748 21016 2752
rect 20952 2692 20956 2748
rect 20956 2692 21012 2748
rect 21012 2692 21016 2748
rect 20952 2688 21016 2692
rect 21032 2748 21096 2752
rect 21032 2692 21036 2748
rect 21036 2692 21092 2748
rect 21092 2692 21096 2748
rect 21032 2688 21096 2692
rect 21112 2748 21176 2752
rect 21112 2692 21116 2748
rect 21116 2692 21172 2748
rect 21172 2692 21176 2748
rect 21112 2688 21176 2692
rect 21192 2748 21256 2752
rect 21192 2692 21196 2748
rect 21196 2692 21252 2748
rect 21252 2692 21256 2748
rect 21192 2688 21256 2692
rect 24900 2620 24964 2684
rect 5952 2204 6016 2208
rect 5952 2148 5956 2204
rect 5956 2148 6012 2204
rect 6012 2148 6016 2204
rect 5952 2144 6016 2148
rect 6032 2204 6096 2208
rect 6032 2148 6036 2204
rect 6036 2148 6092 2204
rect 6092 2148 6096 2204
rect 6032 2144 6096 2148
rect 6112 2204 6176 2208
rect 6112 2148 6116 2204
rect 6116 2148 6172 2204
rect 6172 2148 6176 2204
rect 6112 2144 6176 2148
rect 6192 2204 6256 2208
rect 6192 2148 6196 2204
rect 6196 2148 6252 2204
rect 6252 2148 6256 2204
rect 6192 2144 6256 2148
rect 15952 2204 16016 2208
rect 15952 2148 15956 2204
rect 15956 2148 16012 2204
rect 16012 2148 16016 2204
rect 15952 2144 16016 2148
rect 16032 2204 16096 2208
rect 16032 2148 16036 2204
rect 16036 2148 16092 2204
rect 16092 2148 16096 2204
rect 16032 2144 16096 2148
rect 16112 2204 16176 2208
rect 16112 2148 16116 2204
rect 16116 2148 16172 2204
rect 16172 2148 16176 2204
rect 16112 2144 16176 2148
rect 16192 2204 16256 2208
rect 16192 2148 16196 2204
rect 16196 2148 16252 2204
rect 16252 2148 16256 2204
rect 16192 2144 16256 2148
rect 25952 2204 26016 2208
rect 25952 2148 25956 2204
rect 25956 2148 26012 2204
rect 26012 2148 26016 2204
rect 25952 2144 26016 2148
rect 26032 2204 26096 2208
rect 26032 2148 26036 2204
rect 26036 2148 26092 2204
rect 26092 2148 26096 2204
rect 26032 2144 26096 2148
rect 26112 2204 26176 2208
rect 26112 2148 26116 2204
rect 26116 2148 26172 2204
rect 26172 2148 26176 2204
rect 26112 2144 26176 2148
rect 26192 2204 26256 2208
rect 26192 2148 26196 2204
rect 26196 2148 26252 2204
rect 26252 2148 26256 2204
rect 26192 2144 26256 2148
<< metal4 >>
rect 5944 77280 6264 77840
rect 5944 77216 5952 77280
rect 6016 77216 6032 77280
rect 6096 77216 6112 77280
rect 6176 77216 6192 77280
rect 6256 77216 6264 77280
rect 5944 76192 6264 77216
rect 5944 76128 5952 76192
rect 6016 76128 6032 76192
rect 6096 76128 6112 76192
rect 6176 76128 6192 76192
rect 6256 76128 6264 76192
rect 5944 75104 6264 76128
rect 5944 75040 5952 75104
rect 6016 75040 6032 75104
rect 6096 75040 6112 75104
rect 6176 75040 6192 75104
rect 6256 75040 6264 75104
rect 5944 74016 6264 75040
rect 10944 77824 11264 77840
rect 10944 77760 10952 77824
rect 11016 77760 11032 77824
rect 11096 77760 11112 77824
rect 11176 77760 11192 77824
rect 11256 77760 11264 77824
rect 10944 76736 11264 77760
rect 10944 76672 10952 76736
rect 11016 76672 11032 76736
rect 11096 76672 11112 76736
rect 11176 76672 11192 76736
rect 11256 76672 11264 76736
rect 10944 75648 11264 76672
rect 15944 77280 16264 77840
rect 20944 77824 21264 77840
rect 20944 77760 20952 77824
rect 21016 77760 21032 77824
rect 21096 77760 21112 77824
rect 21176 77760 21192 77824
rect 21256 77760 21264 77824
rect 20667 77484 20733 77485
rect 20667 77420 20668 77484
rect 20732 77420 20733 77484
rect 20667 77419 20733 77420
rect 15944 77216 15952 77280
rect 16016 77216 16032 77280
rect 16096 77216 16112 77280
rect 16176 77216 16192 77280
rect 16256 77216 16264 77280
rect 15944 76192 16264 77216
rect 15944 76128 15952 76192
rect 16016 76128 16032 76192
rect 16096 76128 16112 76192
rect 16176 76128 16192 76192
rect 16256 76128 16264 76192
rect 11835 75716 11901 75717
rect 11835 75652 11836 75716
rect 11900 75652 11901 75716
rect 11835 75651 11901 75652
rect 10944 75584 10952 75648
rect 11016 75584 11032 75648
rect 11096 75584 11112 75648
rect 11176 75584 11192 75648
rect 11256 75584 11264 75648
rect 9995 74764 10061 74765
rect 9995 74700 9996 74764
rect 10060 74700 10061 74764
rect 9995 74699 10061 74700
rect 5944 73952 5952 74016
rect 6016 73952 6032 74016
rect 6096 73952 6112 74016
rect 6176 73952 6192 74016
rect 6256 73952 6264 74016
rect 5944 72928 6264 73952
rect 5944 72864 5952 72928
rect 6016 72864 6032 72928
rect 6096 72864 6112 72928
rect 6176 72864 6192 72928
rect 6256 72864 6264 72928
rect 5944 71840 6264 72864
rect 5944 71776 5952 71840
rect 6016 71776 6032 71840
rect 6096 71776 6112 71840
rect 6176 71776 6192 71840
rect 6256 71776 6264 71840
rect 5944 70752 6264 71776
rect 5944 70688 5952 70752
rect 6016 70688 6032 70752
rect 6096 70688 6112 70752
rect 6176 70688 6192 70752
rect 6256 70688 6264 70752
rect 5944 69664 6264 70688
rect 5944 69600 5952 69664
rect 6016 69600 6032 69664
rect 6096 69600 6112 69664
rect 6176 69600 6192 69664
rect 6256 69600 6264 69664
rect 5944 68912 6264 69600
rect 5944 68676 5986 68912
rect 6222 68676 6264 68912
rect 5944 68576 6264 68676
rect 5944 68512 5952 68576
rect 6016 68512 6032 68576
rect 6096 68512 6112 68576
rect 6176 68512 6192 68576
rect 6256 68512 6264 68576
rect 5944 67488 6264 68512
rect 5944 67424 5952 67488
rect 6016 67424 6032 67488
rect 6096 67424 6112 67488
rect 6176 67424 6192 67488
rect 6256 67424 6264 67488
rect 5944 66400 6264 67424
rect 5944 66336 5952 66400
rect 6016 66336 6032 66400
rect 6096 66336 6112 66400
rect 6176 66336 6192 66400
rect 6256 66336 6264 66400
rect 5944 65312 6264 66336
rect 5944 65248 5952 65312
rect 6016 65248 6032 65312
rect 6096 65248 6112 65312
rect 6176 65248 6192 65312
rect 6256 65248 6264 65312
rect 5944 64224 6264 65248
rect 5944 64160 5952 64224
rect 6016 64160 6032 64224
rect 6096 64160 6112 64224
rect 6176 64160 6192 64224
rect 6256 64160 6264 64224
rect 5944 63136 6264 64160
rect 5944 63072 5952 63136
rect 6016 63072 6032 63136
rect 6096 63072 6112 63136
rect 6176 63072 6192 63136
rect 6256 63072 6264 63136
rect 5944 62048 6264 63072
rect 5944 61984 5952 62048
rect 6016 61984 6032 62048
rect 6096 61984 6112 62048
rect 6176 61984 6192 62048
rect 6256 61984 6264 62048
rect 5944 60960 6264 61984
rect 5944 60896 5952 60960
rect 6016 60896 6032 60960
rect 6096 60896 6112 60960
rect 6176 60896 6192 60960
rect 6256 60896 6264 60960
rect 5944 59872 6264 60896
rect 5944 59808 5952 59872
rect 6016 59808 6032 59872
rect 6096 59808 6112 59872
rect 6176 59808 6192 59872
rect 6256 59808 6264 59872
rect 5944 58784 6264 59808
rect 5944 58720 5952 58784
rect 6016 58720 6032 58784
rect 6096 58720 6112 58784
rect 6176 58720 6192 58784
rect 6256 58720 6264 58784
rect 5944 57696 6264 58720
rect 5944 57632 5952 57696
rect 6016 57632 6032 57696
rect 6096 57632 6112 57696
rect 6176 57632 6192 57696
rect 6256 57632 6264 57696
rect 5944 56608 6264 57632
rect 5944 56544 5952 56608
rect 6016 56544 6032 56608
rect 6096 56544 6112 56608
rect 6176 56544 6192 56608
rect 6256 56544 6264 56608
rect 5944 55520 6264 56544
rect 5944 55456 5952 55520
rect 6016 55456 6032 55520
rect 6096 55456 6112 55520
rect 6176 55456 6192 55520
rect 6256 55456 6264 55520
rect 5944 54432 6264 55456
rect 5944 54368 5952 54432
rect 6016 54368 6032 54432
rect 6096 54368 6112 54432
rect 6176 54368 6192 54432
rect 6256 54368 6264 54432
rect 5944 53344 6264 54368
rect 5944 53280 5952 53344
rect 6016 53280 6032 53344
rect 6096 53280 6112 53344
rect 6176 53280 6192 53344
rect 6256 53280 6264 53344
rect 5944 52256 6264 53280
rect 5944 52192 5952 52256
rect 6016 52192 6032 52256
rect 6096 52192 6112 52256
rect 6176 52192 6192 52256
rect 6256 52192 6264 52256
rect 5944 51168 6264 52192
rect 5944 51104 5952 51168
rect 6016 51104 6032 51168
rect 6096 51104 6112 51168
rect 6176 51104 6192 51168
rect 6256 51104 6264 51168
rect 5944 50080 6264 51104
rect 5944 50016 5952 50080
rect 6016 50016 6032 50080
rect 6096 50016 6112 50080
rect 6176 50016 6192 50080
rect 6256 50016 6264 50080
rect 5944 48992 6264 50016
rect 5944 48928 5952 48992
rect 6016 48928 6032 48992
rect 6096 48928 6112 48992
rect 6176 48928 6192 48992
rect 6256 48928 6264 48992
rect 5944 47904 6264 48928
rect 5944 47840 5952 47904
rect 6016 47840 6032 47904
rect 6096 47840 6112 47904
rect 6176 47840 6192 47904
rect 6256 47840 6264 47904
rect 5944 46816 6264 47840
rect 9627 47020 9693 47021
rect 9627 46956 9628 47020
rect 9692 46956 9693 47020
rect 9627 46955 9693 46956
rect 5944 46752 5952 46816
rect 6016 46752 6032 46816
rect 6096 46752 6112 46816
rect 6176 46752 6192 46816
rect 6256 46752 6264 46816
rect 5944 45728 6264 46752
rect 5944 45664 5952 45728
rect 6016 45664 6032 45728
rect 6096 45664 6112 45728
rect 6176 45664 6192 45728
rect 6256 45664 6264 45728
rect 5944 44640 6264 45664
rect 5944 44576 5952 44640
rect 6016 44576 6032 44640
rect 6096 44576 6112 44640
rect 6176 44576 6192 44640
rect 6256 44576 6264 44640
rect 5944 43552 6264 44576
rect 5944 43488 5952 43552
rect 6016 43488 6032 43552
rect 6096 43488 6112 43552
rect 6176 43488 6192 43552
rect 6256 43488 6264 43552
rect 5944 42464 6264 43488
rect 5944 42400 5952 42464
rect 6016 42400 6032 42464
rect 6096 42400 6112 42464
rect 6176 42400 6192 42464
rect 6256 42400 6264 42464
rect 5944 42246 6264 42400
rect 5944 42010 5986 42246
rect 6222 42010 6264 42246
rect 5944 41376 6264 42010
rect 5944 41312 5952 41376
rect 6016 41312 6032 41376
rect 6096 41312 6112 41376
rect 6176 41312 6192 41376
rect 6256 41312 6264 41376
rect 5944 40288 6264 41312
rect 5944 40224 5952 40288
rect 6016 40224 6032 40288
rect 6096 40224 6112 40288
rect 6176 40224 6192 40288
rect 6256 40224 6264 40288
rect 5944 39200 6264 40224
rect 5944 39136 5952 39200
rect 6016 39136 6032 39200
rect 6096 39136 6112 39200
rect 6176 39136 6192 39200
rect 6256 39136 6264 39200
rect 3374 32061 3434 37622
rect 3742 35733 3802 36942
rect 3739 35732 3805 35733
rect 3739 35668 3740 35732
rect 3804 35668 3805 35732
rect 3739 35667 3805 35668
rect 5582 33013 5642 38982
rect 5944 38112 6264 39136
rect 5944 38048 5952 38112
rect 6016 38048 6032 38112
rect 6096 38048 6112 38112
rect 6176 38048 6192 38112
rect 6256 38048 6264 38112
rect 5944 37024 6264 38048
rect 9630 37365 9690 46955
rect 9811 37636 9877 37637
rect 9811 37572 9812 37636
rect 9876 37572 9877 37636
rect 9811 37571 9877 37572
rect 9627 37364 9693 37365
rect 9627 37300 9628 37364
rect 9692 37300 9693 37364
rect 9627 37299 9693 37300
rect 5944 36960 5952 37024
rect 6016 36960 6032 37024
rect 6096 36960 6112 37024
rect 6176 36960 6192 37024
rect 6256 36960 6264 37024
rect 5944 35936 6264 36960
rect 9627 36004 9693 36005
rect 9627 35940 9628 36004
rect 9692 35940 9693 36004
rect 9627 35939 9693 35940
rect 5944 35872 5952 35936
rect 6016 35872 6032 35936
rect 6096 35872 6112 35936
rect 6176 35872 6192 35936
rect 6256 35872 6264 35936
rect 5944 34848 6264 35872
rect 9259 35732 9325 35733
rect 9259 35668 9260 35732
rect 9324 35668 9325 35732
rect 9259 35667 9325 35668
rect 7419 35324 7485 35325
rect 7419 35260 7420 35324
rect 7484 35260 7485 35324
rect 7419 35259 7485 35260
rect 5944 34784 5952 34848
rect 6016 34784 6032 34848
rect 6096 34784 6112 34848
rect 6176 34784 6192 34848
rect 6256 34784 6264 34848
rect 5944 33760 6264 34784
rect 6683 33964 6749 33965
rect 6683 33900 6684 33964
rect 6748 33900 6749 33964
rect 6683 33899 6749 33900
rect 5944 33696 5952 33760
rect 6016 33696 6032 33760
rect 6096 33696 6112 33760
rect 6176 33696 6192 33760
rect 6256 33696 6264 33760
rect 5579 33012 5645 33013
rect 5579 32948 5580 33012
rect 5644 32948 5645 33012
rect 5579 32947 5645 32948
rect 5944 32672 6264 33696
rect 6686 33098 6746 33899
rect 5944 32608 5952 32672
rect 6016 32608 6032 32672
rect 6096 32608 6112 32672
rect 6176 32608 6192 32672
rect 6256 32608 6264 32672
rect 3371 32060 3437 32061
rect 3371 31996 3372 32060
rect 3436 31996 3437 32060
rect 3371 31995 3437 31996
rect 5944 31584 6264 32608
rect 5944 31520 5952 31584
rect 6016 31520 6032 31584
rect 6096 31520 6112 31584
rect 6176 31520 6192 31584
rect 6256 31520 6264 31584
rect 5944 30496 6264 31520
rect 5944 30432 5952 30496
rect 6016 30432 6032 30496
rect 6096 30432 6112 30496
rect 6176 30432 6192 30496
rect 6256 30432 6264 30496
rect 5944 29408 6264 30432
rect 5944 29344 5952 29408
rect 6016 29344 6032 29408
rect 6096 29344 6112 29408
rect 6176 29344 6192 29408
rect 6256 29344 6264 29408
rect 5944 28320 6264 29344
rect 7422 28933 7482 35259
rect 9075 34916 9141 34917
rect 9075 34852 9076 34916
rect 9140 34852 9141 34916
rect 9075 34851 9141 34852
rect 9078 32061 9138 34851
rect 9262 32741 9322 35667
rect 9443 34372 9509 34373
rect 9443 34308 9444 34372
rect 9508 34308 9509 34372
rect 9443 34307 9509 34308
rect 9259 32740 9325 32741
rect 9259 32676 9260 32740
rect 9324 32676 9325 32740
rect 9259 32675 9325 32676
rect 9075 32060 9141 32061
rect 9075 31996 9076 32060
rect 9140 31996 9141 32060
rect 9075 31995 9141 31996
rect 9262 29477 9322 32675
rect 9446 31653 9506 34307
rect 9443 31652 9509 31653
rect 9443 31588 9444 31652
rect 9508 31588 9509 31652
rect 9443 31587 9509 31588
rect 9259 29476 9325 29477
rect 9259 29412 9260 29476
rect 9324 29412 9325 29476
rect 9259 29411 9325 29412
rect 7419 28932 7485 28933
rect 7419 28868 7420 28932
rect 7484 28868 7485 28932
rect 7419 28867 7485 28868
rect 5944 28256 5952 28320
rect 6016 28256 6032 28320
rect 6096 28256 6112 28320
rect 6176 28256 6192 28320
rect 6256 28256 6264 28320
rect 5944 27232 6264 28256
rect 9630 27845 9690 35939
rect 9814 34781 9874 37571
rect 9811 34780 9877 34781
rect 9811 34716 9812 34780
rect 9876 34716 9877 34780
rect 9811 34715 9877 34716
rect 9811 33964 9877 33965
rect 9811 33900 9812 33964
rect 9876 33900 9877 33964
rect 9811 33899 9877 33900
rect 9627 27844 9693 27845
rect 9627 27780 9628 27844
rect 9692 27780 9693 27844
rect 9627 27779 9693 27780
rect 5944 27168 5952 27232
rect 6016 27168 6032 27232
rect 6096 27168 6112 27232
rect 6176 27168 6192 27232
rect 6256 27168 6264 27232
rect 5944 26144 6264 27168
rect 9814 26893 9874 33899
rect 9811 26892 9877 26893
rect 9811 26828 9812 26892
rect 9876 26828 9877 26892
rect 9811 26827 9877 26828
rect 5944 26080 5952 26144
rect 6016 26080 6032 26144
rect 6096 26080 6112 26144
rect 6176 26080 6192 26144
rect 6256 26080 6264 26144
rect 5944 25056 6264 26080
rect 9627 25668 9693 25669
rect 9627 25604 9628 25668
rect 9692 25604 9693 25668
rect 9627 25603 9693 25604
rect 5944 24992 5952 25056
rect 6016 24992 6032 25056
rect 6096 24992 6112 25056
rect 6176 24992 6192 25056
rect 6256 24992 6264 25056
rect 5944 23968 6264 24992
rect 5944 23904 5952 23968
rect 6016 23904 6032 23968
rect 6096 23904 6112 23968
rect 6176 23904 6192 23968
rect 6256 23904 6264 23968
rect 5944 22880 6264 23904
rect 5944 22816 5952 22880
rect 6016 22816 6032 22880
rect 6096 22816 6112 22880
rect 6176 22816 6192 22880
rect 6256 22816 6264 22880
rect 5944 21792 6264 22816
rect 5944 21728 5952 21792
rect 6016 21728 6032 21792
rect 6096 21728 6112 21792
rect 6176 21728 6192 21792
rect 6256 21728 6264 21792
rect 5944 20704 6264 21728
rect 5944 20640 5952 20704
rect 6016 20640 6032 20704
rect 6096 20640 6112 20704
rect 6176 20640 6192 20704
rect 6256 20640 6264 20704
rect 5944 19616 6264 20640
rect 9630 20229 9690 25603
rect 9998 21997 10058 74699
rect 10944 74560 11264 75584
rect 10944 74496 10952 74560
rect 11016 74496 11032 74560
rect 11096 74496 11112 74560
rect 11176 74496 11192 74560
rect 11256 74496 11264 74560
rect 10944 73472 11264 74496
rect 10944 73408 10952 73472
rect 11016 73408 11032 73472
rect 11096 73408 11112 73472
rect 11176 73408 11192 73472
rect 11256 73408 11264 73472
rect 10944 72384 11264 73408
rect 10944 72320 10952 72384
rect 11016 72320 11032 72384
rect 11096 72320 11112 72384
rect 11176 72320 11192 72384
rect 11256 72320 11264 72384
rect 10944 71296 11264 72320
rect 10944 71232 10952 71296
rect 11016 71232 11032 71296
rect 11096 71232 11112 71296
rect 11176 71232 11192 71296
rect 11256 71232 11264 71296
rect 10944 70208 11264 71232
rect 10944 70144 10952 70208
rect 11016 70144 11032 70208
rect 11096 70144 11112 70208
rect 11176 70144 11192 70208
rect 11256 70144 11264 70208
rect 10944 69120 11264 70144
rect 10944 69056 10952 69120
rect 11016 69056 11032 69120
rect 11096 69056 11112 69120
rect 11176 69056 11192 69120
rect 11256 69056 11264 69120
rect 10944 68032 11264 69056
rect 10944 67968 10952 68032
rect 11016 67968 11032 68032
rect 11096 67968 11112 68032
rect 11176 67968 11192 68032
rect 11256 67968 11264 68032
rect 10944 66944 11264 67968
rect 10944 66880 10952 66944
rect 11016 66880 11032 66944
rect 11096 66880 11112 66944
rect 11176 66880 11192 66944
rect 11256 66880 11264 66944
rect 10944 65856 11264 66880
rect 10944 65792 10952 65856
rect 11016 65792 11032 65856
rect 11096 65792 11112 65856
rect 11176 65792 11192 65856
rect 11256 65792 11264 65856
rect 10944 64768 11264 65792
rect 10944 64704 10952 64768
rect 11016 64704 11032 64768
rect 11096 64704 11112 64768
rect 11176 64704 11192 64768
rect 11256 64704 11264 64768
rect 10944 63680 11264 64704
rect 10944 63616 10952 63680
rect 11016 63616 11032 63680
rect 11096 63616 11112 63680
rect 11176 63616 11192 63680
rect 11256 63616 11264 63680
rect 10944 62592 11264 63616
rect 10944 62528 10952 62592
rect 11016 62528 11032 62592
rect 11096 62528 11112 62592
rect 11176 62528 11192 62592
rect 11256 62528 11264 62592
rect 10944 61504 11264 62528
rect 10944 61440 10952 61504
rect 11016 61440 11032 61504
rect 11096 61440 11112 61504
rect 11176 61440 11192 61504
rect 11256 61440 11264 61504
rect 10944 60416 11264 61440
rect 10944 60352 10952 60416
rect 11016 60352 11032 60416
rect 11096 60352 11112 60416
rect 11176 60352 11192 60416
rect 11256 60352 11264 60416
rect 10944 59328 11264 60352
rect 10944 59264 10952 59328
rect 11016 59264 11032 59328
rect 11096 59264 11112 59328
rect 11176 59264 11192 59328
rect 11256 59264 11264 59328
rect 10944 58240 11264 59264
rect 10944 58176 10952 58240
rect 11016 58176 11032 58240
rect 11096 58176 11112 58240
rect 11176 58176 11192 58240
rect 11256 58176 11264 58240
rect 10944 57152 11264 58176
rect 11467 58036 11533 58037
rect 11467 57972 11468 58036
rect 11532 57972 11533 58036
rect 11467 57971 11533 57972
rect 10944 57088 10952 57152
rect 11016 57088 11032 57152
rect 11096 57088 11112 57152
rect 11176 57088 11192 57152
rect 11256 57088 11264 57152
rect 10944 56064 11264 57088
rect 10944 56000 10952 56064
rect 11016 56000 11032 56064
rect 11096 56000 11112 56064
rect 11176 56000 11192 56064
rect 11256 56000 11264 56064
rect 10944 55579 11264 56000
rect 10944 55343 10986 55579
rect 11222 55343 11264 55579
rect 10944 54976 11264 55343
rect 10944 54912 10952 54976
rect 11016 54912 11032 54976
rect 11096 54912 11112 54976
rect 11176 54912 11192 54976
rect 11256 54912 11264 54976
rect 10944 53888 11264 54912
rect 10944 53824 10952 53888
rect 11016 53824 11032 53888
rect 11096 53824 11112 53888
rect 11176 53824 11192 53888
rect 11256 53824 11264 53888
rect 10944 52800 11264 53824
rect 10944 52736 10952 52800
rect 11016 52736 11032 52800
rect 11096 52736 11112 52800
rect 11176 52736 11192 52800
rect 11256 52736 11264 52800
rect 10944 51712 11264 52736
rect 10944 51648 10952 51712
rect 11016 51648 11032 51712
rect 11096 51648 11112 51712
rect 11176 51648 11192 51712
rect 11256 51648 11264 51712
rect 10944 50624 11264 51648
rect 10944 50560 10952 50624
rect 11016 50560 11032 50624
rect 11096 50560 11112 50624
rect 11176 50560 11192 50624
rect 11256 50560 11264 50624
rect 10944 49536 11264 50560
rect 10944 49472 10952 49536
rect 11016 49472 11032 49536
rect 11096 49472 11112 49536
rect 11176 49472 11192 49536
rect 11256 49472 11264 49536
rect 10944 48448 11264 49472
rect 10944 48384 10952 48448
rect 11016 48384 11032 48448
rect 11096 48384 11112 48448
rect 11176 48384 11192 48448
rect 11256 48384 11264 48448
rect 10944 47360 11264 48384
rect 10944 47296 10952 47360
rect 11016 47296 11032 47360
rect 11096 47296 11112 47360
rect 11176 47296 11192 47360
rect 11256 47296 11264 47360
rect 10944 46272 11264 47296
rect 10944 46208 10952 46272
rect 11016 46208 11032 46272
rect 11096 46208 11112 46272
rect 11176 46208 11192 46272
rect 11256 46208 11264 46272
rect 10944 45184 11264 46208
rect 10944 45120 10952 45184
rect 11016 45120 11032 45184
rect 11096 45120 11112 45184
rect 11176 45120 11192 45184
rect 11256 45120 11264 45184
rect 10944 44096 11264 45120
rect 10944 44032 10952 44096
rect 11016 44032 11032 44096
rect 11096 44032 11112 44096
rect 11176 44032 11192 44096
rect 11256 44032 11264 44096
rect 10944 43008 11264 44032
rect 10944 42944 10952 43008
rect 11016 42944 11032 43008
rect 11096 42944 11112 43008
rect 11176 42944 11192 43008
rect 11256 42944 11264 43008
rect 10944 41920 11264 42944
rect 10944 41856 10952 41920
rect 11016 41856 11032 41920
rect 11096 41856 11112 41920
rect 11176 41856 11192 41920
rect 11256 41856 11264 41920
rect 10944 40832 11264 41856
rect 10944 40768 10952 40832
rect 11016 40768 11032 40832
rect 11096 40768 11112 40832
rect 11176 40768 11192 40832
rect 11256 40768 11264 40832
rect 10944 39744 11264 40768
rect 10944 39680 10952 39744
rect 11016 39680 11032 39744
rect 11096 39680 11112 39744
rect 11176 39680 11192 39744
rect 11256 39680 11264 39744
rect 10944 38656 11264 39680
rect 10944 38592 10952 38656
rect 11016 38592 11032 38656
rect 11096 38592 11112 38656
rect 11176 38592 11192 38656
rect 11256 38592 11264 38656
rect 10363 37772 10429 37773
rect 10363 37708 10364 37772
rect 10428 37708 10429 37772
rect 10363 37707 10429 37708
rect 10179 37364 10245 37365
rect 10179 37300 10180 37364
rect 10244 37300 10245 37364
rect 10179 37299 10245 37300
rect 10182 25941 10242 37299
rect 10366 34373 10426 37707
rect 10944 37568 11264 38592
rect 10944 37504 10952 37568
rect 11016 37504 11032 37568
rect 11096 37504 11112 37568
rect 11176 37504 11192 37568
rect 11256 37504 11264 37568
rect 10547 37092 10613 37093
rect 10547 37028 10548 37092
rect 10612 37028 10613 37092
rect 10547 37027 10613 37028
rect 10550 34781 10610 37027
rect 10944 36480 11264 37504
rect 10944 36416 10952 36480
rect 11016 36416 11032 36480
rect 11096 36416 11112 36480
rect 11176 36416 11192 36480
rect 11256 36416 11264 36480
rect 10731 35460 10797 35461
rect 10731 35396 10732 35460
rect 10796 35396 10797 35460
rect 10731 35395 10797 35396
rect 10547 34780 10613 34781
rect 10547 34716 10548 34780
rect 10612 34716 10613 34780
rect 10547 34715 10613 34716
rect 10363 34372 10429 34373
rect 10363 34308 10364 34372
rect 10428 34308 10429 34372
rect 10363 34307 10429 34308
rect 10363 32196 10429 32197
rect 10363 32132 10364 32196
rect 10428 32132 10429 32196
rect 10363 32131 10429 32132
rect 10366 30021 10426 32131
rect 10550 32061 10610 34715
rect 10547 32060 10613 32061
rect 10547 31996 10548 32060
rect 10612 31996 10613 32060
rect 10547 31995 10613 31996
rect 10734 31786 10794 35395
rect 10550 31726 10794 31786
rect 10944 35392 11264 36416
rect 10944 35328 10952 35392
rect 11016 35328 11032 35392
rect 11096 35328 11112 35392
rect 11176 35328 11192 35392
rect 11256 35328 11264 35392
rect 10944 34304 11264 35328
rect 10944 34240 10952 34304
rect 11016 34240 11032 34304
rect 11096 34240 11112 34304
rect 11176 34240 11192 34304
rect 11256 34240 11264 34304
rect 10944 33216 11264 34240
rect 10944 33152 10952 33216
rect 11016 33152 11032 33216
rect 11096 33152 11112 33216
rect 11176 33152 11192 33216
rect 11256 33152 11264 33216
rect 10944 32128 11264 33152
rect 11470 33013 11530 57971
rect 11651 36004 11717 36005
rect 11651 35940 11652 36004
rect 11716 35940 11717 36004
rect 11651 35939 11717 35940
rect 11654 33829 11714 35939
rect 11651 33828 11717 33829
rect 11651 33764 11652 33828
rect 11716 33764 11717 33828
rect 11651 33763 11717 33764
rect 11654 33421 11714 33763
rect 11651 33420 11717 33421
rect 11651 33356 11652 33420
rect 11716 33356 11717 33420
rect 11651 33355 11717 33356
rect 11467 33012 11533 33013
rect 11467 32948 11468 33012
rect 11532 32948 11533 33012
rect 11467 32947 11533 32948
rect 10944 32064 10952 32128
rect 11016 32064 11032 32128
rect 11096 32064 11112 32128
rect 11176 32064 11192 32128
rect 11256 32064 11264 32128
rect 10363 30020 10429 30021
rect 10363 29956 10364 30020
rect 10428 29956 10429 30020
rect 10363 29955 10429 29956
rect 10550 29749 10610 31726
rect 10731 31652 10797 31653
rect 10731 31588 10732 31652
rect 10796 31588 10797 31652
rect 10731 31587 10797 31588
rect 10547 29748 10613 29749
rect 10547 29684 10548 29748
rect 10612 29684 10613 29748
rect 10547 29683 10613 29684
rect 10547 28116 10613 28117
rect 10547 28052 10548 28116
rect 10612 28052 10613 28116
rect 10547 28051 10613 28052
rect 10179 25940 10245 25941
rect 10179 25876 10180 25940
rect 10244 25876 10245 25940
rect 10179 25875 10245 25876
rect 10550 25669 10610 28051
rect 10734 26349 10794 31587
rect 10944 31040 11264 32064
rect 11467 32060 11533 32061
rect 11467 31996 11468 32060
rect 11532 31996 11533 32060
rect 11467 31995 11533 31996
rect 11470 31381 11530 31995
rect 11654 31653 11714 33355
rect 11651 31652 11717 31653
rect 11651 31588 11652 31652
rect 11716 31588 11717 31652
rect 11651 31587 11717 31588
rect 11651 31516 11717 31517
rect 11651 31452 11652 31516
rect 11716 31452 11717 31516
rect 11651 31451 11717 31452
rect 11467 31380 11533 31381
rect 11467 31316 11468 31380
rect 11532 31316 11533 31380
rect 11467 31315 11533 31316
rect 10944 30976 10952 31040
rect 11016 30976 11032 31040
rect 11096 30976 11112 31040
rect 11176 30976 11192 31040
rect 11256 30976 11264 31040
rect 10944 29952 11264 30976
rect 11654 30157 11714 31451
rect 11651 30156 11717 30157
rect 11651 30092 11652 30156
rect 11716 30092 11717 30156
rect 11651 30091 11717 30092
rect 10944 29888 10952 29952
rect 11016 29888 11032 29952
rect 11096 29888 11112 29952
rect 11176 29888 11192 29952
rect 11256 29888 11264 29952
rect 10944 28912 11264 29888
rect 11651 29748 11717 29749
rect 11651 29684 11652 29748
rect 11716 29684 11717 29748
rect 11651 29683 11717 29684
rect 10944 28864 10986 28912
rect 11222 28864 11264 28912
rect 10944 28800 10952 28864
rect 11256 28800 11264 28864
rect 10944 28676 10986 28800
rect 11222 28676 11264 28800
rect 10944 27776 11264 28676
rect 10944 27712 10952 27776
rect 11016 27712 11032 27776
rect 11096 27712 11112 27776
rect 11176 27712 11192 27776
rect 11256 27712 11264 27776
rect 10944 26688 11264 27712
rect 10944 26624 10952 26688
rect 11016 26624 11032 26688
rect 11096 26624 11112 26688
rect 11176 26624 11192 26688
rect 11256 26624 11264 26688
rect 10731 26348 10797 26349
rect 10731 26284 10732 26348
rect 10796 26284 10797 26348
rect 10731 26283 10797 26284
rect 10547 25668 10613 25669
rect 10547 25604 10548 25668
rect 10612 25604 10613 25668
rect 10547 25603 10613 25604
rect 10731 25668 10797 25669
rect 10731 25604 10732 25668
rect 10796 25604 10797 25668
rect 10731 25603 10797 25604
rect 9995 21996 10061 21997
rect 9995 21932 9996 21996
rect 10060 21932 10061 21996
rect 9995 21931 10061 21932
rect 10734 21725 10794 25603
rect 10944 25600 11264 26624
rect 11467 26348 11533 26349
rect 11467 26284 11468 26348
rect 11532 26284 11533 26348
rect 11467 26283 11533 26284
rect 10944 25536 10952 25600
rect 11016 25536 11032 25600
rect 11096 25536 11112 25600
rect 11176 25536 11192 25600
rect 11256 25536 11264 25600
rect 10944 24512 11264 25536
rect 11470 24581 11530 26283
rect 11467 24580 11533 24581
rect 11467 24516 11468 24580
rect 11532 24516 11533 24580
rect 11467 24515 11533 24516
rect 10944 24448 10952 24512
rect 11016 24448 11032 24512
rect 11096 24448 11112 24512
rect 11176 24448 11192 24512
rect 11256 24448 11264 24512
rect 10944 23424 11264 24448
rect 10944 23360 10952 23424
rect 11016 23360 11032 23424
rect 11096 23360 11112 23424
rect 11176 23360 11192 23424
rect 11256 23360 11264 23424
rect 10944 22336 11264 23360
rect 11467 22676 11533 22677
rect 11467 22612 11468 22676
rect 11532 22612 11533 22676
rect 11467 22611 11533 22612
rect 10944 22272 10952 22336
rect 11016 22272 11032 22336
rect 11096 22272 11112 22336
rect 11176 22272 11192 22336
rect 11256 22272 11264 22336
rect 10731 21724 10797 21725
rect 10731 21660 10732 21724
rect 10796 21660 10797 21724
rect 10731 21659 10797 21660
rect 10944 21248 11264 22272
rect 10944 21184 10952 21248
rect 11016 21184 11032 21248
rect 11096 21184 11112 21248
rect 11176 21184 11192 21248
rect 11256 21184 11264 21248
rect 9627 20228 9693 20229
rect 9627 20164 9628 20228
rect 9692 20164 9693 20228
rect 9627 20163 9693 20164
rect 5944 19552 5952 19616
rect 6016 19552 6032 19616
rect 6096 19552 6112 19616
rect 6176 19552 6192 19616
rect 6256 19552 6264 19616
rect 5944 18528 6264 19552
rect 10944 20160 11264 21184
rect 10944 20096 10952 20160
rect 11016 20096 11032 20160
rect 11096 20096 11112 20160
rect 11176 20096 11192 20160
rect 11256 20096 11264 20160
rect 9075 19276 9141 19277
rect 9075 19212 9076 19276
rect 9140 19212 9141 19276
rect 9075 19211 9141 19212
rect 5944 18464 5952 18528
rect 6016 18464 6032 18528
rect 6096 18464 6112 18528
rect 6176 18464 6192 18528
rect 6256 18464 6264 18528
rect 5944 17440 6264 18464
rect 5944 17376 5952 17440
rect 6016 17376 6032 17440
rect 6096 17376 6112 17440
rect 6176 17376 6192 17440
rect 6256 17376 6264 17440
rect 5944 16352 6264 17376
rect 5944 16288 5952 16352
rect 6016 16288 6032 16352
rect 6096 16288 6112 16352
rect 6176 16288 6192 16352
rect 6256 16288 6264 16352
rect 5944 15579 6264 16288
rect 5944 15343 5986 15579
rect 6222 15343 6264 15579
rect 5944 15264 6264 15343
rect 5944 15200 5952 15264
rect 6016 15200 6032 15264
rect 6096 15200 6112 15264
rect 6176 15200 6192 15264
rect 6256 15200 6264 15264
rect 5944 14176 6264 15200
rect 5944 14112 5952 14176
rect 6016 14112 6032 14176
rect 6096 14112 6112 14176
rect 6176 14112 6192 14176
rect 6256 14112 6264 14176
rect 5944 13088 6264 14112
rect 5944 13024 5952 13088
rect 6016 13024 6032 13088
rect 6096 13024 6112 13088
rect 6176 13024 6192 13088
rect 6256 13024 6264 13088
rect 5944 12000 6264 13024
rect 9078 12069 9138 19211
rect 10944 19072 11264 20096
rect 11470 19821 11530 22611
rect 11654 22405 11714 29683
rect 11651 22404 11717 22405
rect 11651 22340 11652 22404
rect 11716 22340 11717 22404
rect 11651 22339 11717 22340
rect 11467 19820 11533 19821
rect 11467 19756 11468 19820
rect 11532 19756 11533 19820
rect 11467 19755 11533 19756
rect 10944 19008 10952 19072
rect 11016 19008 11032 19072
rect 11096 19008 11112 19072
rect 11176 19008 11192 19072
rect 11256 19008 11264 19072
rect 10547 18868 10613 18869
rect 10547 18804 10548 18868
rect 10612 18804 10613 18868
rect 10547 18803 10613 18804
rect 9075 12068 9141 12069
rect 9075 12004 9076 12068
rect 9140 12004 9141 12068
rect 9075 12003 9141 12004
rect 5944 11936 5952 12000
rect 6016 11936 6032 12000
rect 6096 11936 6112 12000
rect 6176 11936 6192 12000
rect 6256 11936 6264 12000
rect 5944 10912 6264 11936
rect 5944 10848 5952 10912
rect 6016 10848 6032 10912
rect 6096 10848 6112 10912
rect 6176 10848 6192 10912
rect 6256 10848 6264 10912
rect 5944 9824 6264 10848
rect 10550 10845 10610 18803
rect 10944 17984 11264 19008
rect 10944 17920 10952 17984
rect 11016 17920 11032 17984
rect 11096 17920 11112 17984
rect 11176 17920 11192 17984
rect 11256 17920 11264 17984
rect 10944 16896 11264 17920
rect 10944 16832 10952 16896
rect 11016 16832 11032 16896
rect 11096 16832 11112 16896
rect 11176 16832 11192 16896
rect 11256 16832 11264 16896
rect 10944 15808 11264 16832
rect 10944 15744 10952 15808
rect 11016 15744 11032 15808
rect 11096 15744 11112 15808
rect 11176 15744 11192 15808
rect 11256 15744 11264 15808
rect 10944 14720 11264 15744
rect 10944 14656 10952 14720
rect 11016 14656 11032 14720
rect 11096 14656 11112 14720
rect 11176 14656 11192 14720
rect 11256 14656 11264 14720
rect 10944 13632 11264 14656
rect 10944 13568 10952 13632
rect 11016 13568 11032 13632
rect 11096 13568 11112 13632
rect 11176 13568 11192 13632
rect 11256 13568 11264 13632
rect 10944 12544 11264 13568
rect 10944 12480 10952 12544
rect 11016 12480 11032 12544
rect 11096 12480 11112 12544
rect 11176 12480 11192 12544
rect 11256 12480 11264 12544
rect 10944 11456 11264 12480
rect 10944 11392 10952 11456
rect 11016 11392 11032 11456
rect 11096 11392 11112 11456
rect 11176 11392 11192 11456
rect 11256 11392 11264 11456
rect 10547 10844 10613 10845
rect 10547 10780 10548 10844
rect 10612 10780 10613 10844
rect 10547 10779 10613 10780
rect 5944 9760 5952 9824
rect 6016 9760 6032 9824
rect 6096 9760 6112 9824
rect 6176 9760 6192 9824
rect 6256 9760 6264 9824
rect 5944 8736 6264 9760
rect 5944 8672 5952 8736
rect 6016 8672 6032 8736
rect 6096 8672 6112 8736
rect 6176 8672 6192 8736
rect 6256 8672 6264 8736
rect 5944 7648 6264 8672
rect 5944 7584 5952 7648
rect 6016 7584 6032 7648
rect 6096 7584 6112 7648
rect 6176 7584 6192 7648
rect 6256 7584 6264 7648
rect 5944 6560 6264 7584
rect 5944 6496 5952 6560
rect 6016 6496 6032 6560
rect 6096 6496 6112 6560
rect 6176 6496 6192 6560
rect 6256 6496 6264 6560
rect 5944 5472 6264 6496
rect 5944 5408 5952 5472
rect 6016 5408 6032 5472
rect 6096 5408 6112 5472
rect 6176 5408 6192 5472
rect 6256 5408 6264 5472
rect 5944 4384 6264 5408
rect 5944 4320 5952 4384
rect 6016 4320 6032 4384
rect 6096 4320 6112 4384
rect 6176 4320 6192 4384
rect 6256 4320 6264 4384
rect 5944 3296 6264 4320
rect 5944 3232 5952 3296
rect 6016 3232 6032 3296
rect 6096 3232 6112 3296
rect 6176 3232 6192 3296
rect 6256 3232 6264 3296
rect 5944 2208 6264 3232
rect 5944 2144 5952 2208
rect 6016 2144 6032 2208
rect 6096 2144 6112 2208
rect 6176 2144 6192 2208
rect 6256 2144 6264 2208
rect 5944 2128 6264 2144
rect 10944 10368 11264 11392
rect 10944 10304 10952 10368
rect 11016 10304 11032 10368
rect 11096 10304 11112 10368
rect 11176 10304 11192 10368
rect 11256 10304 11264 10368
rect 10944 9280 11264 10304
rect 10944 9216 10952 9280
rect 11016 9216 11032 9280
rect 11096 9216 11112 9280
rect 11176 9216 11192 9280
rect 11256 9216 11264 9280
rect 10944 8192 11264 9216
rect 10944 8128 10952 8192
rect 11016 8128 11032 8192
rect 11096 8128 11112 8192
rect 11176 8128 11192 8192
rect 11256 8128 11264 8192
rect 10944 7104 11264 8128
rect 10944 7040 10952 7104
rect 11016 7040 11032 7104
rect 11096 7040 11112 7104
rect 11176 7040 11192 7104
rect 11256 7040 11264 7104
rect 10944 6016 11264 7040
rect 10944 5952 10952 6016
rect 11016 5952 11032 6016
rect 11096 5952 11112 6016
rect 11176 5952 11192 6016
rect 11256 5952 11264 6016
rect 10944 4928 11264 5952
rect 11838 5541 11898 75651
rect 15944 75104 16264 76128
rect 15944 75040 15952 75104
rect 16016 75040 16032 75104
rect 16096 75040 16112 75104
rect 16176 75040 16192 75104
rect 16256 75040 16264 75104
rect 15944 74016 16264 75040
rect 15944 73952 15952 74016
rect 16016 73952 16032 74016
rect 16096 73952 16112 74016
rect 16176 73952 16192 74016
rect 16256 73952 16264 74016
rect 15944 72928 16264 73952
rect 15944 72864 15952 72928
rect 16016 72864 16032 72928
rect 16096 72864 16112 72928
rect 16176 72864 16192 72928
rect 16256 72864 16264 72928
rect 15944 71840 16264 72864
rect 15944 71776 15952 71840
rect 16016 71776 16032 71840
rect 16096 71776 16112 71840
rect 16176 71776 16192 71840
rect 16256 71776 16264 71840
rect 15944 70752 16264 71776
rect 15944 70688 15952 70752
rect 16016 70688 16032 70752
rect 16096 70688 16112 70752
rect 16176 70688 16192 70752
rect 16256 70688 16264 70752
rect 15944 69664 16264 70688
rect 15944 69600 15952 69664
rect 16016 69600 16032 69664
rect 16096 69600 16112 69664
rect 16176 69600 16192 69664
rect 16256 69600 16264 69664
rect 15944 68912 16264 69600
rect 17171 69324 17237 69325
rect 17171 69260 17172 69324
rect 17236 69260 17237 69324
rect 17171 69259 17237 69260
rect 15944 68676 15986 68912
rect 16222 68676 16264 68912
rect 15944 68576 16264 68676
rect 15944 68512 15952 68576
rect 16016 68512 16032 68576
rect 16096 68512 16112 68576
rect 16176 68512 16192 68576
rect 16256 68512 16264 68576
rect 15944 67488 16264 68512
rect 15944 67424 15952 67488
rect 16016 67424 16032 67488
rect 16096 67424 16112 67488
rect 16176 67424 16192 67488
rect 16256 67424 16264 67488
rect 15944 66400 16264 67424
rect 15944 66336 15952 66400
rect 16016 66336 16032 66400
rect 16096 66336 16112 66400
rect 16176 66336 16192 66400
rect 16256 66336 16264 66400
rect 15944 65312 16264 66336
rect 15944 65248 15952 65312
rect 16016 65248 16032 65312
rect 16096 65248 16112 65312
rect 16176 65248 16192 65312
rect 16256 65248 16264 65312
rect 15944 64224 16264 65248
rect 15944 64160 15952 64224
rect 16016 64160 16032 64224
rect 16096 64160 16112 64224
rect 16176 64160 16192 64224
rect 16256 64160 16264 64224
rect 15944 63136 16264 64160
rect 15944 63072 15952 63136
rect 16016 63072 16032 63136
rect 16096 63072 16112 63136
rect 16176 63072 16192 63136
rect 16256 63072 16264 63136
rect 15944 62048 16264 63072
rect 15944 61984 15952 62048
rect 16016 61984 16032 62048
rect 16096 61984 16112 62048
rect 16176 61984 16192 62048
rect 16256 61984 16264 62048
rect 15944 60960 16264 61984
rect 15944 60896 15952 60960
rect 16016 60896 16032 60960
rect 16096 60896 16112 60960
rect 16176 60896 16192 60960
rect 16256 60896 16264 60960
rect 15944 59872 16264 60896
rect 15944 59808 15952 59872
rect 16016 59808 16032 59872
rect 16096 59808 16112 59872
rect 16176 59808 16192 59872
rect 16256 59808 16264 59872
rect 15944 58784 16264 59808
rect 15944 58720 15952 58784
rect 16016 58720 16032 58784
rect 16096 58720 16112 58784
rect 16176 58720 16192 58784
rect 16256 58720 16264 58784
rect 15944 57696 16264 58720
rect 15944 57632 15952 57696
rect 16016 57632 16032 57696
rect 16096 57632 16112 57696
rect 16176 57632 16192 57696
rect 16256 57632 16264 57696
rect 15699 56676 15765 56677
rect 15699 56612 15700 56676
rect 15764 56612 15765 56676
rect 15699 56611 15765 56612
rect 12019 52596 12085 52597
rect 12019 52532 12020 52596
rect 12084 52532 12085 52596
rect 12019 52531 12085 52532
rect 12022 12749 12082 52531
rect 15515 51372 15581 51373
rect 15515 51308 15516 51372
rect 15580 51308 15581 51372
rect 15515 51307 15581 51308
rect 15518 50829 15578 51307
rect 15515 50828 15581 50829
rect 15515 50764 15516 50828
rect 15580 50764 15581 50828
rect 15515 50763 15581 50764
rect 15331 48380 15397 48381
rect 15331 48316 15332 48380
rect 15396 48316 15397 48380
rect 15331 48315 15397 48316
rect 13675 42940 13741 42941
rect 13675 42876 13676 42940
rect 13740 42876 13741 42940
rect 13675 42875 13741 42876
rect 12387 42124 12453 42125
rect 12387 42060 12388 42124
rect 12452 42060 12453 42124
rect 12387 42059 12453 42060
rect 12203 35868 12269 35869
rect 12203 35804 12204 35868
rect 12268 35804 12269 35868
rect 12203 35803 12269 35804
rect 12206 33965 12266 35803
rect 12203 33964 12269 33965
rect 12203 33900 12204 33964
rect 12268 33900 12269 33964
rect 12203 33899 12269 33900
rect 12203 33284 12269 33285
rect 12203 33220 12204 33284
rect 12268 33220 12269 33284
rect 12203 33219 12269 33220
rect 12206 33013 12266 33219
rect 12203 33012 12269 33013
rect 12203 32948 12204 33012
rect 12268 32948 12269 33012
rect 12203 32947 12269 32948
rect 12206 27029 12266 32947
rect 12390 27709 12450 42059
rect 12939 41852 13005 41853
rect 12939 41788 12940 41852
rect 13004 41788 13005 41852
rect 12939 41787 13005 41788
rect 12755 39676 12821 39677
rect 12755 39612 12756 39676
rect 12820 39612 12821 39676
rect 12755 39611 12821 39612
rect 12571 34372 12637 34373
rect 12571 34308 12572 34372
rect 12636 34308 12637 34372
rect 12571 34307 12637 34308
rect 12574 31653 12634 34307
rect 12758 31925 12818 39611
rect 12942 33149 13002 41787
rect 13491 39812 13557 39813
rect 13491 39748 13492 39812
rect 13556 39748 13557 39812
rect 13491 39747 13557 39748
rect 13307 39676 13373 39677
rect 13307 39612 13308 39676
rect 13372 39612 13373 39676
rect 13307 39611 13373 39612
rect 13310 39405 13370 39611
rect 13307 39404 13373 39405
rect 13307 39340 13308 39404
rect 13372 39340 13373 39404
rect 13307 39339 13373 39340
rect 13123 38452 13189 38453
rect 13123 38388 13124 38452
rect 13188 38388 13189 38452
rect 13123 38387 13189 38388
rect 12939 33148 13005 33149
rect 12939 33084 12940 33148
rect 13004 33084 13005 33148
rect 12939 33083 13005 33084
rect 13126 33010 13186 38387
rect 13307 35188 13373 35189
rect 13307 35124 13308 35188
rect 13372 35124 13373 35188
rect 13307 35123 13373 35124
rect 12942 32950 13186 33010
rect 12755 31924 12821 31925
rect 12755 31860 12756 31924
rect 12820 31860 12821 31924
rect 12755 31859 12821 31860
rect 12755 31788 12821 31789
rect 12755 31724 12756 31788
rect 12820 31724 12821 31788
rect 12755 31723 12821 31724
rect 12571 31652 12637 31653
rect 12571 31588 12572 31652
rect 12636 31588 12637 31652
rect 12571 31587 12637 31588
rect 12758 30970 12818 31723
rect 12574 30910 12818 30970
rect 12387 27708 12453 27709
rect 12387 27644 12388 27708
rect 12452 27644 12453 27708
rect 12387 27643 12453 27644
rect 12574 27165 12634 30910
rect 12942 30429 13002 32950
rect 13310 32330 13370 35123
rect 13126 32270 13370 32330
rect 12755 30428 12821 30429
rect 12755 30364 12756 30428
rect 12820 30364 12821 30428
rect 12755 30363 12821 30364
rect 12939 30428 13005 30429
rect 12939 30364 12940 30428
rect 13004 30364 13005 30428
rect 12939 30363 13005 30364
rect 12758 30290 12818 30363
rect 12758 30230 13002 30290
rect 12942 29885 13002 30230
rect 12939 29884 13005 29885
rect 12939 29820 12940 29884
rect 13004 29820 13005 29884
rect 12939 29819 13005 29820
rect 12755 29340 12821 29341
rect 12755 29276 12756 29340
rect 12820 29276 12821 29340
rect 12755 29275 12821 29276
rect 12571 27164 12637 27165
rect 12571 27100 12572 27164
rect 12636 27100 12637 27164
rect 12571 27099 12637 27100
rect 12203 27028 12269 27029
rect 12203 26964 12204 27028
rect 12268 26964 12269 27028
rect 12203 26963 12269 26964
rect 12206 23629 12266 26963
rect 12387 25396 12453 25397
rect 12387 25332 12388 25396
rect 12452 25332 12453 25396
rect 12387 25331 12453 25332
rect 12203 23628 12269 23629
rect 12203 23564 12204 23628
rect 12268 23564 12269 23628
rect 12203 23563 12269 23564
rect 12203 22268 12269 22269
rect 12203 22204 12204 22268
rect 12268 22204 12269 22268
rect 12203 22203 12269 22204
rect 12206 20365 12266 22203
rect 12203 20364 12269 20365
rect 12203 20300 12204 20364
rect 12268 20300 12269 20364
rect 12203 20299 12269 20300
rect 12390 18325 12450 25331
rect 12387 18324 12453 18325
rect 12387 18260 12388 18324
rect 12452 18260 12453 18324
rect 12387 18259 12453 18260
rect 12758 15061 12818 29275
rect 12942 22269 13002 29819
rect 13126 29341 13186 32270
rect 13307 31924 13373 31925
rect 13307 31860 13308 31924
rect 13372 31860 13373 31924
rect 13307 31859 13373 31860
rect 13310 30701 13370 31859
rect 13307 30700 13373 30701
rect 13307 30636 13308 30700
rect 13372 30636 13373 30700
rect 13307 30635 13373 30636
rect 13307 30020 13373 30021
rect 13307 29956 13308 30020
rect 13372 29956 13373 30020
rect 13307 29955 13373 29956
rect 13123 29340 13189 29341
rect 13123 29276 13124 29340
rect 13188 29276 13189 29340
rect 13123 29275 13189 29276
rect 13310 22541 13370 29955
rect 13307 22540 13373 22541
rect 13307 22476 13308 22540
rect 13372 22476 13373 22540
rect 13307 22475 13373 22476
rect 12939 22268 13005 22269
rect 12939 22204 12940 22268
rect 13004 22204 13005 22268
rect 12939 22203 13005 22204
rect 13494 22133 13554 39747
rect 13491 22132 13557 22133
rect 13491 22068 13492 22132
rect 13556 22068 13557 22132
rect 13491 22067 13557 22068
rect 12755 15060 12821 15061
rect 12755 14996 12756 15060
rect 12820 14996 12821 15060
rect 12755 14995 12821 14996
rect 13678 13565 13738 42875
rect 14595 37636 14661 37637
rect 14595 37572 14596 37636
rect 14660 37572 14661 37636
rect 14595 37571 14661 37572
rect 14043 35460 14109 35461
rect 14043 35396 14044 35460
rect 14108 35396 14109 35460
rect 14043 35395 14109 35396
rect 13859 31924 13925 31925
rect 13859 31860 13860 31924
rect 13924 31860 13925 31924
rect 13859 31859 13925 31860
rect 13862 31381 13922 31859
rect 14046 31789 14106 35395
rect 14598 34509 14658 37571
rect 14595 34508 14661 34509
rect 14595 34444 14596 34508
rect 14660 34444 14661 34508
rect 14595 34443 14661 34444
rect 14227 34100 14293 34101
rect 14227 34036 14228 34100
rect 14292 34036 14293 34100
rect 14227 34035 14293 34036
rect 14043 31788 14109 31789
rect 14043 31724 14044 31788
rect 14108 31724 14109 31788
rect 14043 31723 14109 31724
rect 14043 31652 14109 31653
rect 14043 31588 14044 31652
rect 14108 31588 14109 31652
rect 14043 31587 14109 31588
rect 13859 31380 13925 31381
rect 13859 31316 13860 31380
rect 13924 31316 13925 31380
rect 13859 31315 13925 31316
rect 13859 30156 13925 30157
rect 13859 30092 13860 30156
rect 13924 30092 13925 30156
rect 13859 30091 13925 30092
rect 13862 28661 13922 30091
rect 14046 29749 14106 31587
rect 14230 31381 14290 34035
rect 14595 33284 14661 33285
rect 14595 33220 14596 33284
rect 14660 33220 14661 33284
rect 14595 33219 14661 33220
rect 14411 31788 14477 31789
rect 14411 31724 14412 31788
rect 14476 31724 14477 31788
rect 14411 31723 14477 31724
rect 14227 31380 14293 31381
rect 14227 31316 14228 31380
rect 14292 31316 14293 31380
rect 14227 31315 14293 31316
rect 14043 29748 14109 29749
rect 14043 29684 14044 29748
rect 14108 29684 14109 29748
rect 14043 29683 14109 29684
rect 14227 29612 14293 29613
rect 14227 29548 14228 29612
rect 14292 29548 14293 29612
rect 14227 29547 14293 29548
rect 13859 28660 13925 28661
rect 13859 28596 13860 28660
rect 13924 28596 13925 28660
rect 13859 28595 13925 28596
rect 14230 28389 14290 29547
rect 14227 28388 14293 28389
rect 14227 28324 14228 28388
rect 14292 28324 14293 28388
rect 14227 28323 14293 28324
rect 14414 25397 14474 31723
rect 14411 25396 14477 25397
rect 14411 25332 14412 25396
rect 14476 25332 14477 25396
rect 14411 25331 14477 25332
rect 14598 18189 14658 33219
rect 14782 32741 14842 33542
rect 15147 33420 15213 33421
rect 15147 33356 15148 33420
rect 15212 33356 15213 33420
rect 15147 33355 15213 33356
rect 14779 32740 14845 32741
rect 14779 32676 14780 32740
rect 14844 32676 14845 32740
rect 14779 32675 14845 32676
rect 14963 31108 15029 31109
rect 14963 31044 14964 31108
rect 15028 31044 15029 31108
rect 14963 31043 15029 31044
rect 14779 30972 14845 30973
rect 14779 30908 14780 30972
rect 14844 30908 14845 30972
rect 14779 30907 14845 30908
rect 14782 21997 14842 30907
rect 14966 22949 15026 31043
rect 14963 22948 15029 22949
rect 14963 22884 14964 22948
rect 15028 22884 15029 22948
rect 14963 22883 15029 22884
rect 15150 22810 15210 33355
rect 14966 22750 15210 22810
rect 14779 21996 14845 21997
rect 14779 21932 14780 21996
rect 14844 21932 14845 21996
rect 14779 21931 14845 21932
rect 14966 20501 15026 22750
rect 15147 22676 15213 22677
rect 15147 22612 15148 22676
rect 15212 22612 15213 22676
rect 15147 22611 15213 22612
rect 14963 20500 15029 20501
rect 14963 20436 14964 20500
rect 15028 20436 15029 20500
rect 14963 20435 15029 20436
rect 14595 18188 14661 18189
rect 14595 18124 14596 18188
rect 14660 18124 14661 18188
rect 14595 18123 14661 18124
rect 13675 13564 13741 13565
rect 13675 13500 13676 13564
rect 13740 13500 13741 13564
rect 13675 13499 13741 13500
rect 12019 12748 12085 12749
rect 12019 12684 12020 12748
rect 12084 12684 12085 12748
rect 12019 12683 12085 12684
rect 11835 5540 11901 5541
rect 11835 5476 11836 5540
rect 11900 5476 11901 5540
rect 11835 5475 11901 5476
rect 10944 4864 10952 4928
rect 11016 4864 11032 4928
rect 11096 4864 11112 4928
rect 11176 4864 11192 4928
rect 11256 4864 11264 4928
rect 10944 3840 11264 4864
rect 10944 3776 10952 3840
rect 11016 3776 11032 3840
rect 11096 3776 11112 3840
rect 11176 3776 11192 3840
rect 11256 3776 11264 3840
rect 10944 2752 11264 3776
rect 15150 3637 15210 22611
rect 15334 7853 15394 48315
rect 15515 47020 15581 47021
rect 15515 46956 15516 47020
rect 15580 46956 15581 47020
rect 15515 46955 15581 46956
rect 15331 7852 15397 7853
rect 15331 7788 15332 7852
rect 15396 7788 15397 7852
rect 15331 7787 15397 7788
rect 15147 3636 15213 3637
rect 15147 3572 15148 3636
rect 15212 3572 15213 3636
rect 15147 3571 15213 3572
rect 15518 3229 15578 46955
rect 15702 11389 15762 56611
rect 15944 56608 16264 57632
rect 15944 56544 15952 56608
rect 16016 56544 16032 56608
rect 16096 56544 16112 56608
rect 16176 56544 16192 56608
rect 16256 56544 16264 56608
rect 15944 55520 16264 56544
rect 15944 55456 15952 55520
rect 16016 55456 16032 55520
rect 16096 55456 16112 55520
rect 16176 55456 16192 55520
rect 16256 55456 16264 55520
rect 15944 54432 16264 55456
rect 15944 54368 15952 54432
rect 16016 54368 16032 54432
rect 16096 54368 16112 54432
rect 16176 54368 16192 54432
rect 16256 54368 16264 54432
rect 15944 53344 16264 54368
rect 15944 53280 15952 53344
rect 16016 53280 16032 53344
rect 16096 53280 16112 53344
rect 16176 53280 16192 53344
rect 16256 53280 16264 53344
rect 15944 52256 16264 53280
rect 16435 52596 16501 52597
rect 16435 52532 16436 52596
rect 16500 52532 16501 52596
rect 16435 52531 16501 52532
rect 15944 52192 15952 52256
rect 16016 52192 16032 52256
rect 16096 52192 16112 52256
rect 16176 52192 16192 52256
rect 16256 52192 16264 52256
rect 15944 51168 16264 52192
rect 15944 51104 15952 51168
rect 16016 51104 16032 51168
rect 16096 51104 16112 51168
rect 16176 51104 16192 51168
rect 16256 51104 16264 51168
rect 15944 50080 16264 51104
rect 15944 50016 15952 50080
rect 16016 50016 16032 50080
rect 16096 50016 16112 50080
rect 16176 50016 16192 50080
rect 16256 50016 16264 50080
rect 15944 48992 16264 50016
rect 16438 49605 16498 52531
rect 16435 49604 16501 49605
rect 16435 49540 16436 49604
rect 16500 49540 16501 49604
rect 16435 49539 16501 49540
rect 15944 48928 15952 48992
rect 16016 48928 16032 48992
rect 16096 48928 16112 48992
rect 16176 48928 16192 48992
rect 16256 48928 16264 48992
rect 15944 47904 16264 48928
rect 15944 47840 15952 47904
rect 16016 47840 16032 47904
rect 16096 47840 16112 47904
rect 16176 47840 16192 47904
rect 16256 47840 16264 47904
rect 15944 46816 16264 47840
rect 16435 47020 16501 47021
rect 16435 46956 16436 47020
rect 16500 46956 16501 47020
rect 16435 46955 16501 46956
rect 15944 46752 15952 46816
rect 16016 46752 16032 46816
rect 16096 46752 16112 46816
rect 16176 46752 16192 46816
rect 16256 46752 16264 46816
rect 15944 45728 16264 46752
rect 15944 45664 15952 45728
rect 16016 45664 16032 45728
rect 16096 45664 16112 45728
rect 16176 45664 16192 45728
rect 16256 45664 16264 45728
rect 15944 44640 16264 45664
rect 15944 44576 15952 44640
rect 16016 44576 16032 44640
rect 16096 44576 16112 44640
rect 16176 44576 16192 44640
rect 16256 44576 16264 44640
rect 15944 43552 16264 44576
rect 15944 43488 15952 43552
rect 16016 43488 16032 43552
rect 16096 43488 16112 43552
rect 16176 43488 16192 43552
rect 16256 43488 16264 43552
rect 15944 42464 16264 43488
rect 15944 42400 15952 42464
rect 16016 42400 16032 42464
rect 16096 42400 16112 42464
rect 16176 42400 16192 42464
rect 16256 42400 16264 42464
rect 15944 42246 16264 42400
rect 15944 42010 15986 42246
rect 16222 42010 16264 42246
rect 15944 41376 16264 42010
rect 15944 41312 15952 41376
rect 16016 41312 16032 41376
rect 16096 41312 16112 41376
rect 16176 41312 16192 41376
rect 16256 41312 16264 41376
rect 15944 40288 16264 41312
rect 15944 40224 15952 40288
rect 16016 40224 16032 40288
rect 16096 40224 16112 40288
rect 16176 40224 16192 40288
rect 16256 40224 16264 40288
rect 15944 39200 16264 40224
rect 15944 39136 15952 39200
rect 16016 39136 16032 39200
rect 16096 39136 16112 39200
rect 16176 39136 16192 39200
rect 16256 39136 16264 39200
rect 15944 38112 16264 39136
rect 15944 38048 15952 38112
rect 16016 38048 16032 38112
rect 16096 38048 16112 38112
rect 16176 38048 16192 38112
rect 16256 38048 16264 38112
rect 15944 37024 16264 38048
rect 15944 36960 15952 37024
rect 16016 36960 16032 37024
rect 16096 36960 16112 37024
rect 16176 36960 16192 37024
rect 16256 36960 16264 37024
rect 15944 35936 16264 36960
rect 15944 35872 15952 35936
rect 16016 35872 16032 35936
rect 16096 35872 16112 35936
rect 16176 35872 16192 35936
rect 16256 35872 16264 35936
rect 15944 34848 16264 35872
rect 15944 34784 15952 34848
rect 16016 34784 16032 34848
rect 16096 34784 16112 34848
rect 16176 34784 16192 34848
rect 16256 34784 16264 34848
rect 15944 33760 16264 34784
rect 15944 33696 15952 33760
rect 16016 33696 16032 33760
rect 16096 33696 16112 33760
rect 16176 33696 16192 33760
rect 16256 33696 16264 33760
rect 15944 32672 16264 33696
rect 15944 32608 15952 32672
rect 16016 32608 16032 32672
rect 16096 32608 16112 32672
rect 16176 32608 16192 32672
rect 16256 32608 16264 32672
rect 15944 31584 16264 32608
rect 15944 31520 15952 31584
rect 16016 31520 16032 31584
rect 16096 31520 16112 31584
rect 16176 31520 16192 31584
rect 16256 31520 16264 31584
rect 15944 30496 16264 31520
rect 15944 30432 15952 30496
rect 16016 30432 16032 30496
rect 16096 30432 16112 30496
rect 16176 30432 16192 30496
rect 16256 30432 16264 30496
rect 15944 29408 16264 30432
rect 15944 29344 15952 29408
rect 16016 29344 16032 29408
rect 16096 29344 16112 29408
rect 16176 29344 16192 29408
rect 16256 29344 16264 29408
rect 15944 28320 16264 29344
rect 15944 28256 15952 28320
rect 16016 28256 16032 28320
rect 16096 28256 16112 28320
rect 16176 28256 16192 28320
rect 16256 28256 16264 28320
rect 15944 27232 16264 28256
rect 15944 27168 15952 27232
rect 16016 27168 16032 27232
rect 16096 27168 16112 27232
rect 16176 27168 16192 27232
rect 16256 27168 16264 27232
rect 15944 26144 16264 27168
rect 15944 26080 15952 26144
rect 16016 26080 16032 26144
rect 16096 26080 16112 26144
rect 16176 26080 16192 26144
rect 16256 26080 16264 26144
rect 15944 25056 16264 26080
rect 15944 24992 15952 25056
rect 16016 24992 16032 25056
rect 16096 24992 16112 25056
rect 16176 24992 16192 25056
rect 16256 24992 16264 25056
rect 15944 23968 16264 24992
rect 15944 23904 15952 23968
rect 16016 23904 16032 23968
rect 16096 23904 16112 23968
rect 16176 23904 16192 23968
rect 16256 23904 16264 23968
rect 15944 22880 16264 23904
rect 15944 22816 15952 22880
rect 16016 22816 16032 22880
rect 16096 22816 16112 22880
rect 16176 22816 16192 22880
rect 16256 22816 16264 22880
rect 15944 21792 16264 22816
rect 15944 21728 15952 21792
rect 16016 21728 16032 21792
rect 16096 21728 16112 21792
rect 16176 21728 16192 21792
rect 16256 21728 16264 21792
rect 15944 20704 16264 21728
rect 15944 20640 15952 20704
rect 16016 20640 16032 20704
rect 16096 20640 16112 20704
rect 16176 20640 16192 20704
rect 16256 20640 16264 20704
rect 15944 19616 16264 20640
rect 15944 19552 15952 19616
rect 16016 19552 16032 19616
rect 16096 19552 16112 19616
rect 16176 19552 16192 19616
rect 16256 19552 16264 19616
rect 15944 18528 16264 19552
rect 15944 18464 15952 18528
rect 16016 18464 16032 18528
rect 16096 18464 16112 18528
rect 16176 18464 16192 18528
rect 16256 18464 16264 18528
rect 15944 17440 16264 18464
rect 15944 17376 15952 17440
rect 16016 17376 16032 17440
rect 16096 17376 16112 17440
rect 16176 17376 16192 17440
rect 16256 17376 16264 17440
rect 15944 16352 16264 17376
rect 15944 16288 15952 16352
rect 16016 16288 16032 16352
rect 16096 16288 16112 16352
rect 16176 16288 16192 16352
rect 16256 16288 16264 16352
rect 15944 15579 16264 16288
rect 15944 15343 15986 15579
rect 16222 15343 16264 15579
rect 15944 15264 16264 15343
rect 15944 15200 15952 15264
rect 16016 15200 16032 15264
rect 16096 15200 16112 15264
rect 16176 15200 16192 15264
rect 16256 15200 16264 15264
rect 15944 14176 16264 15200
rect 15944 14112 15952 14176
rect 16016 14112 16032 14176
rect 16096 14112 16112 14176
rect 16176 14112 16192 14176
rect 16256 14112 16264 14176
rect 15944 13088 16264 14112
rect 15944 13024 15952 13088
rect 16016 13024 16032 13088
rect 16096 13024 16112 13088
rect 16176 13024 16192 13088
rect 16256 13024 16264 13088
rect 15944 12000 16264 13024
rect 15944 11936 15952 12000
rect 16016 11936 16032 12000
rect 16096 11936 16112 12000
rect 16176 11936 16192 12000
rect 16256 11936 16264 12000
rect 15699 11388 15765 11389
rect 15699 11324 15700 11388
rect 15764 11324 15765 11388
rect 15699 11323 15765 11324
rect 15944 10912 16264 11936
rect 15944 10848 15952 10912
rect 16016 10848 16032 10912
rect 16096 10848 16112 10912
rect 16176 10848 16192 10912
rect 16256 10848 16264 10912
rect 15944 9824 16264 10848
rect 15944 9760 15952 9824
rect 16016 9760 16032 9824
rect 16096 9760 16112 9824
rect 16176 9760 16192 9824
rect 16256 9760 16264 9824
rect 15944 8736 16264 9760
rect 15944 8672 15952 8736
rect 16016 8672 16032 8736
rect 16096 8672 16112 8736
rect 16176 8672 16192 8736
rect 16256 8672 16264 8736
rect 15944 7648 16264 8672
rect 15944 7584 15952 7648
rect 16016 7584 16032 7648
rect 16096 7584 16112 7648
rect 16176 7584 16192 7648
rect 16256 7584 16264 7648
rect 15944 6560 16264 7584
rect 15944 6496 15952 6560
rect 16016 6496 16032 6560
rect 16096 6496 16112 6560
rect 16176 6496 16192 6560
rect 16256 6496 16264 6560
rect 15944 5472 16264 6496
rect 15944 5408 15952 5472
rect 16016 5408 16032 5472
rect 16096 5408 16112 5472
rect 16176 5408 16192 5472
rect 16256 5408 16264 5472
rect 15944 4384 16264 5408
rect 15944 4320 15952 4384
rect 16016 4320 16032 4384
rect 16096 4320 16112 4384
rect 16176 4320 16192 4384
rect 16256 4320 16264 4384
rect 15944 3296 16264 4320
rect 16438 4045 16498 46955
rect 16803 37500 16869 37501
rect 16803 37436 16804 37500
rect 16868 37436 16869 37500
rect 16803 37435 16869 37436
rect 16619 37228 16685 37229
rect 16619 37164 16620 37228
rect 16684 37164 16685 37228
rect 16619 37163 16685 37164
rect 16622 36413 16682 37163
rect 16619 36412 16685 36413
rect 16619 36348 16620 36412
rect 16684 36348 16685 36412
rect 16619 36347 16685 36348
rect 16622 35461 16682 36347
rect 16619 35460 16685 35461
rect 16619 35396 16620 35460
rect 16684 35396 16685 35460
rect 16619 35395 16685 35396
rect 16619 33828 16685 33829
rect 16619 33764 16620 33828
rect 16684 33764 16685 33828
rect 16619 33763 16685 33764
rect 16622 30565 16682 33763
rect 16619 30564 16685 30565
rect 16619 30500 16620 30564
rect 16684 30500 16685 30564
rect 16619 30499 16685 30500
rect 16806 30293 16866 37435
rect 16987 36004 17053 36005
rect 16987 35940 16988 36004
rect 17052 35940 17053 36004
rect 16987 35939 17053 35940
rect 16990 32333 17050 35939
rect 16987 32332 17053 32333
rect 16987 32268 16988 32332
rect 17052 32268 17053 32332
rect 16987 32267 17053 32268
rect 16803 30292 16869 30293
rect 16803 30228 16804 30292
rect 16868 30228 16869 30292
rect 16803 30227 16869 30228
rect 16619 27708 16685 27709
rect 16619 27644 16620 27708
rect 16684 27644 16685 27708
rect 16619 27643 16685 27644
rect 16622 23629 16682 27643
rect 16619 23628 16685 23629
rect 16619 23564 16620 23628
rect 16684 23564 16685 23628
rect 16619 23563 16685 23564
rect 17174 17781 17234 69259
rect 18091 62932 18157 62933
rect 18091 62868 18092 62932
rect 18156 62868 18157 62932
rect 18091 62867 18157 62868
rect 17723 56540 17789 56541
rect 17723 56476 17724 56540
rect 17788 56476 17789 56540
rect 17723 56475 17789 56476
rect 17726 52189 17786 56475
rect 17723 52188 17789 52189
rect 17723 52124 17724 52188
rect 17788 52124 17789 52188
rect 17723 52123 17789 52124
rect 17539 30292 17605 30293
rect 17539 30228 17540 30292
rect 17604 30228 17605 30292
rect 17539 30227 17605 30228
rect 17542 27709 17602 30227
rect 17539 27708 17605 27709
rect 17539 27644 17540 27708
rect 17604 27644 17605 27708
rect 17539 27643 17605 27644
rect 18094 21725 18154 62867
rect 20483 57356 20549 57357
rect 20483 57292 20484 57356
rect 20548 57292 20549 57356
rect 20483 57291 20549 57292
rect 20299 50012 20365 50013
rect 20299 49948 20300 50012
rect 20364 49948 20365 50012
rect 20299 49947 20365 49948
rect 20302 49330 20362 49947
rect 20486 49469 20546 57291
rect 20483 49468 20549 49469
rect 20483 49404 20484 49468
rect 20548 49404 20549 49468
rect 20483 49403 20549 49404
rect 20302 49270 20546 49330
rect 20299 49196 20365 49197
rect 20299 49132 20300 49196
rect 20364 49132 20365 49196
rect 20299 49131 20365 49132
rect 19931 47972 19997 47973
rect 19931 47908 19932 47972
rect 19996 47908 19997 47972
rect 19931 47907 19997 47908
rect 19934 42397 19994 47907
rect 20115 46748 20181 46749
rect 20115 46684 20116 46748
rect 20180 46684 20181 46748
rect 20115 46683 20181 46684
rect 20118 45661 20178 46683
rect 20115 45660 20181 45661
rect 20115 45596 20116 45660
rect 20180 45596 20181 45660
rect 20115 45595 20181 45596
rect 19931 42396 19997 42397
rect 19931 42332 19932 42396
rect 19996 42332 19997 42396
rect 19931 42331 19997 42332
rect 20118 41989 20178 45595
rect 20302 44845 20362 49131
rect 20299 44844 20365 44845
rect 20299 44780 20300 44844
rect 20364 44780 20365 44844
rect 20299 44779 20365 44780
rect 20115 41988 20181 41989
rect 20115 41924 20116 41988
rect 20180 41924 20181 41988
rect 20115 41923 20181 41924
rect 20486 41581 20546 49270
rect 20483 41580 20549 41581
rect 20483 41516 20484 41580
rect 20548 41516 20549 41580
rect 20483 41515 20549 41516
rect 20483 41444 20549 41445
rect 20483 41380 20484 41444
rect 20548 41380 20549 41444
rect 20483 41379 20549 41380
rect 20486 41173 20546 41379
rect 20670 41173 20730 77419
rect 20944 76736 21264 77760
rect 20944 76672 20952 76736
rect 21016 76672 21032 76736
rect 21096 76672 21112 76736
rect 21176 76672 21192 76736
rect 21256 76672 21264 76736
rect 20944 75648 21264 76672
rect 20944 75584 20952 75648
rect 21016 75584 21032 75648
rect 21096 75584 21112 75648
rect 21176 75584 21192 75648
rect 21256 75584 21264 75648
rect 20944 74560 21264 75584
rect 25944 77280 26264 77840
rect 25944 77216 25952 77280
rect 26016 77216 26032 77280
rect 26096 77216 26112 77280
rect 26176 77216 26192 77280
rect 26256 77216 26264 77280
rect 25944 76192 26264 77216
rect 25944 76128 25952 76192
rect 26016 76128 26032 76192
rect 26096 76128 26112 76192
rect 26176 76128 26192 76192
rect 26256 76128 26264 76192
rect 25944 75104 26264 76128
rect 25944 75040 25952 75104
rect 26016 75040 26032 75104
rect 26096 75040 26112 75104
rect 26176 75040 26192 75104
rect 26256 75040 26264 75104
rect 25083 74628 25149 74629
rect 25083 74564 25084 74628
rect 25148 74564 25149 74628
rect 25083 74563 25149 74564
rect 20944 74496 20952 74560
rect 21016 74496 21032 74560
rect 21096 74496 21112 74560
rect 21176 74496 21192 74560
rect 21256 74496 21264 74560
rect 20944 73472 21264 74496
rect 24899 74492 24965 74493
rect 24899 74428 24900 74492
rect 24964 74428 24965 74492
rect 24899 74427 24965 74428
rect 20944 73408 20952 73472
rect 21016 73408 21032 73472
rect 21096 73408 21112 73472
rect 21176 73408 21192 73472
rect 21256 73408 21264 73472
rect 20944 72384 21264 73408
rect 20944 72320 20952 72384
rect 21016 72320 21032 72384
rect 21096 72320 21112 72384
rect 21176 72320 21192 72384
rect 21256 72320 21264 72384
rect 20944 71296 21264 72320
rect 20944 71232 20952 71296
rect 21016 71232 21032 71296
rect 21096 71232 21112 71296
rect 21176 71232 21192 71296
rect 21256 71232 21264 71296
rect 20944 70208 21264 71232
rect 20944 70144 20952 70208
rect 21016 70144 21032 70208
rect 21096 70144 21112 70208
rect 21176 70144 21192 70208
rect 21256 70144 21264 70208
rect 20944 69120 21264 70144
rect 20944 69056 20952 69120
rect 21016 69056 21032 69120
rect 21096 69056 21112 69120
rect 21176 69056 21192 69120
rect 21256 69056 21264 69120
rect 20944 68032 21264 69056
rect 20944 67968 20952 68032
rect 21016 67968 21032 68032
rect 21096 67968 21112 68032
rect 21176 67968 21192 68032
rect 21256 67968 21264 68032
rect 20944 66944 21264 67968
rect 20944 66880 20952 66944
rect 21016 66880 21032 66944
rect 21096 66880 21112 66944
rect 21176 66880 21192 66944
rect 21256 66880 21264 66944
rect 20944 65856 21264 66880
rect 20944 65792 20952 65856
rect 21016 65792 21032 65856
rect 21096 65792 21112 65856
rect 21176 65792 21192 65856
rect 21256 65792 21264 65856
rect 20944 64768 21264 65792
rect 21955 65516 22021 65517
rect 21955 65452 21956 65516
rect 22020 65452 22021 65516
rect 21955 65451 22021 65452
rect 20944 64704 20952 64768
rect 21016 64704 21032 64768
rect 21096 64704 21112 64768
rect 21176 64704 21192 64768
rect 21256 64704 21264 64768
rect 20944 63680 21264 64704
rect 21587 64564 21653 64565
rect 21587 64500 21588 64564
rect 21652 64500 21653 64564
rect 21587 64499 21653 64500
rect 20944 63616 20952 63680
rect 21016 63616 21032 63680
rect 21096 63616 21112 63680
rect 21176 63616 21192 63680
rect 21256 63616 21264 63680
rect 20944 62592 21264 63616
rect 20944 62528 20952 62592
rect 21016 62528 21032 62592
rect 21096 62528 21112 62592
rect 21176 62528 21192 62592
rect 21256 62528 21264 62592
rect 20944 61504 21264 62528
rect 20944 61440 20952 61504
rect 21016 61440 21032 61504
rect 21096 61440 21112 61504
rect 21176 61440 21192 61504
rect 21256 61440 21264 61504
rect 20944 60416 21264 61440
rect 20944 60352 20952 60416
rect 21016 60352 21032 60416
rect 21096 60352 21112 60416
rect 21176 60352 21192 60416
rect 21256 60352 21264 60416
rect 20944 59328 21264 60352
rect 20944 59264 20952 59328
rect 21016 59264 21032 59328
rect 21096 59264 21112 59328
rect 21176 59264 21192 59328
rect 21256 59264 21264 59328
rect 20944 58240 21264 59264
rect 20944 58176 20952 58240
rect 21016 58176 21032 58240
rect 21096 58176 21112 58240
rect 21176 58176 21192 58240
rect 21256 58176 21264 58240
rect 20944 57152 21264 58176
rect 20944 57088 20952 57152
rect 21016 57088 21032 57152
rect 21096 57088 21112 57152
rect 21176 57088 21192 57152
rect 21256 57088 21264 57152
rect 20944 56064 21264 57088
rect 20944 56000 20952 56064
rect 21016 56000 21032 56064
rect 21096 56000 21112 56064
rect 21176 56000 21192 56064
rect 21256 56000 21264 56064
rect 20944 55579 21264 56000
rect 20944 55343 20986 55579
rect 21222 55343 21264 55579
rect 20944 54976 21264 55343
rect 21403 55316 21469 55317
rect 21403 55252 21404 55316
rect 21468 55252 21469 55316
rect 21403 55251 21469 55252
rect 20944 54912 20952 54976
rect 21016 54912 21032 54976
rect 21096 54912 21112 54976
rect 21176 54912 21192 54976
rect 21256 54912 21264 54976
rect 20944 53888 21264 54912
rect 20944 53824 20952 53888
rect 21016 53824 21032 53888
rect 21096 53824 21112 53888
rect 21176 53824 21192 53888
rect 21256 53824 21264 53888
rect 20944 52800 21264 53824
rect 20944 52736 20952 52800
rect 21016 52736 21032 52800
rect 21096 52736 21112 52800
rect 21176 52736 21192 52800
rect 21256 52736 21264 52800
rect 20944 51712 21264 52736
rect 20944 51648 20952 51712
rect 21016 51648 21032 51712
rect 21096 51648 21112 51712
rect 21176 51648 21192 51712
rect 21256 51648 21264 51712
rect 20944 50624 21264 51648
rect 20944 50560 20952 50624
rect 21016 50560 21032 50624
rect 21096 50560 21112 50624
rect 21176 50560 21192 50624
rect 21256 50560 21264 50624
rect 20944 49536 21264 50560
rect 20944 49472 20952 49536
rect 21016 49472 21032 49536
rect 21096 49472 21112 49536
rect 21176 49472 21192 49536
rect 21256 49472 21264 49536
rect 20944 48448 21264 49472
rect 20944 48384 20952 48448
rect 21016 48384 21032 48448
rect 21096 48384 21112 48448
rect 21176 48384 21192 48448
rect 21256 48384 21264 48448
rect 20944 47360 21264 48384
rect 20944 47296 20952 47360
rect 21016 47296 21032 47360
rect 21096 47296 21112 47360
rect 21176 47296 21192 47360
rect 21256 47296 21264 47360
rect 20944 46272 21264 47296
rect 20944 46208 20952 46272
rect 21016 46208 21032 46272
rect 21096 46208 21112 46272
rect 21176 46208 21192 46272
rect 21256 46208 21264 46272
rect 20944 45184 21264 46208
rect 20944 45120 20952 45184
rect 21016 45120 21032 45184
rect 21096 45120 21112 45184
rect 21176 45120 21192 45184
rect 21256 45120 21264 45184
rect 20944 44096 21264 45120
rect 20944 44032 20952 44096
rect 21016 44032 21032 44096
rect 21096 44032 21112 44096
rect 21176 44032 21192 44096
rect 21256 44032 21264 44096
rect 20944 43008 21264 44032
rect 20944 42944 20952 43008
rect 21016 42944 21032 43008
rect 21096 42944 21112 43008
rect 21176 42944 21192 43008
rect 21256 42944 21264 43008
rect 20944 41920 21264 42944
rect 20944 41856 20952 41920
rect 21016 41856 21032 41920
rect 21096 41856 21112 41920
rect 21176 41856 21192 41920
rect 21256 41856 21264 41920
rect 20483 41172 20549 41173
rect 20483 41108 20484 41172
rect 20548 41108 20549 41172
rect 20483 41107 20549 41108
rect 20667 41172 20733 41173
rect 20667 41108 20668 41172
rect 20732 41108 20733 41172
rect 20667 41107 20733 41108
rect 20483 40900 20549 40901
rect 20483 40836 20484 40900
rect 20548 40836 20549 40900
rect 20483 40835 20549 40836
rect 20486 31109 20546 40835
rect 20944 40832 21264 41856
rect 20944 40768 20952 40832
rect 21016 40768 21032 40832
rect 21096 40768 21112 40832
rect 21176 40768 21192 40832
rect 21256 40768 21264 40832
rect 20944 39744 21264 40768
rect 20944 39680 20952 39744
rect 21016 39680 21032 39744
rect 21096 39680 21112 39744
rect 21176 39680 21192 39744
rect 21256 39680 21264 39744
rect 20944 38656 21264 39680
rect 20944 38592 20952 38656
rect 21016 38592 21032 38656
rect 21096 38592 21112 38656
rect 21176 38592 21192 38656
rect 21256 38592 21264 38656
rect 20944 37568 21264 38592
rect 20944 37504 20952 37568
rect 21016 37504 21032 37568
rect 21096 37504 21112 37568
rect 21176 37504 21192 37568
rect 21256 37504 21264 37568
rect 20944 36480 21264 37504
rect 20944 36416 20952 36480
rect 21016 36416 21032 36480
rect 21096 36416 21112 36480
rect 21176 36416 21192 36480
rect 21256 36416 21264 36480
rect 20944 35392 21264 36416
rect 20944 35328 20952 35392
rect 21016 35328 21032 35392
rect 21096 35328 21112 35392
rect 21176 35328 21192 35392
rect 21256 35328 21264 35392
rect 20944 34304 21264 35328
rect 20944 34240 20952 34304
rect 21016 34240 21032 34304
rect 21096 34240 21112 34304
rect 21176 34240 21192 34304
rect 21256 34240 21264 34304
rect 20944 33216 21264 34240
rect 20944 33152 20952 33216
rect 21016 33152 21032 33216
rect 21096 33152 21112 33216
rect 21176 33152 21192 33216
rect 21256 33152 21264 33216
rect 20944 32128 21264 33152
rect 20944 32064 20952 32128
rect 21016 32064 21032 32128
rect 21096 32064 21112 32128
rect 21176 32064 21192 32128
rect 21256 32064 21264 32128
rect 20667 31924 20733 31925
rect 20667 31860 20668 31924
rect 20732 31860 20733 31924
rect 20667 31859 20733 31860
rect 20483 31108 20549 31109
rect 20483 31044 20484 31108
rect 20548 31044 20549 31108
rect 20483 31043 20549 31044
rect 20670 30837 20730 31859
rect 20944 31040 21264 32064
rect 20944 30976 20952 31040
rect 21016 30976 21032 31040
rect 21096 30976 21112 31040
rect 21176 30976 21192 31040
rect 21256 30976 21264 31040
rect 20667 30836 20733 30837
rect 20667 30772 20668 30836
rect 20732 30772 20733 30836
rect 20667 30771 20733 30772
rect 20944 29952 21264 30976
rect 20944 29888 20952 29952
rect 21016 29888 21032 29952
rect 21096 29888 21112 29952
rect 21176 29888 21192 29952
rect 21256 29888 21264 29952
rect 20944 28912 21264 29888
rect 20944 28864 20986 28912
rect 21222 28864 21264 28912
rect 20944 28800 20952 28864
rect 21256 28800 21264 28864
rect 20944 28676 20986 28800
rect 21222 28676 21264 28800
rect 20944 27776 21264 28676
rect 20944 27712 20952 27776
rect 21016 27712 21032 27776
rect 21096 27712 21112 27776
rect 21176 27712 21192 27776
rect 21256 27712 21264 27776
rect 20944 26688 21264 27712
rect 20944 26624 20952 26688
rect 21016 26624 21032 26688
rect 21096 26624 21112 26688
rect 21176 26624 21192 26688
rect 21256 26624 21264 26688
rect 20944 25600 21264 26624
rect 20944 25536 20952 25600
rect 21016 25536 21032 25600
rect 21096 25536 21112 25600
rect 21176 25536 21192 25600
rect 21256 25536 21264 25600
rect 20944 24512 21264 25536
rect 20944 24448 20952 24512
rect 21016 24448 21032 24512
rect 21096 24448 21112 24512
rect 21176 24448 21192 24512
rect 21256 24448 21264 24512
rect 20944 23424 21264 24448
rect 20944 23360 20952 23424
rect 21016 23360 21032 23424
rect 21096 23360 21112 23424
rect 21176 23360 21192 23424
rect 21256 23360 21264 23424
rect 20944 22336 21264 23360
rect 20944 22272 20952 22336
rect 21016 22272 21032 22336
rect 21096 22272 21112 22336
rect 21176 22272 21192 22336
rect 21256 22272 21264 22336
rect 18091 21724 18157 21725
rect 18091 21660 18092 21724
rect 18156 21660 18157 21724
rect 18091 21659 18157 21660
rect 20944 21248 21264 22272
rect 20944 21184 20952 21248
rect 21016 21184 21032 21248
rect 21096 21184 21112 21248
rect 21176 21184 21192 21248
rect 21256 21184 21264 21248
rect 20944 20160 21264 21184
rect 20944 20096 20952 20160
rect 21016 20096 21032 20160
rect 21096 20096 21112 20160
rect 21176 20096 21192 20160
rect 21256 20096 21264 20160
rect 20944 19072 21264 20096
rect 20944 19008 20952 19072
rect 21016 19008 21032 19072
rect 21096 19008 21112 19072
rect 21176 19008 21192 19072
rect 21256 19008 21264 19072
rect 20944 17984 21264 19008
rect 20944 17920 20952 17984
rect 21016 17920 21032 17984
rect 21096 17920 21112 17984
rect 21176 17920 21192 17984
rect 21256 17920 21264 17984
rect 17171 17780 17237 17781
rect 17171 17716 17172 17780
rect 17236 17716 17237 17780
rect 17171 17715 17237 17716
rect 20944 16896 21264 17920
rect 20944 16832 20952 16896
rect 21016 16832 21032 16896
rect 21096 16832 21112 16896
rect 21176 16832 21192 16896
rect 21256 16832 21264 16896
rect 20944 15808 21264 16832
rect 20944 15744 20952 15808
rect 21016 15744 21032 15808
rect 21096 15744 21112 15808
rect 21176 15744 21192 15808
rect 21256 15744 21264 15808
rect 20944 14720 21264 15744
rect 20944 14656 20952 14720
rect 21016 14656 21032 14720
rect 21096 14656 21112 14720
rect 21176 14656 21192 14720
rect 21256 14656 21264 14720
rect 20944 13632 21264 14656
rect 20944 13568 20952 13632
rect 21016 13568 21032 13632
rect 21096 13568 21112 13632
rect 21176 13568 21192 13632
rect 21256 13568 21264 13632
rect 19379 12748 19445 12749
rect 19379 12684 19380 12748
rect 19444 12684 19445 12748
rect 19379 12683 19445 12684
rect 19382 12341 19442 12683
rect 20944 12544 21264 13568
rect 20944 12480 20952 12544
rect 21016 12480 21032 12544
rect 21096 12480 21112 12544
rect 21176 12480 21192 12544
rect 21256 12480 21264 12544
rect 19379 12340 19445 12341
rect 19379 12276 19380 12340
rect 19444 12276 19445 12340
rect 19379 12275 19445 12276
rect 20944 11456 21264 12480
rect 20944 11392 20952 11456
rect 21016 11392 21032 11456
rect 21096 11392 21112 11456
rect 21176 11392 21192 11456
rect 21256 11392 21264 11456
rect 20944 10368 21264 11392
rect 20944 10304 20952 10368
rect 21016 10304 21032 10368
rect 21096 10304 21112 10368
rect 21176 10304 21192 10368
rect 21256 10304 21264 10368
rect 20944 9280 21264 10304
rect 20944 9216 20952 9280
rect 21016 9216 21032 9280
rect 21096 9216 21112 9280
rect 21176 9216 21192 9280
rect 21256 9216 21264 9280
rect 20944 8192 21264 9216
rect 20944 8128 20952 8192
rect 21016 8128 21032 8192
rect 21096 8128 21112 8192
rect 21176 8128 21192 8192
rect 21256 8128 21264 8192
rect 20944 7104 21264 8128
rect 20944 7040 20952 7104
rect 21016 7040 21032 7104
rect 21096 7040 21112 7104
rect 21176 7040 21192 7104
rect 21256 7040 21264 7104
rect 20944 6016 21264 7040
rect 20944 5952 20952 6016
rect 21016 5952 21032 6016
rect 21096 5952 21112 6016
rect 21176 5952 21192 6016
rect 21256 5952 21264 6016
rect 20944 4928 21264 5952
rect 20944 4864 20952 4928
rect 21016 4864 21032 4928
rect 21096 4864 21112 4928
rect 21176 4864 21192 4928
rect 21256 4864 21264 4928
rect 16435 4044 16501 4045
rect 16435 3980 16436 4044
rect 16500 3980 16501 4044
rect 16435 3979 16501 3980
rect 15944 3232 15952 3296
rect 16016 3232 16032 3296
rect 16096 3232 16112 3296
rect 16176 3232 16192 3296
rect 16256 3232 16264 3296
rect 15515 3228 15581 3229
rect 15515 3164 15516 3228
rect 15580 3164 15581 3228
rect 15515 3163 15581 3164
rect 10944 2688 10952 2752
rect 11016 2688 11032 2752
rect 11096 2688 11112 2752
rect 11176 2688 11192 2752
rect 11256 2688 11264 2752
rect 10944 2128 11264 2688
rect 15944 2208 16264 3232
rect 15944 2144 15952 2208
rect 16016 2144 16032 2208
rect 16096 2144 16112 2208
rect 16176 2144 16192 2208
rect 16256 2144 16264 2208
rect 15944 2128 16264 2144
rect 20944 3840 21264 4864
rect 20944 3776 20952 3840
rect 21016 3776 21032 3840
rect 21096 3776 21112 3840
rect 21176 3776 21192 3840
rect 21256 3776 21264 3840
rect 20944 2752 21264 3776
rect 21406 3773 21466 55251
rect 21590 35869 21650 64499
rect 21771 53140 21837 53141
rect 21771 53076 21772 53140
rect 21836 53076 21837 53140
rect 21771 53075 21837 53076
rect 21774 48517 21834 53075
rect 21771 48516 21837 48517
rect 21771 48452 21772 48516
rect 21836 48452 21837 48516
rect 21771 48451 21837 48452
rect 21771 38724 21837 38725
rect 21771 38660 21772 38724
rect 21836 38660 21837 38724
rect 21771 38659 21837 38660
rect 21587 35868 21653 35869
rect 21587 35804 21588 35868
rect 21652 35804 21653 35868
rect 21587 35803 21653 35804
rect 21774 32469 21834 38659
rect 21958 36413 22018 65451
rect 23979 47700 24045 47701
rect 23979 47636 23980 47700
rect 24044 47636 24045 47700
rect 23979 47635 24045 47636
rect 23059 44708 23125 44709
rect 23059 44658 23060 44708
rect 23124 44658 23125 44708
rect 23062 41445 23122 44422
rect 23059 41444 23125 41445
rect 23059 41380 23060 41444
rect 23124 41380 23125 41444
rect 23059 41379 23125 41380
rect 23982 40901 24042 47635
rect 24715 41580 24781 41581
rect 24715 41516 24716 41580
rect 24780 41516 24781 41580
rect 24715 41515 24781 41516
rect 23979 40900 24045 40901
rect 23979 40836 23980 40900
rect 24044 40836 24045 40900
rect 23979 40835 24045 40836
rect 24718 39269 24778 41515
rect 24715 39268 24781 39269
rect 24715 39204 24716 39268
rect 24780 39204 24781 39268
rect 24715 39203 24781 39204
rect 24350 38453 24410 38982
rect 24347 38452 24413 38453
rect 24347 38388 24348 38452
rect 24412 38388 24413 38452
rect 24347 38387 24413 38388
rect 21955 36412 22021 36413
rect 21955 36348 21956 36412
rect 22020 36348 22021 36412
rect 21955 36347 22021 36348
rect 21771 32468 21837 32469
rect 21771 32404 21772 32468
rect 21836 32404 21837 32468
rect 21771 32403 21837 32404
rect 21403 3772 21469 3773
rect 21403 3708 21404 3772
rect 21468 3708 21469 3772
rect 21403 3707 21469 3708
rect 20944 2688 20952 2752
rect 21016 2688 21032 2752
rect 21096 2688 21112 2752
rect 21176 2688 21192 2752
rect 21256 2688 21264 2752
rect 20944 2128 21264 2688
rect 24902 2685 24962 74427
rect 25086 31381 25146 74563
rect 25944 74016 26264 75040
rect 25944 73952 25952 74016
rect 26016 73952 26032 74016
rect 26096 73952 26112 74016
rect 26176 73952 26192 74016
rect 26256 73952 26264 74016
rect 25944 72928 26264 73952
rect 25944 72864 25952 72928
rect 26016 72864 26032 72928
rect 26096 72864 26112 72928
rect 26176 72864 26192 72928
rect 26256 72864 26264 72928
rect 25944 71840 26264 72864
rect 25944 71776 25952 71840
rect 26016 71776 26032 71840
rect 26096 71776 26112 71840
rect 26176 71776 26192 71840
rect 26256 71776 26264 71840
rect 25944 70752 26264 71776
rect 25944 70688 25952 70752
rect 26016 70688 26032 70752
rect 26096 70688 26112 70752
rect 26176 70688 26192 70752
rect 26256 70688 26264 70752
rect 25944 69664 26264 70688
rect 25944 69600 25952 69664
rect 26016 69600 26032 69664
rect 26096 69600 26112 69664
rect 26176 69600 26192 69664
rect 26256 69600 26264 69664
rect 25944 68912 26264 69600
rect 25635 68780 25701 68781
rect 25635 68716 25636 68780
rect 25700 68716 25701 68780
rect 25635 68715 25701 68716
rect 25451 53004 25517 53005
rect 25451 52940 25452 53004
rect 25516 52940 25517 53004
rect 25451 52939 25517 52940
rect 25267 45660 25333 45661
rect 25267 45596 25268 45660
rect 25332 45596 25333 45660
rect 25267 45595 25333 45596
rect 25083 31380 25149 31381
rect 25083 31316 25084 31380
rect 25148 31316 25149 31380
rect 25083 31315 25149 31316
rect 25270 8261 25330 45595
rect 25454 38589 25514 52939
rect 25451 38588 25517 38589
rect 25451 38524 25452 38588
rect 25516 38524 25517 38588
rect 25451 38523 25517 38524
rect 25451 38452 25517 38453
rect 25451 38388 25452 38452
rect 25516 38388 25517 38452
rect 25451 38387 25517 38388
rect 25454 35053 25514 38387
rect 25451 35052 25517 35053
rect 25451 34988 25452 35052
rect 25516 34988 25517 35052
rect 25451 34987 25517 34988
rect 25638 23629 25698 68715
rect 25944 68676 25986 68912
rect 26222 68676 26264 68912
rect 25944 68576 26264 68676
rect 25944 68512 25952 68576
rect 26016 68512 26032 68576
rect 26096 68512 26112 68576
rect 26176 68512 26192 68576
rect 26256 68512 26264 68576
rect 25944 67488 26264 68512
rect 25944 67424 25952 67488
rect 26016 67424 26032 67488
rect 26096 67424 26112 67488
rect 26176 67424 26192 67488
rect 26256 67424 26264 67488
rect 25944 66400 26264 67424
rect 25944 66336 25952 66400
rect 26016 66336 26032 66400
rect 26096 66336 26112 66400
rect 26176 66336 26192 66400
rect 26256 66336 26264 66400
rect 25944 65312 26264 66336
rect 27843 66196 27909 66197
rect 27843 66132 27844 66196
rect 27908 66132 27909 66196
rect 27843 66131 27909 66132
rect 25944 65248 25952 65312
rect 26016 65248 26032 65312
rect 26096 65248 26112 65312
rect 26176 65248 26192 65312
rect 26256 65248 26264 65312
rect 25944 64224 26264 65248
rect 25944 64160 25952 64224
rect 26016 64160 26032 64224
rect 26096 64160 26112 64224
rect 26176 64160 26192 64224
rect 26256 64160 26264 64224
rect 25944 63136 26264 64160
rect 25944 63072 25952 63136
rect 26016 63072 26032 63136
rect 26096 63072 26112 63136
rect 26176 63072 26192 63136
rect 26256 63072 26264 63136
rect 25944 62048 26264 63072
rect 25944 61984 25952 62048
rect 26016 61984 26032 62048
rect 26096 61984 26112 62048
rect 26176 61984 26192 62048
rect 26256 61984 26264 62048
rect 25944 60960 26264 61984
rect 25944 60896 25952 60960
rect 26016 60896 26032 60960
rect 26096 60896 26112 60960
rect 26176 60896 26192 60960
rect 26256 60896 26264 60960
rect 25944 59872 26264 60896
rect 25944 59808 25952 59872
rect 26016 59808 26032 59872
rect 26096 59808 26112 59872
rect 26176 59808 26192 59872
rect 26256 59808 26264 59872
rect 25944 58784 26264 59808
rect 25944 58720 25952 58784
rect 26016 58720 26032 58784
rect 26096 58720 26112 58784
rect 26176 58720 26192 58784
rect 26256 58720 26264 58784
rect 25944 57696 26264 58720
rect 25944 57632 25952 57696
rect 26016 57632 26032 57696
rect 26096 57632 26112 57696
rect 26176 57632 26192 57696
rect 26256 57632 26264 57696
rect 25944 56608 26264 57632
rect 27846 56677 27906 66131
rect 27843 56676 27909 56677
rect 27843 56612 27844 56676
rect 27908 56612 27909 56676
rect 27843 56611 27909 56612
rect 25944 56544 25952 56608
rect 26016 56544 26032 56608
rect 26096 56544 26112 56608
rect 26176 56544 26192 56608
rect 26256 56544 26264 56608
rect 25944 55520 26264 56544
rect 25944 55456 25952 55520
rect 26016 55456 26032 55520
rect 26096 55456 26112 55520
rect 26176 55456 26192 55520
rect 26256 55456 26264 55520
rect 25944 54432 26264 55456
rect 25944 54368 25952 54432
rect 26016 54368 26032 54432
rect 26096 54368 26112 54432
rect 26176 54368 26192 54432
rect 26256 54368 26264 54432
rect 25944 53344 26264 54368
rect 25944 53280 25952 53344
rect 26016 53280 26032 53344
rect 26096 53280 26112 53344
rect 26176 53280 26192 53344
rect 26256 53280 26264 53344
rect 25944 52256 26264 53280
rect 25944 52192 25952 52256
rect 26016 52192 26032 52256
rect 26096 52192 26112 52256
rect 26176 52192 26192 52256
rect 26256 52192 26264 52256
rect 25944 51168 26264 52192
rect 25944 51104 25952 51168
rect 26016 51104 26032 51168
rect 26096 51104 26112 51168
rect 26176 51104 26192 51168
rect 26256 51104 26264 51168
rect 25944 50080 26264 51104
rect 25944 50016 25952 50080
rect 26016 50016 26032 50080
rect 26096 50016 26112 50080
rect 26176 50016 26192 50080
rect 26256 50016 26264 50080
rect 25944 48992 26264 50016
rect 25944 48928 25952 48992
rect 26016 48928 26032 48992
rect 26096 48928 26112 48992
rect 26176 48928 26192 48992
rect 26256 48928 26264 48992
rect 25944 47904 26264 48928
rect 25944 47840 25952 47904
rect 26016 47840 26032 47904
rect 26096 47840 26112 47904
rect 26176 47840 26192 47904
rect 26256 47840 26264 47904
rect 25944 46816 26264 47840
rect 25944 46752 25952 46816
rect 26016 46752 26032 46816
rect 26096 46752 26112 46816
rect 26176 46752 26192 46816
rect 26256 46752 26264 46816
rect 25944 45728 26264 46752
rect 25944 45664 25952 45728
rect 26016 45664 26032 45728
rect 26096 45664 26112 45728
rect 26176 45664 26192 45728
rect 26256 45664 26264 45728
rect 25944 44640 26264 45664
rect 25944 44576 25952 44640
rect 26016 44576 26032 44640
rect 26096 44576 26112 44640
rect 26176 44576 26192 44640
rect 26256 44576 26264 44640
rect 25944 43552 26264 44576
rect 25944 43488 25952 43552
rect 26016 43488 26032 43552
rect 26096 43488 26112 43552
rect 26176 43488 26192 43552
rect 26256 43488 26264 43552
rect 25944 42464 26264 43488
rect 25944 42400 25952 42464
rect 26016 42400 26032 42464
rect 26096 42400 26112 42464
rect 26176 42400 26192 42464
rect 26256 42400 26264 42464
rect 25944 42246 26264 42400
rect 25944 42010 25986 42246
rect 26222 42010 26264 42246
rect 25944 41376 26264 42010
rect 25944 41312 25952 41376
rect 26016 41312 26032 41376
rect 26096 41312 26112 41376
rect 26176 41312 26192 41376
rect 26256 41312 26264 41376
rect 25944 40288 26264 41312
rect 25944 40224 25952 40288
rect 26016 40224 26032 40288
rect 26096 40224 26112 40288
rect 26176 40224 26192 40288
rect 26256 40224 26264 40288
rect 25944 39200 26264 40224
rect 25944 39136 25952 39200
rect 26016 39136 26032 39200
rect 26096 39136 26112 39200
rect 26176 39136 26192 39200
rect 26256 39136 26264 39200
rect 25944 38112 26264 39136
rect 25944 38048 25952 38112
rect 26016 38048 26032 38112
rect 26096 38048 26112 38112
rect 26176 38048 26192 38112
rect 26256 38048 26264 38112
rect 25944 37024 26264 38048
rect 25944 36960 25952 37024
rect 26016 36960 26032 37024
rect 26096 36960 26112 37024
rect 26176 36960 26192 37024
rect 26256 36960 26264 37024
rect 25944 35936 26264 36960
rect 25944 35872 25952 35936
rect 26016 35872 26032 35936
rect 26096 35872 26112 35936
rect 26176 35872 26192 35936
rect 26256 35872 26264 35936
rect 25944 34848 26264 35872
rect 25944 34784 25952 34848
rect 26016 34784 26032 34848
rect 26096 34784 26112 34848
rect 26176 34784 26192 34848
rect 26256 34784 26264 34848
rect 25944 33760 26264 34784
rect 25944 33696 25952 33760
rect 26016 33696 26032 33760
rect 26096 33696 26112 33760
rect 26176 33696 26192 33760
rect 26256 33696 26264 33760
rect 25944 32672 26264 33696
rect 25944 32608 25952 32672
rect 26016 32608 26032 32672
rect 26096 32608 26112 32672
rect 26176 32608 26192 32672
rect 26256 32608 26264 32672
rect 25944 31584 26264 32608
rect 25944 31520 25952 31584
rect 26016 31520 26032 31584
rect 26096 31520 26112 31584
rect 26176 31520 26192 31584
rect 26256 31520 26264 31584
rect 25944 30496 26264 31520
rect 25944 30432 25952 30496
rect 26016 30432 26032 30496
rect 26096 30432 26112 30496
rect 26176 30432 26192 30496
rect 26256 30432 26264 30496
rect 25944 29408 26264 30432
rect 25944 29344 25952 29408
rect 26016 29344 26032 29408
rect 26096 29344 26112 29408
rect 26176 29344 26192 29408
rect 26256 29344 26264 29408
rect 25944 28320 26264 29344
rect 25944 28256 25952 28320
rect 26016 28256 26032 28320
rect 26096 28256 26112 28320
rect 26176 28256 26192 28320
rect 26256 28256 26264 28320
rect 25944 27232 26264 28256
rect 25944 27168 25952 27232
rect 26016 27168 26032 27232
rect 26096 27168 26112 27232
rect 26176 27168 26192 27232
rect 26256 27168 26264 27232
rect 25944 26144 26264 27168
rect 25944 26080 25952 26144
rect 26016 26080 26032 26144
rect 26096 26080 26112 26144
rect 26176 26080 26192 26144
rect 26256 26080 26264 26144
rect 25944 25056 26264 26080
rect 25944 24992 25952 25056
rect 26016 24992 26032 25056
rect 26096 24992 26112 25056
rect 26176 24992 26192 25056
rect 26256 24992 26264 25056
rect 25944 23968 26264 24992
rect 25944 23904 25952 23968
rect 26016 23904 26032 23968
rect 26096 23904 26112 23968
rect 26176 23904 26192 23968
rect 26256 23904 26264 23968
rect 25635 23628 25701 23629
rect 25635 23564 25636 23628
rect 25700 23564 25701 23628
rect 25635 23563 25701 23564
rect 25944 22880 26264 23904
rect 25944 22816 25952 22880
rect 26016 22816 26032 22880
rect 26096 22816 26112 22880
rect 26176 22816 26192 22880
rect 26256 22816 26264 22880
rect 25944 21792 26264 22816
rect 25944 21728 25952 21792
rect 26016 21728 26032 21792
rect 26096 21728 26112 21792
rect 26176 21728 26192 21792
rect 26256 21728 26264 21792
rect 25944 20704 26264 21728
rect 25944 20640 25952 20704
rect 26016 20640 26032 20704
rect 26096 20640 26112 20704
rect 26176 20640 26192 20704
rect 26256 20640 26264 20704
rect 25944 19616 26264 20640
rect 25944 19552 25952 19616
rect 26016 19552 26032 19616
rect 26096 19552 26112 19616
rect 26176 19552 26192 19616
rect 26256 19552 26264 19616
rect 25944 18528 26264 19552
rect 25944 18464 25952 18528
rect 26016 18464 26032 18528
rect 26096 18464 26112 18528
rect 26176 18464 26192 18528
rect 26256 18464 26264 18528
rect 25944 17440 26264 18464
rect 25944 17376 25952 17440
rect 26016 17376 26032 17440
rect 26096 17376 26112 17440
rect 26176 17376 26192 17440
rect 26256 17376 26264 17440
rect 25944 16352 26264 17376
rect 25944 16288 25952 16352
rect 26016 16288 26032 16352
rect 26096 16288 26112 16352
rect 26176 16288 26192 16352
rect 26256 16288 26264 16352
rect 25944 15579 26264 16288
rect 25944 15343 25986 15579
rect 26222 15343 26264 15579
rect 25944 15264 26264 15343
rect 25944 15200 25952 15264
rect 26016 15200 26032 15264
rect 26096 15200 26112 15264
rect 26176 15200 26192 15264
rect 26256 15200 26264 15264
rect 25944 14176 26264 15200
rect 25944 14112 25952 14176
rect 26016 14112 26032 14176
rect 26096 14112 26112 14176
rect 26176 14112 26192 14176
rect 26256 14112 26264 14176
rect 25944 13088 26264 14112
rect 25944 13024 25952 13088
rect 26016 13024 26032 13088
rect 26096 13024 26112 13088
rect 26176 13024 26192 13088
rect 26256 13024 26264 13088
rect 25944 12000 26264 13024
rect 25944 11936 25952 12000
rect 26016 11936 26032 12000
rect 26096 11936 26112 12000
rect 26176 11936 26192 12000
rect 26256 11936 26264 12000
rect 25944 10912 26264 11936
rect 25944 10848 25952 10912
rect 26016 10848 26032 10912
rect 26096 10848 26112 10912
rect 26176 10848 26192 10912
rect 26256 10848 26264 10912
rect 25944 9824 26264 10848
rect 25944 9760 25952 9824
rect 26016 9760 26032 9824
rect 26096 9760 26112 9824
rect 26176 9760 26192 9824
rect 26256 9760 26264 9824
rect 25944 8736 26264 9760
rect 25944 8672 25952 8736
rect 26016 8672 26032 8736
rect 26096 8672 26112 8736
rect 26176 8672 26192 8736
rect 26256 8672 26264 8736
rect 25267 8260 25333 8261
rect 25267 8196 25268 8260
rect 25332 8196 25333 8260
rect 25267 8195 25333 8196
rect 25944 7648 26264 8672
rect 25944 7584 25952 7648
rect 26016 7584 26032 7648
rect 26096 7584 26112 7648
rect 26176 7584 26192 7648
rect 26256 7584 26264 7648
rect 25944 6560 26264 7584
rect 25944 6496 25952 6560
rect 26016 6496 26032 6560
rect 26096 6496 26112 6560
rect 26176 6496 26192 6560
rect 26256 6496 26264 6560
rect 25944 5472 26264 6496
rect 25944 5408 25952 5472
rect 26016 5408 26032 5472
rect 26096 5408 26112 5472
rect 26176 5408 26192 5472
rect 26256 5408 26264 5472
rect 25944 4384 26264 5408
rect 25944 4320 25952 4384
rect 26016 4320 26032 4384
rect 26096 4320 26112 4384
rect 26176 4320 26192 4384
rect 26256 4320 26264 4384
rect 25944 3296 26264 4320
rect 25944 3232 25952 3296
rect 26016 3232 26032 3296
rect 26096 3232 26112 3296
rect 26176 3232 26192 3296
rect 26256 3232 26264 3296
rect 24899 2684 24965 2685
rect 24899 2620 24900 2684
rect 24964 2620 24965 2684
rect 24899 2619 24965 2620
rect 25944 2208 26264 3232
rect 25944 2144 25952 2208
rect 26016 2144 26032 2208
rect 26096 2144 26112 2208
rect 26176 2144 26192 2208
rect 26256 2144 26264 2208
rect 25944 2128 26264 2144
<< via4 >>
rect 5986 68676 6222 68912
rect 3102 44572 3338 44658
rect 3102 44508 3188 44572
rect 3188 44508 3252 44572
rect 3252 44508 3338 44572
rect 3102 44422 3338 44508
rect 5986 42010 6222 42246
rect 5494 38982 5730 39218
rect 3286 37622 3522 37858
rect 3654 36942 3890 37178
rect 6598 32862 6834 33098
rect 10986 55343 11222 55579
rect 10986 28864 11222 28912
rect 10986 28800 11016 28864
rect 11016 28800 11032 28864
rect 11032 28800 11096 28864
rect 11096 28800 11112 28864
rect 11112 28800 11176 28864
rect 11176 28800 11192 28864
rect 11192 28800 11222 28864
rect 10986 28676 11222 28800
rect 5986 15343 6222 15579
rect 15986 68676 16222 68912
rect 14694 33542 14930 33778
rect 15986 42010 16222 42246
rect 15986 15343 16222 15579
rect 20986 55343 21222 55579
rect 19294 37772 19530 37858
rect 19294 37708 19380 37772
rect 19380 37708 19444 37772
rect 19444 37708 19530 37772
rect 19294 37622 19530 37708
rect 20986 28864 21222 28912
rect 20986 28800 21016 28864
rect 21016 28800 21032 28864
rect 21032 28800 21096 28864
rect 21096 28800 21112 28864
rect 21112 28800 21176 28864
rect 21176 28800 21192 28864
rect 21192 28800 21222 28864
rect 20986 28676 21222 28800
rect 22974 44644 23060 44658
rect 23060 44644 23124 44658
rect 23124 44644 23210 44658
rect 22974 44422 23210 44644
rect 24262 38982 24498 39218
rect 23710 37092 23946 37178
rect 23710 37028 23796 37092
rect 23796 37028 23860 37092
rect 23860 37028 23946 37092
rect 23710 36942 23946 37028
rect 25986 68676 26222 68912
rect 25986 42010 26222 42246
rect 25986 15343 26222 15579
<< metal5 >>
rect 1104 68912 28888 68954
rect 1104 68676 5986 68912
rect 6222 68676 15986 68912
rect 16222 68676 25986 68912
rect 26222 68676 28888 68912
rect 1104 68634 28888 68676
rect 1104 55579 28888 55621
rect 1104 55343 10986 55579
rect 11222 55343 20986 55579
rect 21222 55343 28888 55579
rect 1104 55301 28888 55343
rect 3060 44658 23252 44700
rect 3060 44422 3102 44658
rect 3338 44422 22974 44658
rect 23210 44422 23252 44658
rect 3060 44380 23252 44422
rect 1104 42246 28888 42288
rect 1104 42010 5986 42246
rect 6222 42010 15986 42246
rect 16222 42010 25986 42246
rect 26222 42010 28888 42246
rect 1104 41968 28888 42010
rect 5452 39218 24540 39260
rect 5452 38982 5494 39218
rect 5730 38982 24262 39218
rect 24498 38982 24540 39218
rect 5452 38940 24540 38982
rect 3244 37858 19572 37900
rect 3244 37622 3286 37858
rect 3522 37622 19294 37858
rect 19530 37622 19572 37858
rect 3244 37580 19572 37622
rect 3612 37178 23988 37220
rect 3612 36942 3654 37178
rect 3890 36942 23710 37178
rect 23946 36942 23988 37178
rect 3612 36900 23988 36942
rect 13594 33778 14972 33820
rect 13594 33542 14694 33778
rect 14930 33542 14972 33778
rect 13594 33500 14972 33542
rect 13594 33140 13914 33500
rect 6556 33098 13914 33140
rect 6556 32862 6598 33098
rect 6834 32862 13914 33098
rect 6556 32820 13914 32862
rect 1104 28912 28888 28955
rect 1104 28676 10986 28912
rect 11222 28676 20986 28912
rect 21222 28676 28888 28912
rect 1104 28634 28888 28676
rect 1104 15579 28888 15621
rect 1104 15343 5986 15579
rect 6222 15343 15986 15579
rect 16222 15343 25986 15579
rect 26222 15343 28888 15579
rect 1104 15301 28888 15343
use sky130_fd_sc_hd__decap_3  PHY_0 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 1104 0 -1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606120353
transform 1 0 1104 0 1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 1380 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1606120353
transform 1 0 2484 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1606120353
transform 1 0 1380 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1606120353
transform 1 0 2484 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 3956 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 3588 0 -1 2720
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1606120353
transform 1 0 4048 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1606120353
transform 1 0 5152 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1606120353
transform 1 0 3588 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1606120353
transform 1 0 4692 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1606120353
transform 1 0 6808 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1606120353
transform 1 0 6716 0 1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 6256 0 -1 2720
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1606120353
transform 1 0 6900 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 5796 0 1 2720
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 6532 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1606120353
transform 1 0 6808 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1606120353
transform 1 0 8004 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1606120353
transform 1 0 9108 0 -1 2720
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1606120353
transform 1 0 7912 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_1_86
timestamp 1606120353
transform 1 0 9016 0 1 2720
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_1_92 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 9568 0 1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_0_94
timestamp 1606120353
transform 1 0 9752 0 -1 2720
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__D /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 9660 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1606120353
transform 1 0 9660 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_0_107
timestamp 1606120353
transform 1 0 10948 0 -1 2720
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_0_103
timestamp 1606120353
transform 1 0 10580 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_0_100
timestamp 1606120353
transform 1 0 10304 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__CLK
timestamp 1606120353
transform 1 0 10764 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__D
timestamp 1606120353
transform 1 0 10396 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1125_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 9844 0 1 2720
box 0 -48 1748 592
use sky130_fd_sc_hd__dfxtp_4  _1143_
timestamp 1606120353
transform 1 0 12604 0 -1 2720
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1606120353
transform 1 0 12512 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1606120353
transform 1 0 12328 0 1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__D
timestamp 1606120353
transform 1 0 12328 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__CLK
timestamp 1606120353
transform 1 0 11960 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_0_115
timestamp 1606120353
transform 1 0 11684 0 -1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1606120353
transform 1 0 12144 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_1_114
timestamp 1606120353
transform 1 0 11592 0 1 2720
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1606120353
transform 1 0 12420 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_0_144
timestamp 1606120353
transform 1 0 14352 0 -1 2720
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_0_152
timestamp 1606120353
transform 1 0 15088 0 -1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1606120353
transform 1 0 13524 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1606120353
transform 1 0 14628 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1606120353
transform 1 0 15364 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1606120353
transform 1 0 15456 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1606120353
transform 1 0 16560 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1606120353
transform 1 0 15732 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1606120353
transform 1 0 16836 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_1_184
timestamp 1606120353
transform 1 0 18032 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_0_182
timestamp 1606120353
transform 1 0 17848 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__CLK
timestamp 1606120353
transform 1 0 17664 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__D
timestamp 1606120353
transform 1 0 18216 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__D
timestamp 1606120353
transform 1 0 18032 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1606120353
transform 1 0 17940 0 1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1606120353
transform 1 0 18216 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_1_188
timestamp 1606120353
transform 1 0 18400 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__CLK
timestamp 1606120353
transform 1 0 18584 0 1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_1_192
timestamp 1606120353
transform 1 0 18768 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1215_
timestamp 1606120353
transform 1 0 18308 0 -1 2720
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1606120353
transform 1 0 21068 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__D
timestamp 1606120353
transform 1 0 20884 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__CLK
timestamp 1606120353
transform 1 0 20516 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_0_206
timestamp 1606120353
transform 1 0 20056 0 -1 2720
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_0_210
timestamp 1606120353
transform 1 0 20424 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_0_213
timestamp 1606120353
transform 1 0 20700 0 -1 2720
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_0_218
timestamp 1606120353
transform 1 0 21160 0 -1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_1_204
timestamp 1606120353
transform 1 0 19872 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_1_216
timestamp 1606120353
transform 1 0 20976 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1204_
timestamp 1606120353
transform 1 0 21436 0 -1 2720
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_8  FILLER_0_240
timestamp 1606120353
transform 1 0 23184 0 -1 2720
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_1_228
timestamp 1606120353
transform 1 0 22080 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_1_240
timestamp 1606120353
transform 1 0 23184 0 1 2720
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1606120353
transform 1 0 23920 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1606120353
transform 1 0 23552 0 1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_0_249
timestamp 1606120353
transform 1 0 24012 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_0_261
timestamp 1606120353
transform 1 0 25116 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245
timestamp 1606120353
transform 1 0 23644 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_1_257
timestamp 1606120353
transform 1 0 24748 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1606120353
transform 1 0 26772 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1606120353
transform 1 0 26220 0 -1 2720
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_0_280
timestamp 1606120353
transform 1 0 26864 0 -1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_1_269
timestamp 1606120353
transform 1 0 25852 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1606120353
transform 1 0 26956 0 1 2720
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606120353
transform -1 0 28888 0 -1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606120353
transform -1 0 28888 0 1 2720
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_0_292
timestamp 1606120353
transform 1 0 27968 0 -1 2720
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_0_298
timestamp 1606120353
transform 1 0 28520 0 -1 2720
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_1_293
timestamp 1606120353
transform 1 0 28060 0 1 2720
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606120353
transform 1 0 1104 0 -1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1606120353
transform 1 0 1380 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1606120353
transform 1 0 2484 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1606120353
transform 1 0 3956 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1606120353
transform 1 0 3588 0 -1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1606120353
transform 1 0 4048 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1606120353
transform 1 0 5152 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1606120353
transform 1 0 6256 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1606120353
transform 1 0 7360 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1606120353
transform 1 0 8464 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1119_
timestamp 1606120353
transform 1 0 10396 0 -1 3808
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1606120353
transform 1 0 9568 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__CLK
timestamp 1606120353
transform 1 0 9844 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_2_93
timestamp 1606120353
transform 1 0 9660 0 -1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_2_97
timestamp 1606120353
transform 1 0 10028 0 -1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_2_120
timestamp 1606120353
transform 1 0 12144 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_132
timestamp 1606120353
transform 1 0 13248 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1606120353
transform 1 0 15180 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_2_144
timestamp 1606120353
transform 1 0 14352 0 -1 3808
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_2_152
timestamp 1606120353
transform 1 0 15088 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1606120353
transform 1 0 15272 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1606120353
transform 1 0 16376 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1227_
timestamp 1606120353
transform 1 0 17848 0 -1 3808
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_4  FILLER_2_178
timestamp 1606120353
transform 1 0 17480 0 -1 3808
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1606120353
transform 1 0 20792 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_2_201
timestamp 1606120353
transform 1 0 19596 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_2_213
timestamp 1606120353
transform 1 0 20700 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1606120353
transform 1 0 20884 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1606120353
transform 1 0 21988 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1606120353
transform 1 0 23092 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_251
timestamp 1606120353
transform 1 0 24196 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_2_263
timestamp 1606120353
transform 1 0 25300 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1606120353
transform 1 0 26404 0 -1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_2_276
timestamp 1606120353
transform 1 0 26496 0 -1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606120353
transform -1 0 28888 0 -1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_2_288
timestamp 1606120353
transform 1 0 27600 0 -1 3808
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_2_296
timestamp 1606120353
transform 1 0 28336 0 -1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606120353
transform 1 0 1104 0 1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1606120353
transform 1 0 1380 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1606120353
transform 1 0 2484 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1606120353
transform 1 0 3588 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1606120353
transform 1 0 4692 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1606120353
transform 1 0 6716 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1606120353
transform 1 0 5796 0 1 3808
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1606120353
transform 1 0 6532 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1606120353
transform 1 0 6808 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1606120353
transform 1 0 7912 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1606120353
transform 1 0 9016 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__D
timestamp 1606120353
transform 1 0 10948 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_3_98
timestamp 1606120353
transform 1 0 10120 0 1 3808
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_3_106
timestamp 1606120353
transform 1 0 10856 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_3_109
timestamp 1606120353
transform 1 0 11132 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1606120353
transform 1 0 12328 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__CLK
timestamp 1606120353
transform 1 0 11316 0 1 3808
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_3_113
timestamp 1606120353
transform 1 0 11500 0 1 3808
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_3_121
timestamp 1606120353
transform 1 0 12236 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1606120353
transform 1 0 12420 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1606120353
transform 1 0 13524 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1606120353
transform 1 0 14628 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1606120353
transform 1 0 15732 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1606120353
transform 1 0 16836 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1606120353
transform 1 0 17940 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1606120353
transform 1 0 18032 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1606120353
transform 1 0 19136 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1606120353
transform 1 0 20240 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_220
timestamp 1606120353
transform 1 0 21344 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_232
timestamp 1606120353
transform 1 0 22448 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1606120353
transform 1 0 23552 0 1 3808
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1606120353
transform 1 0 23644 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1606120353
transform 1 0 24748 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_269
timestamp 1606120353
transform 1 0 25852 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1606120353
transform 1 0 26956 0 1 3808
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606120353
transform -1 0 28888 0 1 3808
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_3_293
timestamp 1606120353
transform 1 0 28060 0 1 3808
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606120353
transform 1 0 1104 0 -1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1606120353
transform 1 0 1380 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1606120353
transform 1 0 2484 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1606120353
transform 1 0 3956 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1606120353
transform 1 0 3588 0 -1 4896
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1606120353
transform 1 0 4048 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1606120353
transform 1 0 5152 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1606120353
transform 1 0 6256 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1606120353
transform 1 0 7360 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1606120353
transform 1 0 8464 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1131_
timestamp 1606120353
transform 1 0 10948 0 -1 4896
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1606120353
transform 1 0 9568 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1606120353
transform 1 0 9660 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_4_105
timestamp 1606120353
transform 1 0 10764 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__B1
timestamp 1606120353
transform 1 0 13156 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_4_126
timestamp 1606120353
transform 1 0 12696 0 -1 4896
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_4_130
timestamp 1606120353
transform 1 0 13064 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1606120353
transform 1 0 15180 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__B2
timestamp 1606120353
transform 1 0 13524 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__A2
timestamp 1606120353
transform 1 0 13892 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_4_133
timestamp 1606120353
transform 1 0 13340 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_4_137
timestamp 1606120353
transform 1 0 13708 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1606120353
transform 1 0 14076 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_4_154
timestamp 1606120353
transform 1 0 15272 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__A2
timestamp 1606120353
transform 1 0 15456 0 -1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_4_158
timestamp 1606120353
transform 1 0 15640 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_170
timestamp 1606120353
transform 1 0 16744 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_182
timestamp 1606120353
transform 1 0 17848 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_194
timestamp 1606120353
transform 1 0 18952 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1606120353
transform 1 0 20792 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_4_206
timestamp 1606120353
transform 1 0 20056 0 -1 4896
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1606120353
transform 1 0 20884 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1606120353
transform 1 0 21988 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_239
timestamp 1606120353
transform 1 0 23092 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_251
timestamp 1606120353
transform 1 0 24196 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_4_263
timestamp 1606120353
transform 1 0 25300 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1606120353
transform 1 0 26404 0 -1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_4_276
timestamp 1606120353
transform 1 0 26496 0 -1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606120353
transform -1 0 28888 0 -1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_4_288
timestamp 1606120353
transform 1 0 27600 0 -1 4896
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_4_296
timestamp 1606120353
transform 1 0 28336 0 -1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606120353
transform 1 0 1104 0 1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1606120353
transform 1 0 1380 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1606120353
transform 1 0 2484 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1606120353
transform 1 0 3588 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1606120353
transform 1 0 4692 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1606120353
transform 1 0 6716 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1606120353
transform 1 0 5796 0 1 4896
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1606120353
transform 1 0 6532 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1606120353
transform 1 0 6808 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1606120353
transform 1 0 7912 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1606120353
transform 1 0 9016 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1606120353
transform 1 0 10120 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_5_110
timestamp 1606120353
transform 1 0 11224 0 1 4896
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1096_
timestamp 1606120353
transform 1 0 13064 0 1 4896
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1606120353
transform 1 0 12328 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__A1
timestamp 1606120353
transform 1 0 12880 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__D
timestamp 1606120353
transform 1 0 12144 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_5_118
timestamp 1606120353
transform 1 0 11960 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_5_123
timestamp 1606120353
transform 1 0 12420 0 1 4896
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_5_127
timestamp 1606120353
transform 1 0 12788 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__A1
timestamp 1606120353
transform 1 0 15272 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_5_149
timestamp 1606120353
transform 1 0 14812 0 1 4896
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_5_153
timestamp 1606120353
transform 1 0 15180 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__B1
timestamp 1606120353
transform 1 0 15640 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__B2
timestamp 1606120353
transform 1 0 16008 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_5_156
timestamp 1606120353
transform 1 0 15456 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_5_160
timestamp 1606120353
transform 1 0 15824 0 1 4896
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_5_164
timestamp 1606120353
transform 1 0 16192 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_5_176
timestamp 1606120353
transform 1 0 17296 0 1 4896
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1606120353
transform 1 0 17940 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_5_182
timestamp 1606120353
transform 1 0 17848 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1606120353
transform 1 0 18032 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1606120353
transform 1 0 19136 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1606120353
transform 1 0 20240 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_220
timestamp 1606120353
transform 1 0 21344 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_232
timestamp 1606120353
transform 1 0 22448 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1606120353
transform 1 0 23552 0 1 4896
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1606120353
transform 1 0 23644 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_257
timestamp 1606120353
transform 1 0 24748 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_269
timestamp 1606120353
transform 1 0 25852 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1606120353
transform 1 0 26956 0 1 4896
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606120353
transform -1 0 28888 0 1 4896
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_5_293
timestamp 1606120353
transform 1 0 28060 0 1 4896
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606120353
transform 1 0 1104 0 -1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606120353
transform 1 0 1104 0 1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1606120353
transform 1 0 1380 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1606120353
transform 1 0 2484 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1606120353
transform 1 0 1380 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1606120353
transform 1 0 2484 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1606120353
transform 1 0 3956 0 -1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1606120353
transform 1 0 3588 0 -1 5984
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1606120353
transform 1 0 4048 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1606120353
transform 1 0 5152 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1606120353
transform 1 0 3588 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1606120353
transform 1 0 4692 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1606120353
transform 1 0 6716 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1606120353
transform 1 0 6256 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1606120353
transform 1 0 5796 0 1 5984
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1606120353
transform 1 0 6532 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1606120353
transform 1 0 6808 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1606120353
transform 1 0 7360 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1606120353
transform 1 0 8464 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1606120353
transform 1 0 7912 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1606120353
transform 1 0 9016 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1606120353
transform 1 0 9568 0 -1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1606120353
transform 1 0 9660 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1606120353
transform 1 0 10764 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1606120353
transform 1 0 10120 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1606120353
transform 1 0 11224 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__o22a_4  _0794_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 13156 0 -1 5984
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1606120353
transform 1 0 12328 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__CLK
timestamp 1606120353
transform 1 0 12972 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1606120353
transform 1 0 11868 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1606120353
transform 1 0 12420 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__o22a_4  _0796_
timestamp 1606120353
transform 1 0 15272 0 -1 5984
box 0 -48 1288 592
use sky130_fd_sc_hd__dfxtp_4  _1097_
timestamp 1606120353
transform 1 0 14536 0 1 5984
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1606120353
transform 1 0 15180 0 -1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__D
timestamp 1606120353
transform 1 0 14352 0 1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_6_145
timestamp 1606120353
transform 1 0 14444 0 -1 5984
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_7_135
timestamp 1606120353
transform 1 0 13524 0 1 5984
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_7_143
timestamp 1606120353
transform 1 0 14260 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_6_168
timestamp 1606120353
transform 1 0 16560 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_165
timestamp 1606120353
transform 1 0 16284 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1606120353
transform 1 0 17940 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_6_180
timestamp 1606120353
transform 1 0 17664 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_6_192
timestamp 1606120353
transform 1 0 18768 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_7_177
timestamp 1606120353
transform 1 0 17388 0 1 5984
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1606120353
transform 1 0 18032 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1606120353
transform 1 0 19136 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1606120353
transform 1 0 20792 0 -1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_6_204
timestamp 1606120353
transform 1 0 19872 0 -1 5984
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_6_212
timestamp 1606120353
transform 1 0 20608 0 -1 5984
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1606120353
transform 1 0 20884 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1606120353
transform 1 0 20240 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_220
timestamp 1606120353
transform 1 0 21344 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1606120353
transform 1 0 21988 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_6_239
timestamp 1606120353
transform 1 0 23092 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_232
timestamp 1606120353
transform 1 0 22448 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1606120353
transform 1 0 23552 0 1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_6_251
timestamp 1606120353
transform 1 0 24196 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_6_263
timestamp 1606120353
transform 1 0 25300 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1606120353
transform 1 0 23644 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1606120353
transform 1 0 24748 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1606120353
transform 1 0 26404 0 -1 5984
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_6_276
timestamp 1606120353
transform 1 0 26496 0 -1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_269
timestamp 1606120353
transform 1 0 25852 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1606120353
transform 1 0 26956 0 1 5984
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606120353
transform -1 0 28888 0 -1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606120353
transform -1 0 28888 0 1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_6_288
timestamp 1606120353
transform 1 0 27600 0 -1 5984
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_6_296
timestamp 1606120353
transform 1 0 28336 0 -1 5984
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_7_293
timestamp 1606120353
transform 1 0 28060 0 1 5984
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606120353
transform 1 0 1104 0 -1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1606120353
transform 1 0 1380 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1606120353
transform 1 0 2484 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1606120353
transform 1 0 3956 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1606120353
transform 1 0 3588 0 -1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1606120353
transform 1 0 4048 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1606120353
transform 1 0 5152 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1606120353
transform 1 0 6256 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1606120353
transform 1 0 7360 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1606120353
transform 1 0 8464 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1606120353
transform 1 0 9568 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1606120353
transform 1 0 9660 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1606120353
transform 1 0 10764 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__CLK
timestamp 1606120353
transform 1 0 13064 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1606120353
transform 1 0 11868 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_8_129
timestamp 1606120353
transform 1 0 12972 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_8_132
timestamp 1606120353
transform 1 0 13248 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1606120353
transform 1 0 15180 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__CLK
timestamp 1606120353
transform 1 0 14536 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_8_144
timestamp 1606120353
transform 1 0 14352 0 -1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_8_148
timestamp 1606120353
transform 1 0 14720 0 -1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_8_152
timestamp 1606120353
transform 1 0 15088 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1606120353
transform 1 0 15272 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1606120353
transform 1 0 16376 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1606120353
transform 1 0 17480 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_190
timestamp 1606120353
transform 1 0 18584 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1606120353
transform 1 0 20792 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_8_202
timestamp 1606120353
transform 1 0 19688 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1606120353
transform 1 0 20884 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_227
timestamp 1606120353
transform 1 0 21988 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_239
timestamp 1606120353
transform 1 0 23092 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_251
timestamp 1606120353
transform 1 0 24196 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_8_263
timestamp 1606120353
transform 1 0 25300 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1606120353
transform 1 0 26404 0 -1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_8_276
timestamp 1606120353
transform 1 0 26496 0 -1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606120353
transform -1 0 28888 0 -1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_8_288
timestamp 1606120353
transform 1 0 27600 0 -1 7072
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_8_296
timestamp 1606120353
transform 1 0 28336 0 -1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606120353
transform 1 0 1104 0 1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1606120353
transform 1 0 1380 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1606120353
transform 1 0 2484 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1606120353
transform 1 0 3588 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1606120353
transform 1 0 4692 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1606120353
transform 1 0 6716 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1606120353
transform 1 0 5796 0 1 7072
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1606120353
transform 1 0 6532 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1606120353
transform 1 0 6808 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1606120353
transform 1 0 7912 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_9_86
timestamp 1606120353
transform 1 0 9016 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__D
timestamp 1606120353
transform 1 0 11040 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_9_98
timestamp 1606120353
transform 1 0 10120 0 1 7072
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_9_106
timestamp 1606120353
transform 1 0 10856 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_9_110
timestamp 1606120353
transform 1 0 11224 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1094_
timestamp 1606120353
transform 1 0 13064 0 1 7072
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1606120353
transform 1 0 12328 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__D
timestamp 1606120353
transform 1 0 12880 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__CLK
timestamp 1606120353
transform 1 0 11408 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_9_114
timestamp 1606120353
transform 1 0 11592 0 1 7072
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_9_123
timestamp 1606120353
transform 1 0 12420 0 1 7072
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_9_127
timestamp 1606120353
transform 1 0 12788 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1606120353
transform 1 0 14812 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__D
timestamp 1606120353
transform 1 0 16560 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__CLK
timestamp 1606120353
transform 1 0 16928 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1606120353
transform 1 0 15916 0 1 7072
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1606120353
transform 1 0 16468 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_9_170
timestamp 1606120353
transform 1 0 16744 0 1 7072
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_9_174
timestamp 1606120353
transform 1 0 17112 0 1 7072
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1606120353
transform 1 0 17940 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_9_182
timestamp 1606120353
transform 1 0 17848 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1606120353
transform 1 0 18032 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1606120353
transform 1 0 19136 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1606120353
transform 1 0 20240 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_9_220
timestamp 1606120353
transform 1 0 21344 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_9_232
timestamp 1606120353
transform 1 0 22448 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1606120353
transform 1 0 23552 0 1 7072
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1606120353
transform 1 0 23644 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1606120353
transform 1 0 24748 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_9_269
timestamp 1606120353
transform 1 0 25852 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1606120353
transform 1 0 26956 0 1 7072
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606120353
transform -1 0 28888 0 1 7072
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_9_293
timestamp 1606120353
transform 1 0 28060 0 1 7072
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606120353
transform 1 0 1104 0 -1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1606120353
transform 1 0 1380 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1606120353
transform 1 0 2484 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1606120353
transform 1 0 3956 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1606120353
transform 1 0 3588 0 -1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1606120353
transform 1 0 4048 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1606120353
transform 1 0 5152 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1606120353
transform 1 0 6256 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__B1
timestamp 1606120353
transform 1 0 9016 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1606120353
transform 1 0 7360 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_10_80
timestamp 1606120353
transform 1 0 8464 0 -1 8160
box 0 -48 552 592
use sky130_fd_sc_hd__decap_4  FILLER_10_88
timestamp 1606120353
transform 1 0 9200 0 -1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1083_
timestamp 1606120353
transform 1 0 11040 0 -1 8160
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1606120353
transform 1 0 9568 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__CLK
timestamp 1606120353
transform 1 0 9844 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_10_93
timestamp 1606120353
transform 1 0 9660 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_10_97
timestamp 1606120353
transform 1 0 10028 0 -1 8160
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_10_105
timestamp 1606120353
transform 1 0 10764 0 -1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_10_127
timestamp 1606120353
transform 1 0 12788 0 -1 8160
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1606120353
transform 1 0 15180 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__B1
timestamp 1606120353
transform 1 0 13432 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__A2
timestamp 1606120353
transform 1 0 13800 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_10_133
timestamp 1606120353
transform 1 0 13340 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_10_136
timestamp 1606120353
transform 1 0 13616 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_10_140
timestamp 1606120353
transform 1 0 13984 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_10_152
timestamp 1606120353
transform 1 0 15088 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1606120353
transform 1 0 15272 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1210_
timestamp 1606120353
transform 1 0 16560 0 -1 8160
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_2  FILLER_10_166
timestamp 1606120353
transform 1 0 16376 0 -1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_10_187
timestamp 1606120353
transform 1 0 18308 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1606120353
transform 1 0 20792 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_10_199
timestamp 1606120353
transform 1 0 19412 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_10_211
timestamp 1606120353
transform 1 0 20516 0 -1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1606120353
transform 1 0 20884 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1606120353
transform 1 0 21988 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1606120353
transform 1 0 23092 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_10_251
timestamp 1606120353
transform 1 0 24196 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_10_263
timestamp 1606120353
transform 1 0 25300 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1606120353
transform 1 0 26404 0 -1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_10_276
timestamp 1606120353
transform 1 0 26496 0 -1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606120353
transform -1 0 28888 0 -1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_10_288
timestamp 1606120353
transform 1 0 27600 0 -1 8160
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_10_296
timestamp 1606120353
transform 1 0 28336 0 -1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606120353
transform 1 0 1104 0 1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__D
timestamp 1606120353
transform 1 0 1564 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__CLK
timestamp 1606120353
transform 1 0 1932 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_3
timestamp 1606120353
transform 1 0 1380 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_7
timestamp 1606120353
transform 1 0 1748 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_11_11
timestamp 1606120353
transform 1 0 2116 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_11_23
timestamp 1606120353
transform 1 0 3220 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_11_35
timestamp 1606120353
transform 1 0 4324 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1606120353
transform 1 0 6716 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_11_47
timestamp 1606120353
transform 1 0 5428 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1606120353
transform 1 0 6532 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1606120353
transform 1 0 6808 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__o22a_4  _0786_
timestamp 1606120353
transform 1 0 9016 0 1 8160
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__A1
timestamp 1606120353
transform 1 0 8832 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__A2
timestamp 1606120353
transform 1 0 8464 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_11_74
timestamp 1606120353
transform 1 0 7912 0 1 8160
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_11_82
timestamp 1606120353
transform 1 0 8648 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__D
timestamp 1606120353
transform 1 0 10488 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_100
timestamp 1606120353
transform 1 0 10304 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_11_104
timestamp 1606120353
transform 1 0 10672 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1606120353
transform 1 0 12328 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__A1
timestamp 1606120353
transform 1 0 12144 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__B1
timestamp 1606120353
transform 1 0 12604 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__A1
timestamp 1606120353
transform 1 0 13248 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__A2
timestamp 1606120353
transform 1 0 11776 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_118
timestamp 1606120353
transform 1 0 11960 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_123
timestamp 1606120353
transform 1 0 12420 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_11_127
timestamp 1606120353
transform 1 0 12788 0 1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_11_131
timestamp 1606120353
transform 1 0 13156 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _0789_
timestamp 1606120353
transform 1 0 13432 0 1 8160
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILLER_11_148
timestamp 1606120353
transform 1 0 14720 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__A1
timestamp 1606120353
transform 1 0 16192 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__B1
timestamp 1606120353
transform 1 0 16560 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__A2
timestamp 1606120353
transform 1 0 16928 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_11_160
timestamp 1606120353
transform 1 0 15824 0 1 8160
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_11_166
timestamp 1606120353
transform 1 0 16376 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_11_170
timestamp 1606120353
transform 1 0 16744 0 1 8160
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_11_174
timestamp 1606120353
transform 1 0 17112 0 1 8160
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1606120353
transform 1 0 17940 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_11_182
timestamp 1606120353
transform 1 0 17848 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1606120353
transform 1 0 18032 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1606120353
transform 1 0 19136 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1606120353
transform 1 0 20240 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_11_220
timestamp 1606120353
transform 1 0 21344 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_11_232
timestamp 1606120353
transform 1 0 22448 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1606120353
transform 1 0 23552 0 1 8160
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_11_245
timestamp 1606120353
transform 1 0 23644 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_11_257
timestamp 1606120353
transform 1 0 24748 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_11_269
timestamp 1606120353
transform 1 0 25852 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1606120353
transform 1 0 26956 0 1 8160
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606120353
transform -1 0 28888 0 1 8160
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_11_293
timestamp 1606120353
transform 1 0 28060 0 1 8160
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1218_
timestamp 1606120353
transform 1 0 1380 0 -1 9248
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606120353
transform 1 0 1104 0 -1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_12_22
timestamp 1606120353
transform 1 0 3128 0 -1 9248
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1606120353
transform 1 0 3956 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_12_30
timestamp 1606120353
transform 1 0 3864 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1606120353
transform 1 0 4048 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1606120353
transform 1 0 5152 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1606120353
transform 1 0 6256 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__B2
timestamp 1606120353
transform 1 0 9016 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1606120353
transform 1 0 7360 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_12_80
timestamp 1606120353
transform 1 0 8464 0 -1 9248
box 0 -48 552 592
use sky130_fd_sc_hd__decap_4  FILLER_12_88
timestamp 1606120353
transform 1 0 9200 0 -1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1093_
timestamp 1606120353
transform 1 0 9660 0 -1 9248
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1606120353
transform 1 0 9568 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__a21o_4  _0666_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 12144 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_12_112
timestamp 1606120353
transform 1 0 11408 0 -1 9248
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_12_132
timestamp 1606120353
transform 1 0 13248 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1606120353
transform 1 0 15180 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__B2
timestamp 1606120353
transform 1 0 13432 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_12_136
timestamp 1606120353
transform 1 0 13616 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_12_148
timestamp 1606120353
transform 1 0 14720 0 -1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1606120353
transform 1 0 15088 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_12_154
timestamp 1606120353
transform 1 0 15272 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0715_
timestamp 1606120353
transform 1 0 16192 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__CLK
timestamp 1606120353
transform 1 0 15456 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_12_158
timestamp 1606120353
transform 1 0 15640 0 -1 9248
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_12_176
timestamp 1606120353
transform 1 0 17296 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_12_188
timestamp 1606120353
transform 1 0 18400 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1606120353
transform 1 0 20792 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_12_200
timestamp 1606120353
transform 1 0 19504 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_12_212
timestamp 1606120353
transform 1 0 20608 0 -1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1606120353
transform 1 0 20884 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1606120353
transform 1 0 21988 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1606120353
transform 1 0 23092 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_12_251
timestamp 1606120353
transform 1 0 24196 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_12_263
timestamp 1606120353
transform 1 0 25300 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1606120353
transform 1 0 26404 0 -1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_12_276
timestamp 1606120353
transform 1 0 26496 0 -1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606120353
transform -1 0 28888 0 -1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_12_288
timestamp 1606120353
transform 1 0 27600 0 -1 9248
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_12_296
timestamp 1606120353
transform 1 0 28336 0 -1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606120353
transform 1 0 1104 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606120353
transform 1 0 1104 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1606120353
transform 1 0 1380 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1606120353
transform 1 0 2484 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1606120353
transform 1 0 1380 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1606120353
transform 1 0 2484 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1606120353
transform 1 0 3956 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1606120353
transform 1 0 3588 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1606120353
transform 1 0 4692 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1606120353
transform 1 0 3588 0 -1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1606120353
transform 1 0 4048 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1606120353
transform 1 0 5152 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1606120353
transform 1 0 6716 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1606120353
transform 1 0 5796 0 1 9248
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1606120353
transform 1 0 6532 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1606120353
transform 1 0 6808 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1606120353
transform 1 0 6256 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_13_74
timestamp 1606120353
transform 1 0 7912 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_13_86
timestamp 1606120353
transform 1 0 9016 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1606120353
transform 1 0 7360 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1606120353
transform 1 0 8464 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1606120353
transform 1 0 9568 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_13_98
timestamp 1606120353
transform 1 0 10120 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_13_110
timestamp 1606120353
transform 1 0 11224 0 1 9248
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1606120353
transform 1 0 9660 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_14_105
timestamp 1606120353
transform 1 0 10764 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__and2_4  _0665_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 12512 0 1 9248
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1606120353
transform 1 0 12328 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0665__A
timestamp 1606120353
transform 1 0 12144 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_118
timestamp 1606120353
transform 1 0 11960 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_13_123
timestamp 1606120353
transform 1 0 12420 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_13_131
timestamp 1606120353
transform 1 0 13156 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_14_117
timestamp 1606120353
transform 1 0 11868 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_14_129
timestamp 1606120353
transform 1 0 12972 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_13_142
timestamp 1606120353
transform 1 0 14168 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_13_135
timestamp 1606120353
transform 1 0 13524 0 1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0665__B
timestamp 1606120353
transform 1 0 13340 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0779_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 13892 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_14_154
timestamp 1606120353
transform 1 0 15272 0 -1 10336
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_13_150
timestamp 1606120353
transform 1 0 14904 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_13_146
timestamp 1606120353
transform 1 0 14536 0 1 9248
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__D
timestamp 1606120353
transform 1 0 14996 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__A
timestamp 1606120353
transform 1 0 14352 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1606120353
transform 1 0 15180 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1606120353
transform 1 0 14076 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1084_
timestamp 1606120353
transform 1 0 15180 0 1 9248
box 0 -48 1748 592
use sky130_fd_sc_hd__and2_4  _0714_
timestamp 1606120353
transform 1 0 16284 0 -1 10336
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__A
timestamp 1606120353
transform 1 0 17112 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_172
timestamp 1606120353
transform 1 0 16928 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_13_176
timestamp 1606120353
transform 1 0 17296 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_14_162
timestamp 1606120353
transform 1 0 16008 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_14_172
timestamp 1606120353
transform 1 0 16928 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_14_184
timestamp 1606120353
transform 1 0 18032 0 -1 10336
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_13_184
timestamp 1606120353
transform 1 0 18032 0 1 9248
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_13_180
timestamp 1606120353
transform 1 0 17664 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__B
timestamp 1606120353
transform 1 0 17480 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1606120353
transform 1 0 17940 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_14_195
timestamp 1606120353
transform 1 0 19044 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__CLK
timestamp 1606120353
transform 1 0 19228 0 -1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_clk_A
timestamp 1606120353
transform 1 0 18768 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_clk /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 18768 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_13_194
timestamp 1606120353
transform 1 0 18952 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1606120353
transform 1 0 20792 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_13_206
timestamp 1606120353
transform 1 0 20056 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_13_218
timestamp 1606120353
transform 1 0 21160 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_14_199
timestamp 1606120353
transform 1 0 19412 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_14_211
timestamp 1606120353
transform 1 0 20516 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_14_215
timestamp 1606120353
transform 1 0 20884 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_13_230
timestamp 1606120353
transform 1 0 22264 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_13_242
timestamp 1606120353
transform 1 0 23368 0 1 9248
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_14_227
timestamp 1606120353
transform 1 0 21988 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_14_239
timestamp 1606120353
transform 1 0 23092 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1606120353
transform 1 0 23552 0 1 9248
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_13_245
timestamp 1606120353
transform 1 0 23644 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_13_257
timestamp 1606120353
transform 1 0 24748 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_14_251
timestamp 1606120353
transform 1 0 24196 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_14_263
timestamp 1606120353
transform 1 0 25300 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1606120353
transform 1 0 26404 0 -1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_13_269
timestamp 1606120353
transform 1 0 25852 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1606120353
transform 1 0 26956 0 1 9248
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_14_276
timestamp 1606120353
transform 1 0 26496 0 -1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606120353
transform -1 0 28888 0 1 9248
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606120353
transform -1 0 28888 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_13_293
timestamp 1606120353
transform 1 0 28060 0 1 9248
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILLER_14_288
timestamp 1606120353
transform 1 0 27600 0 -1 10336
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_14_296
timestamp 1606120353
transform 1 0 28336 0 -1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606120353
transform 1 0 1104 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1606120353
transform 1 0 1380 0 1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1606120353
transform 1 0 2484 0 1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1606120353
transform 1 0 3588 0 1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1606120353
transform 1 0 4692 0 1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1606120353
transform 1 0 6716 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1606120353
transform 1 0 5796 0 1 10336
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1606120353
transform 1 0 6532 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_15_62
timestamp 1606120353
transform 1 0 6808 0 1 10336
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_clk_A
timestamp 1606120353
transform 1 0 7820 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_15_70
timestamp 1606120353
transform 1 0 7544 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_15_75
timestamp 1606120353
transform 1 0 8004 0 1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_15_87
timestamp 1606120353
transform 1 0 9108 0 1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__B
timestamp 1606120353
transform 1 0 10764 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__A
timestamp 1606120353
transform 1 0 11132 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_15_99
timestamp 1606120353
transform 1 0 10212 0 1 10336
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_15_107
timestamp 1606120353
transform 1 0 10948 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1606120353
transform 1 0 12328 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__A1_N
timestamp 1606120353
transform 1 0 12972 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__B1
timestamp 1606120353
transform 1 0 12604 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_15_111
timestamp 1606120353
transform 1 0 11316 0 1 10336
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_15_119
timestamp 1606120353
transform 1 0 12052 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_15_123
timestamp 1606120353
transform 1 0 12420 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_127
timestamp 1606120353
transform 1 0 12788 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_131
timestamp 1606120353
transform 1 0 13156 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__B2
timestamp 1606120353
transform 1 0 13340 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__A2_N
timestamp 1606120353
transform 1 0 13708 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__D
timestamp 1606120353
transform 1 0 15272 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_135
timestamp 1606120353
transform 1 0 13524 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_15_139
timestamp 1606120353
transform 1 0 13892 0 1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_15_151
timestamp 1606120353
transform 1 0 14996 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__CLK
timestamp 1606120353
transform 1 0 15640 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_15_156
timestamp 1606120353
transform 1 0 15456 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_15_160
timestamp 1606120353
transform 1 0 15824 0 1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_15_172
timestamp 1606120353
transform 1 0 16928 0 1 10336
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1167_
timestamp 1606120353
transform 1 0 19228 0 1 10336
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1606120353
transform 1 0 17940 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__D
timestamp 1606120353
transform 1 0 19044 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_clk_A
timestamp 1606120353
transform 1 0 17756 0 1 10336
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_15_180
timestamp 1606120353
transform 1 0 17664 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_15_184
timestamp 1606120353
transform 1 0 18032 0 1 10336
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_15_192
timestamp 1606120353
transform 1 0 18768 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_15_216
timestamp 1606120353
transform 1 0 20976 0 1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_15_228
timestamp 1606120353
transform 1 0 22080 0 1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_15_240
timestamp 1606120353
transform 1 0 23184 0 1 10336
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1606120353
transform 1 0 23552 0 1 10336
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_15_245
timestamp 1606120353
transform 1 0 23644 0 1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_15_257
timestamp 1606120353
transform 1 0 24748 0 1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_15_269
timestamp 1606120353
transform 1 0 25852 0 1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1606120353
transform 1 0 26956 0 1 10336
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606120353
transform -1 0 28888 0 1 10336
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_15_293
timestamp 1606120353
transform 1 0 28060 0 1 10336
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606120353
transform 1 0 1104 0 -1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1606120353
transform 1 0 1380 0 -1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1606120353
transform 1 0 2484 0 -1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1606120353
transform 1 0 3956 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1606120353
transform 1 0 3588 0 -1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1606120353
transform 1 0 4048 0 -1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1606120353
transform 1 0 5152 0 -1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1606120353
transform 1 0 6256 0 -1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_clk
timestamp 1606120353
transform 1 0 7820 0 -1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_16_68
timestamp 1606120353
transform 1 0 7360 0 -1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_16_72
timestamp 1606120353
transform 1 0 7728 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_16_76
timestamp 1606120353
transform 1 0 8096 0 -1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_16_88
timestamp 1606120353
transform 1 0 9200 0 -1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__and2_4  _0783_
timestamp 1606120353
transform 1 0 10764 0 -1 11424
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1606120353
transform 1 0 9568 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__A2
timestamp 1606120353
transform 1 0 10304 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_16_93
timestamp 1606120353
transform 1 0 9660 0 -1 11424
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_16_99
timestamp 1606120353
transform 1 0 10212 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_16_102
timestamp 1606120353
transform 1 0 10488 0 -1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__a2bb2o_4  _0790_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 12972 0 -1 11424
box 0 -48 1472 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__B1
timestamp 1606120353
transform 1 0 12420 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__A2
timestamp 1606120353
transform 1 0 11592 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__A2_N
timestamp 1606120353
transform 1 0 12788 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__B1
timestamp 1606120353
transform 1 0 11960 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_112
timestamp 1606120353
transform 1 0 11408 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_116
timestamp 1606120353
transform 1 0 11776 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_16_120
timestamp 1606120353
transform 1 0 12144 0 -1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_16_125
timestamp 1606120353
transform 1 0 12604 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1095_
timestamp 1606120353
transform 1 0 15272 0 -1 11424
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1606120353
transform 1 0 15180 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__B1
timestamp 1606120353
transform 1 0 14628 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_16_145
timestamp 1606120353
transform 1 0 14444 0 -1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_16_149
timestamp 1606120353
transform 1 0 14812 0 -1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILLER_16_173
timestamp 1606120353
transform 1 0 17020 0 -1 11424
box 0 -48 736 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_clk
timestamp 1606120353
transform 1 0 17756 0 -1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_16_184
timestamp 1606120353
transform 1 0 18032 0 -1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_16_196
timestamp 1606120353
transform 1 0 19136 0 -1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1606120353
transform 1 0 20792 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_16_208
timestamp 1606120353
transform 1 0 20240 0 -1 11424
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1606120353
transform 1 0 20884 0 -1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_16_227
timestamp 1606120353
transform 1 0 21988 0 -1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_16_239
timestamp 1606120353
transform 1 0 23092 0 -1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_16_251
timestamp 1606120353
transform 1 0 24196 0 -1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_16_263
timestamp 1606120353
transform 1 0 25300 0 -1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1606120353
transform 1 0 26404 0 -1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_16_276
timestamp 1606120353
transform 1 0 26496 0 -1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606120353
transform -1 0 28888 0 -1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_16_288
timestamp 1606120353
transform 1 0 27600 0 -1 11424
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_16_296
timestamp 1606120353
transform 1 0 28336 0 -1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606120353
transform 1 0 1104 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1606120353
transform 1 0 1380 0 1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1606120353
transform 1 0 2484 0 1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1606120353
transform 1 0 3588 0 1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1606120353
transform 1 0 4692 0 1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1606120353
transform 1 0 6716 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1606120353
transform 1 0 5796 0 1 11424
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1606120353
transform 1 0 6532 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1606120353
transform 1 0 6808 0 1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0637__A
timestamp 1606120353
transform 1 0 9108 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_17_74
timestamp 1606120353
transform 1 0 7912 0 1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_17_86
timestamp 1606120353
transform 1 0 9016 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0637_
timestamp 1606120353
transform 1 0 9292 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__a21o_4  _0784_
timestamp 1606120353
transform 1 0 10304 0 1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__A1
timestamp 1606120353
transform 1 0 10120 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__A
timestamp 1606120353
transform 1 0 9752 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_92
timestamp 1606120353
transform 1 0 9568 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_96
timestamp 1606120353
transform 1 0 9936 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__a2bb2o_4  _0788_
timestamp 1606120353
transform 1 0 12420 0 1 11424
box 0 -48 1472 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1606120353
transform 1 0 12328 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__A1_N
timestamp 1606120353
transform 1 0 12144 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__A1
timestamp 1606120353
transform 1 0 11592 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_112
timestamp 1606120353
transform 1 0 11408 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_17_116
timestamp 1606120353
transform 1 0 11776 0 1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__o22a_4  _0791_
timestamp 1606120353
transform 1 0 15088 0 1 11424
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__A1_N
timestamp 1606120353
transform 1 0 14076 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__B2
timestamp 1606120353
transform 1 0 14444 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__A1
timestamp 1606120353
transform 1 0 14904 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_139
timestamp 1606120353
transform 1 0 13892 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_143
timestamp 1606120353
transform 1 0 14260 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_17_147
timestamp 1606120353
transform 1 0 14628 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__A2
timestamp 1606120353
transform 1 0 16560 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_clk_A
timestamp 1606120353
transform 1 0 16928 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_166
timestamp 1606120353
transform 1 0 16376 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_17_170
timestamp 1606120353
transform 1 0 16744 0 1 11424
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_17_174
timestamp 1606120353
transform 1 0 17112 0 1 11424
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1606120353
transform 1 0 17940 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_17_182
timestamp 1606120353
transform 1 0 17848 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1606120353
transform 1 0 18032 0 1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1606120353
transform 1 0 19136 0 1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1606120353
transform 1 0 20240 0 1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_17_220
timestamp 1606120353
transform 1 0 21344 0 1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_17_232
timestamp 1606120353
transform 1 0 22448 0 1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1606120353
transform 1 0 23552 0 1 11424
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_17_245
timestamp 1606120353
transform 1 0 23644 0 1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_17_257
timestamp 1606120353
transform 1 0 24748 0 1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_17_269
timestamp 1606120353
transform 1 0 25852 0 1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1606120353
transform 1 0 26956 0 1 11424
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606120353
transform -1 0 28888 0 1 11424
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_17_293
timestamp 1606120353
transform 1 0 28060 0 1 11424
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606120353
transform 1 0 1104 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1606120353
transform 1 0 1380 0 -1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1606120353
transform 1 0 2484 0 -1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1606120353
transform 1 0 3956 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1606120353
transform 1 0 3588 0 -1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1606120353
transform 1 0 4048 0 -1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1606120353
transform 1 0 5152 0 -1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1606120353
transform 1 0 6256 0 -1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__CLK
timestamp 1606120353
transform 1 0 8648 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1606120353
transform 1 0 7360 0 -1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_18_80
timestamp 1606120353
transform 1 0 8464 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_18_84
timestamp 1606120353
transform 1 0 8832 0 -1 12512
box 0 -48 736 592
use sky130_fd_sc_hd__buf_1  _0785_
timestamp 1606120353
transform 1 0 9752 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__a21o_4  _0793_
timestamp 1606120353
transform 1 0 11132 0 -1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1606120353
transform 1 0 9568 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__B1
timestamp 1606120353
transform 1 0 10304 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_18_93
timestamp 1606120353
transform 1 0 9660 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_18_97
timestamp 1606120353
transform 1 0 10028 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_18_102
timestamp 1606120353
transform 1 0 10488 0 -1 12512
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_18_108
timestamp 1606120353
transform 1 0 11040 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__a2bb2o_4  _0795_
timestamp 1606120353
transform 1 0 12972 0 -1 12512
box 0 -48 1472 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__B2
timestamp 1606120353
transform 1 0 12420 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__A2_N
timestamp 1606120353
transform 1 0 12788 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_121
timestamp 1606120353
transform 1 0 12236 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_125
timestamp 1606120353
transform 1 0 12604 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1606120353
transform 1 0 15180 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_18_145
timestamp 1606120353
transform 1 0 14444 0 -1 12512
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_18_154
timestamp 1606120353
transform 1 0 15272 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_clk
timestamp 1606120353
transform 1 0 16008 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__B1
timestamp 1606120353
transform 1 0 15456 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__B2
timestamp 1606120353
transform 1 0 15824 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_18_158
timestamp 1606120353
transform 1 0 15640 0 -1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1606120353
transform 1 0 16284 0 -1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_18_177
timestamp 1606120353
transform 1 0 17388 0 -1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_18_189
timestamp 1606120353
transform 1 0 18492 0 -1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1606120353
transform 1 0 20792 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_18_201
timestamp 1606120353
transform 1 0 19596 0 -1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_18_213
timestamp 1606120353
transform 1 0 20700 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_18_215
timestamp 1606120353
transform 1 0 20884 0 -1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_18_227
timestamp 1606120353
transform 1 0 21988 0 -1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_18_239
timestamp 1606120353
transform 1 0 23092 0 -1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_18_251
timestamp 1606120353
transform 1 0 24196 0 -1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_18_263
timestamp 1606120353
transform 1 0 25300 0 -1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1606120353
transform 1 0 26404 0 -1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_18_276
timestamp 1606120353
transform 1 0 26496 0 -1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606120353
transform -1 0 28888 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_18_288
timestamp 1606120353
transform 1 0 27600 0 -1 12512
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_18_296
timestamp 1606120353
transform 1 0 28336 0 -1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606120353
transform 1 0 1104 0 1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606120353
transform 1 0 1104 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1606120353
transform 1 0 1380 0 1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1606120353
transform 1 0 2484 0 1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1606120353
transform 1 0 1380 0 -1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1606120353
transform 1 0 2484 0 -1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1606120353
transform 1 0 3956 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1606120353
transform 1 0 3588 0 1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1606120353
transform 1 0 4692 0 1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1606120353
transform 1 0 3588 0 -1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1606120353
transform 1 0 4048 0 -1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1606120353
transform 1 0 5152 0 -1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1606120353
transform 1 0 6716 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1606120353
transform 1 0 5796 0 1 12512
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1606120353
transform 1 0 6532 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_19_62
timestamp 1606120353
transform 1 0 6808 0 1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_19_66
timestamp 1606120353
transform 1 0 7176 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_20_56
timestamp 1606120353
transform 1 0 6256 0 -1 13600
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_20_64
timestamp 1606120353
transform 1 0 6992 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_20_74
timestamp 1606120353
transform 1 0 7912 0 -1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_20_70
timestamp 1606120353
transform 1 0 7544 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_19_77
timestamp 1606120353
transform 1 0 8188 0 1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_19_69
timestamp 1606120353
transform 1 0 7452 0 1 12512
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_clk_A
timestamp 1606120353
transform 1 0 7268 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__B2
timestamp 1606120353
transform 1 0 7728 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_clk
timestamp 1606120353
transform 1 0 7268 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_20_85
timestamp 1606120353
transform 1 0 8924 0 -1 13600
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_20_81
timestamp 1606120353
transform 1 0 8556 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_20_78
timestamp 1606120353
transform 1 0 8280 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__D
timestamp 1606120353
transform 1 0 8464 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__B2
timestamp 1606120353
transform 1 0 8740 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__A1
timestamp 1606120353
transform 1 0 8372 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1109_
timestamp 1606120353
transform 1 0 8648 0 1 12512
box 0 -48 1748 592
use sky130_fd_sc_hd__inv_8  _0494_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 10580 0 -1 13600
box 0 -48 828 592
use sky130_fd_sc_hd__buf_1  _0495_
timestamp 1606120353
transform 1 0 11132 0 1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1606120353
transform 1 0 9568 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0494__A
timestamp 1606120353
transform 1 0 10580 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_101
timestamp 1606120353
transform 1 0 10396 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_19_105
timestamp 1606120353
transform 1 0 10764 0 1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1606120353
transform 1 0 9476 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_20_93
timestamp 1606120353
transform 1 0 9660 0 -1 13600
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_20_101
timestamp 1606120353
transform 1 0 10396 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_20_112
timestamp 1606120353
transform 1 0 11408 0 -1 13600
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_19_116
timestamp 1606120353
transform 1 0 11776 0 1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_19_112
timestamp 1606120353
transform 1 0 11408 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0495__A
timestamp 1606120353
transform 1 0 11592 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_126
timestamp 1606120353
transform 1 0 12696 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__B
timestamp 1606120353
transform 1 0 12144 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1606120353
transform 1 0 12328 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _0792_
timestamp 1606120353
transform 1 0 12144 0 -1 13600
box 0 -48 644 592
use sky130_fd_sc_hd__buf_1  _0787_
timestamp 1606120353
transform 1 0 12420 0 1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_20_131
timestamp 1606120353
transform 1 0 13156 0 -1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_20_127
timestamp 1606120353
transform 1 0 12788 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_19_130
timestamp 1606120353
transform 1 0 13064 0 1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0554__A
timestamp 1606120353
transform 1 0 12972 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__A
timestamp 1606120353
transform 1 0 12880 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_137
timestamp 1606120353
transform 1 0 13708 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_19_134
timestamp 1606120353
transform 1 0 13432 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__A
timestamp 1606120353
transform 1 0 13892 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0667__A
timestamp 1606120353
transform 1 0 13524 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0667_
timestamp 1606120353
transform 1 0 13524 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_20_150
timestamp 1606120353
transform 1 0 14904 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1606120353
transform 1 0 15180 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1606120353
transform 1 0 15272 0 -1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_20_138
timestamp 1606120353
transform 1 0 13800 0 -1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_19_153
timestamp 1606120353
transform 1 0 15180 0 1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_19_141
timestamp 1606120353
transform 1 0 14076 0 1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_19_165
timestamp 1606120353
transform 1 0 16284 0 1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1606120353
transform 1 0 16376 0 -1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1606120353
transform 1 0 17940 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_19_177
timestamp 1606120353
transform 1 0 17388 0 1 12512
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1606120353
transform 1 0 18032 0 1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1606120353
transform 1 0 19136 0 1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1606120353
transform 1 0 17480 0 -1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_20_190
timestamp 1606120353
transform 1 0 18584 0 -1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1144_
timestamp 1606120353
transform 1 0 21160 0 -1 13600
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1606120353
transform 1 0 20792 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__D
timestamp 1606120353
transform 1 0 21160 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_19_208
timestamp 1606120353
transform 1 0 20240 0 1 12512
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_19_216
timestamp 1606120353
transform 1 0 20976 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_19_220
timestamp 1606120353
transform 1 0 21344 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_20_202
timestamp 1606120353
transform 1 0 19688 0 -1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_20_215
timestamp 1606120353
transform 1 0 20884 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__CLK
timestamp 1606120353
transform 1 0 21528 0 1 12512
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_19_224
timestamp 1606120353
transform 1 0 21712 0 1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_19_236
timestamp 1606120353
transform 1 0 22816 0 1 12512
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_20_237
timestamp 1606120353
transform 1 0 22908 0 -1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1606120353
transform 1 0 23552 0 1 12512
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_19_245
timestamp 1606120353
transform 1 0 23644 0 1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_19_257
timestamp 1606120353
transform 1 0 24748 0 1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_20_249
timestamp 1606120353
transform 1 0 24012 0 -1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_20_261
timestamp 1606120353
transform 1 0 25116 0 -1 13600
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1606120353
transform 1 0 26404 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__CLK
timestamp 1606120353
transform 1 0 26128 0 -1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_19_269
timestamp 1606120353
transform 1 0 25852 0 1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1606120353
transform 1 0 26956 0 1 12512
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_20_269
timestamp 1606120353
transform 1 0 25852 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_20_274
timestamp 1606120353
transform 1 0 26312 0 -1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_20_276
timestamp 1606120353
transform 1 0 26496 0 -1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606120353
transform -1 0 28888 0 1 12512
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606120353
transform -1 0 28888 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_19_293
timestamp 1606120353
transform 1 0 28060 0 1 12512
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILLER_20_288
timestamp 1606120353
transform 1 0 27600 0 -1 13600
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_20_296
timestamp 1606120353
transform 1 0 28336 0 -1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606120353
transform 1 0 1104 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1606120353
transform 1 0 1380 0 1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1606120353
transform 1 0 2484 0 1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1606120353
transform 1 0 3588 0 1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1606120353
transform 1 0 4692 0 1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1606120353
transform 1 0 6716 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__A1
timestamp 1606120353
transform 1 0 7176 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1606120353
transform 1 0 5796 0 1 13600
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1606120353
transform 1 0 6532 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_21_62
timestamp 1606120353
transform 1 0 6808 0 1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__o22a_4  _0816_
timestamp 1606120353
transform 1 0 8372 0 1 13600
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__B1
timestamp 1606120353
transform 1 0 8188 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__B1
timestamp 1606120353
transform 1 0 7544 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_68
timestamp 1606120353
transform 1 0 7360 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_21_72
timestamp 1606120353
transform 1 0 7728 0 1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_21_76
timestamp 1606120353
transform 1 0 8096 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0497_
timestamp 1606120353
transform 1 0 10488 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0497__A
timestamp 1606120353
transform 1 0 10948 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__A
timestamp 1606120353
transform 1 0 9936 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_21_93
timestamp 1606120353
transform 1 0 9660 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_21_98
timestamp 1606120353
transform 1 0 10120 0 1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_21_105
timestamp 1606120353
transform 1 0 10764 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_109
timestamp 1606120353
transform 1 0 11132 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0554_
timestamp 1606120353
transform 1 0 12420 0 1 13600
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1606120353
transform 1 0 12328 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__A
timestamp 1606120353
transform 1 0 11316 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0559__A1_N
timestamp 1606120353
transform 1 0 12144 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0559__A2_N
timestamp 1606120353
transform 1 0 11776 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_21_113
timestamp 1606120353
transform 1 0 11500 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_21_118
timestamp 1606120353
transform 1 0 11960 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_132
timestamp 1606120353
transform 1 0 13248 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0604_
timestamp 1606120353
transform 1 0 13984 0 1 13600
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0604__A
timestamp 1606120353
transform 1 0 13800 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0559__B2
timestamp 1606120353
transform 1 0 13432 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_136
timestamp 1606120353
transform 1 0 13616 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_21_149
timestamp 1606120353
transform 1 0 14812 0 1 13600
box 0 -48 552 592
use sky130_fd_sc_hd__inv_8  _0575_
timestamp 1606120353
transform 1 0 15548 0 1 13600
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__A1
timestamp 1606120353
transform 1 0 16652 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__B1
timestamp 1606120353
transform 1 0 17020 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0575__A
timestamp 1606120353
transform 1 0 15364 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_21_166
timestamp 1606120353
transform 1 0 16376 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_21_171
timestamp 1606120353
transform 1 0 16836 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_21_175
timestamp 1606120353
transform 1 0 17204 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1606120353
transform 1 0 17940 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__A2
timestamp 1606120353
transform 1 0 17388 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_21_179
timestamp 1606120353
transform 1 0 17572 0 1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1606120353
transform 1 0 18032 0 1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1606120353
transform 1 0 19136 0 1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1606120353
transform 1 0 20240 0 1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_21_220
timestamp 1606120353
transform 1 0 21344 0 1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_21_232
timestamp 1606120353
transform 1 0 22448 0 1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1606120353
transform 1 0 23552 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_21_245
timestamp 1606120353
transform 1 0 23644 0 1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_21_257
timestamp 1606120353
transform 1 0 24748 0 1 13600
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1166_
timestamp 1606120353
transform 1 0 26128 0 1 13600
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__D
timestamp 1606120353
transform 1 0 25944 0 1 13600
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_21_269
timestamp 1606120353
transform 1 0 25852 0 1 13600
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606120353
transform -1 0 28888 0 1 13600
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_21_291
timestamp 1606120353
transform 1 0 27876 0 1 13600
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606120353
transform 1 0 1104 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1606120353
transform 1 0 1380 0 -1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1606120353
transform 1 0 2484 0 -1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1606120353
transform 1 0 3956 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1606120353
transform 1 0 3588 0 -1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1606120353
transform 1 0 4048 0 -1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1606120353
transform 1 0 5152 0 -1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1606120353
transform 1 0 6256 0 -1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__o22a_4  _0817_
timestamp 1606120353
transform 1 0 7544 0 -1 14688
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__A2
timestamp 1606120353
transform 1 0 9016 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__A2
timestamp 1606120353
transform 1 0 7360 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_84
timestamp 1606120353
transform 1 0 8832 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_22_88
timestamp 1606120353
transform 1 0 9200 0 -1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__buf_1  _0678_
timestamp 1606120353
transform 1 0 9936 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0711_
timestamp 1606120353
transform 1 0 10948 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1606120353
transform 1 0 9568 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_22_93
timestamp 1606120353
transform 1 0 9660 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_22_99
timestamp 1606120353
transform 1 0 10212 0 -1 14688
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_22_110
timestamp 1606120353
transform 1 0 11224 0 -1 14688
box 0 -48 736 592
use sky130_fd_sc_hd__a2bb2o_4  _0559_
timestamp 1606120353
transform 1 0 12420 0 -1 14688
box 0 -48 1472 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0559__B1
timestamp 1606120353
transform 1 0 12236 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_22_118
timestamp 1606120353
transform 1 0 11960 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1606120353
transform 1 0 15180 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0615__A2_N
timestamp 1606120353
transform 1 0 14076 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0615__A1_N
timestamp 1606120353
transform 1 0 14444 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0615__B1
timestamp 1606120353
transform 1 0 14812 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_139
timestamp 1606120353
transform 1 0 13892 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_143
timestamp 1606120353
transform 1 0 14260 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_147
timestamp 1606120353
transform 1 0 14628 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_22_151
timestamp 1606120353
transform 1 0 14996 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_22_154
timestamp 1606120353
transform 1 0 15272 0 -1 14688
box 0 -48 552 592
use sky130_fd_sc_hd__a21o_4  _0756_
timestamp 1606120353
transform 1 0 16652 0 -1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__CLK
timestamp 1606120353
transform 1 0 15916 0 -1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_22_160
timestamp 1606120353
transform 1 0 15824 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_22_163
timestamp 1606120353
transform 1 0 16100 0 -1 14688
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_22_181
timestamp 1606120353
transform 1 0 17756 0 -1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_22_193
timestamp 1606120353
transform 1 0 18860 0 -1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1606120353
transform 1 0 20792 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_22_205
timestamp 1606120353
transform 1 0 19964 0 -1 14688
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_22_213
timestamp 1606120353
transform 1 0 20700 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_22_215
timestamp 1606120353
transform 1 0 20884 0 -1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_22_227
timestamp 1606120353
transform 1 0 21988 0 -1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_22_239
timestamp 1606120353
transform 1 0 23092 0 -1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_22_251
timestamp 1606120353
transform 1 0 24196 0 -1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_22_263
timestamp 1606120353
transform 1 0 25300 0 -1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1606120353
transform 1 0 26404 0 -1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_22_276
timestamp 1606120353
transform 1 0 26496 0 -1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606120353
transform -1 0 28888 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_22_288
timestamp 1606120353
transform 1 0 27600 0 -1 14688
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_22_296
timestamp 1606120353
transform 1 0 28336 0 -1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606120353
transform 1 0 1104 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1606120353
transform 1 0 1380 0 1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1606120353
transform 1 0 2484 0 1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1606120353
transform 1 0 3588 0 1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1606120353
transform 1 0 4692 0 1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1606120353
transform 1 0 6716 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__D
timestamp 1606120353
transform 1 0 6992 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__CLK
timestamp 1606120353
transform 1 0 6532 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1606120353
transform 1 0 5796 0 1 14688
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_23_62
timestamp 1606120353
transform 1 0 6808 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_66
timestamp 1606120353
transform 1 0 7176 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1110_
timestamp 1606120353
transform 1 0 8280 0 1 14688
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__D
timestamp 1606120353
transform 1 0 8096 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_clk_A
timestamp 1606120353
transform 1 0 7360 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__CLK
timestamp 1606120353
transform 1 0 7728 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_70
timestamp 1606120353
transform 1 0 7544 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_74
timestamp 1606120353
transform 1 0 7912 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0663_
timestamp 1606120353
transform 1 0 10764 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0663__A
timestamp 1606120353
transform 1 0 11224 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__A
timestamp 1606120353
transform 1 0 10212 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_97
timestamp 1606120353
transform 1 0 10028 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_23_101
timestamp 1606120353
transform 1 0 10396 0 1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_23_108
timestamp 1606120353
transform 1 0 11040 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0614_
timestamp 1606120353
transform 1 0 12512 0 1 14688
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1606120353
transform 1 0 12328 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0577__B2
timestamp 1606120353
transform 1 0 12144 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0614__A
timestamp 1606120353
transform 1 0 11776 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_23_112
timestamp 1606120353
transform 1 0 11408 0 1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_23_118
timestamp 1606120353
transform 1 0 11960 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_23_123
timestamp 1606120353
transform 1 0 12420 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__a2bb2o_4  _0615_
timestamp 1606120353
transform 1 0 14076 0 1 14688
box 0 -48 1472 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0577__B1
timestamp 1606120353
transform 1 0 13524 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0615__B2
timestamp 1606120353
transform 1 0 13892 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_133
timestamp 1606120353
transform 1 0 13340 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_23_137
timestamp 1606120353
transform 1 0 13708 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0755_
timestamp 1606120353
transform 1 0 16560 0 1 14688
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__B
timestamp 1606120353
transform 1 0 16376 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__D
timestamp 1606120353
transform 1 0 15916 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_23_157
timestamp 1606120353
transform 1 0 15548 0 1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_23_163
timestamp 1606120353
transform 1 0 16100 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_23_175
timestamp 1606120353
transform 1 0 17204 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1606120353
transform 1 0 17940 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__A
timestamp 1606120353
transform 1 0 17388 0 1 14688
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_23_179
timestamp 1606120353
transform 1 0 17572 0 1 14688
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1606120353
transform 1 0 18032 0 1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1606120353
transform 1 0 19136 0 1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1606120353
transform 1 0 20240 0 1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_23_220
timestamp 1606120353
transform 1 0 21344 0 1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_23_232
timestamp 1606120353
transform 1 0 22448 0 1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1606120353
transform 1 0 23552 0 1 14688
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_23_245
timestamp 1606120353
transform 1 0 23644 0 1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_23_257
timestamp 1606120353
transform 1 0 24748 0 1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_23_269
timestamp 1606120353
transform 1 0 25852 0 1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1606120353
transform 1 0 26956 0 1 14688
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606120353
transform -1 0 28888 0 1 14688
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_23_293
timestamp 1606120353
transform 1 0 28060 0 1 14688
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606120353
transform 1 0 1104 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1606120353
transform 1 0 1380 0 -1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_24_15
timestamp 1606120353
transform 1 0 2484 0 -1 15776
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1606120353
transform 1 0 3956 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__CLK
timestamp 1606120353
transform 1 0 3404 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_23
timestamp 1606120353
transform 1 0 3220 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1606120353
transform 1 0 3588 0 -1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1606120353
transform 1 0 4048 0 -1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1606120353
transform 1 0 5152 0 -1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1129_
timestamp 1606120353
transform 1 0 6992 0 -1 15776
box 0 -48 1748 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_clk
timestamp 1606120353
transform 1 0 6624 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_24_56
timestamp 1606120353
transform 1 0 6256 0 -1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_24_63
timestamp 1606120353
transform 1 0 6900 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_24_83
timestamp 1606120353
transform 1 0 8740 0 -1 15776
box 0 -48 736 592
use sky130_fd_sc_hd__buf_1  _0691_
timestamp 1606120353
transform 1 0 9844 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1606120353
transform 1 0 9568 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__A1
timestamp 1606120353
transform 1 0 10304 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1606120353
transform 1 0 9476 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_24_93
timestamp 1606120353
transform 1 0 9660 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_98
timestamp 1606120353
transform 1 0 10120 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_24_102
timestamp 1606120353
transform 1 0 10488 0 -1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__a2bb2o_4  _0577_
timestamp 1606120353
transform 1 0 12972 0 -1 15776
box 0 -48 1472 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0577__A1_N
timestamp 1606120353
transform 1 0 12788 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0577__A2_N
timestamp 1606120353
transform 1 0 12420 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_24_114
timestamp 1606120353
transform 1 0 11592 0 -1 15776
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_24_122
timestamp 1606120353
transform 1 0 12328 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_24_125
timestamp 1606120353
transform 1 0 12604 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1606120353
transform 1 0 15180 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0578__B
timestamp 1606120353
transform 1 0 14628 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0578__D
timestamp 1606120353
transform 1 0 14996 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_145
timestamp 1606120353
transform 1 0 14444 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_149
timestamp 1606120353
transform 1 0 14812 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_24_154
timestamp 1606120353
transform 1 0 15272 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1087_
timestamp 1606120353
transform 1 0 15916 0 -1 15776
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0574__A
timestamp 1606120353
transform 1 0 15456 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_24_158
timestamp 1606120353
transform 1 0 15640 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__CLK
timestamp 1606120353
transform 1 0 18032 0 -1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_24_180
timestamp 1606120353
transform 1 0 17664 0 -1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_24_186
timestamp 1606120353
transform 1 0 18216 0 -1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_24_198
timestamp 1606120353
transform 1 0 19320 0 -1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1606120353
transform 1 0 20792 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_24_210
timestamp 1606120353
transform 1 0 20424 0 -1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_24_215
timestamp 1606120353
transform 1 0 20884 0 -1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_24_227
timestamp 1606120353
transform 1 0 21988 0 -1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_24_239
timestamp 1606120353
transform 1 0 23092 0 -1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_24_251
timestamp 1606120353
transform 1 0 24196 0 -1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_24_263
timestamp 1606120353
transform 1 0 25300 0 -1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1606120353
transform 1 0 26404 0 -1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_24_276
timestamp 1606120353
transform 1 0 26496 0 -1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606120353
transform -1 0 28888 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_24_288
timestamp 1606120353
transform 1 0 27600 0 -1 15776
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_24_296
timestamp 1606120353
transform 1 0 28336 0 -1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606120353
transform 1 0 1104 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1606120353
transform 1 0 1380 0 1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_25_15
timestamp 1606120353
transform 1 0 2484 0 1 15776
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1137_
timestamp 1606120353
transform 1 0 3404 0 1 15776
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__D
timestamp 1606120353
transform 1 0 3220 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_25_44
timestamp 1606120353
transform 1 0 5152 0 1 15776
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1606120353
transform 1 0 6716 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__D
timestamp 1606120353
transform 1 0 6072 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__CLK
timestamp 1606120353
transform 1 0 6440 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_52
timestamp 1606120353
transform 1 0 5888 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_56
timestamp 1606120353
transform 1 0 6256 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_25_60
timestamp 1606120353
transform 1 0 6624 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_25_62
timestamp 1606120353
transform 1 0 6808 0 1 15776
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1112_
timestamp 1606120353
transform 1 0 8280 0 1 15776
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__D
timestamp 1606120353
transform 1 0 8096 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__CLK
timestamp 1606120353
transform 1 0 7728 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_70
timestamp 1606120353
transform 1 0 7544 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_74
timestamp 1606120353
transform 1 0 7912 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0750_
timestamp 1606120353
transform 1 0 10764 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__A2
timestamp 1606120353
transform 1 0 11224 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__B1
timestamp 1606120353
transform 1 0 10580 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__A1
timestamp 1606120353
transform 1 0 10212 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_97
timestamp 1606120353
transform 1 0 10028 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_101
timestamp 1606120353
transform 1 0 10396 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_108
timestamp 1606120353
transform 1 0 11040 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0560_
timestamp 1606120353
transform 1 0 12604 0 1 15776
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1606120353
transform 1 0 12328 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__A
timestamp 1606120353
transform 1 0 11592 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0560__A
timestamp 1606120353
transform 1 0 12144 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_112
timestamp 1606120353
transform 1 0 11408 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_25_116
timestamp 1606120353
transform 1 0 11776 0 1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_25_123
timestamp 1606120353
transform 1 0 12420 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__nor4_4  _0578_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 14628 0 1 15776
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0578__A
timestamp 1606120353
transform 1 0 14444 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0568__A1
timestamp 1606120353
transform 1 0 13616 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0568__A2
timestamp 1606120353
transform 1 0 13984 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_134
timestamp 1606120353
transform 1 0 13432 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_138
timestamp 1606120353
transform 1 0 13800 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_25_142
timestamp 1606120353
transform 1 0 14168 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0557__A
timestamp 1606120353
transform 1 0 17204 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0574__B
timestamp 1606120353
transform 1 0 16376 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0574__C
timestamp 1606120353
transform 1 0 16744 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_164
timestamp 1606120353
transform 1 0 16192 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_25_168
timestamp 1606120353
transform 1 0 16560 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_25_172
timestamp 1606120353
transform 1 0 16928 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1180_
timestamp 1606120353
transform 1 0 18032 0 1 15776
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1606120353
transform 1 0 17940 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__D
timestamp 1606120353
transform 1 0 17756 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_25_177
timestamp 1606120353
transform 1 0 17388 0 1 15776
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_25_203
timestamp 1606120353
transform 1 0 19780 0 1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_25_215
timestamp 1606120353
transform 1 0 20884 0 1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__D
timestamp 1606120353
transform 1 0 22264 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__CLK
timestamp 1606120353
transform 1 0 22632 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_25_227
timestamp 1606120353
transform 1 0 21988 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_25_232
timestamp 1606120353
transform 1 0 22448 0 1 15776
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_25_236
timestamp 1606120353
transform 1 0 22816 0 1 15776
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1606120353
transform 1 0 23552 0 1 15776
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_25_245
timestamp 1606120353
transform 1 0 23644 0 1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_25_257
timestamp 1606120353
transform 1 0 24748 0 1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_25_269
timestamp 1606120353
transform 1 0 25852 0 1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1606120353
transform 1 0 26956 0 1 15776
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606120353
transform -1 0 28888 0 1 15776
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_25_293
timestamp 1606120353
transform 1 0 28060 0 1 15776
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1202_
timestamp 1606120353
transform 1 0 1380 0 1 16864
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606120353
transform 1 0 1104 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606120353
transform 1 0 1104 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__D
timestamp 1606120353
transform 1 0 1564 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__CLK
timestamp 1606120353
transform 1 0 1932 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1606120353
transform 1 0 1380 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_7
timestamp 1606120353
transform 1 0 1748 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_26_11
timestamp 1606120353
transform 1 0 2116 0 -1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_27_22
timestamp 1606120353
transform 1 0 3128 0 1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1606120353
transform 1 0 3956 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_26_23
timestamp 1606120353
transform 1 0 3220 0 -1 16864
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1606120353
transform 1 0 4048 0 -1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_26_44
timestamp 1606120353
transform 1 0 5152 0 -1 16864
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_27_34
timestamp 1606120353
transform 1 0 4232 0 1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1120_
timestamp 1606120353
transform 1 0 6072 0 -1 16864
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1606120353
transform 1 0 6716 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_26_52
timestamp 1606120353
transform 1 0 5888 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_27_46
timestamp 1606120353
transform 1 0 5336 0 1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_27_58
timestamp 1606120353
transform 1 0 6440 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_27_62
timestamp 1606120353
transform 1 0 6808 0 1 16864
box 0 -48 736 592
use sky130_fd_sc_hd__o22a_4  _0819_
timestamp 1606120353
transform 1 0 8188 0 1 16864
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__B1
timestamp 1606120353
transform 1 0 8004 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__A1
timestamp 1606120353
transform 1 0 8188 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__A2
timestamp 1606120353
transform 1 0 7636 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_26_73
timestamp 1606120353
transform 1 0 7820 0 -1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILLER_26_79
timestamp 1606120353
transform 1 0 8372 0 -1 16864
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_26_87
timestamp 1606120353
transform 1 0 9108 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_27_70
timestamp 1606120353
transform 1 0 7544 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_27_73
timestamp 1606120353
transform 1 0 7820 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_96
timestamp 1606120353
transform 1 0 9936 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_27_91
timestamp 1606120353
transform 1 0 9476 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_26_98
timestamp 1606120353
transform 1 0 10120 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_26_93
timestamp 1606120353
transform 1 0 9660 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__A1
timestamp 1606120353
transform 1 0 9384 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__B2
timestamp 1606120353
transform 1 0 9936 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__A2
timestamp 1606120353
transform 1 0 9752 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__A2
timestamp 1606120353
transform 1 0 10120 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1606120353
transform 1 0 9568 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_26_102
timestamp 1606120353
transform 1 0 10488 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__B1
timestamp 1606120353
transform 1 0 10304 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _0754_
timestamp 1606120353
transform 1 0 10304 0 1 16864
box 0 -48 1288 592
use sky130_fd_sc_hd__o21a_4  _0753_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 10672 0 -1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_27_118
timestamp 1606120353
transform 1 0 11960 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_114
timestamp 1606120353
transform 1 0 11592 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_120
timestamp 1606120353
transform 1 0 12144 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_116
timestamp 1606120353
transform 1 0 11776 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0603__A
timestamp 1606120353
transform 1 0 11960 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__B1
timestamp 1606120353
transform 1 0 11776 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__A2_N
timestamp 1606120353
transform 1 0 12144 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_27_123
timestamp 1606120353
transform 1 0 12420 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_26_128
timestamp 1606120353
transform 1 0 12880 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_124
timestamp 1606120353
transform 1 0 12512 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__B2
timestamp 1606120353
transform 1 0 12696 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__A1_N
timestamp 1606120353
transform 1 0 12328 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0568__B1
timestamp 1606120353
transform 1 0 13064 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1606120353
transform 1 0 12328 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _0603_
timestamp 1606120353
transform 1 0 12512 0 1 16864
box 0 -48 828 592
use sky130_fd_sc_hd__o21ai_4  _0568_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 13248 0 -1 16864
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_27_137
timestamp 1606120353
transform 1 0 13708 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_133
timestamp 1606120353
transform 1 0 13340 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__B2
timestamp 1606120353
transform 1 0 13524 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__A2_N
timestamp 1606120353
transform 1 0 13892 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_149
timestamp 1606120353
transform 1 0 14812 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_145
timestamp 1606120353
transform 1 0 14444 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__B1
timestamp 1606120353
transform 1 0 14996 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0578__C
timestamp 1606120353
transform 1 0 14628 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1606120353
transform 1 0 15180 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__a2bb2o_4  _0605_
timestamp 1606120353
transform 1 0 14076 0 1 16864
box 0 -48 1472 592
use sky130_fd_sc_hd__nor3_4  _0574_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 15272 0 -1 16864
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_27_161
timestamp 1606120353
transform 1 0 15916 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_27_157
timestamp 1606120353
transform 1 0 15548 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__A2
timestamp 1606120353
transform 1 0 15732 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_26_167
timestamp 1606120353
transform 1 0 16468 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__B2
timestamp 1606120353
transform 1 0 16100 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0639_
timestamp 1606120353
transform 1 0 16284 0 1 16864
box 0 -48 644 592
use sky130_fd_sc_hd__decap_4  FILLER_27_172
timestamp 1606120353
transform 1 0 16928 0 1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_26_171
timestamp 1606120353
transform 1 0 16836 0 -1 16864
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__B
timestamp 1606120353
transform 1 0 16652 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0557_
timestamp 1606120353
transform 1 0 17204 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__D
timestamp 1606120353
transform 1 0 17296 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1606120353
transform 1 0 17940 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__CLK
timestamp 1606120353
transform 1 0 17664 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1606120353
transform 1 0 17480 0 -1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1606120353
transform 1 0 18584 0 -1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_27_178
timestamp 1606120353
transform 1 0 17480 0 1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_27_182
timestamp 1606120353
transform 1 0 17848 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1606120353
transform 1 0 18032 0 1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1606120353
transform 1 0 19136 0 1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1606120353
transform 1 0 20792 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_26_202
timestamp 1606120353
transform 1 0 19688 0 -1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1606120353
transform 1 0 20884 0 -1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1606120353
transform 1 0 20240 0 1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_27_220
timestamp 1606120353
transform 1 0 21344 0 1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1188_
timestamp 1606120353
transform 1 0 22264 0 -1 16864
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  FILLER_26_227
timestamp 1606120353
transform 1 0 21988 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_27_232
timestamp 1606120353
transform 1 0 22448 0 1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1606120353
transform 1 0 23552 0 1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_26_249
timestamp 1606120353
transform 1 0 24012 0 -1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_26_261
timestamp 1606120353
transform 1 0 25116 0 -1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_27_245
timestamp 1606120353
transform 1 0 23644 0 1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_27_257
timestamp 1606120353
transform 1 0 24748 0 1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1606120353
transform 1 0 26404 0 -1 16864
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_26_273
timestamp 1606120353
transform 1 0 26220 0 -1 16864
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_26_276
timestamp 1606120353
transform 1 0 26496 0 -1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_27_269
timestamp 1606120353
transform 1 0 25852 0 1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1606120353
transform 1 0 26956 0 1 16864
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606120353
transform -1 0 28888 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606120353
transform -1 0 28888 0 1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_26_288
timestamp 1606120353
transform 1 0 27600 0 -1 16864
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_26_296
timestamp 1606120353
transform 1 0 28336 0 -1 16864
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_27_293
timestamp 1606120353
transform 1 0 28060 0 1 16864
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1606120353
transform 1 0 1104 0 -1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__CLK
timestamp 1606120353
transform 1 0 1840 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_28_3
timestamp 1606120353
transform 1 0 1380 0 -1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_28_7
timestamp 1606120353
transform 1 0 1748 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_28_10
timestamp 1606120353
transform 1 0 2024 0 -1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_28_22
timestamp 1606120353
transform 1 0 3128 0 -1 17952
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1606120353
transform 1 0 3956 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_28_30
timestamp 1606120353
transform 1 0 3864 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1606120353
transform 1 0 4048 0 -1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1606120353
transform 1 0 5152 0 -1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1606120353
transform 1 0 6256 0 -1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__B2
timestamp 1606120353
transform 1 0 8188 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A1
timestamp 1606120353
transform 1 0 9016 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_28_68
timestamp 1606120353
transform 1 0 7360 0 -1 17952
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_28_76
timestamp 1606120353
transform 1 0 8096 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_28_79
timestamp 1606120353
transform 1 0 8372 0 -1 17952
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_28_85
timestamp 1606120353
transform 1 0 8924 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_28_88
timestamp 1606120353
transform 1 0 9200 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0767_
timestamp 1606120353
transform 1 0 10304 0 -1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1606120353
transform 1 0 9568 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__B1
timestamp 1606120353
transform 1 0 10120 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__A1
timestamp 1606120353
transform 1 0 9384 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_28_93
timestamp 1606120353
transform 1 0 9660 0 -1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_28_97
timestamp 1606120353
transform 1 0 10028 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__a2bb2o_4  _0765_
timestamp 1606120353
transform 1 0 12328 0 -1 17952
box 0 -48 1472 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__A2
timestamp 1606120353
transform 1 0 12144 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__B1
timestamp 1606120353
transform 1 0 11592 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_112
timestamp 1606120353
transform 1 0 11408 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_28_116
timestamp 1606120353
transform 1 0 11776 0 -1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__o22a_4  _0625_
timestamp 1606120353
transform 1 0 15272 0 -1 17952
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1606120353
transform 1 0 15180 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__B2
timestamp 1606120353
transform 1 0 14536 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__A1_N
timestamp 1606120353
transform 1 0 14076 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__A1
timestamp 1606120353
transform 1 0 14996 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_28_138
timestamp 1606120353
transform 1 0 13800 0 -1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_28_143
timestamp 1606120353
transform 1 0 14260 0 -1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_28_148
timestamp 1606120353
transform 1 0 14720 0 -1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1139_
timestamp 1606120353
transform 1 0 17296 0 -1 17952
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__A
timestamp 1606120353
transform 1 0 16744 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__CLK
timestamp 1606120353
transform 1 0 17112 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_168
timestamp 1606120353
transform 1 0 16560 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_28_172
timestamp 1606120353
transform 1 0 16928 0 -1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_28_195
timestamp 1606120353
transform 1 0 19044 0 -1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1606120353
transform 1 0 20792 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_28_207
timestamp 1606120353
transform 1 0 20148 0 -1 17952
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_28_213
timestamp 1606120353
transform 1 0 20700 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1606120353
transform 1 0 20884 0 -1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1606120353
transform 1 0 21988 0 -1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1606120353
transform 1 0 23092 0 -1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_28_251
timestamp 1606120353
transform 1 0 24196 0 -1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_28_263
timestamp 1606120353
transform 1 0 25300 0 -1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1606120353
transform 1 0 26404 0 -1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_28_276
timestamp 1606120353
transform 1 0 26496 0 -1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1606120353
transform -1 0 28888 0 -1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_28_288
timestamp 1606120353
transform 1 0 27600 0 -1 17952
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_28_296
timestamp 1606120353
transform 1 0 28336 0 -1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1136_
timestamp 1606120353
transform 1 0 1840 0 1 17952
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1606120353
transform 1 0 1104 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__D
timestamp 1606120353
transform 1 0 1656 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_29_3
timestamp 1606120353
transform 1 0 1380 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1606120353
transform 1 0 3588 0 1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1606120353
transform 1 0 4692 0 1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1606120353
transform 1 0 6716 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__D
timestamp 1606120353
transform 1 0 7084 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1606120353
transform 1 0 5796 0 1 17952
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1606120353
transform 1 0 6532 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_29_62
timestamp 1606120353
transform 1 0 6808 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__B1
timestamp 1606120353
transform 1 0 9200 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__B2
timestamp 1606120353
transform 1 0 8832 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__CLK
timestamp 1606120353
transform 1 0 7452 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_67
timestamp 1606120353
transform 1 0 7268 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_29_71
timestamp 1606120353
transform 1 0 7636 0 1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_29_83
timestamp 1606120353
transform 1 0 8740 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_29_86
timestamp 1606120353
transform 1 0 9016 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0760_
timestamp 1606120353
transform 1 0 9752 0 1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A2
timestamp 1606120353
transform 1 0 9568 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__A2
timestamp 1606120353
transform 1 0 11040 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_90
timestamp 1606120353
transform 1 0 9384 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_106
timestamp 1606120353
transform 1 0 10856 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_110
timestamp 1606120353
transform 1 0 11224 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0766_
timestamp 1606120353
transform 1 0 12420 0 1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1606120353
transform 1 0 12328 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__A1
timestamp 1606120353
transform 1 0 12144 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__B1
timestamp 1606120353
transform 1 0 11776 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__A2
timestamp 1606120353
transform 1 0 11408 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_114
timestamp 1606120353
transform 1 0 11592 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_118
timestamp 1606120353
transform 1 0 11960 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__a22oi_4  _0573_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 14536 0 1 17952
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__A2
timestamp 1606120353
transform 1 0 14352 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__B1
timestamp 1606120353
transform 1 0 13708 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_135
timestamp 1606120353
transform 1 0 13524 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_29_139
timestamp 1606120353
transform 1 0 13892 0 1 17952
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_29_143
timestamp 1606120353
transform 1 0 14260 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0571_
timestamp 1606120353
transform 1 0 16836 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0571__A
timestamp 1606120353
transform 1 0 17296 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0572__A
timestamp 1606120353
transform 1 0 16284 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0609__A
timestamp 1606120353
transform 1 0 16652 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_163
timestamp 1606120353
transform 1 0 16100 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_167
timestamp 1606120353
transform 1 0 16468 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_174
timestamp 1606120353
transform 1 0 17112 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1606120353
transform 1 0 17940 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0609__B
timestamp 1606120353
transform 1 0 17664 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_29_178
timestamp 1606120353
transform 1 0 17480 0 1 17952
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_29_182
timestamp 1606120353
transform 1 0 17848 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1606120353
transform 1 0 18032 0 1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1606120353
transform 1 0 19136 0 1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1606120353
transform 1 0 20240 0 1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_29_220
timestamp 1606120353
transform 1 0 21344 0 1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_29_232
timestamp 1606120353
transform 1 0 22448 0 1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1606120353
transform 1 0 23552 0 1 17952
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_29_245
timestamp 1606120353
transform 1 0 23644 0 1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_29_257
timestamp 1606120353
transform 1 0 24748 0 1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_29_269
timestamp 1606120353
transform 1 0 25852 0 1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1606120353
transform 1 0 26956 0 1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1606120353
transform -1 0 28888 0 1 17952
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_29_293
timestamp 1606120353
transform 1 0 28060 0 1 17952
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1606120353
transform 1 0 1104 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1606120353
transform 1 0 1380 0 -1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1606120353
transform 1 0 2484 0 -1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1606120353
transform 1 0 3956 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1606120353
transform 1 0 3588 0 -1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1606120353
transform 1 0 4048 0 -1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1606120353
transform 1 0 5152 0 -1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1111_
timestamp 1606120353
transform 1 0 7084 0 -1 19040
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_8  FILLER_30_56
timestamp 1606120353
transform 1 0 6256 0 -1 19040
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_30_64
timestamp 1606120353
transform 1 0 6992 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_30_84
timestamp 1606120353
transform 1 0 8832 0 -1 19040
box 0 -48 552 592
use sky130_fd_sc_hd__o22a_4  _0768_
timestamp 1606120353
transform 1 0 10672 0 -1 19040
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1606120353
transform 1 0 9568 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A2
timestamp 1606120353
transform 1 0 9844 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__B2
timestamp 1606120353
transform 1 0 10212 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A1
timestamp 1606120353
transform 1 0 9384 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_93
timestamp 1606120353
transform 1 0 9660 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_97
timestamp 1606120353
transform 1 0 10028 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_30_101
timestamp 1606120353
transform 1 0 10396 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__o21a_4  _0752_
timestamp 1606120353
transform 1 0 12696 0 -1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__A1
timestamp 1606120353
transform 1 0 12420 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_30_118
timestamp 1606120353
transform 1 0 11960 0 -1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_30_122
timestamp 1606120353
transform 1 0 12328 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_30_125
timestamp 1606120353
transform 1 0 12604 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _0572_
timestamp 1606120353
transform 1 0 15272 0 -1 19040
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1606120353
transform 1 0 15180 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__A2
timestamp 1606120353
transform 1 0 13984 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__A
timestamp 1606120353
transform 1 0 14352 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__B1
timestamp 1606120353
transform 1 0 14720 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_138
timestamp 1606120353
transform 1 0 13800 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_142
timestamp 1606120353
transform 1 0 14168 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_146
timestamp 1606120353
transform 1 0 14536 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_30_150
timestamp 1606120353
transform 1 0 14904 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__and2_4  _0609_
timestamp 1606120353
transform 1 0 16836 0 -1 19040
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__D
timestamp 1606120353
transform 1 0 16284 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__B1
timestamp 1606120353
transform 1 0 16652 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_163
timestamp 1606120353
transform 1 0 16100 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_167
timestamp 1606120353
transform 1 0 16468 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__B
timestamp 1606120353
transform 1 0 18032 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__CLK
timestamp 1606120353
transform 1 0 17664 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_178
timestamp 1606120353
transform 1 0 17480 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_30_182
timestamp 1606120353
transform 1 0 17848 0 -1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_30_186
timestamp 1606120353
transform 1 0 18216 0 -1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_30_198
timestamp 1606120353
transform 1 0 19320 0 -1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1606120353
transform 1 0 20792 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_30_210
timestamp 1606120353
transform 1 0 20424 0 -1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1606120353
transform 1 0 20884 0 -1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1606120353
transform 1 0 21988 0 -1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_30_239
timestamp 1606120353
transform 1 0 23092 0 -1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_30_251
timestamp 1606120353
transform 1 0 24196 0 -1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_30_263
timestamp 1606120353
transform 1 0 25300 0 -1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1606120353
transform 1 0 26404 0 -1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_30_276
timestamp 1606120353
transform 1 0 26496 0 -1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1606120353
transform -1 0 28888 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_30_288
timestamp 1606120353
transform 1 0 27600 0 -1 19040
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_30_296
timestamp 1606120353
transform 1 0 28336 0 -1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1606120353
transform 1 0 1104 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1606120353
transform 1 0 1380 0 1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1606120353
transform 1 0 2484 0 1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1606120353
transform 1 0 3588 0 1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1606120353
transform 1 0 4692 0 1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1606120353
transform 1 0 6716 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A1
timestamp 1606120353
transform 1 0 7176 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A2
timestamp 1606120353
transform 1 0 6532 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1606120353
transform 1 0 5796 0 1 19040
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_31_62
timestamp 1606120353
transform 1 0 6808 0 1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__o22a_4  _0818_
timestamp 1606120353
transform 1 0 7360 0 1 19040
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__B
timestamp 1606120353
transform 1 0 8832 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__A
timestamp 1606120353
transform 1 0 9200 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_82
timestamp 1606120353
transform 1 0 8648 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_86
timestamp 1606120353
transform 1 0 9016 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _0761_
timestamp 1606120353
transform 1 0 9476 0 1 19040
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__A1
timestamp 1606120353
transform 1 0 10948 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_31_90
timestamp 1606120353
transform 1 0 9384 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_31_105
timestamp 1606120353
transform 1 0 10764 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_109
timestamp 1606120353
transform 1 0 11132 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0751_
timestamp 1606120353
transform 1 0 12420 0 1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1606120353
transform 1 0 12328 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__B
timestamp 1606120353
transform 1 0 12144 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__A1
timestamp 1606120353
transform 1 0 11776 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__B1
timestamp 1606120353
transform 1 0 11316 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_31_113
timestamp 1606120353
transform 1 0 11500 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_31_118
timestamp 1606120353
transform 1 0 11960 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0553_
timestamp 1606120353
transform 1 0 14444 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0553__A
timestamp 1606120353
transform 1 0 14904 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0593__A
timestamp 1606120353
transform 1 0 15272 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0630__A
timestamp 1606120353
transform 1 0 13984 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_31_135
timestamp 1606120353
transform 1 0 13524 0 1 19040
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_31_139
timestamp 1606120353
transform 1 0 13892 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_31_142
timestamp 1606120353
transform 1 0 14168 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_31_148
timestamp 1606120353
transform 1 0 14720 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_152
timestamp 1606120353
transform 1 0 15088 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1103_
timestamp 1606120353
transform 1 0 15456 0 1 19040
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_2  FILLER_31_175
timestamp 1606120353
transform 1 0 17204 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0763_
timestamp 1606120353
transform 1 0 18032 0 1 19040
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1606120353
transform 1 0 17940 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0608__B
timestamp 1606120353
transform 1 0 18952 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__A
timestamp 1606120353
transform 1 0 17756 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0608__A
timestamp 1606120353
transform 1 0 19320 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__D
timestamp 1606120353
transform 1 0 17388 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_31_179
timestamp 1606120353
transform 1 0 17572 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_31_191
timestamp 1606120353
transform 1 0 18676 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_31_196
timestamp 1606120353
transform 1 0 19136 0 1 19040
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_31_200
timestamp 1606120353
transform 1 0 19504 0 1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_31_212
timestamp 1606120353
transform 1 0 20608 0 1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_31_224
timestamp 1606120353
transform 1 0 21712 0 1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_31_236
timestamp 1606120353
transform 1 0 22816 0 1 19040
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1606120353
transform 1 0 23552 0 1 19040
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_31_245
timestamp 1606120353
transform 1 0 23644 0 1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_31_257
timestamp 1606120353
transform 1 0 24748 0 1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_31_269
timestamp 1606120353
transform 1 0 25852 0 1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1606120353
transform 1 0 26956 0 1 19040
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1606120353
transform -1 0 28888 0 1 19040
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_31_293
timestamp 1606120353
transform 1 0 28060 0 1 19040
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1606120353
transform 1 0 1104 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1606120353
transform 1 0 1380 0 -1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1606120353
transform 1 0 2484 0 -1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1606120353
transform 1 0 3956 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1606120353
transform 1 0 3588 0 -1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1606120353
transform 1 0 4048 0 -1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1606120353
transform 1 0 5152 0 -1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1606120353
transform 1 0 6256 0 -1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__and2_4  _0757_
timestamp 1606120353
transform 1 0 8188 0 -1 20128
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__B2
timestamp 1606120353
transform 1 0 7360 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__B1
timestamp 1606120353
transform 1 0 7728 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_70
timestamp 1606120353
transform 1 0 7544 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_32_74
timestamp 1606120353
transform 1 0 7912 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_32_84
timestamp 1606120353
transform 1 0 8832 0 -1 20128
box 0 -48 736 592
use sky130_fd_sc_hd__a21o_4  _0758_
timestamp 1606120353
transform 1 0 10764 0 -1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1606120353
transform 1 0 9568 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__A1
timestamp 1606120353
transform 1 0 10304 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__B1
timestamp 1606120353
transform 1 0 9844 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_93
timestamp 1606120353
transform 1 0 9660 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_32_97
timestamp 1606120353
transform 1 0 10028 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_32_102
timestamp 1606120353
transform 1 0 10488 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__and2_4  _0634_
timestamp 1606120353
transform 1 0 12604 0 -1 20128
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__B1
timestamp 1606120353
transform 1 0 12420 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__B
timestamp 1606120353
transform 1 0 12052 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_117
timestamp 1606120353
transform 1 0 11868 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_121
timestamp 1606120353
transform 1 0 12236 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_132
timestamp 1606120353
transform 1 0 13248 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__B1
timestamp 1606120353
transform 1 0 13432 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_136
timestamp 1606120353
transform 1 0 13616 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__D1
timestamp 1606120353
transform 1 0 13800 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0630_
timestamp 1606120353
transform 1 0 13984 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_32_143
timestamp 1606120353
transform 1 0 14260 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_147
timestamp 1606120353
transform 1 0 14628 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0526__A
timestamp 1606120353
transform 1 0 14444 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__A1
timestamp 1606120353
transform 1 0 14812 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_151
timestamp 1606120353
transform 1 0 14996 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1606120353
transform 1 0 15180 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0593_
timestamp 1606120353
transform 1 0 15272 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1088_
timestamp 1606120353
transform 1 0 16468 0 -1 20128
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__B2
timestamp 1606120353
transform 1 0 15824 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__A2
timestamp 1606120353
transform 1 0 16192 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_32_157
timestamp 1606120353
transform 1 0 15548 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_32_162
timestamp 1606120353
transform 1 0 16008 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_32_166
timestamp 1606120353
transform 1 0 16376 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _0608_
timestamp 1606120353
transform 1 0 18952 0 -1 20128
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__A2
timestamp 1606120353
transform 1 0 18400 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_32_186
timestamp 1606120353
transform 1 0 18216 0 -1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_32_190
timestamp 1606120353
transform 1 0 18584 0 -1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1606120353
transform 1 0 20792 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_32_201
timestamp 1606120353
transform 1 0 19596 0 -1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_32_213
timestamp 1606120353
transform 1 0 20700 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_32_215
timestamp 1606120353
transform 1 0 20884 0 -1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_32_227
timestamp 1606120353
transform 1 0 21988 0 -1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_32_239
timestamp 1606120353
transform 1 0 23092 0 -1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_32_251
timestamp 1606120353
transform 1 0 24196 0 -1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_32_263
timestamp 1606120353
transform 1 0 25300 0 -1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1606120353
transform 1 0 26404 0 -1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_32_276
timestamp 1606120353
transform 1 0 26496 0 -1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1606120353
transform -1 0 28888 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_32_288
timestamp 1606120353
transform 1 0 27600 0 -1 20128
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_32_296
timestamp 1606120353
transform 1 0 28336 0 -1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1140_
timestamp 1606120353
transform 1 0 1472 0 -1 21216
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1606120353
transform 1 0 1104 0 1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1606120353
transform 1 0 1104 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__D
timestamp 1606120353
transform 1 0 1564 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__CLK
timestamp 1606120353
transform 1 0 1932 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_3
timestamp 1606120353
transform 1 0 1380 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_7
timestamp 1606120353
transform 1 0 1748 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_33_11
timestamp 1606120353
transform 1 0 2116 0 1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_34_3
timestamp 1606120353
transform 1 0 1380 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1606120353
transform 1 0 3956 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_33_23
timestamp 1606120353
transform 1 0 3220 0 1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_33_35
timestamp 1606120353
transform 1 0 4324 0 1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_34_23
timestamp 1606120353
transform 1 0 3220 0 -1 21216
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1606120353
transform 1 0 4048 0 -1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_34_44
timestamp 1606120353
transform 1 0 5152 0 -1 21216
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_34_52
timestamp 1606120353
transform 1 0 5888 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__CLK
timestamp 1606120353
transform 1 0 6072 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_34_65
timestamp 1606120353
transform 1 0 7084 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_34_62
timestamp 1606120353
transform 1 0 6808 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_34_56
timestamp 1606120353
transform 1 0 6256 0 -1 21216
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1606120353
transform 1 0 6532 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__B2
timestamp 1606120353
transform 1 0 6900 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1606120353
transform 1 0 6716 0 1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1606120353
transform 1 0 6808 0 1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_33_47
timestamp 1606120353
transform 1 0 5428 0 1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__A2
timestamp 1606120353
transform 1 0 7268 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__A
timestamp 1606120353
transform 1 0 8924 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_33_74
timestamp 1606120353
transform 1 0 7912 0 1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_33_86
timestamp 1606120353
transform 1 0 9016 0 1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_34_69
timestamp 1606120353
transform 1 0 7452 0 -1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_34_81
timestamp 1606120353
transform 1 0 8556 0 -1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_34_87
timestamp 1606120353
transform 1 0 9108 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_34_96
timestamp 1606120353
transform 1 0 9936 0 -1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_33_95
timestamp 1606120353
transform 1 0 9844 0 1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_33_91
timestamp 1606120353
transform 1 0 9476 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_clk_A
timestamp 1606120353
transform 1 0 9384 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0532__A
timestamp 1606120353
transform 1 0 9292 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__B1
timestamp 1606120353
transform 1 0 10120 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__A
timestamp 1606120353
transform 1 0 9660 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1606120353
transform 1 0 9568 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0762_
timestamp 1606120353
transform 1 0 9660 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_34_107
timestamp 1606120353
transform 1 0 10948 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_34_102
timestamp 1606120353
transform 1 0 10488 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__A2
timestamp 1606120353
transform 1 0 10764 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__A2
timestamp 1606120353
transform 1 0 10304 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0532_
timestamp 1606120353
transform 1 0 11040 0 -1 21216
box 0 -48 644 592
use sky130_fd_sc_hd__o21a_4  _0759_
timestamp 1606120353
transform 1 0 10304 0 1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_34_121
timestamp 1606120353
transform 1 0 12236 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_34_115
timestamp 1606120353
transform 1 0 11684 0 -1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_33_116
timestamp 1606120353
transform 1 0 11776 0 1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_33_112
timestamp 1606120353
transform 1 0 11408 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__A1
timestamp 1606120353
transform 1 0 12052 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__A
timestamp 1606120353
transform 1 0 12144 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0532__B
timestamp 1606120353
transform 1 0 11592 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_34_125
timestamp 1606120353
transform 1 0 12604 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_33_123
timestamp 1606120353
transform 1 0 12420 0 1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0635__B
timestamp 1606120353
transform 1 0 12420 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__A2
timestamp 1606120353
transform 1 0 12788 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1606120353
transform 1 0 12328 0 1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _0688_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 12788 0 -1 21216
box 0 -48 644 592
use sky130_fd_sc_hd__a2111oi_4  _0610_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 12972 0 1 20128
box 0 -48 2024 592
use sky130_fd_sc_hd__fill_2  FILLER_34_134
timestamp 1606120353
transform 1 0 13432 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__C1
timestamp 1606120353
transform 1 0 13616 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_34_138
timestamp 1606120353
transform 1 0 13800 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0633__A
timestamp 1606120353
transform 1 0 13984 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0526_
timestamp 1606120353
transform 1 0 14168 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_34_145
timestamp 1606120353
transform 1 0 14444 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__CLK
timestamp 1606120353
transform 1 0 14628 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_34_149
timestamp 1606120353
transform 1 0 14812 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_33_151
timestamp 1606120353
transform 1 0 14996 0 1 20128
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__D
timestamp 1606120353
transform 1 0 14996 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_34_154
timestamp 1606120353
transform 1 0 15272 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1606120353
transform 1 0 15180 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_34_162
timestamp 1606120353
transform 1 0 16008 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_34_158
timestamp 1606120353
transform 1 0 15640 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_33_157
timestamp 1606120353
transform 1 0 15548 0 1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__B1
timestamp 1606120353
transform 1 0 16192 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__A1
timestamp 1606120353
transform 1 0 15824 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0528__A
timestamp 1606120353
transform 1 0 15364 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0528_
timestamp 1606120353
transform 1 0 15364 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_33_174
timestamp 1606120353
transform 1 0 17112 0 1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1089_
timestamp 1606120353
transform 1 0 16376 0 -1 21216
box 0 -48 1748 592
use sky130_fd_sc_hd__o22a_4  _0807_
timestamp 1606120353
transform 1 0 15824 0 1 20128
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_34_185
timestamp 1606120353
transform 1 0 18124 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_33_179
timestamp 1606120353
transform 1 0 17572 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__A1
timestamp 1606120353
transform 1 0 18308 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__B1
timestamp 1606120353
transform 1 0 17388 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__A1
timestamp 1606120353
transform 1 0 17756 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1606120353
transform 1 0 17940 0 1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_34_193
timestamp 1606120353
transform 1 0 18860 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_34_189
timestamp 1606120353
transform 1 0 18492 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__B1
timestamp 1606120353
transform 1 0 19044 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__B2
timestamp 1606120353
transform 1 0 18676 0 -1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_34_197
timestamp 1606120353
transform 1 0 19228 0 -1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_33_196
timestamp 1606120353
transform 1 0 19136 0 1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__a21o_4  _0764_
timestamp 1606120353
transform 1 0 18032 0 1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1606120353
transform 1 0 20792 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_33_208
timestamp 1606120353
transform 1 0 20240 0 1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_33_220
timestamp 1606120353
transform 1 0 21344 0 1 20128
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_34_209
timestamp 1606120353
transform 1 0 20332 0 -1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_34_213
timestamp 1606120353
transform 1 0 20700 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1606120353
transform 1 0 20884 0 -1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1133_
timestamp 1606120353
transform 1 0 22356 0 -1 21216
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__D
timestamp 1606120353
transform 1 0 22356 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__CLK
timestamp 1606120353
transform 1 0 22724 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_33_228
timestamp 1606120353
transform 1 0 22080 0 1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_33_233
timestamp 1606120353
transform 1 0 22540 0 1 20128
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_33_237
timestamp 1606120353
transform 1 0 22908 0 1 20128
box 0 -48 552 592
use sky130_fd_sc_hd__decap_4  FILLER_34_227
timestamp 1606120353
transform 1 0 21988 0 -1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1606120353
transform 1 0 23552 0 1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_33_243
timestamp 1606120353
transform 1 0 23460 0 1 20128
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_33_245
timestamp 1606120353
transform 1 0 23644 0 1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_33_257
timestamp 1606120353
transform 1 0 24748 0 1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_34_250
timestamp 1606120353
transform 1 0 24104 0 -1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_34_262
timestamp 1606120353
transform 1 0 25208 0 -1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1606120353
transform 1 0 26404 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_33_269
timestamp 1606120353
transform 1 0 25852 0 1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1606120353
transform 1 0 26956 0 1 20128
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_34_274
timestamp 1606120353
transform 1 0 26312 0 -1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_34_276
timestamp 1606120353
transform 1 0 26496 0 -1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1606120353
transform -1 0 28888 0 1 20128
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1606120353
transform -1 0 28888 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_33_293
timestamp 1606120353
transform 1 0 28060 0 1 20128
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILLER_34_288
timestamp 1606120353
transform 1 0 27600 0 -1 21216
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_34_296
timestamp 1606120353
transform 1 0 28336 0 -1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1606120353
transform 1 0 1104 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1606120353
transform 1 0 1380 0 1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1606120353
transform 1 0 2484 0 1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1606120353
transform 1 0 3588 0 1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1606120353
transform 1 0 4692 0 1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__o22a_4  _0814_
timestamp 1606120353
transform 1 0 6900 0 1 21216
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1606120353
transform 1 0 6716 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__B1
timestamp 1606120353
transform 1 0 6532 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__A1
timestamp 1606120353
transform 1 0 6164 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__D
timestamp 1606120353
transform 1 0 5796 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_53
timestamp 1606120353
transform 1 0 5980 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_57
timestamp 1606120353
transform 1 0 6348 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_35_62
timestamp 1606120353
transform 1 0 6808 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0670_
timestamp 1606120353
transform 1 0 8924 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__A
timestamp 1606120353
transform 1 0 8556 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_35_77
timestamp 1606120353
transform 1 0 8188 0 1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_35_83
timestamp 1606120353
transform 1 0 8740 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_35_88
timestamp 1606120353
transform 1 0 9200 0 1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__and2_4  _0687_
timestamp 1606120353
transform 1 0 10948 0 1 21216
box 0 -48 644 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_clk
timestamp 1606120353
transform 1 0 9936 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__D
timestamp 1606120353
transform 1 0 9660 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__B
timestamp 1606120353
transform 1 0 10764 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__A
timestamp 1606120353
transform 1 0 10396 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_35_92
timestamp 1606120353
transform 1 0 9568 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_35_95
timestamp 1606120353
transform 1 0 9844 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_35_99
timestamp 1606120353
transform 1 0 10212 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_103
timestamp 1606120353
transform 1 0 10580 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__nor3_4  _0635_
timestamp 1606120353
transform 1 0 12420 0 1 21216
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1606120353
transform 1 0 12328 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0635__A
timestamp 1606120353
transform 1 0 12144 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0601__A
timestamp 1606120353
transform 1 0 11776 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_114
timestamp 1606120353
transform 1 0 11592 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_118
timestamp 1606120353
transform 1 0 11960 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0529_
timestamp 1606120353
transform 1 0 14536 0 1 21216
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0529__A
timestamp 1606120353
transform 1 0 14352 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0633__B
timestamp 1606120353
transform 1 0 13800 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_136
timestamp 1606120353
transform 1 0 13616 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_35_140
timestamp 1606120353
transform 1 0 13984 0 1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__and2_4  _0769_
timestamp 1606120353
transform 1 0 16560 0 1 21216
box 0 -48 644 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_clk
timestamp 1606120353
transform 1 0 16284 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0525__B
timestamp 1606120353
transform 1 0 15548 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__A
timestamp 1606120353
transform 1 0 16100 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_155
timestamp 1606120353
transform 1 0 15364 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_35_159
timestamp 1606120353
transform 1 0 15732 0 1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_35_175
timestamp 1606120353
transform 1 0 17204 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0770_
timestamp 1606120353
transform 1 0 18032 0 1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1606120353
transform 1 0 17940 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__A
timestamp 1606120353
transform 1 0 17388 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__A1
timestamp 1606120353
transform 1 0 17756 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__A2
timestamp 1606120353
transform 1 0 19320 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_179
timestamp 1606120353
transform 1 0 17572 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_196
timestamp 1606120353
transform 1 0 19136 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__A2
timestamp 1606120353
transform 1 0 19688 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_35_200
timestamp 1606120353
transform 1 0 19504 0 1 21216
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_35_204
timestamp 1606120353
transform 1 0 19872 0 1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_35_216
timestamp 1606120353
transform 1 0 20976 0 1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_35_228
timestamp 1606120353
transform 1 0 22080 0 1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_35_240
timestamp 1606120353
transform 1 0 23184 0 1 21216
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1606120353
transform 1 0 23552 0 1 21216
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_35_245
timestamp 1606120353
transform 1 0 23644 0 1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_35_257
timestamp 1606120353
transform 1 0 24748 0 1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_35_269
timestamp 1606120353
transform 1 0 25852 0 1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1606120353
transform 1 0 26956 0 1 21216
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1606120353
transform -1 0 28888 0 1 21216
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_35_293
timestamp 1606120353
transform 1 0 28060 0 1 21216
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1606120353
transform 1 0 1104 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1606120353
transform 1 0 1380 0 -1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1606120353
transform 1 0 2484 0 -1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1606120353
transform 1 0 3956 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1606120353
transform 1 0 3588 0 -1 22304
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1606120353
transform 1 0 4048 0 -1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_36_44
timestamp 1606120353
transform 1 0 5152 0 -1 22304
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1108_
timestamp 1606120353
transform 1 0 6072 0 -1 22304
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_2  FILLER_36_52
timestamp 1606120353
transform 1 0 5888 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0813_
timestamp 1606120353
transform 1 0 8556 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_36_73
timestamp 1606120353
transform 1 0 7820 0 -1 22304
box 0 -48 736 592
use sky130_fd_sc_hd__decap_6  FILLER_36_84
timestamp 1606120353
transform 1 0 8832 0 -1 22304
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1214_
timestamp 1606120353
transform 1 0 9660 0 -1 22304
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1606120353
transform 1 0 9568 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__CLK
timestamp 1606120353
transform 1 0 9384 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0601_
timestamp 1606120353
transform 1 0 12144 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__and2_4  _0633_
timestamp 1606120353
transform 1 0 13156 0 -1 22304
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0635__C
timestamp 1606120353
transform 1 0 12604 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__C
timestamp 1606120353
transform 1 0 11960 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0607__A
timestamp 1606120353
transform 1 0 12972 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_36_112
timestamp 1606120353
transform 1 0 11408 0 -1 22304
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_36_123
timestamp 1606120353
transform 1 0 12420 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_127
timestamp 1606120353
transform 1 0 12788 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0525_
timestamp 1606120353
transform 1 0 15272 0 -1 22304
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1606120353
transform 1 0 15180 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0611__B
timestamp 1606120353
transform 1 0 13984 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0611__A
timestamp 1606120353
transform 1 0 14352 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_138
timestamp 1606120353
transform 1 0 13800 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_142
timestamp 1606120353
transform 1 0 14168 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_36_146
timestamp 1606120353
transform 1 0 14536 0 -1 22304
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_36_152
timestamp 1606120353
transform 1 0 15088 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0801_
timestamp 1606120353
transform 1 0 16836 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__B
timestamp 1606120353
transform 1 0 16560 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0525__A
timestamp 1606120353
transform 1 0 16100 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_161
timestamp 1606120353
transform 1 0 15916 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_36_165
timestamp 1606120353
transform 1 0 16284 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_36_170
timestamp 1606120353
transform 1 0 16744 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_36_174
timestamp 1606120353
transform 1 0 17112 0 -1 22304
box 0 -48 736 592
use sky130_fd_sc_hd__o22a_4  _0804_
timestamp 1606120353
transform 1 0 18308 0 -1 22304
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__B1
timestamp 1606120353
transform 1 0 18032 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_36_182
timestamp 1606120353
transform 1 0 17848 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_36_186
timestamp 1606120353
transform 1 0 18216 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1606120353
transform 1 0 20792 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_36_201
timestamp 1606120353
transform 1 0 19596 0 -1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_36_213
timestamp 1606120353
transform 1 0 20700 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_36_215
timestamp 1606120353
transform 1 0 20884 0 -1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_36_227
timestamp 1606120353
transform 1 0 21988 0 -1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_36_239
timestamp 1606120353
transform 1 0 23092 0 -1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_36_251
timestamp 1606120353
transform 1 0 24196 0 -1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_36_263
timestamp 1606120353
transform 1 0 25300 0 -1 22304
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1606120353
transform 1 0 26404 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__CLK
timestamp 1606120353
transform 1 0 26128 0 -1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_36_271
timestamp 1606120353
transform 1 0 26036 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_36_274
timestamp 1606120353
transform 1 0 26312 0 -1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_36_276
timestamp 1606120353
transform 1 0 26496 0 -1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1606120353
transform -1 0 28888 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_36_288
timestamp 1606120353
transform 1 0 27600 0 -1 22304
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_36_296
timestamp 1606120353
transform 1 0 28336 0 -1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1606120353
transform 1 0 1104 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1606120353
transform 1 0 1380 0 1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1606120353
transform 1 0 2484 0 1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1606120353
transform 1 0 3588 0 1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_37_39
timestamp 1606120353
transform 1 0 4692 0 1 22304
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1106_
timestamp 1606120353
transform 1 0 6808 0 1 22304
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1606120353
transform 1 0 6716 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A1
timestamp 1606120353
transform 1 0 6164 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__B2
timestamp 1606120353
transform 1 0 6532 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A2
timestamp 1606120353
transform 1 0 5796 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__B1
timestamp 1606120353
transform 1 0 5428 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_49
timestamp 1606120353
transform 1 0 5612 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_53
timestamp 1606120353
transform 1 0 5980 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1606120353
transform 1 0 6348 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__A
timestamp 1606120353
transform 1 0 9108 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__A
timestamp 1606120353
transform 1 0 8740 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_81
timestamp 1606120353
transform 1 0 8556 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_85
timestamp 1606120353
transform 1 0 8924 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0806_
timestamp 1606120353
transform 1 0 9292 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_37_92
timestamp 1606120353
transform 1 0 9568 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0537__B1
timestamp 1606120353
transform 1 0 9752 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_96
timestamp 1606120353
transform 1 0 9936 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0537__A1
timestamp 1606120353
transform 1 0 10120 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0662_
timestamp 1606120353
transform 1 0 10304 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_37_103
timestamp 1606120353
transform 1 0 10580 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0537__A2
timestamp 1606120353
transform 1 0 10764 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_107
timestamp 1606120353
transform 1 0 10948 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0662__A
timestamp 1606120353
transform 1 0 11132 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0607_
timestamp 1606120353
transform 1 0 12420 0 1 22304
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1606120353
transform 1 0 12328 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0607__B
timestamp 1606120353
transform 1 0 13248 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__A
timestamp 1606120353
transform 1 0 11960 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__B
timestamp 1606120353
transform 1 0 11592 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_37_111
timestamp 1606120353
transform 1 0 11316 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_37_116
timestamp 1606120353
transform 1 0 11776 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_120
timestamp 1606120353
transform 1 0 12144 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_130
timestamp 1606120353
transform 1 0 13064 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__nor3_4  _0611_
timestamp 1606120353
transform 1 0 13800 0 1 22304
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0519__A
timestamp 1606120353
transform 1 0 13616 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__B
timestamp 1606120353
transform 1 0 15272 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_134
timestamp 1606120353
transform 1 0 13432 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_37_151
timestamp 1606120353
transform 1 0 14996 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__A
timestamp 1606120353
transform 1 0 15640 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__C
timestamp 1606120353
transform 1 0 16008 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__D
timestamp 1606120353
transform 1 0 16376 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_clk_A
timestamp 1606120353
transform 1 0 16744 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_156
timestamp 1606120353
transform 1 0 15456 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_160
timestamp 1606120353
transform 1 0 15824 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_164
timestamp 1606120353
transform 1 0 16192 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_37_168
timestamp 1606120353
transform 1 0 16560 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_37_172
timestamp 1606120353
transform 1 0 16928 0 1 22304
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1101_
timestamp 1606120353
transform 1 0 18032 0 1 22304
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1606120353
transform 1 0 17940 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__D
timestamp 1606120353
transform 1 0 17756 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_37_180
timestamp 1606120353
transform 1 0 17664 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_37_203
timestamp 1606120353
transform 1 0 19780 0 1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_37_215
timestamp 1606120353
transform 1 0 20884 0 1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_37_227
timestamp 1606120353
transform 1 0 21988 0 1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_37_239
timestamp 1606120353
transform 1 0 23092 0 1 22304
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1606120353
transform 1 0 23552 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_37_243
timestamp 1606120353
transform 1 0 23460 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_37_245
timestamp 1606120353
transform 1 0 23644 0 1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_37_257
timestamp 1606120353
transform 1 0 24748 0 1 22304
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1142_
timestamp 1606120353
transform 1 0 26128 0 1 22304
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__D
timestamp 1606120353
transform 1 0 25944 0 1 22304
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_37_269
timestamp 1606120353
transform 1 0 25852 0 1 22304
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1606120353
transform -1 0 28888 0 1 22304
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_37_291
timestamp 1606120353
transform 1 0 27876 0 1 22304
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1606120353
transform 1 0 1104 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1606120353
transform 1 0 1380 0 -1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1606120353
transform 1 0 2484 0 -1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1606120353
transform 1 0 3956 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1606120353
transform 1 0 3588 0 -1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1606120353
transform 1 0 4048 0 -1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_38_44
timestamp 1606120353
transform 1 0 5152 0 -1 23392
box 0 -48 736 592
use sky130_fd_sc_hd__o22a_4  _0811_
timestamp 1606120353
transform 1 0 6164 0 -1 23392
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_3  FILLER_38_52
timestamp 1606120353
transform 1 0 5888 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0799_
timestamp 1606120353
transform 1 0 8556 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__D
timestamp 1606120353
transform 1 0 7636 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_69
timestamp 1606120353
transform 1 0 7452 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_38_73
timestamp 1606120353
transform 1 0 7820 0 -1 23392
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_38_84
timestamp 1606120353
transform 1 0 8832 0 -1 23392
box 0 -48 736 592
use sky130_fd_sc_hd__o21a_4  _0537_
timestamp 1606120353
transform 1 0 10120 0 -1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1606120353
transform 1 0 9568 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_38_93
timestamp 1606120353
transform 1 0 9660 0 -1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_38_97
timestamp 1606120353
transform 1 0 10028 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_38_110
timestamp 1606120353
transform 1 0 11224 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__nor3_4  _0636_
timestamp 1606120353
transform 1 0 11960 0 -1 23392
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0638__A
timestamp 1606120353
transform 1 0 11776 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0692__A
timestamp 1606120353
transform 1 0 11408 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_114
timestamp 1606120353
transform 1 0 11592 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_131
timestamp 1606120353
transform 1 0 13156 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_135
timestamp 1606120353
transform 1 0 13524 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0626__C
timestamp 1606120353
transform 1 0 13340 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0611__C
timestamp 1606120353
transform 1 0 13708 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0519_
timestamp 1606120353
transform 1 0 13892 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_38_150
timestamp 1606120353
transform 1 0 14904 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_38_146
timestamp 1606120353
transform 1 0 14536 0 -1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_38_142
timestamp 1606120353
transform 1 0 14168 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0612__C
timestamp 1606120353
transform 1 0 14352 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__B
timestamp 1606120353
transform 1 0 14996 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1606120353
transform 1 0 15180 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _0602_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 15272 0 -1 23392
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__A
timestamp 1606120353
transform 1 0 16284 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_38_163
timestamp 1606120353
transform 1 0 16100 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_38_167
timestamp 1606120353
transform 1 0 16468 0 -1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__CLK
timestamp 1606120353
transform 1 0 18032 0 -1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_38_179
timestamp 1606120353
transform 1 0 17572 0 -1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_38_183
timestamp 1606120353
transform 1 0 17940 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_38_186
timestamp 1606120353
transform 1 0 18216 0 -1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_38_198
timestamp 1606120353
transform 1 0 19320 0 -1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1606120353
transform 1 0 20792 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_38_210
timestamp 1606120353
transform 1 0 20424 0 -1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_38_215
timestamp 1606120353
transform 1 0 20884 0 -1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_38_227
timestamp 1606120353
transform 1 0 21988 0 -1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_38_239
timestamp 1606120353
transform 1 0 23092 0 -1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_38_251
timestamp 1606120353
transform 1 0 24196 0 -1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_38_263
timestamp 1606120353
transform 1 0 25300 0 -1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1606120353
transform 1 0 26404 0 -1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_38_276
timestamp 1606120353
transform 1 0 26496 0 -1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1606120353
transform -1 0 28888 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_38_288
timestamp 1606120353
transform 1 0 27600 0 -1 23392
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_38_296
timestamp 1606120353
transform 1 0 28336 0 -1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1606120353
transform 1 0 1104 0 1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1606120353
transform 1 0 1104 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1606120353
transform 1 0 1380 0 1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1606120353
transform 1 0 2484 0 1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1606120353
transform 1 0 1380 0 -1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1606120353
transform 1 0 2484 0 -1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1606120353
transform 1 0 3956 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1606120353
transform 1 0 3588 0 1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1606120353
transform 1 0 4692 0 1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1606120353
transform 1 0 3588 0 -1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1606120353
transform 1 0 4048 0 -1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1606120353
transform 1 0 5152 0 -1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1606120353
transform 1 0 6716 0 1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__CLK
timestamp 1606120353
transform 1 0 6992 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__CLK
timestamp 1606120353
transform 1 0 6992 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_39_51
timestamp 1606120353
transform 1 0 5796 0 1 23392
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_39_59
timestamp 1606120353
transform 1 0 6532 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_62
timestamp 1606120353
transform 1 0 6808 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_39_66
timestamp 1606120353
transform 1 0 7176 0 1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_40_56
timestamp 1606120353
transform 1 0 6256 0 -1 24480
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_40_66
timestamp 1606120353
transform 1 0 7176 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0661_
timestamp 1606120353
transform 1 0 8648 0 1 23392
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0661__A
timestamp 1606120353
transform 1 0 8464 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__A1
timestamp 1606120353
transform 1 0 7360 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__A2
timestamp 1606120353
transform 1 0 7728 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_78
timestamp 1606120353
transform 1 0 8280 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_70
timestamp 1606120353
transform 1 0 7544 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_40_74
timestamp 1606120353
transform 1 0 7912 0 -1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_40_86
timestamp 1606120353
transform 1 0 9016 0 -1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_40_93
timestamp 1606120353
transform 1 0 9660 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_39_91
timestamp 1606120353
transform 1 0 9476 0 1 23392
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__B2
timestamp 1606120353
transform 1 0 9384 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__B1_N
timestamp 1606120353
transform 1 0 9844 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1606120353
transform 1 0 9568 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_40_103
timestamp 1606120353
transform 1 0 10580 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_40_97
timestamp 1606120353
transform 1 0 10028 0 -1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_39_101
timestamp 1606120353
transform 1 0 10396 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__D
timestamp 1606120353
transform 1 0 10212 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__B1
timestamp 1606120353
transform 1 0 10580 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__A4
timestamp 1606120353
transform 1 0 10396 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_107
timestamp 1606120353
transform 1 0 10948 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_109
timestamp 1606120353
transform 1 0 11132 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_105
timestamp 1606120353
transform 1 0 10764 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__B1
timestamp 1606120353
transform 1 0 10948 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__A3
timestamp 1606120353
transform 1 0 10764 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__A2
timestamp 1606120353
transform 1 0 11132 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_40_118
timestamp 1606120353
transform 1 0 11960 0 -1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_39_118
timestamp 1606120353
transform 1 0 11960 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_39_113
timestamp 1606120353
transform 1 0 11500 0 1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0626__B
timestamp 1606120353
transform 1 0 11776 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0638__B
timestamp 1606120353
transform 1 0 12144 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0692__B
timestamp 1606120353
transform 1 0 11316 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0692_
timestamp 1606120353
transform 1 0 11316 0 -1 24480
box 0 -48 644 592
use sky130_fd_sc_hd__fill_1  FILLER_40_125
timestamp 1606120353
transform 1 0 12604 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_40_122
timestamp 1606120353
transform 1 0 12328 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_39_130
timestamp 1606120353
transform 1 0 13064 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__B1
timestamp 1606120353
transform 1 0 12420 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0626__A
timestamp 1606120353
transform 1 0 13248 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1606120353
transform 1 0 12328 0 1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _0638_
timestamp 1606120353
transform 1 0 12420 0 1 23392
box 0 -48 644 592
use sky130_fd_sc_hd__nor3_4  _0626_
timestamp 1606120353
transform 1 0 12696 0 -1 24480
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_40_143
timestamp 1606120353
transform 1 0 14260 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_139
timestamp 1606120353
transform 1 0 13892 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_39_134
timestamp 1606120353
transform 1 0 13432 0 1 23392
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0612__B
timestamp 1606120353
transform 1 0 14076 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0612__A
timestamp 1606120353
transform 1 0 13800 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_151
timestamp 1606120353
transform 1 0 14996 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_147
timestamp 1606120353
transform 1 0 14628 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__C
timestamp 1606120353
transform 1 0 14812 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0612__D
timestamp 1606120353
transform 1 0 14444 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1606120353
transform 1 0 15180 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _0599_
timestamp 1606120353
transform 1 0 15272 0 -1 24480
box 0 -48 828 592
use sky130_fd_sc_hd__nor4_4  _0612_
timestamp 1606120353
transform 1 0 13984 0 1 23392
box 0 -48 1564 592
use sky130_fd_sc_hd__fill_2  FILLER_39_161
timestamp 1606120353
transform 1 0 15916 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_157
timestamp 1606120353
transform 1 0 15548 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__A
timestamp 1606120353
transform 1 0 15732 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_167
timestamp 1606120353
transform 1 0 16468 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_40_163
timestamp 1606120353
transform 1 0 16100 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_39_168
timestamp 1606120353
transform 1 0 16560 0 1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0543__A
timestamp 1606120353
transform 1 0 16652 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__D
timestamp 1606120353
transform 1 0 16284 0 -1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__C
timestamp 1606120353
transform 1 0 16100 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0808_
timestamp 1606120353
transform 1 0 16284 0 1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_40_174
timestamp 1606120353
transform 1 0 17112 0 -1 24480
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_39_173
timestamp 1606120353
transform 1 0 17020 0 1 23392
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0598__A
timestamp 1606120353
transform 1 0 16836 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0598_
timestamp 1606120353
transform 1 0 16836 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0592_
timestamp 1606120353
transform 1 0 17848 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1606120353
transform 1 0 17940 0 1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0592__A
timestamp 1606120353
transform 1 0 18216 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_181
timestamp 1606120353
transform 1 0 17756 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_39_184
timestamp 1606120353
transform 1 0 18032 0 1 23392
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_39_188
timestamp 1606120353
transform 1 0 18400 0 1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_40_185
timestamp 1606120353
transform 1 0 18124 0 -1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_40_197
timestamp 1606120353
transform 1 0 19228 0 -1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1606120353
transform 1 0 20792 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_39_200
timestamp 1606120353
transform 1 0 19504 0 1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_39_212
timestamp 1606120353
transform 1 0 20608 0 1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_40_209
timestamp 1606120353
transform 1 0 20332 0 -1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_40_213
timestamp 1606120353
transform 1 0 20700 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_40_215
timestamp 1606120353
transform 1 0 20884 0 -1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_39_224
timestamp 1606120353
transform 1 0 21712 0 1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_39_236
timestamp 1606120353
transform 1 0 22816 0 1 23392
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_40_227
timestamp 1606120353
transform 1 0 21988 0 -1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_40_239
timestamp 1606120353
transform 1 0 23092 0 -1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1606120353
transform 1 0 23552 0 1 23392
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_39_245
timestamp 1606120353
transform 1 0 23644 0 1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_39_257
timestamp 1606120353
transform 1 0 24748 0 1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_40_251
timestamp 1606120353
transform 1 0 24196 0 -1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_40_263
timestamp 1606120353
transform 1 0 25300 0 -1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1606120353
transform 1 0 26404 0 -1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_39_269
timestamp 1606120353
transform 1 0 25852 0 1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1606120353
transform 1 0 26956 0 1 23392
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_40_276
timestamp 1606120353
transform 1 0 26496 0 -1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1606120353
transform -1 0 28888 0 1 23392
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1606120353
transform -1 0 28888 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_39_293
timestamp 1606120353
transform 1 0 28060 0 1 23392
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILLER_40_288
timestamp 1606120353
transform 1 0 27600 0 -1 24480
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_40_296
timestamp 1606120353
transform 1 0 28336 0 -1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1606120353
transform 1 0 1104 0 1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0486__B
timestamp 1606120353
transform 1 0 1564 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0486__A
timestamp 1606120353
transform 1 0 1932 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1606120353
transform 1 0 1380 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_7
timestamp 1606120353
transform 1 0 1748 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_41_11
timestamp 1606120353
transform 1 0 2116 0 1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_41_23
timestamp 1606120353
transform 1 0 3220 0 1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_41_35
timestamp 1606120353
transform 1 0 4324 0 1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1606120353
transform 1 0 6716 0 1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__B1
timestamp 1606120353
transform 1 0 7176 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__B2
timestamp 1606120353
transform 1 0 6532 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__D
timestamp 1606120353
transform 1 0 6164 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_41_47
timestamp 1606120353
transform 1 0 5428 0 1 24480
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_41_57
timestamp 1606120353
transform 1 0 6348 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_41_62
timestamp 1606120353
transform 1 0 6808 0 1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__o22a_4  _0780_
timestamp 1606120353
transform 1 0 7360 0 1 24480
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__A2
timestamp 1606120353
transform 1 0 9016 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_41_82
timestamp 1606120353
transform 1 0 8648 0 1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_41_88
timestamp 1606120353
transform 1 0 9200 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0660_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 9568 0 1 24480
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__A1
timestamp 1606120353
transform 1 0 9384 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0496__A
timestamp 1606120353
transform 1 0 10948 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_105
timestamp 1606120353
transform 1 0 10764 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_109
timestamp 1606120353
transform 1 0 11132 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0693_
timestamp 1606120353
transform 1 0 12420 0 1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1606120353
transform 1 0 12328 0 1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__A1
timestamp 1606120353
transform 1 0 11316 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__A2
timestamp 1606120353
transform 1 0 12144 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__C1
timestamp 1606120353
transform 1 0 11776 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_41_113
timestamp 1606120353
transform 1 0 11500 0 1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_41_118
timestamp 1606120353
transform 1 0 11960 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0627_
timestamp 1606120353
transform 1 0 14260 0 1 24480
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0627__A
timestamp 1606120353
transform 1 0 14076 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__A
timestamp 1606120353
transform 1 0 13708 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__B
timestamp 1606120353
transform 1 0 15272 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_135
timestamp 1606120353
transform 1 0 13524 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_139
timestamp 1606120353
transform 1 0 13892 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_152
timestamp 1606120353
transform 1 0 15088 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_156
timestamp 1606120353
transform 1 0 15456 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_160
timestamp 1606120353
transform 1 0 15824 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__A1
timestamp 1606120353
transform 1 0 15640 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0543_
timestamp 1606120353
transform 1 0 16008 0 1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_41_165
timestamp 1606120353
transform 1 0 16284 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_169
timestamp 1606120353
transform 1 0 16652 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__A2
timestamp 1606120353
transform 1 0 16468 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__D
timestamp 1606120353
transform 1 0 16836 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_173
timestamp 1606120353
transform 1 0 17020 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__CLK
timestamp 1606120353
transform 1 0 17204 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0664_
timestamp 1606120353
transform 1 0 18032 0 1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1606120353
transform 1 0 17940 0 1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0664__A
timestamp 1606120353
transform 1 0 18492 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__CLK
timestamp 1606120353
transform 1 0 17572 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_177
timestamp 1606120353
transform 1 0 17388 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_181
timestamp 1606120353
transform 1 0 17756 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_41_187
timestamp 1606120353
transform 1 0 18308 0 1 24480
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_41_191
timestamp 1606120353
transform 1 0 18676 0 1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_41_203
timestamp 1606120353
transform 1 0 19780 0 1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_41_215
timestamp 1606120353
transform 1 0 20884 0 1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_41_227
timestamp 1606120353
transform 1 0 21988 0 1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_41_239
timestamp 1606120353
transform 1 0 23092 0 1 24480
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1606120353
transform 1 0 23552 0 1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_41_243
timestamp 1606120353
transform 1 0 23460 0 1 24480
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_41_245
timestamp 1606120353
transform 1 0 23644 0 1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_41_257
timestamp 1606120353
transform 1 0 24748 0 1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_41_269
timestamp 1606120353
transform 1 0 25852 0 1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1606120353
transform 1 0 26956 0 1 24480
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1606120353
transform -1 0 28888 0 1 24480
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_41_293
timestamp 1606120353
transform 1 0 28060 0 1 24480
box 0 -48 552 592
use sky130_fd_sc_hd__or2_4  _0486_
timestamp 1606120353
transform 1 0 1380 0 -1 25568
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1606120353
transform 1 0 1104 0 -1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_42_10
timestamp 1606120353
transform 1 0 2024 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_42_22
timestamp 1606120353
transform 1 0 3128 0 -1 25568
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1606120353
transform 1 0 3956 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__B2
timestamp 1606120353
transform 1 0 4692 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_42_30
timestamp 1606120353
transform 1 0 3864 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_42_32
timestamp 1606120353
transform 1 0 4048 0 -1 25568
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_42_38
timestamp 1606120353
transform 1 0 4600 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_42_41
timestamp 1606120353
transform 1 0 4876 0 -1 25568
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1091_
timestamp 1606120353
transform 1 0 7084 0 -1 25568
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__D
timestamp 1606120353
transform 1 0 5244 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__CLK
timestamp 1606120353
transform 1 0 5612 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__CLK
timestamp 1606120353
transform 1 0 6900 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_47
timestamp 1606120353
transform 1 0 5428 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_42_51
timestamp 1606120353
transform 1 0 5796 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__B1
timestamp 1606120353
transform 1 0 9016 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_84
timestamp 1606120353
transform 1 0 8832 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_88
timestamp 1606120353
transform 1 0 9200 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_42_97
timestamp 1606120353
transform 1 0 10028 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_42_93
timestamp 1606120353
transform 1 0 9660 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__A2
timestamp 1606120353
transform 1 0 9384 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__A1
timestamp 1606120353
transform 1 0 9844 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1606120353
transform 1 0 9568 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0496_
timestamp 1606120353
transform 1 0 10120 0 -1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_42_107
timestamp 1606120353
transform 1 0 10948 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_42_101
timestamp 1606120353
transform 1 0 10396 0 -1 25568
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__C
timestamp 1606120353
transform 1 0 10764 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__o41a_4  _0649_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 11132 0 -1 25568
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0648__B1
timestamp 1606120353
transform 1 0 12880 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__A2
timestamp 1606120353
transform 1 0 13248 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_126
timestamp 1606120353
transform 1 0 12696 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_130
timestamp 1606120353
transform 1 0 13064 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0647_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 13432 0 -1 25568
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1606120353
transform 1 0 15180 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__A
timestamp 1606120353
transform 1 0 14444 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__D
timestamp 1606120353
transform 1 0 14812 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_143
timestamp 1606120353
transform 1 0 14260 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_147
timestamp 1606120353
transform 1 0 14628 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_151
timestamp 1606120353
transform 1 0 14996 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_42_154
timestamp 1606120353
transform 1 0 15272 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1107_
timestamp 1606120353
transform 1 0 16100 0 -1 25568
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0617__B
timestamp 1606120353
transform 1 0 15456 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__A1
timestamp 1606120353
transform 1 0 15916 0 -1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_42_158
timestamp 1606120353
transform 1 0 15640 0 -1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_42_182
timestamp 1606120353
transform 1 0 17848 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_42_194
timestamp 1606120353
transform 1 0 18952 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1606120353
transform 1 0 20792 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_42_206
timestamp 1606120353
transform 1 0 20056 0 -1 25568
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_42_215
timestamp 1606120353
transform 1 0 20884 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_42_227
timestamp 1606120353
transform 1 0 21988 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_42_239
timestamp 1606120353
transform 1 0 23092 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_42_251
timestamp 1606120353
transform 1 0 24196 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_42_263
timestamp 1606120353
transform 1 0 25300 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1606120353
transform 1 0 26404 0 -1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_42_276
timestamp 1606120353
transform 1 0 26496 0 -1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1606120353
transform -1 0 28888 0 -1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_42_288
timestamp 1606120353
transform 1 0 27600 0 -1 25568
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_42_296
timestamp 1606120353
transform 1 0 28336 0 -1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1606120353
transform 1 0 1104 0 1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__D
timestamp 1606120353
transform 1 0 1564 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__CLK
timestamp 1606120353
transform 1 0 1932 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1606120353
transform 1 0 1380 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_7
timestamp 1606120353
transform 1 0 1748 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_43_11
timestamp 1606120353
transform 1 0 2116 0 1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__o22a_4  _0810_
timestamp 1606120353
transform 1 0 4692 0 1 25568
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__A1
timestamp 1606120353
transform 1 0 4508 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__A2
timestamp 1606120353
transform 1 0 4140 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__B1
timestamp 1606120353
transform 1 0 3772 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_43_23
timestamp 1606120353
transform 1 0 3220 0 1 25568
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_43_31
timestamp 1606120353
transform 1 0 3956 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_35
timestamp 1606120353
transform 1 0 4324 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1606120353
transform 1 0 6716 0 1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__A3
timestamp 1606120353
transform 1 0 7084 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__A2
timestamp 1606120353
transform 1 0 6532 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_43_53
timestamp 1606120353
transform 1 0 5980 0 1 25568
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILLER_43_62
timestamp 1606120353
transform 1 0 6808 0 1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__a2bb2o_4  _0778_
timestamp 1606120353
transform 1 0 8372 0 1 25568
box 0 -48 1472 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__A
timestamp 1606120353
transform 1 0 8188 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__A2_N
timestamp 1606120353
transform 1 0 7820 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__A1_N
timestamp 1606120353
transform 1 0 7452 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_67
timestamp 1606120353
transform 1 0 7268 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_71
timestamp 1606120353
transform 1 0 7636 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_75
timestamp 1606120353
transform 1 0 8004 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0631_
timestamp 1606120353
transform 1 0 10764 0 1 25568
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__B1
timestamp 1606120353
transform 1 0 10028 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__A
timestamp 1606120353
transform 1 0 10580 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_95
timestamp 1606120353
transform 1 0 9844 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_43_99
timestamp 1606120353
transform 1 0 10212 0 1 25568
box 0 -48 368 592
use sky130_fd_sc_hd__a21oi_4  _0648_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 12420 0 1 25568
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1606120353
transform 1 0 12328 0 1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0648__A1
timestamp 1606120353
transform 1 0 12144 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__A1
timestamp 1606120353
transform 1 0 11776 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_114
timestamp 1606120353
transform 1 0 11592 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_118
timestamp 1606120353
transform 1 0 11960 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0613_
timestamp 1606120353
transform 1 0 14352 0 1 25568
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__C
timestamp 1606120353
transform 1 0 14168 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__B
timestamp 1606120353
transform 1 0 13800 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_136
timestamp 1606120353
transform 1 0 13616 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_140
timestamp 1606120353
transform 1 0 13984 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_153
timestamp 1606120353
transform 1 0 15180 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _0812_
timestamp 1606120353
transform 1 0 15916 0 1 25568
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__B1
timestamp 1606120353
transform 1 0 15732 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0617__A
timestamp 1606120353
transform 1 0 15364 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_157
timestamp 1606120353
transform 1 0 15548 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_175
timestamp 1606120353
transform 1 0 17204 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1606120353
transform 1 0 17940 0 1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__A
timestamp 1606120353
transform 1 0 17388 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__B
timestamp 1606120353
transform 1 0 17756 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__D
timestamp 1606120353
transform 1 0 18216 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__CLK
timestamp 1606120353
transform 1 0 18584 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_179
timestamp 1606120353
transform 1 0 17572 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_184
timestamp 1606120353
transform 1 0 18032 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_43_188
timestamp 1606120353
transform 1 0 18400 0 1 25568
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_43_192
timestamp 1606120353
transform 1 0 18768 0 1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_43_204
timestamp 1606120353
transform 1 0 19872 0 1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_43_216
timestamp 1606120353
transform 1 0 20976 0 1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_43_228
timestamp 1606120353
transform 1 0 22080 0 1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_43_240
timestamp 1606120353
transform 1 0 23184 0 1 25568
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1606120353
transform 1 0 23552 0 1 25568
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_43_245
timestamp 1606120353
transform 1 0 23644 0 1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_43_257
timestamp 1606120353
transform 1 0 24748 0 1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_43_269
timestamp 1606120353
transform 1 0 25852 0 1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1606120353
transform 1 0 26956 0 1 25568
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1606120353
transform -1 0 28888 0 1 25568
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_43_293
timestamp 1606120353
transform 1 0 28060 0 1 25568
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1165_
timestamp 1606120353
transform 1 0 1380 0 -1 26656
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1606120353
transform 1 0 1104 0 -1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_44_22
timestamp 1606120353
transform 1 0 3128 0 -1 26656
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1606120353
transform 1 0 3956 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__B2
timestamp 1606120353
transform 1 0 4692 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__D
timestamp 1606120353
transform 1 0 5060 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_44_30
timestamp 1606120353
transform 1 0 3864 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_44_32
timestamp 1606120353
transform 1 0 4048 0 -1 26656
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_44_38
timestamp 1606120353
transform 1 0 4600 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_44_41
timestamp 1606120353
transform 1 0 4876 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1105_
timestamp 1606120353
transform 1 0 5244 0 -1 26656
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  FILLER_44_64
timestamp 1606120353
transform 1 0 6992 0 -1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_44_69
timestamp 1606120353
transform 1 0 7452 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__B1
timestamp 1606120353
transform 1 0 7268 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__B1
timestamp 1606120353
transform 1 0 7636 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_73
timestamp 1606120353
transform 1 0 7820 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__A2
timestamp 1606120353
transform 1 0 8004 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_77
timestamp 1606120353
transform 1 0 8188 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__B2
timestamp 1606120353
transform 1 0 8372 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0815_
timestamp 1606120353
transform 1 0 8556 0 -1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_44_84
timestamp 1606120353
transform 1 0 8832 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__B1
timestamp 1606120353
transform 1 0 9016 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_88
timestamp 1606120353
transform 1 0 9200 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__a32o_4  _0712_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 9844 0 -1 26656
box 0 -48 1564 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1606120353
transform 1 0 9568 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__A2_N
timestamp 1606120353
transform 1 0 9384 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_93
timestamp 1606120353
transform 1 0 9660 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__a211o_4  _0632_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 12420 0 -1 26656
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__C
timestamp 1606120353
transform 1 0 12236 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0648__A2
timestamp 1606120353
transform 1 0 11868 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_44_112
timestamp 1606120353
transform 1 0 11408 0 -1 26656
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_44_116
timestamp 1606120353
transform 1 0 11776 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_44_119
timestamp 1606120353
transform 1 0 12052 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0617_
timestamp 1606120353
transform 1 0 15272 0 -1 26656
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1606120353
transform 1 0 15180 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__A
timestamp 1606120353
transform 1 0 14076 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__C
timestamp 1606120353
transform 1 0 14444 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__B
timestamp 1606120353
transform 1 0 14812 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_44_137
timestamp 1606120353
transform 1 0 13708 0 -1 26656
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_44_143
timestamp 1606120353
transform 1 0 14260 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_147
timestamp 1606120353
transform 1 0 14628 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_151
timestamp 1606120353
transform 1 0 14996 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0776_
timestamp 1606120353
transform 1 0 17296 0 -1 26656
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__C
timestamp 1606120353
transform 1 0 16836 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__D
timestamp 1606120353
transform 1 0 16100 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__B2
timestamp 1606120353
transform 1 0 16468 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_161
timestamp 1606120353
transform 1 0 15916 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_165
timestamp 1606120353
transform 1 0 16284 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_169
timestamp 1606120353
transform 1 0 16652 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_44_173
timestamp 1606120353
transform 1 0 17020 0 -1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0629__A
timestamp 1606120353
transform 1 0 18860 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__D
timestamp 1606120353
transform 1 0 18124 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__D
timestamp 1606120353
transform 1 0 18492 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_183
timestamp 1606120353
transform 1 0 17940 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_187
timestamp 1606120353
transform 1 0 18308 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_44_191
timestamp 1606120353
transform 1 0 18676 0 -1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_44_195
timestamp 1606120353
transform 1 0 19044 0 -1 26656
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1606120353
transform 1 0 20792 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_44_207
timestamp 1606120353
transform 1 0 20148 0 -1 26656
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_44_213
timestamp 1606120353
transform 1 0 20700 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_44_215
timestamp 1606120353
transform 1 0 20884 0 -1 26656
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_44_227
timestamp 1606120353
transform 1 0 21988 0 -1 26656
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_44_239
timestamp 1606120353
transform 1 0 23092 0 -1 26656
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_44_251
timestamp 1606120353
transform 1 0 24196 0 -1 26656
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_44_263
timestamp 1606120353
transform 1 0 25300 0 -1 26656
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1606120353
transform 1 0 26404 0 -1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_44_276
timestamp 1606120353
transform 1 0 26496 0 -1 26656
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1606120353
transform -1 0 28888 0 -1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_44_288
timestamp 1606120353
transform 1 0 27600 0 -1 26656
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_44_296
timestamp 1606120353
transform 1 0 28336 0 -1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1606120353
transform 1 0 1104 0 1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__CLK
timestamp 1606120353
transform 1 0 1564 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1606120353
transform 1 0 1380 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_45_7
timestamp 1606120353
transform 1 0 1748 0 1 26656
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_45_19
timestamp 1606120353
transform 1 0 2852 0 1 26656
box 0 -48 736 592
use sky130_fd_sc_hd__o22a_4  _0809_
timestamp 1606120353
transform 1 0 4692 0 1 26656
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__A1
timestamp 1606120353
transform 1 0 4508 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__A2
timestamp 1606120353
transform 1 0 4140 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__B1
timestamp 1606120353
transform 1 0 3772 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_27
timestamp 1606120353
transform 1 0 3588 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_31
timestamp 1606120353
transform 1 0 3956 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_35
timestamp 1606120353
transform 1 0 4324 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1092_
timestamp 1606120353
transform 1 0 6900 0 1 26656
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1606120353
transform 1 0 6716 0 1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__A1
timestamp 1606120353
transform 1 0 6532 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__D
timestamp 1606120353
transform 1 0 6164 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_53
timestamp 1606120353
transform 1 0 5980 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_57
timestamp 1606120353
transform 1 0 6348 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_45_62
timestamp 1606120353
transform 1 0 6808 0 1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__B2
timestamp 1606120353
transform 1 0 9200 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__A1_N
timestamp 1606120353
transform 1 0 8832 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_82
timestamp 1606120353
transform 1 0 8648 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_86
timestamp 1606120353
transform 1 0 9016 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__a2bb2o_4  _0781_
timestamp 1606120353
transform 1 0 9384 0 1 26656
box 0 -48 1472 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__B
timestamp 1606120353
transform 1 0 11040 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_106
timestamp 1606120353
transform 1 0 10856 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1606120353
transform 1 0 11224 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0686_
timestamp 1606120353
transform 1 0 12420 0 1 26656
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1606120353
transform 1 0 12328 0 1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__A
timestamp 1606120353
transform 1 0 12144 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__B1
timestamp 1606120353
transform 1 0 11776 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__A2
timestamp 1606120353
transform 1 0 11408 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_114
timestamp 1606120353
transform 1 0 11592 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_118
timestamp 1606120353
transform 1 0 11960 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_45_132
timestamp 1606120353
transform 1 0 13248 0 1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__nor4_4  _0618_
timestamp 1606120353
transform 1 0 14076 0 1 26656
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0520__A
timestamp 1606120353
transform 1 0 13892 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__B
timestamp 1606120353
transform 1 0 13524 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_137
timestamp 1606120353
transform 1 0 13708 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0628_
timestamp 1606120353
transform 1 0 16376 0 1 26656
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0628__B
timestamp 1606120353
transform 1 0 17204 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0562__A
timestamp 1606120353
transform 1 0 15824 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0628__A
timestamp 1606120353
transform 1 0 16192 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_158
timestamp 1606120353
transform 1 0 15640 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_162
timestamp 1606120353
transform 1 0 16008 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_173
timestamp 1606120353
transform 1 0 17020 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1135_
timestamp 1606120353
transform 1 0 18032 0 1 26656
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1606120353
transform 1 0 17940 0 1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__D
timestamp 1606120353
transform 1 0 17756 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_45_177
timestamp 1606120353
transform 1 0 17388 0 1 26656
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__D
timestamp 1606120353
transform 1 0 19964 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_45_203
timestamp 1606120353
transform 1 0 19780 0 1 26656
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_45_207
timestamp 1606120353
transform 1 0 20148 0 1 26656
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_45_219
timestamp 1606120353
transform 1 0 21252 0 1 26656
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_45_231
timestamp 1606120353
transform 1 0 22356 0 1 26656
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1606120353
transform 1 0 23552 0 1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_45_243
timestamp 1606120353
transform 1 0 23460 0 1 26656
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_45_245
timestamp 1606120353
transform 1 0 23644 0 1 26656
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_45_257
timestamp 1606120353
transform 1 0 24748 0 1 26656
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_45_269
timestamp 1606120353
transform 1 0 25852 0 1 26656
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1606120353
transform 1 0 26956 0 1 26656
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1606120353
transform -1 0 28888 0 1 26656
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_45_293
timestamp 1606120353
transform 1 0 28060 0 1 26656
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_47_3
timestamp 1606120353
transform 1 0 1380 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_11
timestamp 1606120353
transform 1 0 2116 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_7
timestamp 1606120353
transform 1 0 1748 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1606120353
transform 1 0 1380 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__D
timestamp 1606120353
transform 1 0 1932 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__D
timestamp 1606120353
transform 1 0 1564 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1606120353
transform 1 0 1104 0 1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1606120353
transform 1 0 1104 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__CLK
timestamp 1606120353
transform 1 0 2300 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1606120353
transform 1 0 2484 0 -1 27744
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1124_
timestamp 1606120353
transform 1 0 1564 0 1 27744
box 0 -48 1748 592
use sky130_fd_sc_hd__dfxtp_4  _1104_
timestamp 1606120353
transform 1 0 4784 0 -1 27744
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1606120353
transform 1 0 3956 0 -1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__CLK
timestamp 1606120353
transform 1 0 4600 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_46_27
timestamp 1606120353
transform 1 0 3588 0 -1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__decap_6  FILLER_46_32
timestamp 1606120353
transform 1 0 4048 0 -1 27744
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_47_24
timestamp 1606120353
transform 1 0 3312 0 1 27744
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_47_36
timestamp 1606120353
transform 1 0 4416 0 1 27744
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_clk_A
timestamp 1606120353
transform 1 0 5520 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_47_50
timestamp 1606120353
transform 1 0 5704 0 1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_47_54
timestamp 1606120353
transform 1 0 6072 0 1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__A1
timestamp 1606120353
transform 1 0 6164 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_57
timestamp 1606120353
transform 1 0 6348 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_59
timestamp 1606120353
transform 1 0 6532 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0654__A
timestamp 1606120353
transform 1 0 6532 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_62
timestamp 1606120353
transform 1 0 6808 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_63
timestamp 1606120353
transform 1 0 6900 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__B2
timestamp 1606120353
transform 1 0 6716 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1606120353
transform 1 0 6716 0 1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0654_
timestamp 1606120353
transform 1 0 6992 0 1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__B1
timestamp 1606120353
transform 1 0 7084 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_47_74
timestamp 1606120353
transform 1 0 7912 0 1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_47_71
timestamp 1606120353
transform 1 0 7636 0 1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_47_67
timestamp 1606120353
transform 1 0 7268 0 1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__A2
timestamp 1606120353
transform 1 0 7728 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0709_
timestamp 1606120353
transform 1 0 8004 0 1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_47_82
timestamp 1606120353
transform 1 0 8648 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_78
timestamp 1606120353
transform 1 0 8280 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_88
timestamp 1606120353
transform 1 0 9200 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_46_85
timestamp 1606120353
transform 1 0 8924 0 -1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_46_81
timestamp 1606120353
transform 1 0 8556 0 -1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__A2
timestamp 1606120353
transform 1 0 9016 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__A1
timestamp 1606120353
transform 1 0 8832 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__A
timestamp 1606120353
transform 1 0 8464 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _0782_
timestamp 1606120353
transform 1 0 7268 0 -1 27744
box 0 -48 1288 592
use sky130_fd_sc_hd__o22a_4  _0775_
timestamp 1606120353
transform 1 0 9016 0 1 27744
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_46_93
timestamp 1606120353
transform 1 0 9660 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__A1
timestamp 1606120353
transform 1 0 9844 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__B1
timestamp 1606120353
transform 1 0 9384 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1606120353
transform 1 0 9568 0 -1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_47_107
timestamp 1606120353
transform 1 0 10948 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_47_104
timestamp 1606120353
transform 1 0 10672 0 1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_47_100
timestamp 1606120353
transform 1 0 10304 0 1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_46_110
timestamp 1606120353
transform 1 0 11224 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__C
timestamp 1606120353
transform 1 0 10764 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__D
timestamp 1606120353
transform 1 0 11132 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _0710_
timestamp 1606120353
transform 1 0 10028 0 -1 27744
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_47_118
timestamp 1606120353
transform 1 0 11960 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_114
timestamp 1606120353
transform 1 0 11592 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_114
timestamp 1606120353
transform 1 0 11592 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__A1
timestamp 1606120353
transform 1 0 11408 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__C
timestamp 1606120353
transform 1 0 11776 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0541__A
timestamp 1606120353
transform 1 0 11776 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__A
timestamp 1606120353
transform 1 0 12144 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0541_
timestamp 1606120353
transform 1 0 11316 0 1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_47_132
timestamp 1606120353
transform 1 0 13248 0 1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_46_131
timestamp 1606120353
transform 1 0 13156 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1606120353
transform 1 0 12328 0 1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__and3_4  _0689_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 12420 0 1 27744
box 0 -48 828 592
use sky130_fd_sc_hd__a21oi_4  _0706_
timestamp 1606120353
transform 1 0 11960 0 -1 27744
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_47_138
timestamp 1606120353
transform 1 0 13800 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_142
timestamp 1606120353
transform 1 0 14168 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_135
timestamp 1606120353
transform 1 0 13524 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__B
timestamp 1606120353
transform 1 0 13708 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__A
timestamp 1606120353
transform 1 0 13340 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0534__A
timestamp 1606120353
transform 1 0 13616 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__C
timestamp 1606120353
transform 1 0 13984 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0520_
timestamp 1606120353
transform 1 0 13892 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_46_154
timestamp 1606120353
transform 1 0 15272 0 -1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_46_150
timestamp 1606120353
transform 1 0 14904 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_46_146
timestamp 1606120353
transform 1 0 14536 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__D
timestamp 1606120353
transform 1 0 14720 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__A
timestamp 1606120353
transform 1 0 14352 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1606120353
transform 1 0 15180 0 -1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__nand4_4  _0567_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 14168 0 1 27744
box 0 -48 1564 592
use sky130_fd_sc_hd__fill_2  FILLER_47_163
timestamp 1606120353
transform 1 0 16100 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_159
timestamp 1606120353
transform 1 0 15732 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_162
timestamp 1606120353
transform 1 0 16008 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_158
timestamp 1606120353
transform 1 0 15640 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__B
timestamp 1606120353
transform 1 0 16192 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__B
timestamp 1606120353
transform 1 0 15824 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__C
timestamp 1606120353
transform 1 0 16284 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__A
timestamp 1606120353
transform 1 0 15916 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0562_
timestamp 1606120353
transform 1 0 15364 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_47_174
timestamp 1606120353
transform 1 0 17112 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0595__B
timestamp 1606120353
transform 1 0 17296 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0595_
timestamp 1606120353
transform 1 0 16468 0 1 27744
box 0 -48 644 592
use sky130_fd_sc_hd__dfxtp_4  _1090_
timestamp 1606120353
transform 1 0 16376 0 -1 27744
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_1  FILLER_47_182
timestamp 1606120353
transform 1 0 17848 0 1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_47_178
timestamp 1606120353
transform 1 0 17480 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_46_185
timestamp 1606120353
transform 1 0 18124 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__A
timestamp 1606120353
transform 1 0 17664 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1606120353
transform 1 0 17940 0 1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_47_196
timestamp 1606120353
transform 1 0 19136 0 1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_46_196
timestamp 1606120353
transform 1 0 19136 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_46_190
timestamp 1606120353
transform 1 0 18584 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__A1
timestamp 1606120353
transform 1 0 19320 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0518__A
timestamp 1606120353
transform 1 0 18400 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0629_
timestamp 1606120353
transform 1 0 18860 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__a21o_4  _0777_
timestamp 1606120353
transform 1 0 18032 0 1 27744
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_47_201
timestamp 1606120353
transform 1 0 19596 0 1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_46_204
timestamp 1606120353
transform 1 0 19872 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_200
timestamp 1606120353
transform 1 0 19504 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__B1
timestamp 1606120353
transform 1 0 19688 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0600__A
timestamp 1606120353
transform 1 0 19412 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0624_
timestamp 1606120353
transform 1 0 19872 0 1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_47_207
timestamp 1606120353
transform 1 0 20148 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_46_208
timestamp 1606120353
transform 1 0 20240 0 -1 27744
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__A2
timestamp 1606120353
transform 1 0 20056 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0624__A
timestamp 1606120353
transform 1 0 20332 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_47_211
timestamp 1606120353
transform 1 0 20516 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_46_215
timestamp 1606120353
transform 1 0 20884 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__D
timestamp 1606120353
transform 1 0 20700 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_clk
timestamp 1606120353
transform 1 0 20884 0 1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1606120353
transform 1 0 20792 0 -1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_47_218
timestamp 1606120353
transform 1 0 21160 0 1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_46_219
timestamp 1606120353
transform 1 0 21252 0 -1 27744
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_clk_A
timestamp 1606120353
transform 1 0 21068 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0929_
timestamp 1606120353
transform 1 0 21620 0 1 27744
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__B1_N
timestamp 1606120353
transform 1 0 21436 0 1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__A2
timestamp 1606120353
transform 1 0 21620 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_46_225
timestamp 1606120353
transform 1 0 21804 0 -1 27744
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_46_237
timestamp 1606120353
transform 1 0 22908 0 -1 27744
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_47_236
timestamp 1606120353
transform 1 0 22816 0 1 27744
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1606120353
transform 1 0 23552 0 1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_46_249
timestamp 1606120353
transform 1 0 24012 0 -1 27744
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_46_261
timestamp 1606120353
transform 1 0 25116 0 -1 27744
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_47_245
timestamp 1606120353
transform 1 0 23644 0 1 27744
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_47_257
timestamp 1606120353
transform 1 0 24748 0 1 27744
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1606120353
transform 1 0 26404 0 -1 27744
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_46_273
timestamp 1606120353
transform 1 0 26220 0 -1 27744
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_46_276
timestamp 1606120353
transform 1 0 26496 0 -1 27744
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_47_269
timestamp 1606120353
transform 1 0 25852 0 1 27744
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1606120353
transform 1 0 26956 0 1 27744
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1606120353
transform -1 0 28888 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1606120353
transform -1 0 28888 0 1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_46_288
timestamp 1606120353
transform 1 0 27600 0 -1 27744
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_46_296
timestamp 1606120353
transform 1 0 28336 0 -1 27744
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_47_293
timestamp 1606120353
transform 1 0 28060 0 1 27744
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1216_
timestamp 1606120353
transform 1 0 1380 0 -1 28832
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1606120353
transform 1 0 1104 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_48_22
timestamp 1606120353
transform 1 0 3128 0 -1 28832
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1606120353
transform 1 0 3956 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_48_30
timestamp 1606120353
transform 1 0 3864 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_48_32
timestamp 1606120353
transform 1 0 4048 0 -1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_48_44
timestamp 1606120353
transform 1 0 5152 0 -1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_clk
timestamp 1606120353
transform 1 0 5520 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__A2
timestamp 1606120353
transform 1 0 7176 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__B2
timestamp 1606120353
transform 1 0 6808 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__A1
timestamp 1606120353
transform 1 0 6440 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__A2
timestamp 1606120353
transform 1 0 6072 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_48_51
timestamp 1606120353
transform 1 0 5796 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_48_56
timestamp 1606120353
transform 1 0 6256 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_60
timestamp 1606120353
transform 1 0 6624 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_64
timestamp 1606120353
transform 1 0 6992 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0774_
timestamp 1606120353
transform 1 0 7728 0 -1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__D
timestamp 1606120353
transform 1 0 9016 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__B1
timestamp 1606120353
transform 1 0 7544 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_68
timestamp 1606120353
transform 1 0 7360 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_84
timestamp 1606120353
transform 1 0 8832 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_88
timestamp 1606120353
transform 1 0 9200 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__a21oi_4  _0708_
timestamp 1606120353
transform 1 0 10580 0 -1 28832
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1606120353
transform 1 0 9568 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__A1
timestamp 1606120353
transform 1 0 9844 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__D
timestamp 1606120353
transform 1 0 10304 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__C1
timestamp 1606120353
transform 1 0 9384 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_93
timestamp 1606120353
transform 1 0 9660 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_48_97
timestamp 1606120353
transform 1 0 10028 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_48_102
timestamp 1606120353
transform 1 0 10488 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _0690_
timestamp 1606120353
transform 1 0 12512 0 -1 28832
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__B
timestamp 1606120353
transform 1 0 12328 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__B
timestamp 1606120353
transform 1 0 11960 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_116
timestamp 1606120353
transform 1 0 11776 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_120
timestamp 1606120353
transform 1 0 12144 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_137
timestamp 1606120353
transform 1 0 13708 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_133
timestamp 1606120353
transform 1 0 13340 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__C
timestamp 1606120353
transform 1 0 13892 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__B
timestamp 1606120353
transform 1 0 13524 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0534_
timestamp 1606120353
transform 1 0 14076 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_48_148
timestamp 1606120353
transform 1 0 14720 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_144
timestamp 1606120353
transform 1 0 14352 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__C
timestamp 1606120353
transform 1 0 14904 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__B
timestamp 1606120353
transform 1 0 14536 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_48_152
timestamp 1606120353
transform 1 0 15088 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1606120353
transform 1 0 15180 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _0641_
timestamp 1606120353
transform 1 0 15272 0 -1 28832
box 0 -48 828 592
use sky130_fd_sc_hd__or4_4  _0704_
timestamp 1606120353
transform 1 0 16836 0 -1 28832
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__A
timestamp 1606120353
transform 1 0 16284 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0619__C
timestamp 1606120353
transform 1 0 16652 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_163
timestamp 1606120353
transform 1 0 16100 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_167
timestamp 1606120353
transform 1 0 16468 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0518_
timestamp 1606120353
transform 1 0 18400 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0594__B
timestamp 1606120353
transform 1 0 18032 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__C
timestamp 1606120353
transform 1 0 18860 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__D
timestamp 1606120353
transform 1 0 19228 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_48_180
timestamp 1606120353
transform 1 0 17664 0 -1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_48_186
timestamp 1606120353
transform 1 0 18216 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_191
timestamp 1606120353
transform 1 0 18676 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_195
timestamp 1606120353
transform 1 0 19044 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0600_
timestamp 1606120353
transform 1 0 19412 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1606120353
transform 1 0 20792 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0595__A
timestamp 1606120353
transform 1 0 19872 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_clk_A
timestamp 1606120353
transform 1 0 20240 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_202
timestamp 1606120353
transform 1 0 19688 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_48_206
timestamp 1606120353
transform 1 0 20056 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_48_210
timestamp 1606120353
transform 1 0 20424 0 -1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILLER_48_215
timestamp 1606120353
transform 1 0 20884 0 -1 28832
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__A1
timestamp 1606120353
transform 1 0 21620 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_48_225
timestamp 1606120353
transform 1 0 21804 0 -1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_48_237
timestamp 1606120353
transform 1 0 22908 0 -1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_48_249
timestamp 1606120353
transform 1 0 24012 0 -1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_48_261
timestamp 1606120353
transform 1 0 25116 0 -1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1606120353
transform 1 0 26404 0 -1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_48_273
timestamp 1606120353
transform 1 0 26220 0 -1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_48_276
timestamp 1606120353
transform 1 0 26496 0 -1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1606120353
transform -1 0 28888 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_48_288
timestamp 1606120353
transform 1 0 27600 0 -1 28832
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_48_296
timestamp 1606120353
transform 1 0 28336 0 -1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1606120353
transform 1 0 1104 0 1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1606120353
transform 1 0 1380 0 1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1606120353
transform 1 0 2484 0 1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1606120353
transform 1 0 3588 0 1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_49_39
timestamp 1606120353
transform 1 0 4692 0 1 28832
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__A
timestamp 1606120353
transform 1 0 5428 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_49
timestamp 1606120353
transform 1 0 5612 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__D
timestamp 1606120353
transform 1 0 5796 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_53
timestamp 1606120353
transform 1 0 5980 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__A
timestamp 1606120353
transform 1 0 6164 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_57
timestamp 1606120353
transform 1 0 6348 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__D
timestamp 1606120353
transform 1 0 6532 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_62
timestamp 1606120353
transform 1 0 6808 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0640__A
timestamp 1606120353
transform 1 0 6992 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1606120353
transform 1 0 6716 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_49_66
timestamp 1606120353
transform 1 0 7176 0 1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__and2_4  _0771_
timestamp 1606120353
transform 1 0 8188 0 1 28832
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__B
timestamp 1606120353
transform 1 0 9016 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__B1
timestamp 1606120353
transform 1 0 8004 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__A1
timestamp 1606120353
transform 1 0 7636 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_49_70
timestamp 1606120353
transform 1 0 7544 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_49_73
timestamp 1606120353
transform 1 0 7820 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_84
timestamp 1606120353
transform 1 0 8832 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_88
timestamp 1606120353
transform 1 0 9200 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__a211o_4  _0672_
timestamp 1606120353
transform 1 0 9568 0 1 28832
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__B1
timestamp 1606120353
transform 1 0 9384 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_49_106
timestamp 1606120353
transform 1 0 10856 0 1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_49_110
timestamp 1606120353
transform 1 0 11224 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_49_117
timestamp 1606120353
transform 1 0 11868 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_113
timestamp 1606120353
transform 1 0 11500 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__B
timestamp 1606120353
transform 1 0 11316 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__B
timestamp 1606120353
transform 1 0 11684 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__A
timestamp 1606120353
transform 1 0 12052 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_127
timestamp 1606120353
transform 1 0 12788 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_123
timestamp 1606120353
transform 1 0 12420 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_49_121
timestamp 1606120353
transform 1 0 12236 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__C
timestamp 1606120353
transform 1 0 12604 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1606120353
transform 1 0 12328 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__C
timestamp 1606120353
transform 1 0 12972 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0698_
timestamp 1606120353
transform 1 0 13156 0 1 28832
box 0 -48 828 592
use sky130_fd_sc_hd__and4_4  _0696_
timestamp 1606120353
transform 1 0 14720 0 1 28832
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__A
timestamp 1606120353
transform 1 0 14536 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__B
timestamp 1606120353
transform 1 0 14168 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_140
timestamp 1606120353
transform 1 0 13984 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_144
timestamp 1606120353
transform 1 0 14352 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0703_
timestamp 1606120353
transform 1 0 16284 0 1 28832
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__C
timestamp 1606120353
transform 1 0 15732 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0619__A
timestamp 1606120353
transform 1 0 17296 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0619__B
timestamp 1606120353
transform 1 0 16100 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_157
timestamp 1606120353
transform 1 0 15548 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_161
timestamp 1606120353
transform 1 0 15916 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_174
timestamp 1606120353
transform 1 0 17112 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0594_
timestamp 1606120353
transform 1 0 18032 0 1 28832
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1606120353
transform 1 0 17940 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__A
timestamp 1606120353
transform 1 0 18860 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__B
timestamp 1606120353
transform 1 0 19228 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__C
timestamp 1606120353
transform 1 0 17756 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_49_178
timestamp 1606120353
transform 1 0 17480 0 1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_49_191
timestamp 1606120353
transform 1 0 18676 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_195
timestamp 1606120353
transform 1 0 19044 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_202
timestamp 1606120353
transform 1 0 19688 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0695_
timestamp 1606120353
transform 1 0 19412 0 1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_49_206
timestamp 1606120353
transform 1 0 20056 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__D
timestamp 1606120353
transform 1 0 19872 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_210
timestamp 1606120353
transform 1 0 20424 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0594__A
timestamp 1606120353
transform 1 0 20240 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_49_214
timestamp 1606120353
transform 1 0 20792 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__A
timestamp 1606120353
transform 1 0 20608 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_49_218
timestamp 1606120353
transform 1 0 21160 0 1 28832
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__D
timestamp 1606120353
transform 1 0 20976 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_clk_A
timestamp 1606120353
transform 1 0 21620 0 1 28832
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_49_222
timestamp 1606120353
transform 1 0 21528 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1606120353
transform 1 0 21804 0 1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_49_237
timestamp 1606120353
transform 1 0 22908 0 1 28832
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1606120353
transform 1 0 23552 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_49_243
timestamp 1606120353
transform 1 0 23460 0 1 28832
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_49_245
timestamp 1606120353
transform 1 0 23644 0 1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_49_257
timestamp 1606120353
transform 1 0 24748 0 1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_49_269
timestamp 1606120353
transform 1 0 25852 0 1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1606120353
transform 1 0 26956 0 1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1606120353
transform -1 0 28888 0 1 28832
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_49_293
timestamp 1606120353
transform 1 0 28060 0 1 28832
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1606120353
transform 1 0 1104 0 -1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1606120353
transform 1 0 1380 0 -1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1606120353
transform 1 0 2484 0 -1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1606120353
transform 1 0 3956 0 -1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_50_27
timestamp 1606120353
transform 1 0 3588 0 -1 29920
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_50_32
timestamp 1606120353
transform 1 0 4048 0 -1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_50_44
timestamp 1606120353
transform 1 0 5152 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__CLK
timestamp 1606120353
transform 1 0 5336 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_48
timestamp 1606120353
transform 1 0 5520 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__D
timestamp 1606120353
transform 1 0 5704 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_52
timestamp 1606120353
transform 1 0 5888 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_56
timestamp 1606120353
transform 1 0 6256 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__D
timestamp 1606120353
transform 1 0 6072 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__D
timestamp 1606120353
transform 1 0 6440 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_60
timestamp 1606120353
transform 1 0 6624 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__A1
timestamp 1606120353
transform 1 0 6808 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0640_
timestamp 1606120353
transform 1 0 6992 0 -1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__inv_8  _0673_
timestamp 1606120353
transform 1 0 8004 0 -1 29920
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__A1
timestamp 1606120353
transform 1 0 9016 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__A2
timestamp 1606120353
transform 1 0 7820 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__A2
timestamp 1606120353
transform 1 0 7452 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_67
timestamp 1606120353
transform 1 0 7268 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_71
timestamp 1606120353
transform 1 0 7636 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_84
timestamp 1606120353
transform 1 0 8832 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_88
timestamp 1606120353
transform 1 0 9200 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0773_
timestamp 1606120353
transform 1 0 9660 0 -1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1606120353
transform 1 0 9568 0 -1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__C
timestamp 1606120353
transform 1 0 10948 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__A2
timestamp 1606120353
transform 1 0 9384 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_105
timestamp 1606120353
transform 1 0 10764 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_50_109
timestamp 1606120353
transform 1 0 11132 0 -1 29920
box 0 -48 368 592
use sky130_fd_sc_hd__and4_4  _0694_
timestamp 1606120353
transform 1 0 12052 0 -1 29920
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__A
timestamp 1606120353
transform 1 0 13064 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__B
timestamp 1606120353
transform 1 0 11868 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__B
timestamp 1606120353
transform 1 0 11500 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_115
timestamp 1606120353
transform 1 0 11684 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_128
timestamp 1606120353
transform 1 0 12880 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_132
timestamp 1606120353
transform 1 0 13248 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0699_
timestamp 1606120353
transform 1 0 13616 0 -1 29920
box 0 -48 828 592
use sky130_fd_sc_hd__or4_4  _0705_
timestamp 1606120353
transform 1 0 15272 0 -1 29920
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1606120353
transform 1 0 15180 0 -1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__C1
timestamp 1606120353
transform 1 0 14628 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__B1
timestamp 1606120353
transform 1 0 14996 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__A
timestamp 1606120353
transform 1 0 13432 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_145
timestamp 1606120353
transform 1 0 14444 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_149
timestamp 1606120353
transform 1 0 14812 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__and3_4  _0619_
timestamp 1606120353
transform 1 0 16836 0 -1 29920
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__A
timestamp 1606120353
transform 1 0 16284 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__B
timestamp 1606120353
transform 1 0 16652 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_163
timestamp 1606120353
transform 1 0 16100 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_167
timestamp 1606120353
transform 1 0 16468 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0583_
timestamp 1606120353
transform 1 0 18400 0 -1 29920
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__A
timestamp 1606120353
transform 1 0 17848 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__B
timestamp 1606120353
transform 1 0 18216 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_180
timestamp 1606120353
transform 1 0 17664 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_184
timestamp 1606120353
transform 1 0 18032 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_197
timestamp 1606120353
transform 1 0 19228 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_201
timestamp 1606120353
transform 1 0 19596 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__B1
timestamp 1606120353
transform 1 0 19412 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__D
timestamp 1606120353
transform 1 0 19780 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_clk
timestamp 1606120353
transform 1 0 19964 0 -1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_50_208
timestamp 1606120353
transform 1 0 20240 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0487__A
timestamp 1606120353
transform 1 0 20424 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_50_212
timestamp 1606120353
transform 1 0 20608 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1606120353
transform 1 0 20792 0 -1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_50_215
timestamp 1606120353
transform 1 0 20884 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1102__CLK
timestamp 1606120353
transform 1 0 21068 0 -1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_50_219
timestamp 1606120353
transform 1 0 21252 0 -1 29920
box 0 -48 368 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_clk
timestamp 1606120353
transform 1 0 21620 0 -1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_50_226
timestamp 1606120353
transform 1 0 21896 0 -1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_50_238
timestamp 1606120353
transform 1 0 23000 0 -1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_50_250
timestamp 1606120353
transform 1 0 24104 0 -1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_50_262
timestamp 1606120353
transform 1 0 25208 0 -1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1606120353
transform 1 0 26404 0 -1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_50_274
timestamp 1606120353
transform 1 0 26312 0 -1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_50_276
timestamp 1606120353
transform 1 0 26496 0 -1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1606120353
transform -1 0 28888 0 -1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_50_288
timestamp 1606120353
transform 1 0 27600 0 -1 29920
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_50_296
timestamp 1606120353
transform 1 0 28336 0 -1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1606120353
transform 1 0 1104 0 1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1606120353
transform 1 0 1380 0 1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1606120353
transform 1 0 2484 0 1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_clk
timestamp 1606120353
transform 1 0 4232 0 1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_clk_A
timestamp 1606120353
transform 1 0 5152 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_clk_A
timestamp 1606120353
transform 1 0 4692 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_51_27
timestamp 1606120353
transform 1 0 3588 0 1 29920
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_51_33
timestamp 1606120353
transform 1 0 4140 0 1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_51_37
timestamp 1606120353
transform 1 0 4508 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_51_41
timestamp 1606120353
transform 1 0 4876 0 1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__o22a_4  _0820_
timestamp 1606120353
transform 1 0 6808 0 1 29920
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1606120353
transform 1 0 6716 0 1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_clk
timestamp 1606120353
transform 1 0 6440 0 1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__B2
timestamp 1606120353
transform 1 0 6256 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__A2
timestamp 1606120353
transform 1 0 5888 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__B1
timestamp 1606120353
transform 1 0 5520 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_46
timestamp 1606120353
transform 1 0 5336 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_50
timestamp 1606120353
transform 1 0 5704 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_54
timestamp 1606120353
transform 1 0 6072 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0685_
timestamp 1606120353
transform 1 0 9200 0 1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0536__A
timestamp 1606120353
transform 1 0 8556 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__B1
timestamp 1606120353
transform 1 0 9016 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_51_76
timestamp 1606120353
transform 1 0 8096 0 1 29920
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_51_80
timestamp 1606120353
transform 1 0 8464 0 1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_51_83
timestamp 1606120353
transform 1 0 8740 0 1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__B
timestamp 1606120353
transform 1 0 10488 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__A
timestamp 1606120353
transform 1 0 10856 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_100
timestamp 1606120353
transform 1 0 10304 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_104
timestamp 1606120353
transform 1 0 10672 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_51_108
timestamp 1606120353
transform 1 0 11040 0 1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0491_
timestamp 1606120353
transform 1 0 11316 0 1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__and4_4  _0697_
timestamp 1606120353
transform 1 0 12880 0 1 29920
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1606120353
transform 1 0 12328 0 1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0491__A
timestamp 1606120353
transform 1 0 11776 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__C
timestamp 1606120353
transform 1 0 12696 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__C
timestamp 1606120353
transform 1 0 12144 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_114
timestamp 1606120353
transform 1 0 11592 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_118
timestamp 1606120353
transform 1 0 11960 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_51_123
timestamp 1606120353
transform 1 0 12420 0 1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__a2111oi_4  _0596_
timestamp 1606120353
transform 1 0 14444 0 1 29920
box 0 -48 2024 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0563__A
timestamp 1606120353
transform 1 0 14168 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_51_137
timestamp 1606120353
transform 1 0 13708 0 1 29920
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_51_141
timestamp 1606120353
transform 1 0 14076 0 1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_51_144
timestamp 1606120353
transform 1 0 14352 0 1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__A
timestamp 1606120353
transform 1 0 16652 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__B
timestamp 1606120353
transform 1 0 17020 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_167
timestamp 1606120353
transform 1 0 16468 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_171
timestamp 1606120353
transform 1 0 16836 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_175
timestamp 1606120353
transform 1 0 17204 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _0805_
timestamp 1606120353
transform 1 0 18032 0 1 29920
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1606120353
transform 1 0 17940 0 1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__B1
timestamp 1606120353
transform 1 0 17756 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__D
timestamp 1606120353
transform 1 0 17388 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_179
timestamp 1606120353
transform 1 0 17572 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_198
timestamp 1606120353
transform 1 0 19320 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__A1
timestamp 1606120353
transform 1 0 19504 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_202
timestamp 1606120353
transform 1 0 19688 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__A2
timestamp 1606120353
transform 1 0 19872 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0487_
timestamp 1606120353
transform 1 0 20056 0 1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_51_209
timestamp 1606120353
transform 1 0 20332 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_213
timestamp 1606120353
transform 1 0 20700 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__D
timestamp 1606120353
transform 1 0 20516 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0530__A
timestamp 1606120353
transform 1 0 20884 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_217
timestamp 1606120353
transform 1 0 21068 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1102__D
timestamp 1606120353
transform 1 0 21252 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__A1
timestamp 1606120353
transform 1 0 21620 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_51_221
timestamp 1606120353
transform 1 0 21436 0 1 29920
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1606120353
transform 1 0 21804 0 1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_51_237
timestamp 1606120353
transform 1 0 22908 0 1 29920
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1606120353
transform 1 0 23552 0 1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_51_243
timestamp 1606120353
transform 1 0 23460 0 1 29920
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_51_245
timestamp 1606120353
transform 1 0 23644 0 1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_51_257
timestamp 1606120353
transform 1 0 24748 0 1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_51_269
timestamp 1606120353
transform 1 0 25852 0 1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1606120353
transform 1 0 26956 0 1 29920
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1606120353
transform -1 0 28888 0 1 29920
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_51_293
timestamp 1606120353
transform 1 0 28060 0 1 29920
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1606120353
transform 1 0 1104 0 -1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1606120353
transform 1 0 1104 0 1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__D
timestamp 1606120353
transform 1 0 1564 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__CLK
timestamp 1606120353
transform 1 0 1932 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1606120353
transform 1 0 1380 0 -1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1606120353
transform 1 0 2484 0 -1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1606120353
transform 1 0 1380 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_53_7
timestamp 1606120353
transform 1 0 1748 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_53_11
timestamp 1606120353
transform 1 0 2116 0 1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1606120353
transform 1 0 3956 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__D
timestamp 1606120353
transform 1 0 5060 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__CLK
timestamp 1606120353
transform 1 0 4692 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_52_27
timestamp 1606120353
transform 1 0 3588 0 -1 31008
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_52_32
timestamp 1606120353
transform 1 0 4048 0 -1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_52_44
timestamp 1606120353
transform 1 0 5152 0 -1 31008
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_53_23
timestamp 1606120353
transform 1 0 3220 0 1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_53_35
timestamp 1606120353
transform 1 0 4324 0 1 31008
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_53_41
timestamp 1606120353
transform 1 0 4876 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_53_53
timestamp 1606120353
transform 1 0 5980 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_53_49
timestamp 1606120353
transform 1 0 5612 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_53_45
timestamp 1606120353
transform 1 0 5244 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_50
timestamp 1606120353
transform 1 0 5704 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_clk_A
timestamp 1606120353
transform 1 0 5520 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__D
timestamp 1606120353
transform 1 0 5888 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__A1
timestamp 1606120353
transform 1 0 5428 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0655__A
timestamp 1606120353
transform 1 0 6164 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__D
timestamp 1606120353
transform 1 0 5796 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_53_62
timestamp 1606120353
transform 1 0 6808 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_53_57
timestamp 1606120353
transform 1 0 6348 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__B
timestamp 1606120353
transform 1 0 6532 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1606120353
transform 1 0 6716 0 1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0535_
timestamp 1606120353
transform 1 0 6992 0 1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1113_
timestamp 1606120353
transform 1 0 6072 0 -1 31008
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_2  FILLER_53_71
timestamp 1606120353
transform 1 0 7636 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_53_67
timestamp 1606120353
transform 1 0 7268 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_73
timestamp 1606120353
transform 1 0 7820 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0535__A
timestamp 1606120353
transform 1 0 7452 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0512__A
timestamp 1606120353
transform 1 0 7820 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_77
timestamp 1606120353
transform 1 0 8188 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__A3
timestamp 1606120353
transform 1 0 8004 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__B
timestamp 1606120353
transform 1 0 8372 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0674_
timestamp 1606120353
transform 1 0 8004 0 1 31008
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILLER_53_86
timestamp 1606120353
transform 1 0 9016 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_53_82
timestamp 1606120353
transform 1 0 8648 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_84
timestamp 1606120353
transform 1 0 8832 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__B2
timestamp 1606120353
transform 1 0 9016 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__B
timestamp 1606120353
transform 1 0 8832 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0536_
timestamp 1606120353
transform 1 0 8556 0 -1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_52_88
timestamp 1606120353
transform 1 0 9200 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__B1
timestamp 1606120353
transform 1 0 9200 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__a32o_4  _0671_
timestamp 1606120353
transform 1 0 9384 0 1 31008
box 0 -48 1564 592
use sky130_fd_sc_hd__and4_4  _0676_
timestamp 1606120353
transform 1 0 10304 0 -1 31008
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1606120353
transform 1 0 9568 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__A1
timestamp 1606120353
transform 1 0 9384 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__C
timestamp 1606120353
transform 1 0 9844 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_93
timestamp 1606120353
transform 1 0 9660 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_52_97
timestamp 1606120353
transform 1 0 10028 0 -1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_52_109
timestamp 1606120353
transform 1 0 11132 0 -1 31008
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_53_107
timestamp 1606120353
transform 1 0 10948 0 1 31008
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_53_118
timestamp 1606120353
transform 1 0 11960 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_53_113
timestamp 1606120353
transform 1 0 11500 0 1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_52_116
timestamp 1606120353
transform 1 0 11776 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_52_113
timestamp 1606120353
transform 1 0 11500 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__A
timestamp 1606120353
transform 1 0 11592 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__A
timestamp 1606120353
transform 1 0 11960 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__B2
timestamp 1606120353
transform 1 0 11776 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__B1
timestamp 1606120353
transform 1 0 11316 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_53_123
timestamp 1606120353
transform 1 0 12420 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__B1
timestamp 1606120353
transform 1 0 12144 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0545__B
timestamp 1606120353
transform 1 0 12604 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_clk
timestamp 1606120353
transform 1 0 12144 0 -1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1606120353
transform 1 0 12328 0 1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _0702_
timestamp 1606120353
transform 1 0 12788 0 1 31008
box 0 -48 828 592
use sky130_fd_sc_hd__and4_4  _0700_
timestamp 1606120353
transform 1 0 12420 0 -1 31008
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_52_132
timestamp 1606120353
transform 1 0 13248 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_53_140
timestamp 1606120353
transform 1 0 13984 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_53_136
timestamp 1606120353
transform 1 0 13616 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_140
timestamp 1606120353
transform 1 0 13984 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_136
timestamp 1606120353
transform 1 0 13616 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__C
timestamp 1606120353
transform 1 0 13800 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0545__C
timestamp 1606120353
transform 1 0 13432 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0545__A
timestamp 1606120353
transform 1 0 13800 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_149
timestamp 1606120353
transform 1 0 14812 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_145
timestamp 1606120353
transform 1 0 14444 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__C
timestamp 1606120353
transform 1 0 14168 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__A2
timestamp 1606120353
transform 1 0 14628 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0701_
timestamp 1606120353
transform 1 0 14352 0 1 31008
box 0 -48 828 592
use sky130_fd_sc_hd__buf_1  _0563_
timestamp 1606120353
transform 1 0 14168 0 -1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_53_153
timestamp 1606120353
transform 1 0 15180 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__D1
timestamp 1606120353
transform 1 0 14996 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1606120353
transform 1 0 15180 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__or3_4  _0597_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 15272 0 -1 31008
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_53_157
timestamp 1606120353
transform 1 0 15548 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_163
timestamp 1606120353
transform 1 0 16100 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__B
timestamp 1606120353
transform 1 0 15732 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0538__A
timestamp 1606120353
transform 1 0 15364 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0489_
timestamp 1606120353
transform 1 0 15916 0 1 31008
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_53_170
timestamp 1606120353
transform 1 0 16744 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_171
timestamp 1606120353
transform 1 0 16836 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_167
timestamp 1606120353
transform 1 0 16468 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__B
timestamp 1606120353
transform 1 0 16652 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__D
timestamp 1606120353
transform 1 0 16284 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__A
timestamp 1606120353
transform 1 0 16928 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_53_174
timestamp 1606120353
transform 1 0 17112 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_52_175
timestamp 1606120353
transform 1 0 17204 0 -1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__C
timestamp 1606120353
transform 1 0 17020 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__C
timestamp 1606120353
transform 1 0 17296 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1099_
timestamp 1606120353
transform 1 0 18032 0 1 31008
box 0 -48 1748 592
use sky130_fd_sc_hd__dfxtp_4  _1102_
timestamp 1606120353
transform 1 0 17664 0 -1 31008
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1606120353
transform 1 0 17940 0 1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__D
timestamp 1606120353
transform 1 0 17664 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__B2
timestamp 1606120353
transform 1 0 17480 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_53_178
timestamp 1606120353
transform 1 0 17480 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_53_182
timestamp 1606120353
transform 1 0 17848 0 1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_53_203
timestamp 1606120353
transform 1 0 19780 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_203
timestamp 1606120353
transform 1 0 19780 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_199
timestamp 1606120353
transform 1 0 19412 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__B2
timestamp 1606120353
transform 1 0 19964 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__A1
timestamp 1606120353
transform 1 0 19596 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0524__A
timestamp 1606120353
transform 1 0 19964 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_53_207
timestamp 1606120353
transform 1 0 20148 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_52_211
timestamp 1606120353
transform 1 0 20516 0 -1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_52_207
timestamp 1606120353
transform 1 0 20148 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__D
timestamp 1606120353
transform 1 0 20332 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0527__A
timestamp 1606120353
transform 1 0 20332 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _0527_
timestamp 1606120353
transform 1 0 20516 0 1 31008
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILLER_53_218
timestamp 1606120353
transform 1 0 21160 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_218
timestamp 1606120353
transform 1 0 21160 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1606120353
transform 1 0 20792 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0530_
timestamp 1606120353
transform 1 0 20884 0 -1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0489__A
timestamp 1606120353
transform 1 0 21344 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0527__B
timestamp 1606120353
transform 1 0 21344 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_53_229
timestamp 1606120353
transform 1 0 22172 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1606120353
transform 1 0 21528 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_226
timestamp 1606120353
transform 1 0 21896 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_52_222
timestamp 1606120353
transform 1 0 21528 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__CLK
timestamp 1606120353
transform 1 0 22080 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__CLK
timestamp 1606120353
transform 1 0 21712 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0523__A
timestamp 1606120353
transform 1 0 22356 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0524__B
timestamp 1606120353
transform 1 0 21712 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0523_
timestamp 1606120353
transform 1 0 21896 0 1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_53_241
timestamp 1606120353
transform 1 0 23276 0 1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_53_237
timestamp 1606120353
transform 1 0 22908 0 1 31008
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_53_233
timestamp 1606120353
transform 1 0 22540 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_52_242
timestamp 1606120353
transform 1 0 23368 0 -1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__A
timestamp 1606120353
transform 1 0 22724 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__D
timestamp 1606120353
transform 1 0 23368 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_52_230
timestamp 1606120353
transform 1 0 22264 0 -1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1141_
timestamp 1606120353
transform 1 0 23644 0 1 31008
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1606120353
transform 1 0 23552 0 1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__CLK
timestamp 1606120353
transform 1 0 23644 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_52_247
timestamp 1606120353
transform 1 0 23828 0 -1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_52_259
timestamp 1606120353
transform 1 0 24932 0 -1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_53_264
timestamp 1606120353
transform 1 0 25392 0 1 31008
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1168_
timestamp 1606120353
transform 1 0 26128 0 1 31008
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1606120353
transform 1 0 26404 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1168__D
timestamp 1606120353
transform 1 0 25944 0 1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1168__CLK
timestamp 1606120353
transform 1 0 26128 0 -1 31008
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_52_271
timestamp 1606120353
transform 1 0 26036 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_52_274
timestamp 1606120353
transform 1 0 26312 0 -1 31008
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_52_276
timestamp 1606120353
transform 1 0 26496 0 -1 31008
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1606120353
transform -1 0 28888 0 -1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1606120353
transform -1 0 28888 0 1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_52_288
timestamp 1606120353
transform 1 0 27600 0 -1 31008
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_52_296
timestamp 1606120353
transform 1 0 28336 0 -1 31008
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_53_291
timestamp 1606120353
transform 1 0 27876 0 1 31008
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1205_
timestamp 1606120353
transform 1 0 1472 0 -1 32096
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1606120353
transform 1 0 1104 0 -1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_54_3
timestamp 1606120353
transform 1 0 1380 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1606120353
transform 1 0 3956 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__A3
timestamp 1606120353
transform 1 0 4876 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__A2
timestamp 1606120353
transform 1 0 4508 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_54_23
timestamp 1606120353
transform 1 0 3220 0 -1 32096
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_54_32
timestamp 1606120353
transform 1 0 4048 0 -1 32096
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_54_36
timestamp 1606120353
transform 1 0 4416 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_54_39
timestamp 1606120353
transform 1 0 4692 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_54_43
timestamp 1606120353
transform 1 0 5060 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1123_
timestamp 1606120353
transform 1 0 5796 0 -1 32096
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__C
timestamp 1606120353
transform 1 0 5612 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__D
timestamp 1606120353
transform 1 0 5244 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_54_47
timestamp 1606120353
transform 1 0 5428 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0512_
timestamp 1606120353
transform 1 0 8556 0 -1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0655__B
timestamp 1606120353
transform 1 0 8188 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__B1
timestamp 1606120353
transform 1 0 9016 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__A
timestamp 1606120353
transform 1 0 7820 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_54_70
timestamp 1606120353
transform 1 0 7544 0 -1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_54_75
timestamp 1606120353
transform 1 0 8004 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_54_79
timestamp 1606120353
transform 1 0 8372 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_54_84
timestamp 1606120353
transform 1 0 8832 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_54_88
timestamp 1606120353
transform 1 0 9200 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0677_
timestamp 1606120353
transform 1 0 9752 0 -1 32096
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1606120353
transform 1 0 9568 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__A2
timestamp 1606120353
transform 1 0 11132 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__A
timestamp 1606120353
transform 1 0 9384 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__C1
timestamp 1606120353
transform 1 0 10764 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_54_93
timestamp 1606120353
transform 1 0 9660 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_54_103
timestamp 1606120353
transform 1 0 10580 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_54_107
timestamp 1606120353
transform 1 0 10948 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__or3_4  _0545_
timestamp 1606120353
transform 1 0 13156 0 -1 32096
box 0 -48 828 592
use sky130_fd_sc_hd__a21o_4  _0707_
timestamp 1606120353
transform 1 0 11316 0 -1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__A1
timestamp 1606120353
transform 1 0 12696 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_54_123
timestamp 1606120353
transform 1 0 12420 0 -1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_54_128
timestamp 1606120353
transform 1 0 12880 0 -1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0538_
timestamp 1606120353
transform 1 0 15272 0 -1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1606120353
transform 1 0 15180 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__B
timestamp 1606120353
transform 1 0 14168 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0589__D
timestamp 1606120353
transform 1 0 14812 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_54_140
timestamp 1606120353
transform 1 0 13984 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_54_144
timestamp 1606120353
transform 1 0 14352 0 -1 32096
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_54_148
timestamp 1606120353
transform 1 0 14720 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_54_151
timestamp 1606120353
transform 1 0 14996 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1100_
timestamp 1606120353
transform 1 0 16284 0 -1 32096
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__A
timestamp 1606120353
transform 1 0 15732 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__B
timestamp 1606120353
transform 1 0 16100 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_54_157
timestamp 1606120353
transform 1 0 15548 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_54_161
timestamp 1606120353
transform 1 0 15916 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__o22a_4  _0802_
timestamp 1606120353
transform 1 0 18768 0 -1 32096
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__A1
timestamp 1606120353
transform 1 0 18216 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__B2
timestamp 1606120353
transform 1 0 18584 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_54_184
timestamp 1606120353
transform 1 0 18032 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_54_188
timestamp 1606120353
transform 1 0 18400 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0524_
timestamp 1606120353
transform 1 0 20884 0 -1 32096
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1606120353
transform 1 0 20792 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__A2
timestamp 1606120353
transform 1 0 20240 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__D
timestamp 1606120353
transform 1 0 20608 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_54_206
timestamp 1606120353
transform 1 0 20056 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_54_210
timestamp 1606120353
transform 1 0 20424 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0830_
timestamp 1606120353
transform 1 0 22356 0 -1 32096
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__A2
timestamp 1606120353
transform 1 0 21712 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__B1
timestamp 1606120353
transform 1 0 22080 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__CLK
timestamp 1606120353
transform 1 0 23368 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_54_222
timestamp 1606120353
transform 1 0 21528 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_54_226
timestamp 1606120353
transform 1 0 21896 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_54_230
timestamp 1606120353
transform 1 0 22264 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_54_240
timestamp 1606120353
transform 1 0 23184 0 -1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_54_244
timestamp 1606120353
transform 1 0 23552 0 -1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_54_256
timestamp 1606120353
transform 1 0 24656 0 -1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1606120353
transform 1 0 26404 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_54_268
timestamp 1606120353
transform 1 0 25760 0 -1 32096
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_54_274
timestamp 1606120353
transform 1 0 26312 0 -1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_54_276
timestamp 1606120353
transform 1 0 26496 0 -1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1606120353
transform -1 0 28888 0 -1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_54_288
timestamp 1606120353
transform 1 0 27600 0 -1 32096
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_54_296
timestamp 1606120353
transform 1 0 28336 0 -1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1606120353
transform 1 0 1104 0 1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1606120353
transform 1 0 1380 0 1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_55_15
timestamp 1606120353
transform 1 0 2484 0 1 32096
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_55_23
timestamp 1606120353
transform 1 0 3220 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__CLK
timestamp 1606120353
transform 1 0 3404 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_27
timestamp 1606120353
transform 1 0 3588 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_31
timestamp 1606120353
transform 1 0 3956 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0502__A
timestamp 1606120353
transform 1 0 3772 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0540__D
timestamp 1606120353
transform 1 0 4140 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_35
timestamp 1606120353
transform 1 0 4324 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__D
timestamp 1606120353
transform 1 0 4508 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0606_
timestamp 1606120353
transform 1 0 4692 0 1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_55_42
timestamp 1606120353
transform 1 0 4968 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__A
timestamp 1606120353
transform 1 0 5152 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_53
timestamp 1606120353
transform 1 0 5980 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_46
timestamp 1606120353
transform 1 0 5336 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0606__A
timestamp 1606120353
transform 1 0 5520 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0531_
timestamp 1606120353
transform 1 0 5704 0 1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_55_62
timestamp 1606120353
transform 1 0 6808 0 1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_55_57
timestamp 1606120353
transform 1 0 6348 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0531__A
timestamp 1606120353
transform 1 0 6532 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__D
timestamp 1606120353
transform 1 0 6164 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1606120353
transform 1 0 6716 0 1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _0502_
timestamp 1606120353
transform 1 0 6900 0 1 32096
box 0 -48 828 592
use sky130_fd_sc_hd__and4_4  _0675_
timestamp 1606120353
transform 1 0 8464 0 1 32096
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__C
timestamp 1606120353
transform 1 0 8280 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__A
timestamp 1606120353
transform 1 0 7912 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_72
timestamp 1606120353
transform 1 0 7728 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_76
timestamp 1606120353
transform 1 0 8096 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__nor4_4  _0684_
timestamp 1606120353
transform 1 0 10028 0 1 32096
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__A1
timestamp 1606120353
transform 1 0 9660 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_55_89
timestamp 1606120353
transform 1 0 9292 0 1 32096
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_55_95
timestamp 1606120353
transform 1 0 9844 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0683_
timestamp 1606120353
transform 1 0 12420 0 1 32096
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1606120353
transform 1 0 12328 0 1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__A
timestamp 1606120353
transform 1 0 12144 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__A2
timestamp 1606120353
transform 1 0 11776 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_114
timestamp 1606120353
transform 1 0 11592 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_118
timestamp 1606120353
transform 1 0 11960 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_132
timestamp 1606120353
transform 1 0 13248 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0679_
timestamp 1606120353
transform 1 0 13984 0 1 32096
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__A3
timestamp 1606120353
transform 1 0 13432 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__A
timestamp 1606120353
transform 1 0 13800 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__C
timestamp 1606120353
transform 1 0 15272 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_136
timestamp 1606120353
transform 1 0 13616 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_55_149
timestamp 1606120353
transform 1 0 14812 0 1 32096
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_55_153
timestamp 1606120353
transform 1 0 15180 0 1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__o22a_4  _0803_
timestamp 1606120353
transform 1 0 15916 0 1 32096
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__B1
timestamp 1606120353
transform 1 0 15732 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_55_156
timestamp 1606120353
transform 1 0 15456 0 1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_55_175
timestamp 1606120353
transform 1 0 17204 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_187
timestamp 1606120353
transform 1 0 18308 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_179
timestamp 1606120353
transform 1 0 17572 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__C
timestamp 1606120353
transform 1 0 17756 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__D
timestamp 1606120353
transform 1 0 17388 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1606120353
transform 1 0 17940 0 1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0582_
timestamp 1606120353
transform 1 0 18032 0 1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_55_191
timestamp 1606120353
transform 1 0 18676 0 1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0582__A
timestamp 1606120353
transform 1 0 18492 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__D
timestamp 1606120353
transform 1 0 18952 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1134_
timestamp 1606120353
transform 1 0 19136 0 1 32096
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__D
timestamp 1606120353
transform 1 0 21068 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_215
timestamp 1606120353
transform 1 0 20884 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_219
timestamp 1606120353
transform 1 0 21252 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _0850_
timestamp 1606120353
transform 1 0 21620 0 1 32096
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__A1
timestamp 1606120353
transform 1 0 21436 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__D
timestamp 1606120353
transform 1 0 23000 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__CLK
timestamp 1606120353
transform 1 0 23368 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_236
timestamp 1606120353
transform 1 0 22816 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_240
timestamp 1606120353
transform 1 0 23184 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1606120353
transform 1 0 23552 0 1 32096
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__D
timestamp 1606120353
transform 1 0 23828 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__CLK
timestamp 1606120353
transform 1 0 24196 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__CLK
timestamp 1606120353
transform 1 0 24564 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_245
timestamp 1606120353
transform 1 0 23644 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_249
timestamp 1606120353
transform 1 0 24012 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_55_253
timestamp 1606120353
transform 1 0 24380 0 1 32096
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_55_257
timestamp 1606120353
transform 1 0 24748 0 1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_55_269
timestamp 1606120353
transform 1 0 25852 0 1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1606120353
transform 1 0 26956 0 1 32096
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1606120353
transform -1 0 28888 0 1 32096
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_55_293
timestamp 1606120353
transform 1 0 28060 0 1 32096
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1606120353
transform 1 0 1104 0 -1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1606120353
transform 1 0 1380 0 -1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_56_15
timestamp 1606120353
transform 1 0 2484 0 -1 33184
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_56_23
timestamp 1606120353
transform 1 0 3220 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__CLK
timestamp 1606120353
transform 1 0 3404 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_27
timestamp 1606120353
transform 1 0 3588 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__B2
timestamp 1606120353
transform 1 0 3772 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_56_32
timestamp 1606120353
transform 1 0 4048 0 -1 33184
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1606120353
transform 1 0 3956 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_56_36
timestamp 1606120353
transform 1 0 4416 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__B2
timestamp 1606120353
transform 1 0 4508 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_56_42
timestamp 1606120353
transform 1 0 4968 0 -1 33184
box 0 -48 368 592
use sky130_fd_sc_hd__buf_1  _0669_
timestamp 1606120353
transform 1 0 4692 0 -1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1200_
timestamp 1606120353
transform 1 0 5704 0 -1 33184
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0656__B
timestamp 1606120353
transform 1 0 5336 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_48
timestamp 1606120353
transform 1 0 5520 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0655_
timestamp 1606120353
transform 1 0 8188 0 -1 33184
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__B1
timestamp 1606120353
transform 1 0 9200 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__A1
timestamp 1606120353
transform 1 0 7636 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__B
timestamp 1606120353
transform 1 0 8004 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_69
timestamp 1606120353
transform 1 0 7452 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_73
timestamp 1606120353
transform 1 0 7820 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_56_84
timestamp 1606120353
transform 1 0 8832 0 -1 33184
box 0 -48 368 592
use sky130_fd_sc_hd__a211o_4  _0657_
timestamp 1606120353
transform 1 0 9660 0 -1 33184
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1606120353
transform 1 0 9568 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__A
timestamp 1606120353
transform 1 0 11132 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_90
timestamp 1606120353
transform 1 0 9384 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_107
timestamp 1606120353
transform 1 0 10948 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0566_
timestamp 1606120353
transform 1 0 11684 0 -1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__a32o_4  _0590_
timestamp 1606120353
transform 1 0 12696 0 -1 33184
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__A
timestamp 1606120353
transform 1 0 12420 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0566__A
timestamp 1606120353
transform 1 0 11500 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_111
timestamp 1606120353
transform 1 0 11316 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_56_118
timestamp 1606120353
transform 1 0 11960 0 -1 33184
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_56_122
timestamp 1606120353
transform 1 0 12328 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_56_125
timestamp 1606120353
transform 1 0 12604 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _0645_
timestamp 1606120353
transform 1 0 15272 0 -1 33184
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1606120353
transform 1 0 15180 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__C
timestamp 1606120353
transform 1 0 14444 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0589__A
timestamp 1606120353
transform 1 0 14812 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_143
timestamp 1606120353
transform 1 0 14260 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_147
timestamp 1606120353
transform 1 0 14628 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_151
timestamp 1606120353
transform 1 0 14996 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1211_
timestamp 1606120353
transform 1 0 17204 0 -1 33184
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0589__B
timestamp 1606120353
transform 1 0 16284 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__C
timestamp 1606120353
transform 1 0 16652 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__A
timestamp 1606120353
transform 1 0 17020 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_163
timestamp 1606120353
transform 1 0 16100 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_167
timestamp 1606120353
transform 1 0 16468 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_171
timestamp 1606120353
transform 1 0 16836 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__A2
timestamp 1606120353
transform 1 0 19136 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_194
timestamp 1606120353
transform 1 0 18952 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_198
timestamp 1606120353
transform 1 0 19320 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0490_
timestamp 1606120353
transform 1 0 19688 0 -1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1138_
timestamp 1606120353
transform 1 0 20884 0 -1 33184
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1606120353
transform 1 0 20792 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0490__A
timestamp 1606120353
transform 1 0 20148 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__A
timestamp 1606120353
transform 1 0 20608 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__B1_N
timestamp 1606120353
transform 1 0 19504 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_205
timestamp 1606120353
transform 1 0 19964 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_56_209
timestamp 1606120353
transform 1 0 20332 0 -1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A1
timestamp 1606120353
transform 1 0 22816 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__D
timestamp 1606120353
transform 1 0 23184 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_234
timestamp 1606120353
transform 1 0 22632 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_238
timestamp 1606120353
transform 1 0 23000 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_56_242
timestamp 1606120353
transform 1 0 23368 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1196_
timestamp 1606120353
transform 1 0 23736 0 -1 33184
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0522__A
timestamp 1606120353
transform 1 0 23552 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1606120353
transform 1 0 26404 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__CLK
timestamp 1606120353
transform 1 0 26128 0 -1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_56_265
timestamp 1606120353
transform 1 0 25484 0 -1 33184
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_56_271
timestamp 1606120353
transform 1 0 26036 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_56_274
timestamp 1606120353
transform 1 0 26312 0 -1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_56_276
timestamp 1606120353
transform 1 0 26496 0 -1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1606120353
transform -1 0 28888 0 -1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_56_288
timestamp 1606120353
transform 1 0 27600 0 -1 33184
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_56_296
timestamp 1606120353
transform 1 0 28336 0 -1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1606120353
transform 1 0 1104 0 1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__D
timestamp 1606120353
transform 1 0 3036 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__B1
timestamp 1606120353
transform 1 0 2668 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1606120353
transform 1 0 1380 0 1 33184
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_57_15
timestamp 1606120353
transform 1 0 2484 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_19
timestamp 1606120353
transform 1 0 2852 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_23
timestamp 1606120353
transform 1 0 3220 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__D
timestamp 1606120353
transform 1 0 3404 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_27
timestamp 1606120353
transform 1 0 3588 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_31
timestamp 1606120353
transform 1 0 3956 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__A2
timestamp 1606120353
transform 1 0 3772 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0680__A
timestamp 1606120353
transform 1 0 4140 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0680_
timestamp 1606120353
transform 1 0 4324 0 1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_57_38
timestamp 1606120353
transform 1 0 4600 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__A
timestamp 1606120353
transform 1 0 4784 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_42
timestamp 1606120353
transform 1 0 4968 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0540__C
timestamp 1606120353
transform 1 0 5152 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0656_
timestamp 1606120353
transform 1 0 5336 0 1 33184
box 0 -48 644 592
use sky130_fd_sc_hd__o22a_4  _0821_
timestamp 1606120353
transform 1 0 7176 0 1 33184
box 0 -48 1288 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1606120353
transform 1 0 6716 0 1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0540__B
timestamp 1606120353
transform 1 0 6164 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0540__A
timestamp 1606120353
transform 1 0 6532 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0656__A
timestamp 1606120353
transform 1 0 6992 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_53
timestamp 1606120353
transform 1 0 5980 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_57
timestamp 1606120353
transform 1 0 6348 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_62
timestamp 1606120353
transform 1 0 6808 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__a32o_4  _0772_
timestamp 1606120353
transform 1 0 9200 0 1 33184
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__A1
timestamp 1606120353
transform 1 0 9016 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__A2
timestamp 1606120353
transform 1 0 8648 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_80
timestamp 1606120353
transform 1 0 8464 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_84
timestamp 1606120353
transform 1 0 8832 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__A1
timestamp 1606120353
transform 1 0 10948 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_105
timestamp 1606120353
transform 1 0 10764 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_57_109
timestamp 1606120353
transform 1 0 11132 0 1 33184
box 0 -48 368 592
use sky130_fd_sc_hd__and4_4  _0682_
timestamp 1606120353
transform 1 0 12420 0 1 33184
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1606120353
transform 1 0 12328 0 1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__D
timestamp 1606120353
transform 1 0 11960 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__B
timestamp 1606120353
transform 1 0 11592 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_57_113
timestamp 1606120353
transform 1 0 11500 0 1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_57_116
timestamp 1606120353
transform 1 0 11776 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_120
timestamp 1606120353
transform 1 0 12144 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_57_132
timestamp 1606120353
transform 1 0 13248 0 1 33184
box 0 -48 368 592
use sky130_fd_sc_hd__nor4_4  _0589_
timestamp 1606120353
transform 1 0 14812 0 1 33184
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__A
timestamp 1606120353
transform 1 0 13616 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__C
timestamp 1606120353
transform 1 0 13984 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__C
timestamp 1606120353
transform 1 0 14352 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_138
timestamp 1606120353
transform 1 0 13800 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_142
timestamp 1606120353
transform 1 0 14168 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_57_146
timestamp 1606120353
transform 1 0 14536 0 1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0570__A
timestamp 1606120353
transform 1 0 16836 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0589__C
timestamp 1606120353
transform 1 0 17204 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_57_166
timestamp 1606120353
transform 1 0 16376 0 1 33184
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_57_170
timestamp 1606120353
transform 1 0 16744 0 1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_57_173
timestamp 1606120353
transform 1 0 17020 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0522_
timestamp 1606120353
transform 1 0 18032 0 1 33184
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1606120353
transform 1 0 17940 0 1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__D
timestamp 1606120353
transform 1 0 19044 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__B
timestamp 1606120353
transform 1 0 17572 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_177
timestamp 1606120353
transform 1 0 17388 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_181
timestamp 1606120353
transform 1 0 17756 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_193
timestamp 1606120353
transform 1 0 18860 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_197
timestamp 1606120353
transform 1 0 19228 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0915_
timestamp 1606120353
transform 1 0 19872 0 1 33184
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__C
timestamp 1606120353
transform 1 0 21252 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__D
timestamp 1606120353
transform 1 0 19412 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_57_201
timestamp 1606120353
transform 1 0 19596 0 1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_57_217
timestamp 1606120353
transform 1 0 21068 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0579_
timestamp 1606120353
transform 1 0 21804 0 1 33184
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__B
timestamp 1606120353
transform 1 0 21620 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__B1_N
timestamp 1606120353
transform 1 0 22816 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A2
timestamp 1606120353
transform 1 0 23184 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_221
timestamp 1606120353
transform 1 0 21436 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_234
timestamp 1606120353
transform 1 0 22632 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_238
timestamp 1606120353
transform 1 0 23000 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_242
timestamp 1606120353
transform 1 0 23368 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_245
timestamp 1606120353
transform 1 0 23644 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__D
timestamp 1606120353
transform 1 0 23828 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1606120353
transform 1 0 23552 0 1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_57_249
timestamp 1606120353
transform 1 0 24012 0 1 33184
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__A1
timestamp 1606120353
transform 1 0 24380 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_259
timestamp 1606120353
transform 1 0 24932 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_57_255
timestamp 1606120353
transform 1 0 24564 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__A2
timestamp 1606120353
transform 1 0 24748 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_57_263
timestamp 1606120353
transform 1 0 25300 0 1 33184
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__B1
timestamp 1606120353
transform 1 0 25116 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1116_
timestamp 1606120353
transform 1 0 26128 0 1 33184
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__D
timestamp 1606120353
transform 1 0 25944 0 1 33184
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_57_269
timestamp 1606120353
transform 1 0 25852 0 1 33184
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1606120353
transform -1 0 28888 0 1 33184
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_57_291
timestamp 1606120353
transform 1 0 27876 0 1 33184
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1606120353
transform 1 0 1104 0 -1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__D
timestamp 1606120353
transform 1 0 1564 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_58_3
timestamp 1606120353
transform 1 0 1380 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_58_7
timestamp 1606120353
transform 1 0 1748 0 -1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_58_19
timestamp 1606120353
transform 1 0 2852 0 -1 34272
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__D
timestamp 1606120353
transform 1 0 3404 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_58_27
timestamp 1606120353
transform 1 0 3588 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__A1
timestamp 1606120353
transform 1 0 3772 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1606120353
transform 1 0 3956 0 -1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_58_32
timestamp 1606120353
transform 1 0 4048 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__B2
timestamp 1606120353
transform 1 0 4232 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0713_
timestamp 1606120353
transform 1 0 4416 0 -1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_58_39
timestamp 1606120353
transform 1 0 4692 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_58_43
timestamp 1606120353
transform 1 0 5060 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__C
timestamp 1606120353
transform 1 0 4876 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0540_
timestamp 1606120353
transform 1 0 5428 0 -1 34272
box 0 -48 828 592
use sky130_fd_sc_hd__dfxtp_4  _1114_
timestamp 1606120353
transform 1 0 6992 0 -1 34272
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__C
timestamp 1606120353
transform 1 0 6808 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__A3
timestamp 1606120353
transform 1 0 6440 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__B1
timestamp 1606120353
transform 1 0 5244 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_58_56
timestamp 1606120353
transform 1 0 6256 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_58_60
timestamp 1606120353
transform 1 0 6624 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__A2
timestamp 1606120353
transform 1 0 9016 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_58_83
timestamp 1606120353
transform 1 0 8740 0 -1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_58_88
timestamp 1606120353
transform 1 0 9200 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__a32o_4  _0735_
timestamp 1606120353
transform 1 0 9660 0 -1 34272
box 0 -48 1564 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1606120353
transform 1 0 9568 0 -1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__B2
timestamp 1606120353
transform 1 0 9384 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_58_110
timestamp 1606120353
transform 1 0 11224 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0681_
timestamp 1606120353
transform 1 0 11960 0 -1 34272
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__B
timestamp 1606120353
transform 1 0 12972 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__A
timestamp 1606120353
transform 1 0 11776 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__A
timestamp 1606120353
transform 1 0 11408 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_58_114
timestamp 1606120353
transform 1 0 11592 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_58_127
timestamp 1606120353
transform 1 0 12788 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_58_131
timestamp 1606120353
transform 1 0 13156 0 -1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__and4_4  _0643_
timestamp 1606120353
transform 1 0 13616 0 -1 34272
box 0 -48 828 592
use sky130_fd_sc_hd__or4_4  _0646_
timestamp 1606120353
transform 1 0 15272 0 -1 34272
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1606120353
transform 1 0 15180 0 -1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0644__B
timestamp 1606120353
transform 1 0 14628 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__B
timestamp 1606120353
transform 1 0 13432 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__B
timestamp 1606120353
transform 1 0 14996 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_58_145
timestamp 1606120353
transform 1 0 14444 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_58_149
timestamp 1606120353
transform 1 0 14812 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _0570_
timestamp 1606120353
transform 1 0 16836 0 -1 34272
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__A
timestamp 1606120353
transform 1 0 16284 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0542__C
timestamp 1606120353
transform 1 0 16652 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_58_163
timestamp 1606120353
transform 1 0 16100 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_58_167
timestamp 1606120353
transform 1 0 16468 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1132_
timestamp 1606120353
transform 1 0 18216 0 -1 34272
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0542__A
timestamp 1606120353
transform 1 0 17664 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0561__B
timestamp 1606120353
transform 1 0 18032 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_58_178
timestamp 1606120353
transform 1 0 17480 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_58_182
timestamp 1606120353
transform 1 0 17848 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0580_
timestamp 1606120353
transform 1 0 20884 0 -1 34272
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1606120353
transform 1 0 20792 0 -1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__B
timestamp 1606120353
transform 1 0 20608 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A2
timestamp 1606120353
transform 1 0 20148 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_58_205
timestamp 1606120353
transform 1 0 19964 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_58_209
timestamp 1606120353
transform 1 0 20332 0 -1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__a21bo_4  _0924_
timestamp 1606120353
transform 1 0 22448 0 -1 34272
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__A
timestamp 1606120353
transform 1 0 21896 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__C
timestamp 1606120353
transform 1 0 22264 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_58_224
timestamp 1606120353
transform 1 0 21712 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_58_228
timestamp 1606120353
transform 1 0 22080 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0849_
timestamp 1606120353
transform 1 0 24380 0 -1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__CLK
timestamp 1606120353
transform 1 0 23828 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__CLK
timestamp 1606120353
transform 1 0 24196 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_58_245
timestamp 1606120353
transform 1 0 23644 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_58_249
timestamp 1606120353
transform 1 0 24012 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1606120353
transform 1 0 26404 0 -1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__CLK
timestamp 1606120353
transform 1 0 26128 0 -1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_58_265
timestamp 1606120353
transform 1 0 25484 0 -1 34272
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_58_271
timestamp 1606120353
transform 1 0 26036 0 -1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_58_274
timestamp 1606120353
transform 1 0 26312 0 -1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_58_276
timestamp 1606120353
transform 1 0 26496 0 -1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1606120353
transform -1 0 28888 0 -1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_58_288
timestamp 1606120353
transform 1 0 27600 0 -1 34272
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_58_296
timestamp 1606120353
transform 1 0 28336 0 -1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1164_
timestamp 1606120353
transform 1 0 1380 0 1 34272
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1606120353
transform 1 0 1104 0 1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1606120353
transform 1 0 1104 0 -1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__CLK
timestamp 1606120353
transform 1 0 1564 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_59_22
timestamp 1606120353
transform 1 0 3128 0 1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_60_3
timestamp 1606120353
transform 1 0 1380 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_60_7
timestamp 1606120353
transform 1 0 1748 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_60_19
timestamp 1606120353
transform 1 0 2852 0 -1 35360
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__A2
timestamp 1606120353
transform 1 0 3404 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__B1
timestamp 1606120353
transform 1 0 3404 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_60_27
timestamp 1606120353
transform 1 0 3588 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_59_27
timestamp 1606120353
transform 1 0 3588 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__A
timestamp 1606120353
transform 1 0 3772 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__B1
timestamp 1606120353
transform 1 0 3772 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_60_32
timestamp 1606120353
transform 1 0 4048 0 -1 35360
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_59_31
timestamp 1606120353
transform 1 0 3956 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0652__A
timestamp 1606120353
transform 1 0 4140 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1606120353
transform 1 0 3956 0 -1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_60_36
timestamp 1606120353
transform 1 0 4416 0 -1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_59_38
timestamp 1606120353
transform 1 0 4600 0 1 34272
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__A2
timestamp 1606120353
transform 1 0 4508 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0652_
timestamp 1606120353
transform 1 0 4324 0 1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_60_39
timestamp 1606120353
transform 1 0 4692 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_59_42
timestamp 1606120353
transform 1 0 4968 0 1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__D
timestamp 1606120353
transform 1 0 4876 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0539__A
timestamp 1606120353
transform 1 0 5060 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0539_
timestamp 1606120353
transform 1 0 5060 0 -1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_60_50
timestamp 1606120353
transform 1 0 5704 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_60_46
timestamp 1606120353
transform 1 0 5336 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_59_53
timestamp 1606120353
transform 1 0 5980 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_59_45
timestamp 1606120353
transform 1 0 5244 0 1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__B
timestamp 1606120353
transform 1 0 5520 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__A
timestamp 1606120353
transform 1 0 5888 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__B
timestamp 1606120353
transform 1 0 6164 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0797_
timestamp 1606120353
transform 1 0 5336 0 1 34272
box 0 -48 644 592
use sky130_fd_sc_hd__buf_1  _0514_
timestamp 1606120353
transform 1 0 6072 0 -1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_60_61
timestamp 1606120353
transform 1 0 6716 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_60_57
timestamp 1606120353
transform 1 0 6348 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_59_62
timestamp 1606120353
transform 1 0 6808 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_59_57
timestamp 1606120353
transform 1 0 6348 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__A1
timestamp 1606120353
transform 1 0 6532 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__D
timestamp 1606120353
transform 1 0 6900 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0514__A
timestamp 1606120353
transform 1 0 6532 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1606120353
transform 1 0 6716 0 1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0515_
timestamp 1606120353
transform 1 0 6992 0 1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1098_
timestamp 1606120353
transform 1 0 7084 0 -1 35360
box 0 -48 1748 592
use sky130_fd_sc_hd__o22a_4  _0800_
timestamp 1606120353
transform 1 0 8004 0 1 34272
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0515__A
timestamp 1606120353
transform 1 0 7452 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__A
timestamp 1606120353
transform 1 0 9016 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__C
timestamp 1606120353
transform 1 0 7820 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_59_67
timestamp 1606120353
transform 1 0 7268 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_59_71
timestamp 1606120353
transform 1 0 7636 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_60_84
timestamp 1606120353
transform 1 0 8832 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_60_88
timestamp 1606120353
transform 1 0 9200 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_59_95
timestamp 1606120353
transform 1 0 9844 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_59_89
timestamp 1606120353
transform 1 0 9292 0 1 34272
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0546__C
timestamp 1606120353
transform 1 0 9384 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__B
timestamp 1606120353
transform 1 0 9660 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1606120353
transform 1 0 9568 0 -1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _0739_
timestamp 1606120353
transform 1 0 9660 0 -1 35360
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_60_106
timestamp 1606120353
transform 1 0 10856 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_60_102
timestamp 1606120353
transform 1 0 10488 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_59_109
timestamp 1606120353
transform 1 0 11132 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__A
timestamp 1606120353
transform 1 0 11040 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0546__B
timestamp 1606120353
transform 1 0 10672 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0744_
timestamp 1606120353
transform 1 0 11224 0 -1 35360
box 0 -48 828 592
use sky130_fd_sc_hd__a21o_4  _0798_
timestamp 1606120353
transform 1 0 10028 0 1 34272
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_60_119
timestamp 1606120353
transform 1 0 12052 0 -1 35360
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_59_118
timestamp 1606120353
transform 1 0 11960 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_59_113
timestamp 1606120353
transform 1 0 11500 0 1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__C
timestamp 1606120353
transform 1 0 11776 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__A
timestamp 1606120353
transform 1 0 11316 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_60_126
timestamp 1606120353
transform 1 0 12696 0 -1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_60_123
timestamp 1606120353
transform 1 0 12420 0 -1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_59_123
timestamp 1606120353
transform 1 0 12420 0 1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__B
timestamp 1606120353
transform 1 0 12512 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__A
timestamp 1606120353
transform 1 0 12144 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1606120353
transform 1 0 12328 0 1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__or4_4  _0743_
timestamp 1606120353
transform 1 0 12788 0 -1 35360
box 0 -48 828 592
use sky130_fd_sc_hd__and4_4  _0741_
timestamp 1606120353
transform 1 0 12512 0 1 34272
box 0 -48 828 592
use sky130_fd_sc_hd__decap_4  FILLER_60_136
timestamp 1606120353
transform 1 0 13616 0 -1 35360
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_59_137
timestamp 1606120353
transform 1 0 13708 0 1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_59_133
timestamp 1606120353
transform 1 0 13340 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0644__A
timestamp 1606120353
transform 1 0 13984 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__C
timestamp 1606120353
transform 1 0 13984 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__B
timestamp 1606120353
transform 1 0 13524 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_60_150
timestamp 1606120353
transform 1 0 14904 0 -1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_60_146
timestamp 1606120353
transform 1 0 14536 0 -1 35360
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_60_142
timestamp 1606120353
transform 1 0 14168 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__A
timestamp 1606120353
transform 1 0 14352 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0644_
timestamp 1606120353
transform 1 0 14168 0 1 34272
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  FILLER_59_151
timestamp 1606120353
transform 1 0 14996 0 1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__C
timestamp 1606120353
transform 1 0 14996 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__A
timestamp 1606120353
transform 1 0 15272 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1606120353
transform 1 0 15180 0 -1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _0724_
timestamp 1606120353
transform 1 0 15272 0 -1 35360
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_60_163
timestamp 1606120353
transform 1 0 16100 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_59_156
timestamp 1606120353
transform 1 0 15456 0 1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__and4_4  _0642_
timestamp 1606120353
transform 1 0 15732 0 1 34272
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_60_167
timestamp 1606120353
transform 1 0 16468 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_59_172
timestamp 1606120353
transform 1 0 16928 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_59_168
timestamp 1606120353
transform 1 0 16560 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0586__C
timestamp 1606120353
transform 1 0 16652 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0556__D
timestamp 1606120353
transform 1 0 16284 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__B
timestamp 1606120353
transform 1 0 16744 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0542_
timestamp 1606120353
transform 1 0 16836 0 -1 35360
box 0 -48 828 592
use sky130_fd_sc_hd__decap_4  FILLER_59_176
timestamp 1606120353
transform 1 0 17296 0 1 34272
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0542__B
timestamp 1606120353
transform 1 0 17112 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_60_180
timestamp 1606120353
transform 1 0 17664 0 -1 35360
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_59_180
timestamp 1606120353
transform 1 0 17664 0 1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__B
timestamp 1606120353
transform 1 0 18032 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0561__A
timestamp 1606120353
transform 1 0 17756 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1606120353
transform 1 0 17940 0 1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__or4_4  _0561_
timestamp 1606120353
transform 1 0 18032 0 1 34272
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_60_186
timestamp 1606120353
transform 1 0 18216 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_59_193
timestamp 1606120353
transform 1 0 18860 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0516_
timestamp 1606120353
transform 1 0 18400 0 -1 35360
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_60_197
timestamp 1606120353
transform 1 0 19228 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_59_197
timestamp 1606120353
transform 1 0 19228 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__C
timestamp 1606120353
transform 1 0 19044 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_60_206
timestamp 1606120353
transform 1 0 20056 0 -1 35360
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_60_201
timestamp 1606120353
transform 1 0 19596 0 -1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_59_206
timestamp 1606120353
transform 1 0 20056 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_59_201
timestamp 1606120353
transform 1 0 19596 0 1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0644__D
timestamp 1606120353
transform 1 0 19412 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A1
timestamp 1606120353
transform 1 0 19872 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__B1
timestamp 1606120353
transform 1 0 19872 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__A2
timestamp 1606120353
transform 1 0 20240 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__D
timestamp 1606120353
transform 1 0 19412 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_60_215
timestamp 1606120353
transform 1 0 20884 0 -1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_60_212
timestamp 1606120353
transform 1 0 20608 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__A1
timestamp 1606120353
transform 1 0 20424 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1606120353
transform 1 0 20792 0 -1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__o21ai_4  _0871_
timestamp 1606120353
transform 1 0 20424 0 1 34272
box 0 -48 1196 592
use sky130_fd_sc_hd__o21a_4  _0870_
timestamp 1606120353
transform 1 0 21160 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_60_230
timestamp 1606120353
transform 1 0 22264 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_59_231
timestamp 1606120353
transform 1 0 22356 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_59_227
timestamp 1606120353
transform 1 0 21988 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_59_223
timestamp 1606120353
transform 1 0 21620 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__B1
timestamp 1606120353
transform 1 0 22172 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A2
timestamp 1606120353
transform 1 0 21804 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_60_234
timestamp 1606120353
transform 1 0 22632 0 -1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_59_240
timestamp 1606120353
transform 1 0 23184 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_59_235
timestamp 1606120353
transform 1 0 22724 0 1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__CLK
timestamp 1606120353
transform 1 0 22908 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0561__D
timestamp 1606120353
transform 1 0 22448 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A1
timestamp 1606120353
transform 1 0 22540 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__D
timestamp 1606120353
transform 1 0 23000 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__D
timestamp 1606120353
transform 1 0 23368 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1130_
timestamp 1606120353
transform 1 0 23092 0 -1 35360
box 0 -48 1748 592
use sky130_fd_sc_hd__dfxtp_4  _1184_
timestamp 1606120353
transform 1 0 23644 0 1 34272
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1606120353
transform 1 0 23552 0 1 34272
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_59_264
timestamp 1606120353
transform 1 0 25392 0 1 34272
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_60_258
timestamp 1606120353
transform 1 0 24840 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1152_
timestamp 1606120353
transform 1 0 26128 0 1 34272
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1606120353
transform 1 0 26404 0 -1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__D
timestamp 1606120353
transform 1 0 25944 0 1 34272
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__CLK
timestamp 1606120353
transform 1 0 26128 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_60_270
timestamp 1606120353
transform 1 0 25944 0 -1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_60_274
timestamp 1606120353
transform 1 0 26312 0 -1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_60_276
timestamp 1606120353
transform 1 0 26496 0 -1 35360
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1606120353
transform -1 0 28888 0 1 34272
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1606120353
transform -1 0 28888 0 -1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_59_291
timestamp 1606120353
transform 1 0 27876 0 1 34272
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_60_288
timestamp 1606120353
transform 1 0 27600 0 -1 35360
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_60_296
timestamp 1606120353
transform 1 0 28336 0 -1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__or2_4  _1082_
timestamp 1606120353
transform 1 0 2300 0 1 35360
box 0 -48 644 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1606120353
transform 1 0 1104 0 1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__A
timestamp 1606120353
transform 1 0 3128 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__B
timestamp 1606120353
transform 1 0 2116 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__CLK
timestamp 1606120353
transform 1 0 1564 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_3
timestamp 1606120353
transform 1 0 1380 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_61_7
timestamp 1606120353
transform 1 0 1748 0 1 35360
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_61_20
timestamp 1606120353
transform 1 0 2944 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0653_
timestamp 1606120353
transform 1 0 4692 0 1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__D
timestamp 1606120353
transform 1 0 5152 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0521__D
timestamp 1606120353
transform 1 0 4508 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__CLK
timestamp 1606120353
transform 1 0 4140 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_61_24
timestamp 1606120353
transform 1 0 3312 0 1 35360
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_61_32
timestamp 1606120353
transform 1 0 4048 0 1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_61_35
timestamp 1606120353
transform 1 0 4324 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_42
timestamp 1606120353
transform 1 0 4968 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_46
timestamp 1606120353
transform 1 0 5336 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0653__A
timestamp 1606120353
transform 1 0 5520 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0511_
timestamp 1606120353
transform 1 0 5704 0 1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_61_53
timestamp 1606120353
transform 1 0 5980 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0511__A
timestamp 1606120353
transform 1 0 6164 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_57
timestamp 1606120353
transform 1 0 6348 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__A
timestamp 1606120353
transform 1 0 6532 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_62
timestamp 1606120353
transform 1 0 6808 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1606120353
transform 1 0 6716 0 1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__C
timestamp 1606120353
transform 1 0 6992 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_66
timestamp 1606120353
transform 1 0 7176 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0721_
timestamp 1606120353
transform 1 0 7544 0 1 35360
box 0 -48 828 592
use sky130_fd_sc_hd__and4_4  _0723_
timestamp 1606120353
transform 1 0 9108 0 1 35360
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0521__A
timestamp 1606120353
transform 1 0 8556 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__B
timestamp 1606120353
transform 1 0 8924 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__B
timestamp 1606120353
transform 1 0 7360 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_79
timestamp 1606120353
transform 1 0 8372 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_83
timestamp 1606120353
transform 1 0 8740 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0740_
timestamp 1606120353
transform 1 0 10672 0 1 35360
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0546__A
timestamp 1606120353
transform 1 0 10120 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__B
timestamp 1606120353
transform 1 0 10488 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_96
timestamp 1606120353
transform 1 0 9936 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_100
timestamp 1606120353
transform 1 0 10304 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0726_
timestamp 1606120353
transform 1 0 12420 0 1 35360
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1606120353
transform 1 0 12328 0 1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__A
timestamp 1606120353
transform 1 0 12144 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__C
timestamp 1606120353
transform 1 0 11776 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_61_113
timestamp 1606120353
transform 1 0 11500 0 1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_61_118
timestamp 1606120353
transform 1 0 11960 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_132
timestamp 1606120353
transform 1 0 13248 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0738_
timestamp 1606120353
transform 1 0 13984 0 1 35360
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__B
timestamp 1606120353
transform 1 0 13432 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__B
timestamp 1606120353
transform 1 0 13800 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0556__A
timestamp 1606120353
transform 1 0 14996 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_136
timestamp 1606120353
transform 1 0 13616 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_149
timestamp 1606120353
transform 1 0 14812 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_153
timestamp 1606120353
transform 1 0 15180 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0556_
timestamp 1606120353
transform 1 0 15548 0 1 35360
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0556__B
timestamp 1606120353
transform 1 0 15364 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0586__A
timestamp 1606120353
transform 1 0 16836 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0586__B
timestamp 1606120353
transform 1 0 17204 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_61_166
timestamp 1606120353
transform 1 0 16376 0 1 35360
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_61_170
timestamp 1606120353
transform 1 0 16744 0 1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_61_173
timestamp 1606120353
transform 1 0 17020 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0585_
timestamp 1606120353
transform 1 0 18032 0 1 35360
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1606120353
transform 1 0 17940 0 1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__A
timestamp 1606120353
transform 1 0 17756 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0581__A
timestamp 1606120353
transform 1 0 19044 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_61_177
timestamp 1606120353
transform 1 0 17388 0 1 35360
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_61_193
timestamp 1606120353
transform 1 0 18860 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_61_197
timestamp 1606120353
transform 1 0 19228 0 1 35360
box 0 -48 368 592
use sky130_fd_sc_hd__inv_8  _0848_
timestamp 1606120353
transform 1 0 21344 0 1 35360
box 0 -48 828 592
use sky130_fd_sc_hd__inv_8  _0869_
timestamp 1606120353
transform 1 0 19780 0 1 35360
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__A
timestamp 1606120353
transform 1 0 21160 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__B1_N
timestamp 1606120353
transform 1 0 20792 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__A
timestamp 1606120353
transform 1 0 19596 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_212
timestamp 1606120353
transform 1 0 20608 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_216
timestamp 1606120353
transform 1 0 20976 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A2
timestamp 1606120353
transform 1 0 22356 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1160__D
timestamp 1606120353
transform 1 0 23368 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A1
timestamp 1606120353
transform 1 0 22724 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_229
timestamp 1606120353
transform 1 0 22172 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_61_233
timestamp 1606120353
transform 1 0 22540 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_61_237
timestamp 1606120353
transform 1 0 22908 0 1 35360
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_61_241
timestamp 1606120353
transform 1 0 23276 0 1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1160_
timestamp 1606120353
transform 1 0 23644 0 1 35360
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1606120353
transform 1 0 23552 0 1 35360
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_61_264
timestamp 1606120353
transform 1 0 25392 0 1 35360
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1151_
timestamp 1606120353
transform 1 0 26128 0 1 35360
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__D
timestamp 1606120353
transform 1 0 25944 0 1 35360
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1606120353
transform -1 0 28888 0 1 35360
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_61_291
timestamp 1606120353
transform 1 0 27876 0 1 35360
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1606120353
transform 1 0 1104 0 -1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__D
timestamp 1606120353
transform 1 0 1840 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__CLK
timestamp 1606120353
transform 1 0 2208 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_62_3
timestamp 1606120353
transform 1 0 1380 0 -1 36448
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_62_7
timestamp 1606120353
transform 1 0 1748 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_62_10
timestamp 1606120353
transform 1 0 2024 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_62_14
timestamp 1606120353
transform 1 0 2392 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1146_
timestamp 1606120353
transform 1 0 4600 0 -1 36448
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1606120353
transform 1 0 3956 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_62_26
timestamp 1606120353
transform 1 0 3496 0 -1 36448
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_62_30
timestamp 1606120353
transform 1 0 3864 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_62_32
timestamp 1606120353
transform 1 0 4048 0 -1 36448
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__D
timestamp 1606120353
transform 1 0 6808 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_62_57
timestamp 1606120353
transform 1 0 6348 0 -1 36448
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_62_61
timestamp 1606120353
transform 1 0 6716 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_62_64
timestamp 1606120353
transform 1 0 6992 0 -1 36448
box 0 -48 368 592
use sky130_fd_sc_hd__and4_4  _0521_
timestamp 1606120353
transform 1 0 8004 0 -1 36448
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0521__B
timestamp 1606120353
transform 1 0 7820 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0521__C
timestamp 1606120353
transform 1 0 7452 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__C
timestamp 1606120353
transform 1 0 9016 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_62_68
timestamp 1606120353
transform 1 0 7360 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_62_71
timestamp 1606120353
transform 1 0 7636 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_62_84
timestamp 1606120353
transform 1 0 8832 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_62_88
timestamp 1606120353
transform 1 0 9200 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__nor4_4  _0546_
timestamp 1606120353
transform 1 0 9844 0 -1 36448
box 0 -48 1564 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1606120353
transform 1 0 9568 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0546__D
timestamp 1606120353
transform 1 0 9384 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_62_93
timestamp 1606120353
transform 1 0 9660 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0742_
timestamp 1606120353
transform 1 0 12880 0 -1 36448
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__B
timestamp 1606120353
transform 1 0 12420 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__D
timestamp 1606120353
transform 1 0 12052 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__D
timestamp 1606120353
transform 1 0 11592 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_62_112
timestamp 1606120353
transform 1 0 11408 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_62_116
timestamp 1606120353
transform 1 0 11776 0 -1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_62_121
timestamp 1606120353
transform 1 0 12236 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_62_125
timestamp 1606120353
transform 1 0 12604 0 -1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__inv_8  _0555_
timestamp 1606120353
transform 1 0 15272 0 -1 36448
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1606120353
transform 1 0 15180 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__A
timestamp 1606120353
transform 1 0 14444 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__A
timestamp 1606120353
transform 1 0 13892 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0644__C
timestamp 1606120353
transform 1 0 14812 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_62_137
timestamp 1606120353
transform 1 0 13708 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_62_141
timestamp 1606120353
transform 1 0 14076 0 -1 36448
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_62_147
timestamp 1606120353
transform 1 0 14628 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_62_151
timestamp 1606120353
transform 1 0 14996 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0586_
timestamp 1606120353
transform 1 0 16836 0 -1 36448
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0576__B
timestamp 1606120353
transform 1 0 16652 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__B
timestamp 1606120353
transform 1 0 16284 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_62_163
timestamp 1606120353
transform 1 0 16100 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_62_167
timestamp 1606120353
transform 1 0 16468 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0581_
timestamp 1606120353
transform 1 0 18400 0 -1 36448
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__C
timestamp 1606120353
transform 1 0 18032 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__D
timestamp 1606120353
transform 1 0 19228 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_62_180
timestamp 1606120353
transform 1 0 17664 0 -1 36448
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_62_186
timestamp 1606120353
transform 1 0 18216 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_62_195
timestamp 1606120353
transform 1 0 19044 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_62_199
timestamp 1606120353
transform 1 0 19412 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__C
timestamp 1606120353
transform 1 0 19596 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_62_206
timestamp 1606120353
transform 1 0 20056 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0504_
timestamp 1606120353
transform 1 0 19780 0 -1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_62_210
timestamp 1606120353
transform 1 0 20424 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__D
timestamp 1606120353
transform 1 0 20240 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__B
timestamp 1606120353
transform 1 0 20608 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1606120353
transform 1 0 20792 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_62_215
timestamp 1606120353
transform 1 0 20884 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0504__A
timestamp 1606120353
transform 1 0 21068 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_62_219
timestamp 1606120353
transform 1 0 21252 0 -1 36448
box 0 -48 368 592
use sky130_fd_sc_hd__a21bo_4  _0938_
timestamp 1606120353
transform 1 0 21620 0 -1 36448
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_8  FILLER_62_236
timestamp 1606120353
transform 1 0 22816 0 -1 36448
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1160__CLK
timestamp 1606120353
transform 1 0 23644 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_62_244
timestamp 1606120353
transform 1 0 23552 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_62_247
timestamp 1606120353
transform 1 0 23828 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_62_259
timestamp 1606120353
transform 1 0 24932 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_565
timestamp 1606120353
transform 1 0 26404 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__CLK
timestamp 1606120353
transform 1 0 26128 0 -1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_62_271
timestamp 1606120353
transform 1 0 26036 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_62_274
timestamp 1606120353
transform 1 0 26312 0 -1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_62_276
timestamp 1606120353
transform 1 0 26496 0 -1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1606120353
transform -1 0 28888 0 -1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_62_288
timestamp 1606120353
transform 1 0 27600 0 -1 36448
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_62_296
timestamp 1606120353
transform 1 0 28336 0 -1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1145_
timestamp 1606120353
transform 1 0 1840 0 1 36448
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1606120353
transform 1 0 1104 0 1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__D
timestamp 1606120353
transform 1 0 1564 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_3
timestamp 1606120353
transform 1 0 1380 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_63_7
timestamp 1606120353
transform 1 0 1748 0 1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1606120353
transform 1 0 3588 0 1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_63_39
timestamp 1606120353
transform 1 0 4692 0 1 36448
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1122_
timestamp 1606120353
transform 1 0 6808 0 1 36448
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_566
timestamp 1606120353
transform 1 0 6716 0 1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__D
timestamp 1606120353
transform 1 0 6532 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__B
timestamp 1606120353
transform 1 0 6164 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__D
timestamp 1606120353
transform 1 0 5796 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__CLK
timestamp 1606120353
transform 1 0 5428 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_49
timestamp 1606120353
transform 1 0 5612 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_53
timestamp 1606120353
transform 1 0 5980 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_57
timestamp 1606120353
transform 1 0 6348 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__B
timestamp 1606120353
transform 1 0 9200 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__A
timestamp 1606120353
transform 1 0 8832 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_63_81
timestamp 1606120353
transform 1 0 8556 0 1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_63_86
timestamp 1606120353
transform 1 0 9016 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _0659_
timestamp 1606120353
transform 1 0 9384 0 1 36448
box 0 -48 644 592
use sky130_fd_sc_hd__or4_4  _0728_
timestamp 1606120353
transform 1 0 10764 0 1 36448
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0659__A
timestamp 1606120353
transform 1 0 10212 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__A
timestamp 1606120353
transform 1 0 10580 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_97
timestamp 1606120353
transform 1 0 10028 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_101
timestamp 1606120353
transform 1 0 10396 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0727_
timestamp 1606120353
transform 1 0 12880 0 1 36448
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_567
timestamp 1606120353
transform 1 0 12328 0 1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__B
timestamp 1606120353
transform 1 0 11776 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__A
timestamp 1606120353
transform 1 0 12696 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__C
timestamp 1606120353
transform 1 0 12144 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_114
timestamp 1606120353
transform 1 0 11592 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_118
timestamp 1606120353
transform 1 0 11960 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_63_123
timestamp 1606120353
transform 1 0 12420 0 1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__and4_4  _0558_
timestamp 1606120353
transform 1 0 14444 0 1 36448
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__B
timestamp 1606120353
transform 1 0 13892 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__D
timestamp 1606120353
transform 1 0 14260 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_137
timestamp 1606120353
transform 1 0 13708 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_141
timestamp 1606120353
transform 1 0 14076 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_154
timestamp 1606120353
transform 1 0 15272 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0587_
timestamp 1606120353
transform 1 0 16008 0 1 36448
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0576__D
timestamp 1606120353
transform 1 0 17020 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__A
timestamp 1606120353
transform 1 0 15824 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__C
timestamp 1606120353
transform 1 0 15456 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_158
timestamp 1606120353
transform 1 0 15640 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_171
timestamp 1606120353
transform 1 0 16836 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_175
timestamp 1606120353
transform 1 0 17204 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_179
timestamp 1606120353
transform 1 0 17572 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0576__A
timestamp 1606120353
transform 1 0 17388 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0576__C
timestamp 1606120353
transform 1 0 17756 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_568
timestamp 1606120353
transform 1 0 17940 0 1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0564_
timestamp 1606120353
transform 1 0 18032 0 1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_63_187
timestamp 1606120353
transform 1 0 18308 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_191
timestamp 1606120353
transform 1 0 18676 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0517__A
timestamp 1606120353
transform 1 0 18492 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0564__A
timestamp 1606120353
transform 1 0 18860 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0503_
timestamp 1606120353
transform 1 0 19044 0 1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_63_198
timestamp 1606120353
transform 1 0 19320 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _0914_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 20608 0 1 36448
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__A
timestamp 1606120353
transform 1 0 20424 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0570__B
timestamp 1606120353
transform 1 0 19504 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0503__A
timestamp 1606120353
transform 1 0 19872 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_202
timestamp 1606120353
transform 1 0 19688 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_63_206
timestamp 1606120353
transform 1 0 20056 0 1 36448
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__A2
timestamp 1606120353
transform 1 0 21804 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__B1_N
timestamp 1606120353
transform 1 0 22172 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__A1
timestamp 1606120353
transform 1 0 22540 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_63_221
timestamp 1606120353
transform 1 0 21436 0 1 36448
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_63_227
timestamp 1606120353
transform 1 0 21988 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_63_231
timestamp 1606120353
transform 1 0 22356 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_63_235
timestamp 1606120353
transform 1 0 22724 0 1 36448
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_569
timestamp 1606120353
transform 1 0 23552 0 1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__D
timestamp 1606120353
transform 1 0 23920 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__CLK
timestamp 1606120353
transform 1 0 24288 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_63_243
timestamp 1606120353
transform 1 0 23460 0 1 36448
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_63_245
timestamp 1606120353
transform 1 0 23644 0 1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_63_250
timestamp 1606120353
transform 1 0 24104 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_63_254
timestamp 1606120353
transform 1 0 24472 0 1 36448
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1223_
timestamp 1606120353
transform 1 0 26128 0 1 36448
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__D
timestamp 1606120353
transform 1 0 25944 0 1 36448
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_63_266
timestamp 1606120353
transform 1 0 25576 0 1 36448
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1606120353
transform -1 0 28888 0 1 36448
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_63_291
timestamp 1606120353
transform 1 0 27876 0 1 36448
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1190_
timestamp 1606120353
transform 1 0 1380 0 -1 37536
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1606120353
transform 1 0 1104 0 -1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_64_22
timestamp 1606120353
transform 1 0 3128 0 -1 37536
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_570
timestamp 1606120353
transform 1 0 3956 0 -1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_64_30
timestamp 1606120353
transform 1 0 3864 0 -1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_64_32
timestamp 1606120353
transform 1 0 4048 0 -1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_64_44
timestamp 1606120353
transform 1 0 5152 0 -1 37536
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1126_
timestamp 1606120353
transform 1 0 6992 0 -1 37536
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__D
timestamp 1606120353
transform 1 0 6808 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__CLK
timestamp 1606120353
transform 1 0 6440 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__CLK
timestamp 1606120353
transform 1 0 6072 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_52
timestamp 1606120353
transform 1 0 5888 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_56
timestamp 1606120353
transform 1 0 6256 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_60
timestamp 1606120353
transform 1 0 6624 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__C
timestamp 1606120353
transform 1 0 9016 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_64_83
timestamp 1606120353
transform 1 0 8740 0 -1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_64_88
timestamp 1606120353
transform 1 0 9200 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0717_
timestamp 1606120353
transform 1 0 9752 0 -1 37536
box 0 -48 644 592
use sky130_fd_sc_hd__and4_4  _0722_
timestamp 1606120353
transform 1 0 11132 0 -1 37536
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_571
timestamp 1606120353
transform 1 0 9568 0 -1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__A
timestamp 1606120353
transform 1 0 10764 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0659__B
timestamp 1606120353
transform 1 0 9384 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_64_93
timestamp 1606120353
transform 1 0 9660 0 -1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_64_101
timestamp 1606120353
transform 1 0 10396 0 -1 37536
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_64_107
timestamp 1606120353
transform 1 0 10948 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0725_
timestamp 1606120353
transform 1 0 13064 0 -1 37536
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0507__A
timestamp 1606120353
transform 1 0 12512 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__A
timestamp 1606120353
transform 1 0 12880 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__C
timestamp 1606120353
transform 1 0 12144 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_118
timestamp 1606120353
transform 1 0 11960 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_122
timestamp 1606120353
transform 1 0 12328 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_126
timestamp 1606120353
transform 1 0 12696 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0588_
timestamp 1606120353
transform 1 0 15272 0 -1 37536
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_572
timestamp 1606120353
transform 1 0 15180 0 -1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__C
timestamp 1606120353
transform 1 0 14444 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__A
timestamp 1606120353
transform 1 0 14996 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__D
timestamp 1606120353
transform 1 0 14076 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_139
timestamp 1606120353
transform 1 0 13892 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_143
timestamp 1606120353
transform 1 0 14260 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_64_147
timestamp 1606120353
transform 1 0 14628 0 -1 37536
box 0 -48 368 592
use sky130_fd_sc_hd__or4_4  _0576_
timestamp 1606120353
transform 1 0 16836 0 -1 37536
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__C
timestamp 1606120353
transform 1 0 16284 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__D
timestamp 1606120353
transform 1 0 16652 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_163
timestamp 1606120353
transform 1 0 16100 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_167
timestamp 1606120353
transform 1 0 16468 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0517_
timestamp 1606120353
transform 1 0 18400 0 -1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__D
timestamp 1606120353
transform 1 0 17848 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0586__D
timestamp 1606120353
transform 1 0 18216 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0581__B
timestamp 1606120353
transform 1 0 18860 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0516__A
timestamp 1606120353
transform 1 0 19228 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_180
timestamp 1606120353
transform 1 0 17664 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_184
timestamp 1606120353
transform 1 0 18032 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_191
timestamp 1606120353
transform 1 0 18676 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_195
timestamp 1606120353
transform 1 0 19044 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_573
timestamp 1606120353
transform 1 0 20792 0 -1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__B1_N
timestamp 1606120353
transform 1 0 20148 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0555__A
timestamp 1606120353
transform 1 0 19596 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_64_199
timestamp 1606120353
transform 1 0 19412 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_64_203
timestamp 1606120353
transform 1 0 19780 0 -1 37536
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_64_209
timestamp 1606120353
transform 1 0 20332 0 -1 37536
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_64_213
timestamp 1606120353
transform 1 0 20700 0 -1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_64_215
timestamp 1606120353
transform 1 0 20884 0 -1 37536
box 0 -48 736 592
use sky130_fd_sc_hd__a21bo_4  _0939_
timestamp 1606120353
transform 1 0 21804 0 -1 37536
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_64_223
timestamp 1606120353
transform 1 0 21620 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_64_238
timestamp 1606120353
transform 1 0 23000 0 -1 37536
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1163_
timestamp 1606120353
transform 1 0 23920 0 -1 37536
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__A2
timestamp 1606120353
transform 1 0 23644 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_64_244
timestamp 1606120353
transform 1 0 23552 0 -1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_64_247
timestamp 1606120353
transform 1 0 23828 0 -1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_574
timestamp 1606120353
transform 1 0 26404 0 -1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__CLK
timestamp 1606120353
transform 1 0 26128 0 -1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_64_267
timestamp 1606120353
transform 1 0 25668 0 -1 37536
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_64_271
timestamp 1606120353
transform 1 0 26036 0 -1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_64_274
timestamp 1606120353
transform 1 0 26312 0 -1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_64_276
timestamp 1606120353
transform 1 0 26496 0 -1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1606120353
transform -1 0 28888 0 -1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_64_288
timestamp 1606120353
transform 1 0 27600 0 -1 37536
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_64_296
timestamp 1606120353
transform 1 0 28336 0 -1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1606120353
transform 1 0 1104 0 1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1606120353
transform 1 0 1380 0 1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1606120353
transform 1 0 2484 0 1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1606120353
transform 1 0 3588 0 1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1606120353
transform 1 0 4692 0 1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_575
timestamp 1606120353
transform 1 0 6716 0 1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__D
timestamp 1606120353
transform 1 0 7084 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_65_51
timestamp 1606120353
transform 1 0 5796 0 1 37536
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_65_59
timestamp 1606120353
transform 1 0 6532 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_65_62
timestamp 1606120353
transform 1 0 6808 0 1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_65_67
timestamp 1606120353
transform 1 0 7268 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__A2
timestamp 1606120353
transform 1 0 7452 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_71
timestamp 1606120353
transform 1 0 7636 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_75
timestamp 1606120353
transform 1 0 8004 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__C1
timestamp 1606120353
transform 1 0 7820 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__A
timestamp 1606120353
transform 1 0 8188 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0508_
timestamp 1606120353
transform 1 0 8372 0 1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_65_82
timestamp 1606120353
transform 1 0 8648 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0508__A
timestamp 1606120353
transform 1 0 8832 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_86
timestamp 1606120353
transform 1 0 9016 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__A
timestamp 1606120353
transform 1 0 9200 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0716_
timestamp 1606120353
transform 1 0 9384 0 1 37536
box 0 -48 644 592
use sky130_fd_sc_hd__or4_4  _0718_
timestamp 1606120353
transform 1 0 10764 0 1 37536
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__B1
timestamp 1606120353
transform 1 0 10212 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__C
timestamp 1606120353
transform 1 0 10580 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_97
timestamp 1606120353
transform 1 0 10028 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_101
timestamp 1606120353
transform 1 0 10396 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0544_
timestamp 1606120353
transform 1 0 12420 0 1 37536
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_576
timestamp 1606120353
transform 1 0 12328 0 1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0544__B
timestamp 1606120353
transform 1 0 12144 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0544__A
timestamp 1606120353
transform 1 0 11776 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_114
timestamp 1606120353
transform 1 0 11592 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_118
timestamp 1606120353
transform 1 0 11960 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_132
timestamp 1606120353
transform 1 0 13248 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0616_
timestamp 1606120353
transform 1 0 13984 0 1 37536
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__B
timestamp 1606120353
transform 1 0 13800 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0544__C
timestamp 1606120353
transform 1 0 13432 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__B
timestamp 1606120353
transform 1 0 14996 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_136
timestamp 1606120353
transform 1 0 13616 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_149
timestamp 1606120353
transform 1 0 14812 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_153
timestamp 1606120353
transform 1 0 15180 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0584_
timestamp 1606120353
transform 1 0 15548 0 1 37536
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__A
timestamp 1606120353
transform 1 0 15364 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0506__A
timestamp 1606120353
transform 1 0 16560 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__D
timestamp 1606120353
transform 1 0 16928 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__D
timestamp 1606120353
transform 1 0 17296 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_166
timestamp 1606120353
transform 1 0 16376 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_170
timestamp 1606120353
transform 1 0 16744 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_174
timestamp 1606120353
transform 1 0 17112 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_184
timestamp 1606120353
transform 1 0 18032 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_65_182
timestamp 1606120353
transform 1 0 17848 0 1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_65_178
timestamp 1606120353
transform 1 0 17480 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0542__D
timestamp 1606120353
transform 1 0 17664 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_577
timestamp 1606120353
transform 1 0 17940 0 1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_65_192
timestamp 1606120353
transform 1 0 18768 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_65_188
timestamp 1606120353
transform 1 0 18400 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__B
timestamp 1606120353
transform 1 0 18584 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0561__C
timestamp 1606120353
transform 1 0 18216 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_65_196
timestamp 1606120353
transform 1 0 19136 0 1 37536
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__B
timestamp 1606120353
transform 1 0 18952 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0919_
timestamp 1606120353
transform 1 0 20148 0 1 37536
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__A2
timestamp 1606120353
transform 1 0 19964 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_65_204
timestamp 1606120353
transform 1 0 19872 0 1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_65_220
timestamp 1606120353
transform 1 0 21344 0 1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__B1_N
timestamp 1606120353
transform 1 0 23368 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_65_232
timestamp 1606120353
transform 1 0 22448 0 1 37536
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_65_240
timestamp 1606120353
transform 1 0 23184 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0931_
timestamp 1606120353
transform 1 0 23644 0 1 37536
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_578
timestamp 1606120353
transform 1 0 23552 0 1 37536
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_65_258
timestamp 1606120353
transform 1 0 24840 0 1 37536
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1121_
timestamp 1606120353
transform 1 0 26128 0 1 37536
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__D
timestamp 1606120353
transform 1 0 25944 0 1 37536
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1606120353
transform -1 0 28888 0 1 37536
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_65_291
timestamp 1606120353
transform 1 0 27876 0 1 37536
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1115_
timestamp 1606120353
transform 1 0 1564 0 1 38624
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1606120353
transform 1 0 1104 0 -1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1606120353
transform 1 0 1104 0 1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__D
timestamp 1606120353
transform 1 0 1564 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__CLK
timestamp 1606120353
transform 1 0 1932 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_66_3
timestamp 1606120353
transform 1 0 1380 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_66_7
timestamp 1606120353
transform 1 0 1748 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_66_11
timestamp 1606120353
transform 1 0 2116 0 -1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_67_3
timestamp 1606120353
transform 1 0 1380 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_579
timestamp 1606120353
transform 1 0 3956 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_66_23
timestamp 1606120353
transform 1 0 3220 0 -1 38624
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_66_32
timestamp 1606120353
transform 1 0 4048 0 -1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_66_44
timestamp 1606120353
transform 1 0 5152 0 -1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_67_24
timestamp 1606120353
transform 1 0 3312 0 1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_67_36
timestamp 1606120353
transform 1 0 4416 0 1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_584
timestamp 1606120353
transform 1 0 6716 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_66_56
timestamp 1606120353
transform 1 0 6256 0 -1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_67_48
timestamp 1606120353
transform 1 0 5520 0 1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_67_60
timestamp 1606120353
transform 1 0 6624 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_67_62
timestamp 1606120353
transform 1 0 6808 0 1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_67_74
timestamp 1606120353
transform 1 0 7912 0 1 38624
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_66_74
timestamp 1606120353
transform 1 0 7912 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_66_68
timestamp 1606120353
transform 1 0 7360 0 -1 38624
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_66_77
timestamp 1606120353
transform 1 0 8188 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__B
timestamp 1606120353
transform 1 0 8004 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__A
timestamp 1606120353
transform 1 0 8648 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__D
timestamp 1606120353
transform 1 0 8372 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0668_
timestamp 1606120353
transform 1 0 8556 0 -1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_67_88
timestamp 1606120353
transform 1 0 9200 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_67_84
timestamp 1606120353
transform 1 0 8832 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_66_88
timestamp 1606120353
transform 1 0 9200 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_66_84
timestamp 1606120353
transform 1 0 8832 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__C
timestamp 1606120353
transform 1 0 9016 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__A
timestamp 1606120353
transform 1 0 9016 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_67_99
timestamp 1606120353
transform 1 0 10212 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__A1
timestamp 1606120353
transform 1 0 9384 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0509__B
timestamp 1606120353
transform 1 0 9384 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_580
timestamp 1606120353
transform 1 0 9568 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _0509_
timestamp 1606120353
transform 1 0 9568 0 1 38624
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILLER_67_103
timestamp 1606120353
transform 1 0 10580 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_66_107
timestamp 1606120353
transform 1 0 10948 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__B2
timestamp 1606120353
transform 1 0 11132 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__A1
timestamp 1606120353
transform 1 0 10764 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0509__A
timestamp 1606120353
transform 1 0 10396 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _0720_
timestamp 1606120353
transform 1 0 10948 0 1 38624
box 0 -48 644 592
use sky130_fd_sc_hd__a211o_4  _0736_
timestamp 1606120353
transform 1 0 9660 0 -1 38624
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_67_118
timestamp 1606120353
transform 1 0 11960 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_67_114
timestamp 1606120353
transform 1 0 11592 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_66_115
timestamp 1606120353
transform 1 0 11684 0 -1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_66_111
timestamp 1606120353
transform 1 0 11316 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__B
timestamp 1606120353
transform 1 0 11500 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__A
timestamp 1606120353
transform 1 0 11960 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__B
timestamp 1606120353
transform 1 0 11776 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_66_120
timestamp 1606120353
transform 1 0 12144 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__A
timestamp 1606120353
transform 1 0 12144 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0544__D
timestamp 1606120353
transform 1 0 12328 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_585
timestamp 1606120353
transform 1 0 12328 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__and3_4  _0729_
timestamp 1606120353
transform 1 0 12420 0 1 38624
box 0 -48 828 592
use sky130_fd_sc_hd__inv_8  _0507_
timestamp 1606120353
transform 1 0 12512 0 -1 38624
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_67_132
timestamp 1606120353
transform 1 0 13248 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_67_136
timestamp 1606120353
transform 1 0 13616 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_66_137
timestamp 1606120353
transform 1 0 13708 0 -1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_66_133
timestamp 1606120353
transform 1 0 13340 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__B
timestamp 1606120353
transform 1 0 13524 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__B
timestamp 1606120353
transform 1 0 13432 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0505__B
timestamp 1606120353
transform 1 0 13800 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_66_145
timestamp 1606120353
transform 1 0 14444 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__D
timestamp 1606120353
transform 1 0 13984 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0565_
timestamp 1606120353
transform 1 0 14168 0 -1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__or2_4  _0505_
timestamp 1606120353
transform 1 0 13984 0 1 38624
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILLER_67_151
timestamp 1606120353
transform 1 0 14996 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_67_147
timestamp 1606120353
transform 1 0 14628 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_66_149
timestamp 1606120353
transform 1 0 14812 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__B
timestamp 1606120353
transform 1 0 15180 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__C
timestamp 1606120353
transform 1 0 14996 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0565__A
timestamp 1606120353
transform 1 0 14628 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0505__A
timestamp 1606120353
transform 1 0 14812 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_581
timestamp 1606120353
transform 1 0 15180 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0569_
timestamp 1606120353
transform 1 0 15272 0 -1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_66_157
timestamp 1606120353
transform 1 0 15548 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0510_
timestamp 1606120353
transform 1 0 15364 0 1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_67_158
timestamp 1606120353
transform 1 0 15640 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__C
timestamp 1606120353
transform 1 0 15732 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0533__A
timestamp 1606120353
transform 1 0 15824 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_67_162
timestamp 1606120353
transform 1 0 16008 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_66_161
timestamp 1606120353
transform 1 0 15916 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__D
timestamp 1606120353
transform 1 0 16100 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_67_166
timestamp 1606120353
transform 1 0 16376 0 1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__C
timestamp 1606120353
transform 1 0 16192 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0506_
timestamp 1606120353
transform 1 0 16284 0 -1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_66_168
timestamp 1606120353
transform 1 0 16560 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__A
timestamp 1606120353
transform 1 0 16652 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_67_171
timestamp 1606120353
transform 1 0 16836 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_66_172
timestamp 1606120353
transform 1 0 16928 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__D
timestamp 1606120353
transform 1 0 16744 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_67_175
timestamp 1606120353
transform 1 0 17204 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__A
timestamp 1606120353
transform 1 0 17112 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__B
timestamp 1606120353
transform 1 0 17020 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_66_176
timestamp 1606120353
transform 1 0 17296 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_67_179
timestamp 1606120353
transform 1 0 17572 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_66_186
timestamp 1606120353
transform 1 0 18216 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_66_180
timestamp 1606120353
transform 1 0 17664 0 -1 38624
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__CLK
timestamp 1606120353
transform 1 0 17388 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0556__C
timestamp 1606120353
transform 1 0 17480 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__D
timestamp 1606120353
transform 1 0 18032 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1156__D
timestamp 1606120353
transform 1 0 17756 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_586
timestamp 1606120353
transform 1 0 17940 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1156__CLK
timestamp 1606120353
transform 1 0 18400 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_66_190
timestamp 1606120353
transform 1 0 18584 0 -1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1156_
timestamp 1606120353
transform 1 0 18032 0 1 38624
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_4  FILLER_66_209
timestamp 1606120353
transform 1 0 20332 0 -1 38624
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_66_206
timestamp 1606120353
transform 1 0 20056 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_66_202
timestamp 1606120353
transform 1 0 19688 0 -1 38624
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__A1
timestamp 1606120353
transform 1 0 20148 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_67_219
timestamp 1606120353
transform 1 0 21252 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_67_215
timestamp 1606120353
transform 1 0 20884 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_66_213
timestamp 1606120353
transform 1 0 20700 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__A
timestamp 1606120353
transform 1 0 21068 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_582
timestamp 1606120353
transform 1 0 20792 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_67_203
timestamp 1606120353
transform 1 0 19780 0 1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_66_215
timestamp 1606120353
transform 1 0 20884 0 -1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__and2_4  _0844_
timestamp 1606120353
transform 1 0 21988 0 1 38624
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__A
timestamp 1606120353
transform 1 0 22816 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__B
timestamp 1606120353
transform 1 0 21804 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__B
timestamp 1606120353
transform 1 0 21436 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_66_227
timestamp 1606120353
transform 1 0 21988 0 -1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_66_239
timestamp 1606120353
transform 1 0 23092 0 -1 38624
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_67_223
timestamp 1606120353
transform 1 0 21620 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_67_234
timestamp 1606120353
transform 1 0 22632 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_67_238
timestamp 1606120353
transform 1 0 23000 0 1 38624
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_587
timestamp 1606120353
transform 1 0 23552 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A
timestamp 1606120353
transform 1 0 23828 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__A
timestamp 1606120353
transform 1 0 24564 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__A1
timestamp 1606120353
transform 1 0 23644 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_66_247
timestamp 1606120353
transform 1 0 23828 0 -1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_66_259
timestamp 1606120353
transform 1 0 24932 0 -1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_67_245
timestamp 1606120353
transform 1 0 23644 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_67_249
timestamp 1606120353
transform 1 0 24012 0 1 38624
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_67_257
timestamp 1606120353
transform 1 0 24748 0 1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1118_
timestamp 1606120353
transform 1 0 26128 0 1 38624
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_583
timestamp 1606120353
transform 1 0 26404 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__D
timestamp 1606120353
transform 1 0 25944 0 1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__CLK
timestamp 1606120353
transform 1 0 26128 0 -1 38624
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_66_271
timestamp 1606120353
transform 1 0 26036 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_66_274
timestamp 1606120353
transform 1 0 26312 0 -1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_66_276
timestamp 1606120353
transform 1 0 26496 0 -1 38624
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_67_269
timestamp 1606120353
transform 1 0 25852 0 1 38624
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1606120353
transform -1 0 28888 0 -1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1606120353
transform -1 0 28888 0 1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_66_288
timestamp 1606120353
transform 1 0 27600 0 -1 38624
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_66_296
timestamp 1606120353
transform 1 0 28336 0 -1 38624
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_67_291
timestamp 1606120353
transform 1 0 27876 0 1 38624
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1606120353
transform 1 0 1104 0 -1 39712
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__D
timestamp 1606120353
transform 1 0 1564 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_68_3
timestamp 1606120353
transform 1 0 1380 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_68_7
timestamp 1606120353
transform 1 0 1748 0 -1 39712
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_68_19
timestamp 1606120353
transform 1 0 2852 0 -1 39712
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_588
timestamp 1606120353
transform 1 0 3956 0 -1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_68_32
timestamp 1606120353
transform 1 0 4048 0 -1 39712
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_68_44
timestamp 1606120353
transform 1 0 5152 0 -1 39712
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_68_56
timestamp 1606120353
transform 1 0 6256 0 -1 39712
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__B1
timestamp 1606120353
transform 1 0 9016 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_68_68
timestamp 1606120353
transform 1 0 7360 0 -1 39712
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_68_80
timestamp 1606120353
transform 1 0 8464 0 -1 39712
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_68_88
timestamp 1606120353
transform 1 0 9200 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_68_98
timestamp 1606120353
transform 1 0 10120 0 -1 39712
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_68_93
timestamp 1606120353
transform 1 0 9660 0 -1 39712
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__A3
timestamp 1606120353
transform 1 0 9384 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__A1
timestamp 1606120353
transform 1 0 9936 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_589
timestamp 1606120353
transform 1 0 9568 0 -1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_68_107
timestamp 1606120353
transform 1 0 10948 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_68_103
timestamp 1606120353
transform 1 0 10580 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__D
timestamp 1606120353
transform 1 0 10764 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__A
timestamp 1606120353
transform 1 0 10396 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__a32o_4  _0731_
timestamp 1606120353
transform 1 0 11132 0 -1 39712
box 0 -48 1564 592
use sky130_fd_sc_hd__and3_4  _0745_
timestamp 1606120353
transform 1 0 12696 0 -1 39712
box 0 -48 828 592
use sky130_fd_sc_hd__buf_1  _0533_
timestamp 1606120353
transform 1 0 15272 0 -1 39712
box 0 -48 276 592
use sky130_fd_sc_hd__or2_4  _0737_
timestamp 1606120353
transform 1 0 13524 0 -1 39712
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_590
timestamp 1606120353
transform 1 0 15180 0 -1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__D
timestamp 1606120353
transform 1 0 14352 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__A
timestamp 1606120353
transform 1 0 14720 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_68_142
timestamp 1606120353
transform 1 0 14168 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_68_146
timestamp 1606120353
transform 1 0 14536 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_68_150
timestamp 1606120353
transform 1 0 14904 0 -1 39712
box 0 -48 276 592
use sky130_fd_sc_hd__and2_4  _0748_
timestamp 1606120353
transform 1 0 16652 0 -1 39712
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__D
timestamp 1606120353
transform 1 0 15732 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0510__A
timestamp 1606120353
transform 1 0 16100 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0569__A
timestamp 1606120353
transform 1 0 16468 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_68_157
timestamp 1606120353
transform 1 0 15548 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_68_161
timestamp 1606120353
transform 1 0 15916 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_68_165
timestamp 1606120353
transform 1 0 16284 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_68_176
timestamp 1606120353
transform 1 0 17296 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1148_
timestamp 1606120353
transform 1 0 18032 0 -1 39712
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__CLK
timestamp 1606120353
transform 1 0 17480 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_68_180
timestamp 1606120353
transform 1 0 17664 0 -1 39712
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_591
timestamp 1606120353
transform 1 0 20792 0 -1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__A
timestamp 1606120353
transform 1 0 21344 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_68_203
timestamp 1606120353
transform 1 0 19780 0 -1 39712
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_68_211
timestamp 1606120353
transform 1 0 20516 0 -1 39712
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_68_215
timestamp 1606120353
transform 1 0 20884 0 -1 39712
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_68_219
timestamp 1606120353
transform 1 0 21252 0 -1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _0828_
timestamp 1606120353
transform 1 0 21528 0 -1 39712
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0880__B
timestamp 1606120353
transform 1 0 22356 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_68_229
timestamp 1606120353
transform 1 0 22172 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_68_233
timestamp 1606120353
transform 1 0 22540 0 -1 39712
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_68_241
timestamp 1606120353
transform 1 0 23276 0 -1 39712
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0876_
timestamp 1606120353
transform 1 0 23552 0 -1 39712
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0877_
timestamp 1606120353
transform 1 0 24564 0 -1 39712
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__A2
timestamp 1606120353
transform 1 0 24012 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__C1
timestamp 1606120353
transform 1 0 24380 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_68_247
timestamp 1606120353
transform 1 0 23828 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_68_251
timestamp 1606120353
transform 1 0 24196 0 -1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_68_258
timestamp 1606120353
transform 1 0 24840 0 -1 39712
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_592
timestamp 1606120353
transform 1 0 26404 0 -1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_68_270
timestamp 1606120353
transform 1 0 25944 0 -1 39712
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_68_274
timestamp 1606120353
transform 1 0 26312 0 -1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_68_276
timestamp 1606120353
transform 1 0 26496 0 -1 39712
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1606120353
transform -1 0 28888 0 -1 39712
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_68_288
timestamp 1606120353
transform 1 0 27600 0 -1 39712
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_68_296
timestamp 1606120353
transform 1 0 28336 0 -1 39712
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1197_
timestamp 1606120353
transform 1 0 1472 0 1 39712
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1606120353
transform 1 0 1104 0 1 39712
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_69_3
timestamp 1606120353
transform 1 0 1380 0 1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_69_23
timestamp 1606120353
transform 1 0 3220 0 1 39712
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_69_35
timestamp 1606120353
transform 1 0 4324 0 1 39712
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_593
timestamp 1606120353
transform 1 0 6716 0 1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_69_47
timestamp 1606120353
transform 1 0 5428 0 1 39712
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_69_59
timestamp 1606120353
transform 1 0 6532 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_69_62
timestamp 1606120353
transform 1 0 6808 0 1 39712
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__A3
timestamp 1606120353
transform 1 0 9016 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_69_74
timestamp 1606120353
transform 1 0 7912 0 1 39712
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_69_88
timestamp 1606120353
transform 1 0 9200 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__a32o_4  _0747_
timestamp 1606120353
transform 1 0 9936 0 1 39712
box 0 -48 1564 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__B2
timestamp 1606120353
transform 1 0 9752 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__A2
timestamp 1606120353
transform 1 0 9384 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_69_92
timestamp 1606120353
transform 1 0 9568 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_69_113
timestamp 1606120353
transform 1 0 11500 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_69_117
timestamp 1606120353
transform 1 0 11868 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__A2
timestamp 1606120353
transform 1 0 11684 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_69_121
timestamp 1606120353
transform 1 0 12236 0 1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__B1
timestamp 1606120353
transform 1 0 12052 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_594
timestamp 1606120353
transform 1 0 12328 0 1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_69_123
timestamp 1606120353
transform 1 0 12420 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__B
timestamp 1606120353
transform 1 0 12604 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_69_127
timestamp 1606120353
transform 1 0 12788 0 1 39712
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_69_131
timestamp 1606120353
transform 1 0 13156 0 1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0513__A
timestamp 1606120353
transform 1 0 13248 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 13800 0 1 39712
box 0 -48 1840 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1606120353
transform 1 0 13616 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_69_134
timestamp 1606120353
transform 1 0 13432 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1086_
timestamp 1606120353
transform 1 0 15640 0 1 39712
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_595
timestamp 1606120353
transform 1 0 17940 0 1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__D
timestamp 1606120353
transform 1 0 17572 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_69_177
timestamp 1606120353
transform 1 0 17388 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_69_181
timestamp 1606120353
transform 1 0 17756 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_69_184
timestamp 1606120353
transform 1 0 18032 0 1 39712
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_69_196
timestamp 1606120353
transform 1 0 19136 0 1 39712
box 0 -48 1104 592
use sky130_fd_sc_hd__inv_8  _0827_
timestamp 1606120353
transform 1 0 21344 0 1 39712
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__A
timestamp 1606120353
transform 1 0 20976 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_69_208
timestamp 1606120353
transform 1 0 20240 0 1 39712
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_69_218
timestamp 1606120353
transform 1 0 21160 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0880__A
timestamp 1606120353
transform 1 0 22356 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__A
timestamp 1606120353
transform 1 0 23368 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__B1
timestamp 1606120353
transform 1 0 23000 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_69_229
timestamp 1606120353
transform 1 0 22172 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_69_233
timestamp 1606120353
transform 1 0 22540 0 1 39712
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_69_237
timestamp 1606120353
transform 1 0 22908 0 1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_69_240
timestamp 1606120353
transform 1 0 23184 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0907_
timestamp 1606120353
transform 1 0 25208 0 1 39712
box 0 -48 276 592
use sky130_fd_sc_hd__nor2_4  _0922_
timestamp 1606120353
transform 1 0 23644 0 1 39712
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_596
timestamp 1606120353
transform 1 0 23552 0 1 39712
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__B
timestamp 1606120353
transform 1 0 24656 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__A1
timestamp 1606120353
transform 1 0 25024 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_69_254
timestamp 1606120353
transform 1 0 24472 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_69_258
timestamp 1606120353
transform 1 0 24840 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__A
timestamp 1606120353
transform 1 0 25668 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_69_265
timestamp 1606120353
transform 1 0 25484 0 1 39712
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_69_269
timestamp 1606120353
transform 1 0 25852 0 1 39712
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_69_281
timestamp 1606120353
transform 1 0 26956 0 1 39712
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1606120353
transform -1 0 28888 0 1 39712
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_69_293
timestamp 1606120353
transform 1 0 28060 0 1 39712
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1606120353
transform 1 0 1104 0 -1 40800
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__CLK
timestamp 1606120353
transform 1 0 1564 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_70_3
timestamp 1606120353
transform 1 0 1380 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_70_7
timestamp 1606120353
transform 1 0 1748 0 -1 40800
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_70_19
timestamp 1606120353
transform 1 0 2852 0 -1 40800
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_597
timestamp 1606120353
transform 1 0 3956 0 -1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_70_32
timestamp 1606120353
transform 1 0 4048 0 -1 40800
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_70_44
timestamp 1606120353
transform 1 0 5152 0 -1 40800
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_70_56
timestamp 1606120353
transform 1 0 6256 0 -1 40800
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_70_68
timestamp 1606120353
transform 1 0 7360 0 -1 40800
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_70_80
timestamp 1606120353
transform 1 0 8464 0 -1 40800
box 0 -48 1104 592
use sky130_fd_sc_hd__buf_1  _0719_
timestamp 1606120353
transform 1 0 10396 0 -1 40800
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_598
timestamp 1606120353
transform 1 0 9568 0 -1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__B1
timestamp 1606120353
transform 1 0 10856 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__B1
timestamp 1606120353
transform 1 0 9936 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__A2
timestamp 1606120353
transform 1 0 11224 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_70_93
timestamp 1606120353
transform 1 0 9660 0 -1 40800
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_70_98
timestamp 1606120353
transform 1 0 10120 0 -1 40800
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_70_104
timestamp 1606120353
transform 1 0 10672 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_70_108
timestamp 1606120353
transform 1 0 11040 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__a211o_4  _0730_
timestamp 1606120353
transform 1 0 11408 0 -1 40800
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__C
timestamp 1606120353
transform 1 0 12880 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__C
timestamp 1606120353
transform 1 0 13248 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_70_126
timestamp 1606120353
transform 1 0 12696 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_70_130
timestamp 1606120353
transform 1 0 13064 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0513_
timestamp 1606120353
transform 1 0 13984 0 -1 40800
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_599
timestamp 1606120353
transform 1 0 15180 0 -1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_70_134
timestamp 1606120353
transform 1 0 13432 0 -1 40800
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILLER_70_143
timestamp 1606120353
transform 1 0 14260 0 -1 40800
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_70_151
timestamp 1606120353
transform 1 0 14996 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_70_154
timestamp 1606120353
transform 1 0 15272 0 -1 40800
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1117_
timestamp 1606120353
transform 1 0 16744 0 -1 40800
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__B1
timestamp 1606120353
transform 1 0 16100 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__D
timestamp 1606120353
transform 1 0 15640 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__CLK
timestamp 1606120353
transform 1 0 16468 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_70_160
timestamp 1606120353
transform 1 0 15824 0 -1 40800
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_70_165
timestamp 1606120353
transform 1 0 16284 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_70_169
timestamp 1606120353
transform 1 0 16652 0 -1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_70_189
timestamp 1606120353
transform 1 0 18492 0 -1 40800
box 0 -48 1104 592
use sky130_fd_sc_hd__buf_1  _0822_
timestamp 1606120353
transform 1 0 20976 0 -1 40800
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_600
timestamp 1606120353
transform 1 0 20792 0 -1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__A
timestamp 1606120353
transform 1 0 20608 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_70_201
timestamp 1606120353
transform 1 0 19596 0 -1 40800
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_70_209
timestamp 1606120353
transform 1 0 20332 0 -1 40800
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_70_215
timestamp 1606120353
transform 1 0 20884 0 -1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_70_219
timestamp 1606120353
transform 1 0 21252 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0880_
timestamp 1606120353
transform 1 0 21988 0 -1 40800
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__B1_N
timestamp 1606120353
transform 1 0 21436 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__A
timestamp 1606120353
transform 1 0 22816 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__B
timestamp 1606120353
transform 1 0 21804 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__A1
timestamp 1606120353
transform 1 0 23368 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_70_223
timestamp 1606120353
transform 1 0 21620 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_70_234
timestamp 1606120353
transform 1 0 22632 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_70_238
timestamp 1606120353
transform 1 0 23000 0 -1 40800
box 0 -48 368 592
use sky130_fd_sc_hd__a211o_4  _0923_
timestamp 1606120353
transform 1 0 23552 0 -1 40800
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__B1_N
timestamp 1606120353
transform 1 0 25024 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__CLK
timestamp 1606120353
transform 1 0 25392 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_70_258
timestamp 1606120353
transform 1 0 24840 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_70_262
timestamp 1606120353
transform 1 0 25208 0 -1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_601
timestamp 1606120353
transform 1 0 26404 0 -1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_70_266
timestamp 1606120353
transform 1 0 25576 0 -1 40800
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_70_274
timestamp 1606120353
transform 1 0 26312 0 -1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_70_276
timestamp 1606120353
transform 1 0 26496 0 -1 40800
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1606120353
transform -1 0 28888 0 -1 40800
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_70_288
timestamp 1606120353
transform 1 0 27600 0 -1 40800
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_70_296
timestamp 1606120353
transform 1 0 28336 0 -1 40800
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1606120353
transform 1 0 1104 0 1 40800
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1606120353
transform 1 0 1380 0 1 40800
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_71_15
timestamp 1606120353
transform 1 0 2484 0 1 40800
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_71_27
timestamp 1606120353
transform 1 0 3588 0 1 40800
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_71_39
timestamp 1606120353
transform 1 0 4692 0 1 40800
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_602
timestamp 1606120353
transform 1 0 6716 0 1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_71_51
timestamp 1606120353
transform 1 0 5796 0 1 40800
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_71_59
timestamp 1606120353
transform 1 0 6532 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_71_62
timestamp 1606120353
transform 1 0 6808 0 1 40800
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_71_74
timestamp 1606120353
transform 1 0 7912 0 1 40800
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_71_86
timestamp 1606120353
transform 1 0 9016 0 1 40800
box 0 -48 736 592
use sky130_fd_sc_hd__o21ai_4  _0551_
timestamp 1606120353
transform 1 0 10304 0 1 40800
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0551__A1
timestamp 1606120353
transform 1 0 10120 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0551__B1
timestamp 1606120353
transform 1 0 9752 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_71_96
timestamp 1606120353
transform 1 0 9936 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_71_121
timestamp 1606120353
transform 1 0 12236 0 1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_71_117
timestamp 1606120353
transform 1 0 11868 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_71_113
timestamp 1606120353
transform 1 0 11500 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__C1
timestamp 1606120353
transform 1 0 12052 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__A2
timestamp 1606120353
transform 1 0 11684 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_71_127
timestamp 1606120353
transform 1 0 12788 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_71_123
timestamp 1606120353
transform 1 0 12420 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__A1
timestamp 1606120353
transform 1 0 12972 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__C1
timestamp 1606120353
transform 1 0 12604 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_603
timestamp 1606120353
transform 1 0 12328 0 1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_71_131
timestamp 1606120353
transform 1 0 13156 0 1 40800
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_71_143
timestamp 1606120353
transform 1 0 14260 0 1 40800
box 0 -48 1104 592
use sky130_fd_sc_hd__a21o_4  _0749_
timestamp 1606120353
transform 1 0 16100 0 1 40800
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A1
timestamp 1606120353
transform 1 0 15916 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_71_155
timestamp 1606120353
transform 1 0 15364 0 1 40800
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILLER_71_175
timestamp 1606120353
transform 1 0 17204 0 1 40800
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_604
timestamp 1606120353
transform 1 0 17940 0 1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_71_184
timestamp 1606120353
transform 1 0 18032 0 1 40800
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_71_196
timestamp 1606120353
transform 1 0 19136 0 1 40800
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0825_
timestamp 1606120353
transform 1 0 19596 0 1 40800
box 0 -48 276 592
use sky130_fd_sc_hd__a21bo_4  _0829_
timestamp 1606120353
transform 1 0 20976 0 1 40800
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__A1
timestamp 1606120353
transform 1 0 20792 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__A
timestamp 1606120353
transform 1 0 20056 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__A2
timestamp 1606120353
transform 1 0 20424 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__A
timestamp 1606120353
transform 1 0 19412 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_71_204
timestamp 1606120353
transform 1 0 19872 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_71_208
timestamp 1606120353
transform 1 0 20240 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_71_212
timestamp 1606120353
transform 1 0 20608 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__B
timestamp 1606120353
transform 1 0 22356 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__C
timestamp 1606120353
transform 1 0 22724 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__A2
timestamp 1606120353
transform 1 0 23368 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_71_229
timestamp 1606120353
transform 1 0 22172 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_71_233
timestamp 1606120353
transform 1 0 22540 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_71_237
timestamp 1606120353
transform 1 0 22908 0 1 40800
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_71_241
timestamp 1606120353
transform 1 0 23276 0 1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0926_
timestamp 1606120353
transform 1 0 23736 0 1 40800
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1176_
timestamp 1606120353
transform 1 0 24748 0 1 40800
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_605
timestamp 1606120353
transform 1 0 23552 0 1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__D
timestamp 1606120353
transform 1 0 24564 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__A
timestamp 1606120353
transform 1 0 24196 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_71_245
timestamp 1606120353
transform 1 0 23644 0 1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_71_249
timestamp 1606120353
transform 1 0 24012 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_71_253
timestamp 1606120353
transform 1 0 24380 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0552__A
timestamp 1606120353
transform 1 0 26680 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_71_276
timestamp 1606120353
transform 1 0 26496 0 1 40800
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_71_280
timestamp 1606120353
transform 1 0 26864 0 1 40800
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1606120353
transform -1 0 28888 0 1 40800
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_71_292
timestamp 1606120353
transform 1 0 27968 0 1 40800
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_71_298
timestamp 1606120353
transform 1 0 28520 0 1 40800
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1606120353
transform 1 0 1104 0 -1 41888
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1606120353
transform 1 0 1104 0 1 41888
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__CLK
timestamp 1606120353
transform 1 0 1564 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1606120353
transform 1 0 1380 0 -1 41888
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_72_15
timestamp 1606120353
transform 1 0 2484 0 -1 41888
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_73_3
timestamp 1606120353
transform 1 0 1380 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_73_7
timestamp 1606120353
transform 1 0 1748 0 1 41888
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_73_19
timestamp 1606120353
transform 1 0 2852 0 1 41888
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_606
timestamp 1606120353
transform 1 0 3956 0 -1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_72_27
timestamp 1606120353
transform 1 0 3588 0 -1 41888
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_72_32
timestamp 1606120353
transform 1 0 4048 0 -1 41888
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_72_44
timestamp 1606120353
transform 1 0 5152 0 -1 41888
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_73_31
timestamp 1606120353
transform 1 0 3956 0 1 41888
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_73_43
timestamp 1606120353
transform 1 0 5060 0 1 41888
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_611
timestamp 1606120353
transform 1 0 6716 0 1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_72_56
timestamp 1606120353
transform 1 0 6256 0 -1 41888
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_73_55
timestamp 1606120353
transform 1 0 6164 0 1 41888
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_73_62
timestamp 1606120353
transform 1 0 6808 0 1 41888
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_73_77
timestamp 1606120353
transform 1 0 8188 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_73_74
timestamp 1606120353
transform 1 0 7912 0 1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__B1
timestamp 1606120353
transform 1 0 8004 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_72_87
timestamp 1606120353
transform 1 0 9108 0 -1 41888
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_72_83
timestamp 1606120353
transform 1 0 8740 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_72_80
timestamp 1606120353
transform 1 0 8464 0 -1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__B2
timestamp 1606120353
transform 1 0 8924 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__A2
timestamp 1606120353
transform 1 0 8556 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__A1
timestamp 1606120353
transform 1 0 8372 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_72_68
timestamp 1606120353
transform 1 0 7360 0 -1 41888
box 0 -48 1104 592
use sky130_fd_sc_hd__a32oi_4  _0658_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 8556 0 1 41888
box 0 -48 2024 592
use sky130_fd_sc_hd__fill_1  FILLER_72_99
timestamp 1606120353
transform 1 0 10212 0 -1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_72_93
timestamp 1606120353
transform 1 0 9660 0 -1 41888
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_72_91
timestamp 1606120353
transform 1 0 9476 0 -1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_607
timestamp 1606120353
transform 1 0 9568 0 -1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_73_107
timestamp 1606120353
transform 1 0 10948 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_73_103
timestamp 1606120353
transform 1 0 10580 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_72_102
timestamp 1606120353
transform 1 0 10488 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__A1
timestamp 1606120353
transform 1 0 10672 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__A2
timestamp 1606120353
transform 1 0 10764 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__A1
timestamp 1606120353
transform 1 0 11132 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0551__A2
timestamp 1606120353
transform 1 0 10304 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__a211o_4  _0746_
timestamp 1606120353
transform 1 0 10856 0 -1 41888
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_73_118
timestamp 1606120353
transform 1 0 11960 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_73_114
timestamp 1606120353
transform 1 0 11592 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0550__A
timestamp 1606120353
transform 1 0 12144 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__B1
timestamp 1606120353
transform 1 0 11776 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0550_
timestamp 1606120353
transform 1 0 11316 0 1 41888
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_73_123
timestamp 1606120353
transform 1 0 12420 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__C1
timestamp 1606120353
transform 1 0 12604 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_612
timestamp 1606120353
transform 1 0 12328 0 1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_73_127
timestamp 1606120353
transform 1 0 12788 0 1 41888
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_72_132
timestamp 1606120353
transform 1 0 13248 0 -1 41888
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_72_120
timestamp 1606120353
transform 1 0 12144 0 -1 41888
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_73_139
timestamp 1606120353
transform 1 0 13892 0 1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0591__B
timestamp 1606120353
transform 1 0 13984 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0591_
timestamp 1606120353
transform 1 0 14168 0 1 41888
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILLER_73_149
timestamp 1606120353
transform 1 0 14812 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_72_154
timestamp 1606120353
transform 1 0 15272 0 -1 41888
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_72_152
timestamp 1606120353
transform 1 0 15088 0 -1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_72_144
timestamp 1606120353
transform 1 0 14352 0 -1 41888
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0591__A
timestamp 1606120353
transform 1 0 14996 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_608
timestamp 1606120353
transform 1 0 15180 0 -1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_73_153
timestamp 1606120353
transform 1 0 15180 0 1 41888
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A2
timestamp 1606120353
transform 1 0 16100 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__CLK
timestamp 1606120353
transform 1 0 17296 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_72_162
timestamp 1606120353
transform 1 0 16008 0 -1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1606120353
transform 1 0 16284 0 -1 41888
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_73_165
timestamp 1606120353
transform 1 0 16284 0 1 41888
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_73_173
timestamp 1606120353
transform 1 0 17020 0 1 41888
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__CLK
timestamp 1606120353
transform 1 0 17572 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_72_177
timestamp 1606120353
transform 1 0 17388 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_73_178
timestamp 1606120353
transform 1 0 17480 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__B
timestamp 1606120353
transform 1 0 17664 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_72_181
timestamp 1606120353
transform 1 0 17756 0 -1 41888
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_73_182
timestamp 1606120353
transform 1 0 17848 0 1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_613
timestamp 1606120353
transform 1 0 17940 0 1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__D
timestamp 1606120353
transform 1 0 18032 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_73_184
timestamp 1606120353
transform 1 0 18032 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__D
timestamp 1606120353
transform 1 0 18216 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_73_198
timestamp 1606120353
transform 1 0 19320 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_73_194
timestamp 1606120353
transform 1 0 18952 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_73_188
timestamp 1606120353
transform 1 0 18400 0 1 41888
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_72_198
timestamp 1606120353
transform 1 0 19320 0 -1 41888
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__A
timestamp 1606120353
transform 1 0 19136 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0832_
timestamp 1606120353
transform 1 0 18676 0 1 41888
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_72_186
timestamp 1606120353
transform 1 0 18216 0 -1 41888
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_72_206
timestamp 1606120353
transform 1 0 20056 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A1
timestamp 1606120353
transform 1 0 19596 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__D
timestamp 1606120353
transform 1 0 20240 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A2
timestamp 1606120353
transform 1 0 19504 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0881_
timestamp 1606120353
transform 1 0 19780 0 -1 41888
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_73_218
timestamp 1606120353
transform 1 0 21160 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_73_214
timestamp 1606120353
transform 1 0 20792 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_72_210
timestamp 1606120353
transform 1 0 20424 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__A1
timestamp 1606120353
transform 1 0 20608 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__A1
timestamp 1606120353
transform 1 0 20976 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__B1
timestamp 1606120353
transform 1 0 21344 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_609
timestamp 1606120353
transform 1 0 20792 0 -1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__or2_4  _0859_
timestamp 1606120353
transform 1 0 20884 0 -1 41888
box 0 -48 644 592
use sky130_fd_sc_hd__a21o_4  _0913_
timestamp 1606120353
transform 1 0 19688 0 1 41888
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_72_226
timestamp 1606120353
transform 1 0 21896 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_72_222
timestamp 1606120353
transform 1 0 21528 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__A2
timestamp 1606120353
transform 1 0 22080 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__A1
timestamp 1606120353
transform 1 0 21712 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_73_238
timestamp 1606120353
transform 1 0 23000 0 1 41888
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_73_234
timestamp 1606120353
transform 1 0 22632 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__B1
timestamp 1606120353
transform 1 0 22816 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__A1
timestamp 1606120353
transform 1 0 23368 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__nor3_4  _0888_
timestamp 1606120353
transform 1 0 22264 0 -1 41888
box 0 -48 1196 592
use sky130_fd_sc_hd__o21a_4  _0860_
timestamp 1606120353
transform 1 0 21528 0 1 41888
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_72_250
timestamp 1606120353
transform 1 0 24104 0 -1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_72_247
timestamp 1606120353
transform 1 0 23828 0 -1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_72_243
timestamp 1606120353
transform 1 0 23460 0 -1 41888
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__D
timestamp 1606120353
transform 1 0 23920 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_614
timestamp 1606120353
transform 1 0 23552 0 1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_73_261
timestamp 1606120353
transform 1 0 25116 0 1 41888
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_73_257
timestamp 1606120353
transform 1 0 24748 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_72_264
timestamp 1606120353
transform 1 0 25392 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__B1
timestamp 1606120353
transform 1 0 24932 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0921_
timestamp 1606120353
transform 1 0 23644 0 1 41888
box 0 -48 1104 592
use sky130_fd_sc_hd__a21bo_4  _0889_
timestamp 1606120353
transform 1 0 24196 0 -1 41888
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_73_268
timestamp 1606120353
transform 1 0 25760 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_73_265
timestamp 1606120353
transform 1 0 25484 0 1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_72_274
timestamp 1606120353
transform 1 0 26312 0 -1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_72_268
timestamp 1606120353
transform 1 0 25760 0 -1 41888
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__CLK
timestamp 1606120353
transform 1 0 25576 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__D
timestamp 1606120353
transform 1 0 26128 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__A
timestamp 1606120353
transform 1 0 25576 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__B
timestamp 1606120353
transform 1 0 25944 0 1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_610
timestamp 1606120353
transform 1 0 26404 0 -1 41888
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_72_285
timestamp 1606120353
transform 1 0 27324 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0552_
timestamp 1606120353
transform 1 0 26496 0 -1 41888
box 0 -48 828 592
use sky130_fd_sc_hd__dfxtp_4  _1154_
timestamp 1606120353
transform 1 0 26128 0 1 41888
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1606120353
transform -1 0 28888 0 -1 41888
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1606120353
transform -1 0 28888 0 1 41888
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__CLK
timestamp 1606120353
transform 1 0 27508 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_72_289
timestamp 1606120353
transform 1 0 27692 0 -1 41888
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_72_297
timestamp 1606120353
transform 1 0 28428 0 -1 41888
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_73_291
timestamp 1606120353
transform 1 0 27876 0 1 41888
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1606120353
transform 1 0 1104 0 -1 42976
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1172__D
timestamp 1606120353
transform 1 0 1564 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__D
timestamp 1606120353
transform 1 0 1932 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1172__CLK
timestamp 1606120353
transform 1 0 2300 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_74_3
timestamp 1606120353
transform 1 0 1380 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_74_7
timestamp 1606120353
transform 1 0 1748 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_74_11
timestamp 1606120353
transform 1 0 2116 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1606120353
transform 1 0 2484 0 -1 42976
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_615
timestamp 1606120353
transform 1 0 3956 0 -1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_74_27
timestamp 1606120353
transform 1 0 3588 0 -1 42976
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_74_32
timestamp 1606120353
transform 1 0 4048 0 -1 42976
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_74_44
timestamp 1606120353
transform 1 0 5152 0 -1 42976
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_74_56
timestamp 1606120353
transform 1 0 6256 0 -1 42976
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__A3
timestamp 1606120353
transform 1 0 8556 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_74_68
timestamp 1606120353
transform 1 0 7360 0 -1 42976
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_74_80
timestamp 1606120353
transform 1 0 8464 0 -1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_74_83
timestamp 1606120353
transform 1 0 8740 0 -1 42976
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_616
timestamp 1606120353
transform 1 0 9568 0 -1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0623__B1
timestamp 1606120353
transform 1 0 11224 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_74_91
timestamp 1606120353
transform 1 0 9476 0 -1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_74_93
timestamp 1606120353
transform 1 0 9660 0 -1 42976
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_74_105
timestamp 1606120353
transform 1 0 10764 0 -1 42976
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_74_109
timestamp 1606120353
transform 1 0 11132 0 -1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__a211o_4  _0650_
timestamp 1606120353
transform 1 0 11408 0 -1 42976
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0621__A1
timestamp 1606120353
transform 1 0 12880 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_74_126
timestamp 1606120353
transform 1 0 12696 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_74_130
timestamp 1606120353
transform 1 0 13064 0 -1 42976
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_617
timestamp 1606120353
transform 1 0 15180 0 -1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_74_142
timestamp 1606120353
transform 1 0 14168 0 -1 42976
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_74_150
timestamp 1606120353
transform 1 0 14904 0 -1 42976
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_74_154
timestamp 1606120353
transform 1 0 15272 0 -1 42976
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__A
timestamp 1606120353
transform 1 0 16928 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_74_166
timestamp 1606120353
transform 1 0 16376 0 -1 42976
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILLER_74_174
timestamp 1606120353
transform 1 0 17112 0 -1 42976
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1157_
timestamp 1606120353
transform 1 0 17572 0 -1 42976
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__A
timestamp 1606120353
transform 1 0 17388 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_74_198
timestamp 1606120353
transform 1 0 19320 0 -1 42976
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_74_204
timestamp 1606120353
transform 1 0 19872 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__B1
timestamp 1606120353
transform 1 0 19688 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A
timestamp 1606120353
transform 1 0 20056 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_74_208
timestamp 1606120353
transform 1 0 20240 0 -1 42976
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_74_213
timestamp 1606120353
transform 1 0 20700 0 -1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__A2
timestamp 1606120353
transform 1 0 20516 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_74_215
timestamp 1606120353
transform 1 0 20884 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_618
timestamp 1606120353
transform 1 0 20792 0 -1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_74_219
timestamp 1606120353
transform 1 0 21252 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__A2
timestamp 1606120353
transform 1 0 21068 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__a211o_4  _0847_
timestamp 1606120353
transform 1 0 21620 0 -1 42976
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__C1
timestamp 1606120353
transform 1 0 21436 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__A1
timestamp 1606120353
transform 1 0 23092 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_74_237
timestamp 1606120353
transform 1 0 22908 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_74_241
timestamp 1606120353
transform 1 0 23276 0 -1 42976
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1183_
timestamp 1606120353
transform 1 0 23920 0 -1 42976
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__A2
timestamp 1606120353
transform 1 0 23644 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_74_247
timestamp 1606120353
transform 1 0 23828 0 -1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _0920_
timestamp 1606120353
transform 1 0 26496 0 -1 42976
box 0 -48 644 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_619
timestamp 1606120353
transform 1 0 26404 0 -1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__C
timestamp 1606120353
transform 1 0 27324 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__CLK
timestamp 1606120353
transform 1 0 25852 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__CLK
timestamp 1606120353
transform 1 0 26220 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_74_267
timestamp 1606120353
transform 1 0 25668 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_74_271
timestamp 1606120353
transform 1 0 26036 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_74_283
timestamp 1606120353
transform 1 0 27140 0 -1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1606120353
transform -1 0 28888 0 -1 42976
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_74_287
timestamp 1606120353
transform 1 0 27508 0 -1 42976
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1172_
timestamp 1606120353
transform 1 0 1472 0 1 42976
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1606120353
transform 1 0 1104 0 1 42976
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_75_3
timestamp 1606120353
transform 1 0 1380 0 1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_75_23
timestamp 1606120353
transform 1 0 3220 0 1 42976
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_75_35
timestamp 1606120353
transform 1 0 4324 0 1 42976
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_620
timestamp 1606120353
transform 1 0 6716 0 1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_75_47
timestamp 1606120353
transform 1 0 5428 0 1 42976
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_75_59
timestamp 1606120353
transform 1 0 6532 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_75_62
timestamp 1606120353
transform 1 0 6808 0 1 42976
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__B1_N
timestamp 1606120353
transform 1 0 7636 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__A2
timestamp 1606120353
transform 1 0 8004 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__A1
timestamp 1606120353
transform 1 0 8372 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_75_70
timestamp 1606120353
transform 1 0 7544 0 1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_75_73
timestamp 1606120353
transform 1 0 7820 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_77
timestamp 1606120353
transform 1 0 8188 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1606120353
transform 1 0 8556 0 1 42976
box 0 -48 1104 592
use sky130_fd_sc_hd__buf_1  _0501_
timestamp 1606120353
transform 1 0 10764 0 1 42976
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0501__A
timestamp 1606120353
transform 1 0 11224 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0623__A1
timestamp 1606120353
transform 1 0 10580 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_75_93
timestamp 1606120353
transform 1 0 9660 0 1 42976
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_75_101
timestamp 1606120353
transform 1 0 10396 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_108
timestamp 1606120353
transform 1 0 11040 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _0621_
timestamp 1606120353
transform 1 0 12880 0 1 42976
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_621
timestamp 1606120353
transform 1 0 12328 0 1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0493__A
timestamp 1606120353
transform 1 0 12696 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0623__A2
timestamp 1606120353
transform 1 0 11592 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0621__B1
timestamp 1606120353
transform 1 0 12144 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_112
timestamp 1606120353
transform 1 0 11408 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_75_116
timestamp 1606120353
transform 1 0 11776 0 1 42976
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_75_123
timestamp 1606120353
transform 1 0 12420 0 1 42976
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_75_141
timestamp 1606120353
transform 1 0 14076 0 1 42976
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_75_153
timestamp 1606120353
transform 1 0 15180 0 1 42976
box 0 -48 552 592
use sky130_fd_sc_hd__buf_1  _0824_
timestamp 1606120353
transform 1 0 16928 0 1 42976
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__A
timestamp 1606120353
transform 1 0 16100 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__B
timestamp 1606120353
transform 1 0 16468 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__C
timestamp 1606120353
transform 1 0 15732 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_161
timestamp 1606120353
transform 1 0 15916 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_165
timestamp 1606120353
transform 1 0 16284 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_75_169
timestamp 1606120353
transform 1 0 16652 0 1 42976
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_75_175
timestamp 1606120353
transform 1 0 17204 0 1 42976
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1149_
timestamp 1606120353
transform 1 0 18032 0 1 42976
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_622
timestamp 1606120353
transform 1 0 17940 0 1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__C
timestamp 1606120353
transform 1 0 17664 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_75_179
timestamp 1606120353
transform 1 0 17572 0 1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_75_182
timestamp 1606120353
transform 1 0 17848 0 1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__o21a_4  _0826_
timestamp 1606120353
transform 1 0 20516 0 1 42976
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__A1
timestamp 1606120353
transform 1 0 20332 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__C
timestamp 1606120353
transform 1 0 19964 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_203
timestamp 1606120353
transform 1 0 19780 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_207
timestamp 1606120353
transform 1 0 20148 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_223
timestamp 1606120353
transform 1 0 21620 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__A
timestamp 1606120353
transform 1 0 21804 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_227
timestamp 1606120353
transform 1 0 21988 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__A2
timestamp 1606120353
transform 1 0 22172 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_231
timestamp 1606120353
transform 1 0 22356 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0932_
timestamp 1606120353
transform 1 0 22540 0 1 42976
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_75_236
timestamp 1606120353
transform 1 0 22816 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__A
timestamp 1606120353
transform 1 0 23000 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_240
timestamp 1606120353
transform 1 0 23184 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__B1
timestamp 1606120353
transform 1 0 23368 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1169_
timestamp 1606120353
transform 1 0 24564 0 1 42976
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_623
timestamp 1606120353
transform 1 0 23552 0 1 42976
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__D
timestamp 1606120353
transform 1 0 24380 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__D
timestamp 1606120353
transform 1 0 23920 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_75_245
timestamp 1606120353
transform 1 0 23644 0 1 42976
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_75_250
timestamp 1606120353
transform 1 0 24104 0 1 42976
box 0 -48 276 592
use sky130_fd_sc_hd__and2_4  _0846_
timestamp 1606120353
transform 1 0 27048 0 1 42976
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__A
timestamp 1606120353
transform 1 0 26496 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__B
timestamp 1606120353
transform 1 0 26864 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_274
timestamp 1606120353
transform 1 0 26312 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_278
timestamp 1606120353
transform 1 0 26680 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1606120353
transform -1 0 28888 0 1 42976
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__B
timestamp 1606120353
transform 1 0 27876 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__D
timestamp 1606120353
transform 1 0 28244 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_289
timestamp 1606120353
transform 1 0 27692 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_293
timestamp 1606120353
transform 1 0 28060 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_75_297
timestamp 1606120353
transform 1 0 28428 0 1 42976
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1175_
timestamp 1606120353
transform 1 0 1472 0 -1 44064
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1606120353
transform 1 0 1104 0 -1 44064
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_76_3
timestamp 1606120353
transform 1 0 1380 0 -1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_624
timestamp 1606120353
transform 1 0 3956 0 -1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_76_23
timestamp 1606120353
transform 1 0 3220 0 -1 44064
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_76_32
timestamp 1606120353
transform 1 0 4048 0 -1 44064
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_76_44
timestamp 1606120353
transform 1 0 5152 0 -1 44064
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_76_56
timestamp 1606120353
transform 1 0 6256 0 -1 44064
box 0 -48 1104 592
use sky130_fd_sc_hd__a21bo_4  _0934_
timestamp 1606120353
transform 1 0 7636 0 -1 44064
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_3  FILLER_76_68
timestamp 1606120353
transform 1 0 7360 0 -1 44064
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_76_84
timestamp 1606120353
transform 1 0 8832 0 -1 44064
box 0 -48 736 592
use sky130_fd_sc_hd__o21a_4  _0623_
timestamp 1606120353
transform 1 0 11224 0 -1 44064
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_625
timestamp 1606120353
transform 1 0 9568 0 -1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_76_93
timestamp 1606120353
transform 1 0 9660 0 -1 44064
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_76_105
timestamp 1606120353
transform 1 0 10764 0 -1 44064
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_76_109
timestamp 1606120353
transform 1 0 11132 0 -1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0493_
timestamp 1606120353
transform 1 0 13064 0 -1 44064
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0492__C
timestamp 1606120353
transform 1 0 12512 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0621__A2
timestamp 1606120353
transform 1 0 12880 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_76_122
timestamp 1606120353
transform 1 0 12328 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_76_126
timestamp 1606120353
transform 1 0 12696 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_626
timestamp 1606120353
transform 1 0 15180 0 -1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_76_133
timestamp 1606120353
transform 1 0 13340 0 -1 44064
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_76_145
timestamp 1606120353
transform 1 0 14444 0 -1 44064
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_76_154
timestamp 1606120353
transform 1 0 15272 0 -1 44064
box 0 -48 736 592
use sky130_fd_sc_hd__and3_4  _0845_
timestamp 1606120353
transform 1 0 16100 0 -1 44064
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__A
timestamp 1606120353
transform 1 0 17112 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_76_162
timestamp 1606120353
transform 1 0 16008 0 -1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_76_172
timestamp 1606120353
transform 1 0 16928 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_76_176
timestamp 1606120353
transform 1 0 17296 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__or3_4  _0831_
timestamp 1606120353
transform 1 0 17664 0 -1 44064
box 0 -48 828 592
use sky130_fd_sc_hd__inv_8  _0840_
timestamp 1606120353
transform 1 0 19228 0 -1 44064
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__C
timestamp 1606120353
transform 1 0 19044 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__D
timestamp 1606120353
transform 1 0 18676 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__D
timestamp 1606120353
transform 1 0 17480 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_76_189
timestamp 1606120353
transform 1 0 18492 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_76_193
timestamp 1606120353
transform 1 0 18860 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0858_
timestamp 1606120353
transform 1 0 21068 0 -1 44064
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_627
timestamp 1606120353
transform 1 0 20792 0 -1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__B1
timestamp 1606120353
transform 1 0 20516 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_76_206
timestamp 1606120353
transform 1 0 20056 0 -1 44064
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_76_210
timestamp 1606120353
transform 1 0 20424 0 -1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_76_213
timestamp 1606120353
transform 1 0 20700 0 -1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_76_215
timestamp 1606120353
transform 1 0 20884 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_76_220
timestamp 1606120353
transform 1 0 21344 0 -1 44064
box 0 -48 368 592
use sky130_fd_sc_hd__a21o_4  _0896_
timestamp 1606120353
transform 1 0 22080 0 -1 44064
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__B1
timestamp 1606120353
transform 1 0 21712 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__A1
timestamp 1606120353
transform 1 0 23368 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_76_226
timestamp 1606120353
transform 1 0 21896 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_76_240
timestamp 1606120353
transform 1 0 23184 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1162_
timestamp 1606120353
transform 1 0 23920 0 -1 44064
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__B1_N
timestamp 1606120353
transform 1 0 23736 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_76_244
timestamp 1606120353
transform 1 0 23552 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0895_
timestamp 1606120353
transform 1 0 26496 0 -1 44064
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_628
timestamp 1606120353
transform 1 0 26404 0 -1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0884__A
timestamp 1606120353
transform 1 0 25852 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__C
timestamp 1606120353
transform 1 0 26220 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_76_267
timestamp 1606120353
transform 1 0 25668 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_76_271
timestamp 1606120353
transform 1 0 26036 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_76_285
timestamp 1606120353
transform 1 0 27324 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1606120353
transform -1 0 28888 0 -1 44064
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__A
timestamp 1606120353
transform 1 0 27508 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_76_289
timestamp 1606120353
transform 1 0 27692 0 -1 44064
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_76_297
timestamp 1606120353
transform 1 0 28428 0 -1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1174_
timestamp 1606120353
transform 1 0 1380 0 1 44064
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1606120353
transform 1 0 1104 0 1 44064
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_77_22
timestamp 1606120353
transform 1 0 3128 0 1 44064
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_77_34
timestamp 1606120353
transform 1 0 4232 0 1 44064
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_629
timestamp 1606120353
transform 1 0 6716 0 1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_77_46
timestamp 1606120353
transform 1 0 5336 0 1 44064
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_77_58
timestamp 1606120353
transform 1 0 6440 0 1 44064
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_77_62
timestamp 1606120353
transform 1 0 6808 0 1 44064
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_77_74
timestamp 1606120353
transform 1 0 7912 0 1 44064
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_77_86
timestamp 1606120353
transform 1 0 9016 0 1 44064
box 0 -48 1104 592
use sky130_fd_sc_hd__inv_8  _0651_
timestamp 1606120353
transform 1 0 10304 0 1 44064
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0651__A
timestamp 1606120353
transform 1 0 10120 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_77_109
timestamp 1606120353
transform 1 0 11132 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0492_
timestamp 1606120353
transform 1 0 12420 0 1 44064
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_630
timestamp 1606120353
transform 1 0 12328 0 1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0492__B
timestamp 1606120353
transform 1 0 12144 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0549__A
timestamp 1606120353
transform 1 0 11316 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0492__D
timestamp 1606120353
transform 1 0 11776 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_77_113
timestamp 1606120353
transform 1 0 11500 0 1 44064
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_77_118
timestamp 1606120353
transform 1 0 11960 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_77_132
timestamp 1606120353
transform 1 0 13248 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0548_
timestamp 1606120353
transform 1 0 13984 0 1 44064
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0548__A
timestamp 1606120353
transform 1 0 14444 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0498__A
timestamp 1606120353
transform 1 0 13432 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0492__A
timestamp 1606120353
transform 1 0 13800 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_77_136
timestamp 1606120353
transform 1 0 13616 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_77_143
timestamp 1606120353
transform 1 0 14260 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_77_147
timestamp 1606120353
transform 1 0 14628 0 1 44064
box 0 -48 1104 592
use sky130_fd_sc_hd__buf_1  _0823_
timestamp 1606120353
transform 1 0 15916 0 1 44064
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0885_
timestamp 1606120353
transform 1 0 16928 0 1 44064
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__A
timestamp 1606120353
transform 1 0 16652 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__A
timestamp 1606120353
transform 1 0 15732 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_77_164
timestamp 1606120353
transform 1 0 16192 0 1 44064
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_77_168
timestamp 1606120353
transform 1 0 16560 0 1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_77_171
timestamp 1606120353
transform 1 0 16836 0 1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_77_175
timestamp 1606120353
transform 1 0 17204 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0836_
timestamp 1606120353
transform 1 0 18584 0 1 44064
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_631
timestamp 1606120353
transform 1 0 17940 0 1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__A
timestamp 1606120353
transform 1 0 18400 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__A
timestamp 1606120353
transform 1 0 17388 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__C
timestamp 1606120353
transform 1 0 17756 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_77_179
timestamp 1606120353
transform 1 0 17572 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_77_184
timestamp 1606120353
transform 1 0 18032 0 1 44064
box 0 -48 368 592
use sky130_fd_sc_hd__and4_4  _0912_
timestamp 1606120353
transform 1 0 20148 0 1 44064
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__B
timestamp 1606120353
transform 1 0 19596 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__A
timestamp 1606120353
transform 1 0 19964 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__B1
timestamp 1606120353
transform 1 0 21160 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_77_199
timestamp 1606120353
transform 1 0 19412 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_77_203
timestamp 1606120353
transform 1 0 19780 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_77_216
timestamp 1606120353
transform 1 0 20976 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_77_220
timestamp 1606120353
transform 1 0 21344 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0865_
timestamp 1606120353
transform 1 0 21712 0 1 44064
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__A
timestamp 1606120353
transform 1 0 23368 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__A2
timestamp 1606120353
transform 1 0 21528 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__C1
timestamp 1606120353
transform 1 0 23000 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_77_236
timestamp 1606120353
transform 1 0 22816 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_77_240
timestamp 1606120353
transform 1 0 23184 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0898_
timestamp 1606120353
transform 1 0 23828 0 1 44064
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_632
timestamp 1606120353
transform 1 0 23552 0 1 44064
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__A2
timestamp 1606120353
transform 1 0 25208 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_77_245
timestamp 1606120353
transform 1 0 23644 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_77_260
timestamp 1606120353
transform 1 0 25024 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_77_264
timestamp 1606120353
transform 1 0 25392 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1228_
timestamp 1606120353
transform 1 0 26128 0 1 44064
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__D
timestamp 1606120353
transform 1 0 25944 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__A
timestamp 1606120353
transform 1 0 25576 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_77_268
timestamp 1606120353
transform 1 0 25760 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1606120353
transform -1 0 28888 0 1 44064
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__B
timestamp 1606120353
transform 1 0 28060 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_77_291
timestamp 1606120353
transform 1 0 27876 0 1 44064
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_77_295
timestamp 1606120353
transform 1 0 28244 0 1 44064
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1606120353
transform 1 0 1104 0 -1 45152
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__D
timestamp 1606120353
transform 1 0 1564 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__D
timestamp 1606120353
transform 1 0 1932 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__CLK
timestamp 1606120353
transform 1 0 2300 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_3
timestamp 1606120353
transform 1 0 1380 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_7
timestamp 1606120353
transform 1 0 1748 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_11
timestamp 1606120353
transform 1 0 2116 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_78_15
timestamp 1606120353
transform 1 0 2484 0 -1 45152
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_633
timestamp 1606120353
transform 1 0 3956 0 -1 45152
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_78_27
timestamp 1606120353
transform 1 0 3588 0 -1 45152
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_78_32
timestamp 1606120353
transform 1 0 4048 0 -1 45152
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_78_44
timestamp 1606120353
transform 1 0 5152 0 -1 45152
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_78_56
timestamp 1606120353
transform 1 0 6256 0 -1 45152
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_78_68
timestamp 1606120353
transform 1 0 7360 0 -1 45152
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_78_80
timestamp 1606120353
transform 1 0 8464 0 -1 45152
box 0 -48 1104 592
use sky130_fd_sc_hd__inv_8  _0549_
timestamp 1606120353
transform 1 0 11132 0 -1 45152
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_634
timestamp 1606120353
transform 1 0 9568 0 -1 45152
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_78_93
timestamp 1606120353
transform 1 0 9660 0 -1 45152
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_78_105
timestamp 1606120353
transform 1 0 10764 0 -1 45152
box 0 -48 368 592
use sky130_fd_sc_hd__inv_8  _0498_
timestamp 1606120353
transform 1 0 12880 0 -1 45152
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0547__B
timestamp 1606120353
transform 1 0 12420 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_78_118
timestamp 1606120353
transform 1 0 11960 0 -1 45152
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_78_122
timestamp 1606120353
transform 1 0 12328 0 -1 45152
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_78_125
timestamp 1606120353
transform 1 0 12604 0 -1 45152
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_635
timestamp 1606120353
transform 1 0 15180 0 -1 45152
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__B
timestamp 1606120353
transform 1 0 14444 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_78_137
timestamp 1606120353
transform 1 0 13708 0 -1 45152
box 0 -48 736 592
use sky130_fd_sc_hd__decap_6  FILLER_78_147
timestamp 1606120353
transform 1 0 14628 0 -1 45152
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_78_154
timestamp 1606120353
transform 1 0 15272 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0833_
timestamp 1606120353
transform 1 0 16652 0 -1 45152
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__A
timestamp 1606120353
transform 1 0 17204 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__B1
timestamp 1606120353
transform 1 0 15456 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__B1
timestamp 1606120353
transform 1 0 16008 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__B
timestamp 1606120353
transform 1 0 16468 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_78_158
timestamp 1606120353
transform 1 0 15640 0 -1 45152
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_78_164
timestamp 1606120353
transform 1 0 16192 0 -1 45152
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_78_172
timestamp 1606120353
transform 1 0 16928 0 -1 45152
box 0 -48 276 592
use sky130_fd_sc_hd__or3_4  _0841_
timestamp 1606120353
transform 1 0 17664 0 -1 45152
box 0 -48 828 592
use sky130_fd_sc_hd__or4_4  _0943_
timestamp 1606120353
transform 1 0 19228 0 -1 45152
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__C
timestamp 1606120353
transform 1 0 19044 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__B
timestamp 1606120353
transform 1 0 18676 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_78_177
timestamp 1606120353
transform 1 0 17388 0 -1 45152
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_78_189
timestamp 1606120353
transform 1 0 18492 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_193
timestamp 1606120353
transform 1 0 18860 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_636
timestamp 1606120353
transform 1 0 20792 0 -1 45152
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__C
timestamp 1606120353
transform 1 0 20240 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__A
timestamp 1606120353
transform 1 0 20608 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__B
timestamp 1606120353
transform 1 0 21068 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_206
timestamp 1606120353
transform 1 0 20056 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_210
timestamp 1606120353
transform 1 0 20424 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_215
timestamp 1606120353
transform 1 0 20884 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_78_219
timestamp 1606120353
transform 1 0 21252 0 -1 45152
box 0 -48 368 592
use sky130_fd_sc_hd__a211o_4  _0853_
timestamp 1606120353
transform 1 0 21804 0 -1 45152
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__A2
timestamp 1606120353
transform 1 0 21620 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__B1
timestamp 1606120353
transform 1 0 23276 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_239
timestamp 1606120353
transform 1 0 23092 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0875_
timestamp 1606120353
transform 1 0 23828 0 -1 45152
box 0 -48 828 592
use sky130_fd_sc_hd__buf_1  _0884_
timestamp 1606120353
transform 1 0 25392 0 -1 45152
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__B
timestamp 1606120353
transform 1 0 24840 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__B1_N
timestamp 1606120353
transform 1 0 23644 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__A1
timestamp 1606120353
transform 1 0 25208 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_243
timestamp 1606120353
transform 1 0 23460 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_256
timestamp 1606120353
transform 1 0 24656 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_260
timestamp 1606120353
transform 1 0 25024 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0887_
timestamp 1606120353
transform 1 0 26496 0 -1 45152
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_637
timestamp 1606120353
transform 1 0 26404 0 -1 45152
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__C
timestamp 1606120353
transform 1 0 25852 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__A1
timestamp 1606120353
transform 1 0 26220 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_267
timestamp 1606120353
transform 1 0 25668 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_271
timestamp 1606120353
transform 1 0 26036 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_78_285
timestamp 1606120353
transform 1 0 27324 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1606120353
transform -1 0 28888 0 -1 45152
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__CLK
timestamp 1606120353
transform 1 0 27508 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_78_289
timestamp 1606120353
transform 1 0 27692 0 -1 45152
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_78_297
timestamp 1606120353
transform 1 0 28428 0 -1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1192_
timestamp 1606120353
transform 1 0 1380 0 1 45152
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1606120353
transform 1 0 1104 0 1 45152
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1606120353
transform 1 0 1104 0 -1 46240
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__CLK
timestamp 1606120353
transform 1 0 1564 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_79_22
timestamp 1606120353
transform 1 0 3128 0 1 45152
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_80_3
timestamp 1606120353
transform 1 0 1380 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_80_7
timestamp 1606120353
transform 1 0 1748 0 -1 46240
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_80_19
timestamp 1606120353
transform 1 0 2852 0 -1 46240
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_642
timestamp 1606120353
transform 1 0 3956 0 -1 46240
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_79_34
timestamp 1606120353
transform 1 0 4232 0 1 45152
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_80_32
timestamp 1606120353
transform 1 0 4048 0 -1 46240
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_80_44
timestamp 1606120353
transform 1 0 5152 0 -1 46240
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_638
timestamp 1606120353
transform 1 0 6716 0 1 45152
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_79_46
timestamp 1606120353
transform 1 0 5336 0 1 45152
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_79_58
timestamp 1606120353
transform 1 0 6440 0 1 45152
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_79_62
timestamp 1606120353
transform 1 0 6808 0 1 45152
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_80_56
timestamp 1606120353
transform 1 0 6256 0 -1 46240
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_79_74
timestamp 1606120353
transform 1 0 7912 0 1 45152
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_79_86
timestamp 1606120353
transform 1 0 9016 0 1 45152
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_80_68
timestamp 1606120353
transform 1 0 7360 0 -1 46240
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_80_80
timestamp 1606120353
transform 1 0 8464 0 -1 46240
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_643
timestamp 1606120353
transform 1 0 9568 0 -1 46240
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0500__A
timestamp 1606120353
transform 1 0 11132 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_79_98
timestamp 1606120353
transform 1 0 10120 0 1 45152
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_79_106
timestamp 1606120353
transform 1 0 10856 0 1 45152
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_80_93
timestamp 1606120353
transform 1 0 9660 0 -1 46240
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_80_105
timestamp 1606120353
transform 1 0 10764 0 -1 46240
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_80_119
timestamp 1606120353
transform 1 0 12052 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_79_118
timestamp 1606120353
transform 1 0 11960 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_79_114
timestamp 1606120353
transform 1 0 11592 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0547__A
timestamp 1606120353
transform 1 0 11868 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0622__A
timestamp 1606120353
transform 1 0 12236 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0622__C
timestamp 1606120353
transform 1 0 11776 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0622__B
timestamp 1606120353
transform 1 0 12144 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0500_
timestamp 1606120353
transform 1 0 11316 0 1 45152
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_639
timestamp 1606120353
transform 1 0 12328 0 1 45152
box 0 -48 92 592
use sky130_fd_sc_hd__or3_4  _0547_
timestamp 1606120353
transform 1 0 12420 0 -1 46240
box 0 -48 828 592
use sky130_fd_sc_hd__decap_12  FILLER_80_132
timestamp 1606120353
transform 1 0 13248 0 -1 46240
box 0 -48 1104 592
use sky130_fd_sc_hd__nand3_4  _0622_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/maglef
timestamp 1606120353
transform 1 0 12420 0 1 45152
box 0 -48 1288 592
use sky130_fd_sc_hd__fill_2  FILLER_79_141
timestamp 1606120353
transform 1 0 14076 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_79_137
timestamp 1606120353
transform 1 0 13708 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0547__C
timestamp 1606120353
transform 1 0 13892 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__C
timestamp 1606120353
transform 1 0 14260 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_80_147
timestamp 1606120353
transform 1 0 14628 0 -1 46240
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_80_144
timestamp 1606120353
transform 1 0 14352 0 -1 46240
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_79_154
timestamp 1606120353
transform 1 0 15272 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__A
timestamp 1606120353
transform 1 0 14444 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__A2
timestamp 1606120353
transform 1 0 14996 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_644
timestamp 1606120353
transform 1 0 15180 0 -1 46240
box 0 -48 92 592
use sky130_fd_sc_hd__and3_4  _0620_
timestamp 1606120353
transform 1 0 14444 0 1 45152
box 0 -48 828 592
use sky130_fd_sc_hd__o21ai_4  _1081_
timestamp 1606120353
transform 1 0 15272 0 -1 46240
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_4  FILLER_79_162
timestamp 1606120353
transform 1 0 16008 0 1 45152
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_79_158
timestamp 1606120353
transform 1 0 15640 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__A2
timestamp 1606120353
transform 1 0 15824 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__A1
timestamp 1606120353
transform 1 0 15456 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_80_171
timestamp 1606120353
transform 1 0 16836 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_80_167
timestamp 1606120353
transform 1 0 16468 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_79_168
timestamp 1606120353
transform 1 0 16560 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__A1
timestamp 1606120353
transform 1 0 16652 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__B
timestamp 1606120353
transform 1 0 16376 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__A
timestamp 1606120353
transform 1 0 16744 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0882_
timestamp 1606120353
transform 1 0 16928 0 1 45152
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_79_175
timestamp 1606120353
transform 1 0 17204 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__A1
timestamp 1606120353
transform 1 0 17020 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _1036_
timestamp 1606120353
transform 1 0 17204 0 -1 46240
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_80_184
timestamp 1606120353
transform 1 0 18032 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_79_179
timestamp 1606120353
transform 1 0 17572 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__C
timestamp 1606120353
transform 1 0 17388 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__B
timestamp 1606120353
transform 1 0 17756 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_640
timestamp 1606120353
transform 1 0 17940 0 1 45152
box 0 -48 92 592
use sky130_fd_sc_hd__or3_4  _0837_
timestamp 1606120353
transform 1 0 18032 0 1 45152
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  FILLER_80_192
timestamp 1606120353
transform 1 0 18768 0 -1 46240
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_80_188
timestamp 1606120353
transform 1 0 18400 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_79_193
timestamp 1606120353
transform 1 0 18860 0 1 45152
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__B
timestamp 1606120353
transform 1 0 18584 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__A
timestamp 1606120353
transform 1 0 18216 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__B
timestamp 1606120353
transform 1 0 19044 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__A
timestamp 1606120353
transform 1 0 19228 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__or3_4  _0835_
timestamp 1606120353
transform 1 0 19228 0 -1 46240
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_80_206
timestamp 1606120353
transform 1 0 20056 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_79_199
timestamp 1606120353
transform 1 0 19412 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__A
timestamp 1606120353
transform 1 0 20240 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_80_210
timestamp 1606120353
transform 1 0 20424 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_79_218
timestamp 1606120353
transform 1 0 21160 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__B1
timestamp 1606120353
transform 1 0 20608 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__A
timestamp 1606120353
transform 1 0 21344 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_645
timestamp 1606120353
transform 1 0 20792 0 -1 46240
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _0834_
timestamp 1606120353
transform 1 0 20884 0 -1 46240
box 0 -48 828 592
use sky130_fd_sc_hd__nand4_4  _1042_
timestamp 1606120353
transform 1 0 19596 0 1 45152
box 0 -48 1564 592
use sky130_fd_sc_hd__decap_3  FILLER_80_229
timestamp 1606120353
transform 1 0 22172 0 -1 46240
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_80_224
timestamp 1606120353
transform 1 0 21712 0 -1 46240
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_79_222
timestamp 1606120353
transform 1 0 21528 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__A
timestamp 1606120353
transform 1 0 21988 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__A
timestamp 1606120353
transform 1 0 21712 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _0897_
timestamp 1606120353
transform 1 0 21896 0 1 45152
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  FILLER_79_239
timestamp 1606120353
transform 1 0 23092 0 1 45152
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_79_235
timestamp 1606120353
transform 1 0 22724 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__A2
timestamp 1606120353
transform 1 0 22908 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__A2
timestamp 1606120353
transform 1 0 23368 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0892_
timestamp 1606120353
transform 1 0 22448 0 -1 46240
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1606120353
transform 1 0 24196 0 -1 46240
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_80_248
timestamp 1606120353
transform 1 0 23920 0 -1 46240
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_80_244
timestamp 1606120353
transform 1 0 23552 0 -1 46240
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__A1
timestamp 1606120353
transform 1 0 24012 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_641
timestamp 1606120353
transform 1 0 23552 0 1 45152
box 0 -48 92 592
use sky130_fd_sc_hd__nor2_4  _0893_
timestamp 1606120353
transform 1 0 24288 0 -1 46240
box 0 -48 828 592
use sky130_fd_sc_hd__decap_4  FILLER_80_261
timestamp 1606120353
transform 1 0 25116 0 -1 46240
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_79_262
timestamp 1606120353
transform 1 0 25208 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_79_258
timestamp 1606120353
transform 1 0 24840 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__A
timestamp 1606120353
transform 1 0 25392 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__A
timestamp 1606120353
transform 1 0 25024 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0894_
timestamp 1606120353
transform 1 0 23644 0 1 45152
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_3  FILLER_80_272
timestamp 1606120353
transform 1 0 26128 0 -1 46240
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_80_268
timestamp 1606120353
transform 1 0 25760 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_80_265
timestamp 1606120353
transform 1 0 25484 0 -1 46240
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_79_275
timestamp 1606120353
transform 1 0 26404 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__A1
timestamp 1606120353
transform 1 0 25944 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__B
timestamp 1606120353
transform 1 0 25576 0 -1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_646
timestamp 1606120353
transform 1 0 26404 0 -1 46240
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _0891_
timestamp 1606120353
transform 1 0 25576 0 1 45152
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_79_283
timestamp 1606120353
transform 1 0 27140 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_79_279
timestamp 1606120353
transform 1 0 26772 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__D
timestamp 1606120353
transform 1 0 27324 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__A1
timestamp 1606120353
transform 1 0 26956 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__D
timestamp 1606120353
transform 1 0 26588 0 1 45152
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_80_276
timestamp 1606120353
transform 1 0 26496 0 -1 46240
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1606120353
transform -1 0 28888 0 1 45152
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1606120353
transform -1 0 28888 0 -1 46240
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_79_287
timestamp 1606120353
transform 1 0 27508 0 1 45152
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_80_288
timestamp 1606120353
transform 1 0 27600 0 -1 46240
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_80_296
timestamp 1606120353
transform 1 0 28336 0 -1 46240
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1606120353
transform 1 0 1104 0 1 46240
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_81_3
timestamp 1606120353
transform 1 0 1380 0 1 46240
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_81_15
timestamp 1606120353
transform 1 0 2484 0 1 46240
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_81_27
timestamp 1606120353
transform 1 0 3588 0 1 46240
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_81_39
timestamp 1606120353
transform 1 0 4692 0 1 46240
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_647
timestamp 1606120353
transform 1 0 6716 0 1 46240
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_81_51
timestamp 1606120353
transform 1 0 5796 0 1 46240
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_81_59
timestamp 1606120353
transform 1 0 6532 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_81_62
timestamp 1606120353
transform 1 0 6808 0 1 46240
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_81_74
timestamp 1606120353
transform 1 0 7912 0 1 46240
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_81_86
timestamp 1606120353
transform 1 0 9016 0 1 46240
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_81_98
timestamp 1606120353
transform 1 0 10120 0 1 46240
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_81_110
timestamp 1606120353
transform 1 0 11224 0 1 46240
box 0 -48 552 592
use sky130_fd_sc_hd__or3_4  _0499_
timestamp 1606120353
transform 1 0 12420 0 1 46240
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_648
timestamp 1606120353
transform 1 0 12328 0 1 46240
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0499__C
timestamp 1606120353
transform 1 0 12144 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0499__A
timestamp 1606120353
transform 1 0 11776 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_118
timestamp 1606120353
transform 1 0 11960 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_132
timestamp 1606120353
transform 1 0 13248 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_81_136
timestamp 1606120353
transform 1 0 13616 0 1 46240
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0488__A
timestamp 1606120353
transform 1 0 13432 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_81_140
timestamp 1606120353
transform 1 0 13984 0 1 46240
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_81_143
timestamp 1606120353
transform 1 0 14260 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__A
timestamp 1606120353
transform 1 0 14076 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_147
timestamp 1606120353
transform 1 0 14628 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__A2
timestamp 1606120353
transform 1 0 14444 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__B1
timestamp 1606120353
transform 1 0 14812 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0842_
timestamp 1606120353
transform 1 0 14996 0 1 46240
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_81_154
timestamp 1606120353
transform 1 0 15272 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1080_
timestamp 1606120353
transform 1 0 16008 0 1 46240
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__A
timestamp 1606120353
transform 1 0 15456 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__A1
timestamp 1606120353
transform 1 0 15824 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_158
timestamp 1606120353
transform 1 0 15640 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_175
timestamp 1606120353
transform 1 0 17204 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__and3_4  _1065_
timestamp 1606120353
transform 1 0 18032 0 1 46240
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_649
timestamp 1606120353
transform 1 0 17940 0 1 46240
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__A1
timestamp 1606120353
transform 1 0 19136 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__A2
timestamp 1606120353
transform 1 0 17756 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__A
timestamp 1606120353
transform 1 0 17388 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_179
timestamp 1606120353
transform 1 0 17572 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_81_193
timestamp 1606120353
transform 1 0 18860 0 1 46240
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_81_198
timestamp 1606120353
transform 1 0 19320 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0958_
timestamp 1606120353
transform 1 0 19688 0 1 46240
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__B1
timestamp 1606120353
transform 1 0 19504 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A
timestamp 1606120353
transform 1 0 20976 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__B
timestamp 1606120353
transform 1 0 21344 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_214
timestamp 1606120353
transform 1 0 20792 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_218
timestamp 1606120353
transform 1 0 21160 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0899_
timestamp 1606120353
transform 1 0 21988 0 1 46240
box 0 -48 828 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_clk
timestamp 1606120353
transform 1 0 21528 0 1 46240
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__C
timestamp 1606120353
transform 1 0 23000 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__A2
timestamp 1606120353
transform 1 0 23368 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_225
timestamp 1606120353
transform 1 0 21804 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_236
timestamp 1606120353
transform 1 0 22816 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_240
timestamp 1606120353
transform 1 0 23184 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _0874_
timestamp 1606120353
transform 1 0 24012 0 1 46240
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_650
timestamp 1606120353
transform 1 0 23552 0 1 46240
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__A2
timestamp 1606120353
transform 1 0 23828 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__B1_N
timestamp 1606120353
transform 1 0 25392 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_245
timestamp 1606120353
transform 1 0 23644 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_262
timestamp 1606120353
transform 1 0 25208 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0852_
timestamp 1606120353
transform 1 0 25944 0 1 46240
box 0 -48 644 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__A
timestamp 1606120353
transform 1 0 26772 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__B
timestamp 1606120353
transform 1 0 25760 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_clk_A
timestamp 1606120353
transform 1 0 27140 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_266
timestamp 1606120353
transform 1 0 25576 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_277
timestamp 1606120353
transform 1 0 26588 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_81_281
timestamp 1606120353
transform 1 0 26956 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_81_285
timestamp 1606120353
transform 1 0 27324 0 1 46240
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1606120353
transform -1 0 28888 0 1 46240
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_81_297
timestamp 1606120353
transform 1 0 28428 0 1 46240
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1606120353
transform 1 0 1104 0 -1 47328
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_82_3
timestamp 1606120353
transform 1 0 1380 0 -1 47328
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_82_15
timestamp 1606120353
transform 1 0 2484 0 -1 47328
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_651
timestamp 1606120353
transform 1 0 3956 0 -1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_82_27
timestamp 1606120353
transform 1 0 3588 0 -1 47328
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_82_32
timestamp 1606120353
transform 1 0 4048 0 -1 47328
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_82_44
timestamp 1606120353
transform 1 0 5152 0 -1 47328
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_82_56
timestamp 1606120353
transform 1 0 6256 0 -1 47328
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__CLK
timestamp 1606120353
transform 1 0 8188 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_82_68
timestamp 1606120353
transform 1 0 7360 0 -1 47328
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_82_76
timestamp 1606120353
transform 1 0 8096 0 -1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_82_79
timestamp 1606120353
transform 1 0 8372 0 -1 47328
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_652
timestamp 1606120353
transform 1 0 9568 0 -1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_82_91
timestamp 1606120353
transform 1 0 9476 0 -1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_82_93
timestamp 1606120353
transform 1 0 9660 0 -1 47328
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_82_105
timestamp 1606120353
transform 1 0 10764 0 -1 47328
box 0 -48 1104 592
use sky130_fd_sc_hd__inv_8  _0488_
timestamp 1606120353
transform 1 0 12604 0 -1 47328
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0499__B
timestamp 1606120353
transform 1 0 12420 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_82_117
timestamp 1606120353
transform 1 0 11868 0 -1 47328
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_82_138
timestamp 1606120353
transform 1 0 13800 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_82_134
timestamp 1606120353
transform 1 0 13432 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__B1
timestamp 1606120353
transform 1 0 13616 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__A
timestamp 1606120353
transform 1 0 13984 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1070_
timestamp 1606120353
transform 1 0 14168 0 -1 47328
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_82_149
timestamp 1606120353
transform 1 0 14812 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_82_145
timestamp 1606120353
transform 1 0 14444 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__C
timestamp 1606120353
transform 1 0 14628 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__B1
timestamp 1606120353
transform 1 0 14996 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_653
timestamp 1606120353
transform 1 0 15180 0 -1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__o21ai_4  _1041_
timestamp 1606120353
transform 1 0 15272 0 -1 47328
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__A
timestamp 1606120353
transform 1 0 17204 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__B1
timestamp 1606120353
transform 1 0 16836 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_82_167
timestamp 1606120353
transform 1 0 16468 0 -1 47328
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_82_173
timestamp 1606120353
transform 1 0 17020 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0986_
timestamp 1606120353
transform 1 0 17388 0 -1 47328
box 0 -48 276 592
use sky130_fd_sc_hd__o21ai_4  _1047_
timestamp 1606120353
transform 1 0 18400 0 -1 47328
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__C
timestamp 1606120353
transform 1 0 18032 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_82_180
timestamp 1606120353
transform 1 0 17664 0 -1 47328
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_82_186
timestamp 1606120353
transform 1 0 18216 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0878_
timestamp 1606120353
transform 1 0 20884 0 -1 47328
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_654
timestamp 1606120353
transform 1 0 20792 0 -1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__A2
timestamp 1606120353
transform 1 0 19780 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__B
timestamp 1606120353
transform 1 0 20608 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__B1
timestamp 1606120353
transform 1 0 20148 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_82_201
timestamp 1606120353
transform 1 0 19596 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_82_205
timestamp 1606120353
transform 1 0 19964 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_82_209
timestamp 1606120353
transform 1 0 20332 0 -1 47328
box 0 -48 276 592
use sky130_fd_sc_hd__a21o_4  _0900_
timestamp 1606120353
transform 1 0 22448 0 -1 47328
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__A2
timestamp 1606120353
transform 1 0 22264 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__B
timestamp 1606120353
transform 1 0 21896 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_82_224
timestamp 1606120353
transform 1 0 21712 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_82_228
timestamp 1606120353
transform 1 0 22080 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0930_
timestamp 1606120353
transform 1 0 24380 0 -1 47328
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__B1
timestamp 1606120353
transform 1 0 23736 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__B1
timestamp 1606120353
transform 1 0 24104 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_82_244
timestamp 1606120353
transform 1 0 23552 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_82_248
timestamp 1606120353
transform 1 0 23920 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_82_252
timestamp 1606120353
transform 1 0 24288 0 -1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0839_
timestamp 1606120353
transform 1 0 26496 0 -1 47328
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_655
timestamp 1606120353
transform 1 0 26404 0 -1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__A2
timestamp 1606120353
transform 1 0 25760 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__A
timestamp 1606120353
transform 1 0 26128 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_82_266
timestamp 1606120353
transform 1 0 25576 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_82_270
timestamp 1606120353
transform 1 0 25944 0 -1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_82_274
timestamp 1606120353
transform 1 0 26312 0 -1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_82_279
timestamp 1606120353
transform 1 0 26772 0 -1 47328
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1606120353
transform -1 0 28888 0 -1 47328
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_82_291
timestamp 1606120353
transform 1 0 27876 0 -1 47328
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1606120353
transform 1 0 1104 0 1 47328
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_83_3
timestamp 1606120353
transform 1 0 1380 0 1 47328
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_83_15
timestamp 1606120353
transform 1 0 2484 0 1 47328
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_83_27
timestamp 1606120353
transform 1 0 3588 0 1 47328
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_83_39
timestamp 1606120353
transform 1 0 4692 0 1 47328
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_656
timestamp 1606120353
transform 1 0 6716 0 1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_83_51
timestamp 1606120353
transform 1 0 5796 0 1 47328
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_83_59
timestamp 1606120353
transform 1 0 6532 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_83_62
timestamp 1606120353
transform 1 0 6808 0 1 47328
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1127_
timestamp 1606120353
transform 1 0 8188 0 1 47328
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__D
timestamp 1606120353
transform 1 0 8004 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_83_74
timestamp 1606120353
transform 1 0 7912 0 1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_83_96
timestamp 1606120353
transform 1 0 9936 0 1 47328
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_83_108
timestamp 1606120353
transform 1 0 11040 0 1 47328
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_657
timestamp 1606120353
transform 1 0 12328 0 1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__B
timestamp 1606120353
transform 1 0 12972 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__B1
timestamp 1606120353
transform 1 0 12604 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_clk_A
timestamp 1606120353
transform 1 0 12144 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_123
timestamp 1606120353
transform 1 0 12420 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_127
timestamp 1606120353
transform 1 0 12788 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_131
timestamp 1606120353
transform 1 0 13156 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_135
timestamp 1606120353
transform 1 0 13524 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__A1
timestamp 1606120353
transform 1 0 13340 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_83_139
timestamp 1606120353
transform 1 0 13892 0 1 47328
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__A2
timestamp 1606120353
transform 1 0 13708 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__A2
timestamp 1606120353
transform 1 0 14260 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_148
timestamp 1606120353
transform 1 0 14720 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0984_
timestamp 1606120353
transform 1 0 14444 0 1 47328
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_83_152
timestamp 1606120353
transform 1 0 15088 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__A
timestamp 1606120353
transform 1 0 14904 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A1
timestamp 1606120353
transform 1 0 15272 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1038_
timestamp 1606120353
transform 1 0 15456 0 1 47328
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__A1
timestamp 1606120353
transform 1 0 16836 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A2
timestamp 1606120353
transform 1 0 17204 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_169
timestamp 1606120353
transform 1 0 16652 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_173
timestamp 1606120353
transform 1 0 17020 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _0959_
timestamp 1606120353
transform 1 0 18400 0 1 47328
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_658
timestamp 1606120353
transform 1 0 17940 0 1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_clk
timestamp 1606120353
transform 1 0 17388 0 1 47328
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__A2
timestamp 1606120353
transform 1 0 18216 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_83_180
timestamp 1606120353
transform 1 0 17664 0 1 47328
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_83_184
timestamp 1606120353
transform 1 0 18032 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_201
timestamp 1606120353
transform 1 0 19596 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__A
timestamp 1606120353
transform 1 0 19780 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_205
timestamp 1606120353
transform 1 0 19964 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__B
timestamp 1606120353
transform 1 0 20148 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_83_209
timestamp 1606120353
transform 1 0 20332 0 1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0883_
timestamp 1606120353
transform 1 0 20424 0 1 47328
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_83_213
timestamp 1606120353
transform 1 0 20700 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0883__A
timestamp 1606120353
transform 1 0 20884 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_217
timestamp 1606120353
transform 1 0 21068 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__A
timestamp 1606120353
transform 1 0 21252 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _0918_
timestamp 1606120353
transform 1 0 21436 0 1 47328
box 0 -48 828 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_clk
timestamp 1606120353
transform 1 0 23276 0 1 47328
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A2
timestamp 1606120353
transform 1 0 23092 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A1
timestamp 1606120353
transform 1 0 22724 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_83_230
timestamp 1606120353
transform 1 0 22264 0 1 47328
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_83_234
timestamp 1606120353
transform 1 0 22632 0 1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_83_237
timestamp 1606120353
transform 1 0 22908 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0873_
timestamp 1606120353
transform 1 0 23644 0 1 47328
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_659
timestamp 1606120353
transform 1 0 23552 0 1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__A
timestamp 1606120353
transform 1 0 24932 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__A1
timestamp 1606120353
transform 1 0 25300 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_257
timestamp 1606120353
transform 1 0 24748 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_83_261
timestamp 1606120353
transform 1 0 25116 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1212_
timestamp 1606120353
transform 1 0 26128 0 1 47328
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__D
timestamp 1606120353
transform 1 0 25944 0 1 47328
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_83_265
timestamp 1606120353
transform 1 0 25484 0 1 47328
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_83_269
timestamp 1606120353
transform 1 0 25852 0 1 47328
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1606120353
transform -1 0 28888 0 1 47328
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_83_291
timestamp 1606120353
transform 1 0 27876 0 1 47328
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1606120353
transform 1 0 1104 0 -1 48416
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_84_3
timestamp 1606120353
transform 1 0 1380 0 -1 48416
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_84_15
timestamp 1606120353
transform 1 0 2484 0 -1 48416
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_660
timestamp 1606120353
transform 1 0 3956 0 -1 48416
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_84_27
timestamp 1606120353
transform 1 0 3588 0 -1 48416
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_84_32
timestamp 1606120353
transform 1 0 4048 0 -1 48416
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_84_44
timestamp 1606120353
transform 1 0 5152 0 -1 48416
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_84_56
timestamp 1606120353
transform 1 0 6256 0 -1 48416
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_84_68
timestamp 1606120353
transform 1 0 7360 0 -1 48416
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_84_80
timestamp 1606120353
transform 1 0 8464 0 -1 48416
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_661
timestamp 1606120353
transform 1 0 9568 0 -1 48416
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_84_93
timestamp 1606120353
transform 1 0 9660 0 -1 48416
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_84_105
timestamp 1606120353
transform 1 0 10764 0 -1 48416
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__A
timestamp 1606120353
transform 1 0 13156 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__A
timestamp 1606120353
transform 1 0 12788 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__CLK
timestamp 1606120353
transform 1 0 12420 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_84_117
timestamp 1606120353
transform 1 0 11868 0 -1 48416
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_84_125
timestamp 1606120353
transform 1 0 12604 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_129
timestamp 1606120353
transform 1 0 12972 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _1076_
timestamp 1606120353
transform 1 0 13340 0 -1 48416
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_662
timestamp 1606120353
transform 1 0 15180 0 -1 48416
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A2
timestamp 1606120353
transform 1 0 14628 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__A2
timestamp 1606120353
transform 1 0 14996 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_145
timestamp 1606120353
transform 1 0 14444 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_149
timestamp 1606120353
transform 1 0 14812 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_84_154
timestamp 1606120353
transform 1 0 15272 0 -1 48416
box 0 -48 276 592
use sky130_fd_sc_hd__o21a_4  _1079_
timestamp 1606120353
transform 1 0 15548 0 -1 48416
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__B
timestamp 1606120353
transform 1 0 17204 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__C
timestamp 1606120353
transform 1 0 16836 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_169
timestamp 1606120353
transform 1 0 16652 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_173
timestamp 1606120353
transform 1 0 17020 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__nor3_4  _1075_
timestamp 1606120353
transform 1 0 17388 0 -1 48416
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__A1
timestamp 1606120353
transform 1 0 18768 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__B1
timestamp 1606120353
transform 1 0 19136 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_190
timestamp 1606120353
transform 1 0 18584 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_194
timestamp 1606120353
transform 1 0 18952 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_84_198
timestamp 1606120353
transform 1 0 19320 0 -1 48416
box 0 -48 92 592
use sky130_fd_sc_hd__and2_4  _0838_
timestamp 1606120353
transform 1 0 19412 0 -1 48416
box 0 -48 644 592
use sky130_fd_sc_hd__and4_4  _1074_
timestamp 1606120353
transform 1 0 20884 0 -1 48416
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_663
timestamp 1606120353
transform 1 0 20792 0 -1 48416
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__B
timestamp 1606120353
transform 1 0 20608 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__C
timestamp 1606120353
transform 1 0 20240 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_206
timestamp 1606120353
transform 1 0 20056 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_210
timestamp 1606120353
transform 1 0 20424 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0902_
timestamp 1606120353
transform 1 0 22724 0 -1 48416
box 0 -48 1196 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_clk
timestamp 1606120353
transform 1 0 22448 0 -1 48416
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A2
timestamp 1606120353
transform 1 0 21896 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__B1_N
timestamp 1606120353
transform 1 0 22264 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_224
timestamp 1606120353
transform 1 0 21712 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_228
timestamp 1606120353
transform 1 0 22080 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0890_
timestamp 1606120353
transform 1 0 24656 0 -1 48416
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__A1
timestamp 1606120353
transform 1 0 24104 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__D
timestamp 1606120353
transform 1 0 24472 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_clk_A
timestamp 1606120353
transform 1 0 25116 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_248
timestamp 1606120353
transform 1 0 23920 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_252
timestamp 1606120353
transform 1 0 24288 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_84_259
timestamp 1606120353
transform 1 0 24932 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_84_263
timestamp 1606120353
transform 1 0 25300 0 -1 48416
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_664
timestamp 1606120353
transform 1 0 26404 0 -1 48416
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__CLK
timestamp 1606120353
transform 1 0 26128 0 -1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_84_271
timestamp 1606120353
transform 1 0 26036 0 -1 48416
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_84_274
timestamp 1606120353
transform 1 0 26312 0 -1 48416
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_84_276
timestamp 1606120353
transform 1 0 26496 0 -1 48416
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1606120353
transform -1 0 28888 0 -1 48416
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_84_288
timestamp 1606120353
transform 1 0 27600 0 -1 48416
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_84_296
timestamp 1606120353
transform 1 0 28336 0 -1 48416
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1606120353
transform 1 0 1104 0 1 48416
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1606120353
transform 1 0 1104 0 -1 49504
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_85_3
timestamp 1606120353
transform 1 0 1380 0 1 48416
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_85_15
timestamp 1606120353
transform 1 0 2484 0 1 48416
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_86_3
timestamp 1606120353
transform 1 0 1380 0 -1 49504
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_86_15
timestamp 1606120353
transform 1 0 2484 0 -1 49504
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_669
timestamp 1606120353
transform 1 0 3956 0 -1 49504
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_85_27
timestamp 1606120353
transform 1 0 3588 0 1 48416
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_85_39
timestamp 1606120353
transform 1 0 4692 0 1 48416
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_86_27
timestamp 1606120353
transform 1 0 3588 0 -1 49504
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_86_32
timestamp 1606120353
transform 1 0 4048 0 -1 49504
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_86_44
timestamp 1606120353
transform 1 0 5152 0 -1 49504
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_665
timestamp 1606120353
transform 1 0 6716 0 1 48416
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_85_51
timestamp 1606120353
transform 1 0 5796 0 1 48416
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_85_59
timestamp 1606120353
transform 1 0 6532 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_85_62
timestamp 1606120353
transform 1 0 6808 0 1 48416
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_86_56
timestamp 1606120353
transform 1 0 6256 0 -1 49504
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__CLK
timestamp 1606120353
transform 1 0 7360 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_85_74
timestamp 1606120353
transform 1 0 7912 0 1 48416
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_85_86
timestamp 1606120353
transform 1 0 9016 0 1 48416
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_86_70
timestamp 1606120353
transform 1 0 7544 0 -1 49504
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_86_82
timestamp 1606120353
transform 1 0 8648 0 -1 49504
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_86_99
timestamp 1606120353
transform 1 0 10212 0 -1 49504
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_86_93
timestamp 1606120353
transform 1 0 9660 0 -1 49504
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_86_90
timestamp 1606120353
transform 1 0 9384 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_670
timestamp 1606120353
transform 1 0 9568 0 -1 49504
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_86_110
timestamp 1606120353
transform 1 0 11224 0 -1 49504
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_86_106
timestamp 1606120353
transform 1 0 10856 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_86_102
timestamp 1606120353
transform 1 0 10488 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_85_110
timestamp 1606120353
transform 1 0 11224 0 1 48416
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__CLK
timestamp 1606120353
transform 1 0 11040 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__A2
timestamp 1606120353
transform 1 0 10672 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__B1
timestamp 1606120353
transform 1 0 10304 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_85_98
timestamp 1606120353
transform 1 0 10120 0 1 48416
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_86_118
timestamp 1606120353
transform 1 0 11960 0 -1 49504
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  FILLER_85_117
timestamp 1606120353
transform 1 0 11868 0 1 48416
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_85_113
timestamp 1606120353
transform 1 0 11500 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__B
timestamp 1606120353
transform 1 0 11684 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__D
timestamp 1606120353
transform 1 0 12144 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__A
timestamp 1606120353
transform 1 0 11316 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0733_
timestamp 1606120353
transform 1 0 11316 0 -1 49504
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILLER_85_132
timestamp 1606120353
transform 1 0 13248 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_85_128
timestamp 1606120353
transform 1 0 12880 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_85_123
timestamp 1606120353
transform 1 0 12420 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__D
timestamp 1606120353
transform 1 0 12512 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__A
timestamp 1606120353
transform 1 0 13064 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_666
timestamp 1606120353
transform 1 0 12328 0 1 48416
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0732_
timestamp 1606120353
transform 1 0 12604 0 1 48416
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1147_
timestamp 1606120353
transform 1 0 12696 0 -1 49504
box 0 -48 1748 592
use sky130_fd_sc_hd__fill_2  FILLER_85_143
timestamp 1606120353
transform 1 0 14260 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_85_139
timestamp 1606120353
transform 1 0 13892 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__A
timestamp 1606120353
transform 1 0 13432 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__B1
timestamp 1606120353
transform 1 0 14076 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1040_
timestamp 1606120353
transform 1 0 13616 0 1 48416
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_86_154
timestamp 1606120353
transform 1 0 15272 0 -1 49504
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_86_149
timestamp 1606120353
transform 1 0 14812 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_86_145
timestamp 1606120353
transform 1 0 14444 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__B1
timestamp 1606120353
transform 1 0 14628 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__B
timestamp 1606120353
transform 1 0 14996 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A1
timestamp 1606120353
transform 1 0 14444 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_671
timestamp 1606120353
transform 1 0 15180 0 -1 49504
box 0 -48 92 592
use sky130_fd_sc_hd__o21ai_4  _1030_
timestamp 1606120353
transform 1 0 14628 0 1 48416
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_86_162
timestamp 1606120353
transform 1 0 16008 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_86_158
timestamp 1606120353
transform 1 0 15640 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_85_164
timestamp 1606120353
transform 1 0 16192 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_85_160
timestamp 1606120353
transform 1 0 15824 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__B
timestamp 1606120353
transform 1 0 16008 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__A
timestamp 1606120353
transform 1 0 16192 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__A
timestamp 1606120353
transform 1 0 15824 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1035_
timestamp 1606120353
transform 1 0 15364 0 -1 49504
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_85_175
timestamp 1606120353
transform 1 0 17204 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_85_168
timestamp 1606120353
transform 1 0 16560 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__A
timestamp 1606120353
transform 1 0 16744 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__A
timestamp 1606120353
transform 1 0 16376 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0879_
timestamp 1606120353
transform 1 0 16928 0 1 48416
box 0 -48 276 592
use sky130_fd_sc_hd__nor3_4  _1029_
timestamp 1606120353
transform 1 0 16376 0 -1 49504
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_86_183
timestamp 1606120353
transform 1 0 17940 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_86_179
timestamp 1606120353
transform 1 0 17572 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_85_179
timestamp 1606120353
transform 1 0 17572 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__A1
timestamp 1606120353
transform 1 0 17756 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__B1
timestamp 1606120353
transform 1 0 18124 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__A1
timestamp 1606120353
transform 1 0 17756 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__A
timestamp 1606120353
transform 1 0 17388 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_667
timestamp 1606120353
transform 1 0 17940 0 1 48416
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_85_197
timestamp 1606120353
transform 1 0 19228 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__nor3_4  _1066_
timestamp 1606120353
transform 1 0 18032 0 1 48416
box 0 -48 1196 592
use sky130_fd_sc_hd__o21a_4  _1037_
timestamp 1606120353
transform 1 0 18308 0 -1 49504
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_86_207
timestamp 1606120353
transform 1 0 20148 0 -1 49504
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_86_203
timestamp 1606120353
transform 1 0 19780 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_86_199
timestamp 1606120353
transform 1 0 19412 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_85_201
timestamp 1606120353
transform 1 0 19596 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__A2
timestamp 1606120353
transform 1 0 19596 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__A2
timestamp 1606120353
transform 1 0 19412 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__C
timestamp 1606120353
transform 1 0 19964 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__D
timestamp 1606120353
transform 1 0 19780 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _1064_
timestamp 1606120353
transform 1 0 19964 0 1 48416
box 0 -48 828 592
use sky130_fd_sc_hd__fill_1  FILLER_86_211
timestamp 1606120353
transform 1 0 20516 0 -1 49504
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_85_214
timestamp 1606120353
transform 1 0 20792 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__A
timestamp 1606120353
transform 1 0 20608 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__A
timestamp 1606120353
transform 1 0 20976 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_672
timestamp 1606120353
transform 1 0 20792 0 -1 49504
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0886_
timestamp 1606120353
transform 1 0 20884 0 -1 49504
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_86_218
timestamp 1606120353
transform 1 0 21160 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_85_218
timestamp 1606120353
transform 1 0 21160 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__B
timestamp 1606120353
transform 1 0 21344 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__C
timestamp 1606120353
transform 1 0 21344 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_86_222
timestamp 1606120353
transform 1 0 21528 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_85_222
timestamp 1606120353
transform 1 0 21528 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__D
timestamp 1606120353
transform 1 0 21712 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__A
timestamp 1606120353
transform 1 0 21712 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _0901_
timestamp 1606120353
transform 1 0 21896 0 1 48416
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_86_242
timestamp 1606120353
transform 1 0 23368 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_86_238
timestamp 1606120353
transform 1 0 23000 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_85_239
timestamp 1606120353
transform 1 0 23092 0 1 48416
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_85_235
timestamp 1606120353
transform 1 0 22724 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__D
timestamp 1606120353
transform 1 0 23184 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__B1
timestamp 1606120353
transform 1 0 22908 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A
timestamp 1606120353
transform 1 0 23368 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0917_
timestamp 1606120353
transform 1 0 21896 0 -1 49504
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_86_246
timestamp 1606120353
transform 1 0 23736 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_clk_A
timestamp 1606120353
transform 1 0 23920 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A1
timestamp 1606120353
transform 1 0 23552 0 -1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_668
timestamp 1606120353
transform 1 0 23552 0 1 48416
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _0872_
timestamp 1606120353
transform 1 0 24104 0 -1 49504
box 0 -48 828 592
use sky130_fd_sc_hd__inv_8  _0854_
timestamp 1606120353
transform 1 0 23644 0 1 48416
box 0 -48 828 592
use sky130_fd_sc_hd__decap_4  FILLER_85_258
timestamp 1606120353
transform 1 0 24840 0 1 48416
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_85_254
timestamp 1606120353
transform 1 0 24472 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__A
timestamp 1606120353
transform 1 0 24656 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0944_
timestamp 1606120353
transform 1 0 25208 0 1 48416
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_86_259
timestamp 1606120353
transform 1 0 24932 0 -1 49504
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_673
timestamp 1606120353
transform 1 0 26404 0 -1 49504
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0944__A
timestamp 1606120353
transform 1 0 25668 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_85_265
timestamp 1606120353
transform 1 0 25484 0 1 48416
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_85_269
timestamp 1606120353
transform 1 0 25852 0 1 48416
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_85_281
timestamp 1606120353
transform 1 0 26956 0 1 48416
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_86_271
timestamp 1606120353
transform 1 0 26036 0 -1 49504
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_86_276
timestamp 1606120353
transform 1 0 26496 0 -1 49504
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1606120353
transform -1 0 28888 0 1 48416
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1606120353
transform -1 0 28888 0 -1 49504
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_85_293
timestamp 1606120353
transform 1 0 28060 0 1 48416
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILLER_86_288
timestamp 1606120353
transform 1 0 27600 0 -1 49504
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_86_296
timestamp 1606120353
transform 1 0 28336 0 -1 49504
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1606120353
transform 1 0 1104 0 1 49504
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_87_3
timestamp 1606120353
transform 1 0 1380 0 1 49504
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_87_15
timestamp 1606120353
transform 1 0 2484 0 1 49504
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_87_27
timestamp 1606120353
transform 1 0 3588 0 1 49504
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_87_39
timestamp 1606120353
transform 1 0 4692 0 1 49504
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_674
timestamp 1606120353
transform 1 0 6716 0 1 49504
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__D
timestamp 1606120353
transform 1 0 7176 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_87_51
timestamp 1606120353
transform 1 0 5796 0 1 49504
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_87_59
timestamp 1606120353
transform 1 0 6532 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_87_62
timestamp 1606120353
transform 1 0 6808 0 1 49504
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1179_
timestamp 1606120353
transform 1 0 7360 0 1 49504
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_6  FILLER_87_87
timestamp 1606120353
transform 1 0 9108 0 1 49504
box 0 -48 552 592
use sky130_fd_sc_hd__a21o_4  _0734_
timestamp 1606120353
transform 1 0 10304 0 1 49504
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__A1
timestamp 1606120353
transform 1 0 10120 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__D
timestamp 1606120353
transform 1 0 9752 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_87_93
timestamp 1606120353
transform 1 0 9660 0 1 49504
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_87_96
timestamp 1606120353
transform 1 0 9936 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1155_
timestamp 1606120353
transform 1 0 12972 0 1 49504
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_675
timestamp 1606120353
transform 1 0 12328 0 1 49504
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__A
timestamp 1606120353
transform 1 0 12788 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__B
timestamp 1606120353
transform 1 0 12144 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__CLK
timestamp 1606120353
transform 1 0 11776 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_87_112
timestamp 1606120353
transform 1 0 11408 0 1 49504
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_87_118
timestamp 1606120353
transform 1 0 11960 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_87_123
timestamp 1606120353
transform 1 0 12420 0 1 49504
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__C
timestamp 1606120353
transform 1 0 15272 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__A1
timestamp 1606120353
transform 1 0 14904 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_87_148
timestamp 1606120353
transform 1 0 14720 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_87_152
timestamp 1606120353
transform 1 0 15088 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1033_
timestamp 1606120353
transform 1 0 15456 0 1 49504
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__C
timestamp 1606120353
transform 1 0 17020 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_87_169
timestamp 1606120353
transform 1 0 16652 0 1 49504
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_87_175
timestamp 1606120353
transform 1 0 17204 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1002_
timestamp 1606120353
transform 1 0 18492 0 1 49504
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_676
timestamp 1606120353
transform 1 0 17940 0 1 49504
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__A1
timestamp 1606120353
transform 1 0 18308 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__D
timestamp 1606120353
transform 1 0 17388 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__A2
timestamp 1606120353
transform 1 0 17756 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_87_179
timestamp 1606120353
transform 1 0 17572 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_87_184
timestamp 1606120353
transform 1 0 18032 0 1 49504
box 0 -48 276 592
use sky130_fd_sc_hd__and4_4  _0916_
timestamp 1606120353
transform 1 0 21068 0 1 49504
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__A
timestamp 1606120353
transform 1 0 20884 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__B
timestamp 1606120353
transform 1 0 20516 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__A
timestamp 1606120353
transform 1 0 20148 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_87_202
timestamp 1606120353
transform 1 0 19688 0 1 49504
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_87_206
timestamp 1606120353
transform 1 0 20056 0 1 49504
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_87_209
timestamp 1606120353
transform 1 0 20332 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_87_213
timestamp 1606120353
transform 1 0 20700 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__A
timestamp 1606120353
transform 1 0 23368 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__A
timestamp 1606120353
transform 1 0 22448 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__C
timestamp 1606120353
transform 1 0 22816 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__B
timestamp 1606120353
transform 1 0 22080 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_87_226
timestamp 1606120353
transform 1 0 21896 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_87_230
timestamp 1606120353
transform 1 0 22264 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_87_234
timestamp 1606120353
transform 1 0 22632 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_87_238
timestamp 1606120353
transform 1 0 23000 0 1 49504
box 0 -48 368 592
use sky130_fd_sc_hd__inv_8  _0843_
timestamp 1606120353
transform 1 0 23644 0 1 49504
box 0 -48 828 592
use sky130_fd_sc_hd__buf_1  _0998_
timestamp 1606120353
transform 1 0 25208 0 1 49504
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_677
timestamp 1606120353
transform 1 0 23552 0 1 49504
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__A
timestamp 1606120353
transform 1 0 24656 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_87_254
timestamp 1606120353
transform 1 0 24472 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_87_258
timestamp 1606120353
transform 1 0 24840 0 1 49504
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__A
timestamp 1606120353
transform 1 0 25668 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_87_265
timestamp 1606120353
transform 1 0 25484 0 1 49504
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_87_269
timestamp 1606120353
transform 1 0 25852 0 1 49504
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_87_281
timestamp 1606120353
transform 1 0 26956 0 1 49504
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1606120353
transform -1 0 28888 0 1 49504
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_87_293
timestamp 1606120353
transform 1 0 28060 0 1 49504
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1606120353
transform 1 0 1104 0 -1 50592
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_88_3
timestamp 1606120353
transform 1 0 1380 0 -1 50592
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_88_15
timestamp 1606120353
transform 1 0 2484 0 -1 50592
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_678
timestamp 1606120353
transform 1 0 3956 0 -1 50592
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_88_27
timestamp 1606120353
transform 1 0 3588 0 -1 50592
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_88_32
timestamp 1606120353
transform 1 0 4048 0 -1 50592
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_88_44
timestamp 1606120353
transform 1 0 5152 0 -1 50592
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_88_56
timestamp 1606120353
transform 1 0 6256 0 -1 50592
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_88_68
timestamp 1606120353
transform 1 0 7360 0 -1 50592
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_88_80
timestamp 1606120353
transform 1 0 8464 0 -1 50592
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1085_
timestamp 1606120353
transform 1 0 10396 0 -1 50592
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_679
timestamp 1606120353
transform 1 0 9568 0 -1 50592
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_88_93
timestamp 1606120353
transform 1 0 9660 0 -1 50592
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__C
timestamp 1606120353
transform 1 0 13248 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__A
timestamp 1606120353
transform 1 0 12880 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__A
timestamp 1606120353
transform 1 0 12512 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_88_120
timestamp 1606120353
transform 1 0 12144 0 -1 50592
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_88_126
timestamp 1606120353
transform 1 0 12696 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_88_130
timestamp 1606120353
transform 1 0 13064 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _1026_
timestamp 1606120353
transform 1 0 13616 0 -1 50592
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_680
timestamp 1606120353
transform 1 0 15180 0 -1 50592
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__B
timestamp 1606120353
transform 1 0 14812 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_88_134
timestamp 1606120353
transform 1 0 13432 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_88_145
timestamp 1606120353
transform 1 0 14444 0 -1 50592
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_88_151
timestamp 1606120353
transform 1 0 14996 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_88_154
timestamp 1606120353
transform 1 0 15272 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _1009_
timestamp 1606120353
transform 1 0 17020 0 -1 50592
box 0 -48 828 592
use sky130_fd_sc_hd__and3_4  _1046_
timestamp 1606120353
transform 1 0 15456 0 -1 50592
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__A
timestamp 1606120353
transform 1 0 16468 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__C
timestamp 1606120353
transform 1 0 16836 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_88_165
timestamp 1606120353
transform 1 0 16284 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_88_169
timestamp 1606120353
transform 1 0 16652 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _0997_
timestamp 1606120353
transform 1 0 18584 0 -1 50592
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__B1
timestamp 1606120353
transform 1 0 18400 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__B1
timestamp 1606120353
transform 1 0 18032 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_88_182
timestamp 1606120353
transform 1 0 17848 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_88_186
timestamp 1606120353
transform 1 0 18216 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0945_
timestamp 1606120353
transform 1 0 20884 0 -1 50592
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_681
timestamp 1606120353
transform 1 0 20792 0 -1 50592
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__A2
timestamp 1606120353
transform 1 0 20608 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__B1
timestamp 1606120353
transform 1 0 20240 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_88_203
timestamp 1606120353
transform 1 0 19780 0 -1 50592
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_88_207
timestamp 1606120353
transform 1 0 20148 0 -1 50592
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_88_210
timestamp 1606120353
transform 1 0 20424 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0987_
timestamp 1606120353
transform 1 0 22448 0 -1 50592
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__C
timestamp 1606120353
transform 1 0 21896 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__B
timestamp 1606120353
transform 1 0 22264 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_88_224
timestamp 1606120353
transform 1 0 21712 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_88_228
timestamp 1606120353
transform 1 0 22080 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_88_241
timestamp 1606120353
transform 1 0 23276 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0851_
timestamp 1606120353
transform 1 0 24012 0 -1 50592
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__D
timestamp 1606120353
transform 1 0 23460 0 -1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_88_245
timestamp 1606120353
transform 1 0 23644 0 -1 50592
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_88_258
timestamp 1606120353
transform 1 0 24840 0 -1 50592
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_682
timestamp 1606120353
transform 1 0 26404 0 -1 50592
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_88_270
timestamp 1606120353
transform 1 0 25944 0 -1 50592
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_88_274
timestamp 1606120353
transform 1 0 26312 0 -1 50592
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_88_276
timestamp 1606120353
transform 1 0 26496 0 -1 50592
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1606120353
transform -1 0 28888 0 -1 50592
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_88_288
timestamp 1606120353
transform 1 0 27600 0 -1 50592
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_88_296
timestamp 1606120353
transform 1 0 28336 0 -1 50592
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1606120353
transform 1 0 1104 0 1 50592
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_89_3
timestamp 1606120353
transform 1 0 1380 0 1 50592
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_89_15
timestamp 1606120353
transform 1 0 2484 0 1 50592
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_89_27
timestamp 1606120353
transform 1 0 3588 0 1 50592
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_89_39
timestamp 1606120353
transform 1 0 4692 0 1 50592
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_683
timestamp 1606120353
transform 1 0 6716 0 1 50592
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_clk_A
timestamp 1606120353
transform 1 0 5888 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_89_51
timestamp 1606120353
transform 1 0 5796 0 1 50592
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_89_54
timestamp 1606120353
transform 1 0 6072 0 1 50592
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_89_60
timestamp 1606120353
transform 1 0 6624 0 1 50592
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_89_62
timestamp 1606120353
transform 1 0 6808 0 1 50592
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_89_74
timestamp 1606120353
transform 1 0 7912 0 1 50592
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_89_86
timestamp 1606120353
transform 1 0 9016 0 1 50592
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__D
timestamp 1606120353
transform 1 0 11132 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_clk_A
timestamp 1606120353
transform 1 0 10396 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_89_98
timestamp 1606120353
transform 1 0 10120 0 1 50592
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_89_103
timestamp 1606120353
transform 1 0 10580 0 1 50592
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_89_118
timestamp 1606120353
transform 1 0 11960 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_114
timestamp 1606120353
transform 1 0 11592 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__A
timestamp 1606120353
transform 1 0 11776 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0957_
timestamp 1606120353
transform 1 0 11316 0 1 50592
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_89_128
timestamp 1606120353
transform 1 0 12880 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_89_123
timestamp 1606120353
transform 1 0 12420 0 1 50592
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__A
timestamp 1606120353
transform 1 0 12144 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__B
timestamp 1606120353
transform 1 0 12696 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_684
timestamp 1606120353
transform 1 0 12328 0 1 50592
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__D
timestamp 1606120353
transform 1 0 13064 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _1027_
timestamp 1606120353
transform 1 0 13248 0 1 50592
box 0 -48 828 592
use sky130_fd_sc_hd__or4_4  _1039_
timestamp 1606120353
transform 1 0 14812 0 1 50592
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__A
timestamp 1606120353
transform 1 0 14628 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__A
timestamp 1606120353
transform 1 0 14260 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_141
timestamp 1606120353
transform 1 0 14076 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_145
timestamp 1606120353
transform 1 0 14444 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__and3_4  _1010_
timestamp 1606120353
transform 1 0 16376 0 1 50592
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__C
timestamp 1606120353
transform 1 0 16192 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__A
timestamp 1606120353
transform 1 0 15824 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_158
timestamp 1606120353
transform 1 0 15640 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_162
timestamp 1606120353
transform 1 0 16008 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_175
timestamp 1606120353
transform 1 0 17204 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0996_
timestamp 1606120353
transform 1 0 18860 0 1 50592
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_685
timestamp 1606120353
transform 1 0 17940 0 1 50592
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__A
timestamp 1606120353
transform 1 0 18676 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__B
timestamp 1606120353
transform 1 0 17388 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__B
timestamp 1606120353
transform 1 0 17756 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__C
timestamp 1606120353
transform 1 0 18216 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_179
timestamp 1606120353
transform 1 0 17572 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_184
timestamp 1606120353
transform 1 0 18032 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_89_188
timestamp 1606120353
transform 1 0 18400 0 1 50592
box 0 -48 276 592
use sky130_fd_sc_hd__and4_4  _0908_
timestamp 1606120353
transform 1 0 21160 0 1 50592
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__A
timestamp 1606120353
transform 1 0 20976 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__B
timestamp 1606120353
transform 1 0 20608 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__C
timestamp 1606120353
transform 1 0 20240 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_89_205
timestamp 1606120353
transform 1 0 19964 0 1 50592
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_89_210
timestamp 1606120353
transform 1 0 20424 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_214
timestamp 1606120353
transform 1 0 20792 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__A2
timestamp 1606120353
transform 1 0 23184 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__B1
timestamp 1606120353
transform 1 0 22816 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__A1
timestamp 1606120353
transform 1 0 22172 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_227
timestamp 1606120353
transform 1 0 21988 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_89_231
timestamp 1606120353
transform 1 0 22356 0 1 50592
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_89_235
timestamp 1606120353
transform 1 0 22724 0 1 50592
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_89_238
timestamp 1606120353
transform 1 0 23000 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_242
timestamp 1606120353
transform 1 0 23368 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1173_
timestamp 1606120353
transform 1 0 24380 0 1 50592
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_686
timestamp 1606120353
transform 1 0 23552 0 1 50592
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__D
timestamp 1606120353
transform 1 0 24196 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__A1
timestamp 1606120353
transform 1 0 23828 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_245
timestamp 1606120353
transform 1 0 23644 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_89_249
timestamp 1606120353
transform 1 0 24012 0 1 50592
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_89_272
timestamp 1606120353
transform 1 0 26128 0 1 50592
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_89_284
timestamp 1606120353
transform 1 0 27232 0 1 50592
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1606120353
transform -1 0 28888 0 1 50592
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_89_296
timestamp 1606120353
transform 1 0 28336 0 1 50592
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1606120353
transform 1 0 1104 0 -1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_90_3
timestamp 1606120353
transform 1 0 1380 0 -1 51680
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_90_15
timestamp 1606120353
transform 1 0 2484 0 -1 51680
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_687
timestamp 1606120353
transform 1 0 3956 0 -1 51680
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_90_27
timestamp 1606120353
transform 1 0 3588 0 -1 51680
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_90_32
timestamp 1606120353
transform 1 0 4048 0 -1 51680
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_90_44
timestamp 1606120353
transform 1 0 5152 0 -1 51680
box 0 -48 736 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_clk
timestamp 1606120353
transform 1 0 5888 0 -1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_90_55
timestamp 1606120353
transform 1 0 6164 0 -1 51680
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_90_67
timestamp 1606120353
transform 1 0 7268 0 -1 51680
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_90_79
timestamp 1606120353
transform 1 0 8372 0 -1 51680
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_688
timestamp 1606120353
transform 1 0 9568 0 -1 51680
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_clk
timestamp 1606120353
transform 1 0 10396 0 -1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__CLK
timestamp 1606120353
transform 1 0 11040 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_90_91
timestamp 1606120353
transform 1 0 9476 0 -1 51680
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_90_93
timestamp 1606120353
transform 1 0 9660 0 -1 51680
box 0 -48 736 592
use sky130_fd_sc_hd__decap_4  FILLER_90_104
timestamp 1606120353
transform 1 0 10672 0 -1 51680
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_90_110
timestamp 1606120353
transform 1 0 11224 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__A
timestamp 1606120353
transform 1 0 11408 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1007_
timestamp 1606120353
transform 1 0 11592 0 -1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_90_117
timestamp 1606120353
transform 1 0 11868 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__D
timestamp 1606120353
transform 1 0 12052 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_90_121
timestamp 1606120353
transform 1 0 12236 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__C
timestamp 1606120353
transform 1 0 12420 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0995_
timestamp 1606120353
transform 1 0 12604 0 -1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_90_128
timestamp 1606120353
transform 1 0 12880 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__A
timestamp 1606120353
transform 1 0 13064 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_90_132
timestamp 1606120353
transform 1 0 13248 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _1034_
timestamp 1606120353
transform 1 0 13616 0 -1 51680
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_689
timestamp 1606120353
transform 1 0 15180 0 -1 51680
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__B
timestamp 1606120353
transform 1 0 13432 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__C
timestamp 1606120353
transform 1 0 14812 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_90_145
timestamp 1606120353
transform 1 0 14444 0 -1 51680
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_90_151
timestamp 1606120353
transform 1 0 14996 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_90_154
timestamp 1606120353
transform 1 0 15272 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0994_
timestamp 1606120353
transform 1 0 16008 0 -1 51680
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__D
timestamp 1606120353
transform 1 0 15456 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__B
timestamp 1606120353
transform 1 0 17020 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__B
timestamp 1606120353
transform 1 0 15824 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_90_158
timestamp 1606120353
transform 1 0 15640 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_90_171
timestamp 1606120353
transform 1 0 16836 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_90_175
timestamp 1606120353
transform 1 0 17204 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__nor3_4  _1011_
timestamp 1606120353
transform 1 0 17572 0 -1 51680
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__A2
timestamp 1606120353
transform 1 0 18952 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__A1
timestamp 1606120353
transform 1 0 19320 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__A
timestamp 1606120353
transform 1 0 17388 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_90_192
timestamp 1606120353
transform 1 0 18768 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_90_196
timestamp 1606120353
transform 1 0 19136 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__a211o_4  _0961_
timestamp 1606120353
transform 1 0 20884 0 -1 51680
box 0 -48 1288 592
use sky130_fd_sc_hd__buf_1  _0968_
timestamp 1606120353
transform 1 0 19504 0 -1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_690
timestamp 1606120353
transform 1 0 20792 0 -1 51680
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__A1
timestamp 1606120353
transform 1 0 20332 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__C1
timestamp 1606120353
transform 1 0 19964 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_90_203
timestamp 1606120353
transform 1 0 19780 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_90_207
timestamp 1606120353
transform 1 0 20148 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_90_211
timestamp 1606120353
transform 1 0 20516 0 -1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__o21a_4  _0855_
timestamp 1606120353
transform 1 0 23184 0 -1 51680
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__B1
timestamp 1606120353
transform 1 0 22908 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__D
timestamp 1606120353
transform 1 0 22356 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_90_229
timestamp 1606120353
transform 1 0 22172 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_90_233
timestamp 1606120353
transform 1 0 22540 0 -1 51680
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_90_239
timestamp 1606120353
transform 1 0 23092 0 -1 51680
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__C
timestamp 1606120353
transform 1 0 24472 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__CLK
timestamp 1606120353
transform 1 0 24840 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_90_252
timestamp 1606120353
transform 1 0 24288 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_90_256
timestamp 1606120353
transform 1 0 24656 0 -1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_90_260
timestamp 1606120353
transform 1 0 25024 0 -1 51680
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_691
timestamp 1606120353
transform 1 0 26404 0 -1 51680
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_90_272
timestamp 1606120353
transform 1 0 26128 0 -1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_90_276
timestamp 1606120353
transform 1 0 26496 0 -1 51680
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1606120353
transform -1 0 28888 0 -1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_90_288
timestamp 1606120353
transform 1 0 27600 0 -1 51680
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_90_296
timestamp 1606120353
transform 1 0 28336 0 -1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1606120353
transform 1 0 1104 0 1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__D
timestamp 1606120353
transform 1 0 1564 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__CLK
timestamp 1606120353
transform 1 0 1932 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_3
timestamp 1606120353
transform 1 0 1380 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_7
timestamp 1606120353
transform 1 0 1748 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_91_11
timestamp 1606120353
transform 1 0 2116 0 1 51680
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_91_23
timestamp 1606120353
transform 1 0 3220 0 1 51680
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_91_35
timestamp 1606120353
transform 1 0 4324 0 1 51680
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_692
timestamp 1606120353
transform 1 0 6716 0 1 51680
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_91_47
timestamp 1606120353
transform 1 0 5428 0 1 51680
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_91_59
timestamp 1606120353
transform 1 0 6532 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_91_62
timestamp 1606120353
transform 1 0 6808 0 1 51680
box 0 -48 736 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_clk
timestamp 1606120353
transform 1 0 7820 0 1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_clk_A
timestamp 1606120353
transform 1 0 8280 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_91_70
timestamp 1606120353
transform 1 0 7544 0 1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_91_76
timestamp 1606120353
transform 1 0 8096 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_91_80
timestamp 1606120353
transform 1 0 8464 0 1 51680
box 0 -48 1104 592
use sky130_fd_sc_hd__buf_1  _0954_
timestamp 1606120353
transform 1 0 10304 0 1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__A
timestamp 1606120353
transform 1 0 10764 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__A
timestamp 1606120353
transform 1 0 11132 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_91_92
timestamp 1606120353
transform 1 0 9568 0 1 51680
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_91_103
timestamp 1606120353
transform 1 0 10580 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_107
timestamp 1606120353
transform 1 0 10948 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1008_
timestamp 1606120353
transform 1 0 11316 0 1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1209_
timestamp 1606120353
transform 1 0 12788 0 1 51680
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_693
timestamp 1606120353
transform 1 0 12328 0 1 51680
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__D
timestamp 1606120353
transform 1 0 12604 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A
timestamp 1606120353
transform 1 0 11776 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__A
timestamp 1606120353
transform 1 0 12144 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_114
timestamp 1606120353
transform 1 0 11592 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_118
timestamp 1606120353
transform 1 0 11960 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_123
timestamp 1606120353
transform 1 0 12420 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0953_
timestamp 1606120353
transform 1 0 15272 0 1 51680
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__A
timestamp 1606120353
transform 1 0 14720 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__B
timestamp 1606120353
transform 1 0 15088 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_146
timestamp 1606120353
transform 1 0 14536 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_150
timestamp 1606120353
transform 1 0 14904 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0971_
timestamp 1606120353
transform 1 0 16836 0 1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__A
timestamp 1606120353
transform 1 0 16652 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__B
timestamp 1606120353
transform 1 0 16284 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_163
timestamp 1606120353
transform 1 0 16100 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_167
timestamp 1606120353
transform 1 0 16468 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_91_174
timestamp 1606120353
transform 1 0 17112 0 1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__nor3_4  _0988_
timestamp 1606120353
transform 1 0 18400 0 1 51680
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_694
timestamp 1606120353
transform 1 0 17940 0 1 51680
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__A
timestamp 1606120353
transform 1 0 18216 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__C
timestamp 1606120353
transform 1 0 17756 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__B
timestamp 1606120353
transform 1 0 17388 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_179
timestamp 1606120353
transform 1 0 17572 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_184
timestamp 1606120353
transform 1 0 18032 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__a211o_4  _0967_
timestamp 1606120353
transform 1 0 20332 0 1 51680
box 0 -48 1288 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A1
timestamp 1606120353
transform 1 0 20148 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__C1
timestamp 1606120353
transform 1 0 19780 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_201
timestamp 1606120353
transform 1 0 19596 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_205
timestamp 1606120353
transform 1 0 19964 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0949_
timestamp 1606120353
transform 1 0 22356 0 1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__A2
timestamp 1606120353
transform 1 0 22908 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__A1
timestamp 1606120353
transform 1 0 23276 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__A
timestamp 1606120353
transform 1 0 22172 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__B1
timestamp 1606120353
transform 1 0 21804 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_223
timestamp 1606120353
transform 1 0 21620 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_227
timestamp 1606120353
transform 1 0 21988 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_91_234
timestamp 1606120353
transform 1 0 22632 0 1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_91_239
timestamp 1606120353
transform 1 0 23092 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _0903_
timestamp 1606120353
transform 1 0 23644 0 1 51680
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_695
timestamp 1606120353
transform 1 0 23552 0 1 51680
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__A
timestamp 1606120353
transform 1 0 24656 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__D
timestamp 1606120353
transform 1 0 25024 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_91_243
timestamp 1606120353
transform 1 0 23460 0 1 51680
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_91_254
timestamp 1606120353
transform 1 0 24472 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_91_258
timestamp 1606120353
transform 1 0 24840 0 1 51680
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_91_262
timestamp 1606120353
transform 1 0 25208 0 1 51680
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_91_274
timestamp 1606120353
transform 1 0 26312 0 1 51680
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_91_286
timestamp 1606120353
transform 1 0 27416 0 1 51680
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1606120353
transform -1 0 28888 0 1 51680
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_91_298
timestamp 1606120353
transform 1 0 28520 0 1 51680
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1206_
timestamp 1606120353
transform 1 0 1380 0 -1 52768
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1606120353
transform 1 0 1104 0 -1 52768
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1606120353
transform 1 0 1104 0 1 52768
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_92_22
timestamp 1606120353
transform 1 0 3128 0 -1 52768
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_93_3
timestamp 1606120353
transform 1 0 1380 0 1 52768
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_93_15
timestamp 1606120353
transform 1 0 2484 0 1 52768
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_696
timestamp 1606120353
transform 1 0 3956 0 -1 52768
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_92_30
timestamp 1606120353
transform 1 0 3864 0 -1 52768
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_92_32
timestamp 1606120353
transform 1 0 4048 0 -1 52768
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_92_44
timestamp 1606120353
transform 1 0 5152 0 -1 52768
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_93_27
timestamp 1606120353
transform 1 0 3588 0 1 52768
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_93_39
timestamp 1606120353
transform 1 0 4692 0 1 52768
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_701
timestamp 1606120353
transform 1 0 6716 0 1 52768
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_92_56
timestamp 1606120353
transform 1 0 6256 0 -1 52768
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_93_51
timestamp 1606120353
transform 1 0 5796 0 1 52768
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_93_59
timestamp 1606120353
transform 1 0 6532 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_93_62
timestamp 1606120353
transform 1 0 6808 0 1 52768
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_92_68
timestamp 1606120353
transform 1 0 7360 0 -1 52768
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_92_80
timestamp 1606120353
transform 1 0 8464 0 -1 52768
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_93_74
timestamp 1606120353
transform 1 0 7912 0 1 52768
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_93_86
timestamp 1606120353
transform 1 0 9016 0 1 52768
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_92_93
timestamp 1606120353
transform 1 0 9660 0 -1 52768
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_697
timestamp 1606120353
transform 1 0 9568 0 -1 52768
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_93_103
timestamp 1606120353
transform 1 0 10580 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_93_98
timestamp 1606120353
transform 1 0 10120 0 1 52768
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_92_101
timestamp 1606120353
transform 1 0 10396 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__CLK
timestamp 1606120353
transform 1 0 10396 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0956_
timestamp 1606120353
transform 1 0 10580 0 -1 52768
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_93_107
timestamp 1606120353
transform 1 0 10948 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_92_106
timestamp 1606120353
transform 1 0 10856 0 -1 52768
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__CLK
timestamp 1606120353
transform 1 0 10764 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__A
timestamp 1606120353
transform 1 0 11132 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0948_
timestamp 1606120353
transform 1 0 11316 0 1 52768
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__A
timestamp 1606120353
transform 1 0 11408 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0951_
timestamp 1606120353
transform 1 0 11592 0 -1 52768
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__A
timestamp 1606120353
transform 1 0 11776 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_93_114
timestamp 1606120353
transform 1 0 11592 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__A
timestamp 1606120353
transform 1 0 12052 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_92_117
timestamp 1606120353
transform 1 0 11868 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_93_118
timestamp 1606120353
transform 1 0 11960 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__D
timestamp 1606120353
transform 1 0 12144 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_92_121
timestamp 1606120353
transform 1 0 12236 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_92_132
timestamp 1606120353
transform 1 0 13248 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_92_128
timestamp 1606120353
transform 1 0 12880 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__D
timestamp 1606120353
transform 1 0 13064 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__D
timestamp 1606120353
transform 1 0 12420 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_702
timestamp 1606120353
transform 1 0 12328 0 1 52768
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _0999_
timestamp 1606120353
transform 1 0 12604 0 -1 52768
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1207_
timestamp 1606120353
transform 1 0 12420 0 1 52768
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__C
timestamp 1606120353
transform 1 0 13432 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__and4_4  _1055_
timestamp 1606120353
transform 1 0 13616 0 -1 52768
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_93_146
timestamp 1606120353
transform 1 0 14536 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_93_142
timestamp 1606120353
transform 1 0 14168 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_92_149
timestamp 1606120353
transform 1 0 14812 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_92_145
timestamp 1606120353
transform 1 0 14444 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__B
timestamp 1606120353
transform 1 0 14352 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1048__C
timestamp 1606120353
transform 1 0 14628 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__A
timestamp 1606120353
transform 1 0 14720 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0950_
timestamp 1606120353
transform 1 0 14904 0 1 52768
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1048__B
timestamp 1606120353
transform 1 0 14996 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_698
timestamp 1606120353
transform 1 0 15180 0 -1 52768
box 0 -48 92 592
use sky130_fd_sc_hd__inv_8  _1003_
timestamp 1606120353
transform 1 0 15272 0 -1 52768
box 0 -48 828 592
use sky130_fd_sc_hd__decap_4  FILLER_93_159
timestamp 1606120353
transform 1 0 15732 0 1 52768
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_93_166
timestamp 1606120353
transform 1 0 16376 0 1 52768
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_93_163
timestamp 1606120353
transform 1 0 16100 0 1 52768
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_92_163
timestamp 1606120353
transform 1 0 16100 0 -1 52768
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__A
timestamp 1606120353
transform 1 0 16468 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__A
timestamp 1606120353
transform 1 0 16192 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1032_
timestamp 1606120353
transform 1 0 16468 0 1 52768
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_93_174
timestamp 1606120353
transform 1 0 17112 0 1 52768
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_93_170
timestamp 1606120353
transform 1 0 16744 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_92_169
timestamp 1606120353
transform 1 0 16652 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__B
timestamp 1606120353
transform 1 0 16928 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__or2_4  _1028_
timestamp 1606120353
transform 1 0 16836 0 -1 52768
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILLER_93_179
timestamp 1606120353
transform 1 0 17572 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_92_182
timestamp 1606120353
transform 1 0 17848 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_92_178
timestamp 1606120353
transform 1 0 17480 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__B
timestamp 1606120353
transform 1 0 17664 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__D
timestamp 1606120353
transform 1 0 17388 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__C
timestamp 1606120353
transform 1 0 18032 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__A
timestamp 1606120353
transform 1 0 17756 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_703
timestamp 1606120353
transform 1 0 17940 0 1 52768
box 0 -48 92 592
use sky130_fd_sc_hd__and4_4  _1045_
timestamp 1606120353
transform 1 0 18032 0 1 52768
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_93_198
timestamp 1606120353
transform 1 0 19320 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_93_193
timestamp 1606120353
transform 1 0 18860 0 1 52768
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__A1
timestamp 1606120353
transform 1 0 19136 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__nor3_4  _1048_
timestamp 1606120353
transform 1 0 18216 0 -1 52768
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_92_207
timestamp 1606120353
transform 1 0 20148 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_92_203
timestamp 1606120353
transform 1 0 19780 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_92_199
timestamp 1606120353
transform 1 0 19412 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__A2
timestamp 1606120353
transform 1 0 19596 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__C
timestamp 1606120353
transform 1 0 19964 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__B1
timestamp 1606120353
transform 1 0 20332 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1044__A
timestamp 1606120353
transform 1 0 19504 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_93_219
timestamp 1606120353
transform 1 0 21252 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_93_215
timestamp 1606120353
transform 1 0 20884 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_92_211
timestamp 1606120353
transform 1 0 20516 0 -1 52768
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__A
timestamp 1606120353
transform 1 0 21068 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_699
timestamp 1606120353
transform 1 0 20792 0 -1 52768
box 0 -48 92 592
use sky130_fd_sc_hd__o21ai_4  _0980_
timestamp 1606120353
transform 1 0 19688 0 1 52768
box 0 -48 1196 592
use sky130_fd_sc_hd__a21oi_4  _0975_
timestamp 1606120353
transform 1 0 20884 0 -1 52768
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_93_230
timestamp 1606120353
transform 1 0 22264 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_92_228
timestamp 1606120353
transform 1 0 22080 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A2
timestamp 1606120353
transform 1 0 22264 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__B
timestamp 1606120353
transform 1 0 21436 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__and2_4  _0946_
timestamp 1606120353
transform 1 0 21620 0 1 52768
box 0 -48 644 592
use sky130_fd_sc_hd__fill_2  FILLER_93_240
timestamp 1606120353
transform 1 0 23184 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_93_234
timestamp 1606120353
transform 1 0 22632 0 1 52768
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_92_232
timestamp 1606120353
transform 1 0 22448 0 -1 52768
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__A1
timestamp 1606120353
transform 1 0 22724 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__A2
timestamp 1606120353
transform 1 0 23368 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__B1_N
timestamp 1606120353
transform 1 0 23000 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__A
timestamp 1606120353
transform 1 0 22448 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _0856_
timestamp 1606120353
transform 1 0 22908 0 -1 52768
box 0 -48 1196 592
use sky130_fd_sc_hd__dfxtp_4  _1194_
timestamp 1606120353
transform 1 0 24196 0 1 52768
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_704
timestamp 1606120353
transform 1 0 23552 0 1 52768
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__D
timestamp 1606120353
transform 1 0 24012 0 1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__B
timestamp 1606120353
transform 1 0 24288 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_92_250
timestamp 1606120353
transform 1 0 24104 0 -1 52768
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_92_254
timestamp 1606120353
transform 1 0 24472 0 -1 52768
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_93_245
timestamp 1606120353
transform 1 0 23644 0 1 52768
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_700
timestamp 1606120353
transform 1 0 26404 0 -1 52768
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_92_266
timestamp 1606120353
transform 1 0 25576 0 -1 52768
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_92_274
timestamp 1606120353
transform 1 0 26312 0 -1 52768
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_92_276
timestamp 1606120353
transform 1 0 26496 0 -1 52768
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_93_270
timestamp 1606120353
transform 1 0 25944 0 1 52768
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_93_282
timestamp 1606120353
transform 1 0 27048 0 1 52768
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1606120353
transform -1 0 28888 0 -1 52768
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1606120353
transform -1 0 28888 0 1 52768
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_92_288
timestamp 1606120353
transform 1 0 27600 0 -1 52768
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_92_296
timestamp 1606120353
transform 1 0 28336 0 -1 52768
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_93_294
timestamp 1606120353
transform 1 0 28152 0 1 52768
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_93_298
timestamp 1606120353
transform 1 0 28520 0 1 52768
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1606120353
transform 1 0 1104 0 -1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_94_3
timestamp 1606120353
transform 1 0 1380 0 -1 53856
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_94_15
timestamp 1606120353
transform 1 0 2484 0 -1 53856
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_705
timestamp 1606120353
transform 1 0 3956 0 -1 53856
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_94_27
timestamp 1606120353
transform 1 0 3588 0 -1 53856
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_94_32
timestamp 1606120353
transform 1 0 4048 0 -1 53856
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_94_44
timestamp 1606120353
transform 1 0 5152 0 -1 53856
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_94_56
timestamp 1606120353
transform 1 0 6256 0 -1 53856
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_94_68
timestamp 1606120353
transform 1 0 7360 0 -1 53856
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_94_80
timestamp 1606120353
transform 1 0 8464 0 -1 53856
box 0 -48 1104 592
use sky130_fd_sc_hd__buf_1  _0963_
timestamp 1606120353
transform 1 0 11224 0 -1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_706
timestamp 1606120353
transform 1 0 9568 0 -1 53856
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_94_93
timestamp 1606120353
transform 1 0 9660 0 -1 53856
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_94_105
timestamp 1606120353
transform 1 0 10764 0 -1 53856
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_94_109
timestamp 1606120353
transform 1 0 11132 0 -1 53856
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1208_
timestamp 1606120353
transform 1 0 12236 0 -1 53856
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__C
timestamp 1606120353
transform 1 0 12052 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__D
timestamp 1606120353
transform 1 0 11684 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_94_113
timestamp 1606120353
transform 1 0 11500 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_94_117
timestamp 1606120353
transform 1 0 11868 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_707
timestamp 1606120353
transform 1 0 15180 0 -1 53856
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__C
timestamp 1606120353
transform 1 0 14996 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__A
timestamp 1606120353
transform 1 0 14628 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__B
timestamp 1606120353
transform 1 0 14260 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_94_140
timestamp 1606120353
transform 1 0 13984 0 -1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_94_145
timestamp 1606120353
transform 1 0 14444 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_94_149
timestamp 1606120353
transform 1 0 14812 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_94_154
timestamp 1606120353
transform 1 0 15272 0 -1 53856
box 0 -48 368 592
use sky130_fd_sc_hd__or4_4  _0964_
timestamp 1606120353
transform 1 0 16192 0 -1 53856
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__B
timestamp 1606120353
transform 1 0 15640 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__D
timestamp 1606120353
transform 1 0 16008 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1048__A
timestamp 1606120353
transform 1 0 17204 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_94_160
timestamp 1606120353
transform 1 0 15824 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_94_173
timestamp 1606120353
transform 1 0 17020 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__nor3_4  _1056_
timestamp 1606120353
transform 1 0 17756 0 -1 53856
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__C
timestamp 1606120353
transform 1 0 17572 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__A2
timestamp 1606120353
transform 1 0 19136 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_94_177
timestamp 1606120353
transform 1 0 17388 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_94_194
timestamp 1606120353
transform 1 0 18952 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_94_198
timestamp 1606120353
transform 1 0 19320 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__or3_4  _0960_
timestamp 1606120353
transform 1 0 20884 0 -1 53856
box 0 -48 828 592
use sky130_fd_sc_hd__buf_1  _1044_
timestamp 1606120353
transform 1 0 19688 0 -1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_708
timestamp 1606120353
transform 1 0 20792 0 -1 53856
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__B1_N
timestamp 1606120353
transform 1 0 20608 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__B
timestamp 1606120353
transform 1 0 20240 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__B1
timestamp 1606120353
transform 1 0 19504 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_94_205
timestamp 1606120353
transform 1 0 19964 0 -1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_94_210
timestamp 1606120353
transform 1 0 20424 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0936_
timestamp 1606120353
transform 1 0 23000 0 -1 53856
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__B1_N
timestamp 1606120353
transform 1 0 22816 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A1
timestamp 1606120353
transform 1 0 21896 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__A1
timestamp 1606120353
transform 1 0 22264 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_94_224
timestamp 1606120353
transform 1 0 21712 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_94_228
timestamp 1606120353
transform 1 0 22080 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_94_232
timestamp 1606120353
transform 1 0 22448 0 -1 53856
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__CLK
timestamp 1606120353
transform 1 0 24380 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_94_251
timestamp 1606120353
transform 1 0 24196 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_94_255
timestamp 1606120353
transform 1 0 24564 0 -1 53856
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_709
timestamp 1606120353
transform 1 0 26404 0 -1 53856
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__B1_N
timestamp 1606120353
transform 1 0 26680 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__A2
timestamp 1606120353
transform 1 0 27048 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__CLK
timestamp 1606120353
transform 1 0 25944 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_94_267
timestamp 1606120353
transform 1 0 25668 0 -1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_94_272
timestamp 1606120353
transform 1 0 26128 0 -1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_94_276
timestamp 1606120353
transform 1 0 26496 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_94_280
timestamp 1606120353
transform 1 0 26864 0 -1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_94_284
timestamp 1606120353
transform 1 0 27232 0 -1 53856
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1606120353
transform -1 0 28888 0 -1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_94_296
timestamp 1606120353
transform 1 0 28336 0 -1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1606120353
transform 1 0 1104 0 1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_95_3
timestamp 1606120353
transform 1 0 1380 0 1 53856
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_95_15
timestamp 1606120353
transform 1 0 2484 0 1 53856
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_95_27
timestamp 1606120353
transform 1 0 3588 0 1 53856
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_95_39
timestamp 1606120353
transform 1 0 4692 0 1 53856
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_710
timestamp 1606120353
transform 1 0 6716 0 1 53856
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_95_51
timestamp 1606120353
transform 1 0 5796 0 1 53856
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_95_59
timestamp 1606120353
transform 1 0 6532 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_95_62
timestamp 1606120353
transform 1 0 6808 0 1 53856
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_95_74
timestamp 1606120353
transform 1 0 7912 0 1 53856
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_95_86
timestamp 1606120353
transform 1 0 9016 0 1 53856
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_95_98
timestamp 1606120353
transform 1 0 10120 0 1 53856
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_95_110
timestamp 1606120353
transform 1 0 11224 0 1 53856
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_95_114
timestamp 1606120353
transform 1 0 11592 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0941_
timestamp 1606120353
transform 1 0 11316 0 1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_95_118
timestamp 1606120353
transform 1 0 11960 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0941__A
timestamp 1606120353
transform 1 0 11776 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__A
timestamp 1606120353
transform 1 0 12144 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_711
timestamp 1606120353
transform 1 0 12328 0 1 53856
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_95_123
timestamp 1606120353
transform 1 0 12420 0 1 53856
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__A
timestamp 1606120353
transform 1 0 12788 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0981_
timestamp 1606120353
transform 1 0 12972 0 1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_95_132
timestamp 1606120353
transform 1 0 13248 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0947_
timestamp 1606120353
transform 1 0 13984 0 1 53856
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__A
timestamp 1606120353
transform 1 0 13432 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__C
timestamp 1606120353
transform 1 0 14996 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__A
timestamp 1606120353
transform 1 0 13800 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_136
timestamp 1606120353
transform 1 0 13616 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_149
timestamp 1606120353
transform 1 0 14812 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_153
timestamp 1606120353
transform 1 0 15180 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0940_
timestamp 1606120353
transform 1 0 15548 0 1 53856
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A
timestamp 1606120353
transform 1 0 17020 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__A
timestamp 1606120353
transform 1 0 15364 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__D
timestamp 1606120353
transform 1 0 16560 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_166
timestamp 1606120353
transform 1 0 16376 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_95_170
timestamp 1606120353
transform 1 0 16744 0 1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_95_175
timestamp 1606120353
transform 1 0 17204 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__and3_4  _0952_
timestamp 1606120353
transform 1 0 18032 0 1 53856
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_712
timestamp 1606120353
transform 1 0 17940 0 1 53856
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__D
timestamp 1606120353
transform 1 0 17756 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__C
timestamp 1606120353
transform 1 0 17388 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__A
timestamp 1606120353
transform 1 0 19044 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_179
timestamp 1606120353
transform 1 0 17572 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_193
timestamp 1606120353
transform 1 0 18860 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_95_197
timestamp 1606120353
transform 1 0 19228 0 1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__inv_8  _0942_
timestamp 1606120353
transform 1 0 19688 0 1 53856
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__B1
timestamp 1606120353
transform 1 0 21160 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A2
timestamp 1606120353
transform 1 0 20792 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__A
timestamp 1606120353
transform 1 0 19504 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_95_211
timestamp 1606120353
transform 1 0 20516 0 1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_95_216
timestamp 1606120353
transform 1 0 20976 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_220
timestamp 1606120353
transform 1 0 21344 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0904_
timestamp 1606120353
transform 1 0 21712 0 1 53856
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__A
timestamp 1606120353
transform 1 0 23368 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__A2
timestamp 1606120353
transform 1 0 23000 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__A2
timestamp 1606120353
transform 1 0 21528 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_236
timestamp 1606120353
transform 1 0 22816 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_240
timestamp 1606120353
transform 1 0 23184 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _0905_
timestamp 1606120353
transform 1 0 23644 0 1 53856
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_713
timestamp 1606120353
transform 1 0 23552 0 1 53856
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__B
timestamp 1606120353
transform 1 0 24656 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_254
timestamp 1606120353
transform 1 0 24472 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_95_258
timestamp 1606120353
transform 1 0 24840 0 1 53856
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1189_
timestamp 1606120353
transform 1 0 25944 0 1 53856
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__D
timestamp 1606120353
transform 1 0 25760 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_266
timestamp 1606120353
transform 1 0 25576 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1606120353
transform -1 0 28888 0 1 53856
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__A1
timestamp 1606120353
transform 1 0 27876 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_95_289
timestamp 1606120353
transform 1 0 27692 0 1 53856
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_95_293
timestamp 1606120353
transform 1 0 28060 0 1 53856
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1606120353
transform 1 0 1104 0 -1 54944
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_96_3
timestamp 1606120353
transform 1 0 1380 0 -1 54944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_96_15
timestamp 1606120353
transform 1 0 2484 0 -1 54944
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_714
timestamp 1606120353
transform 1 0 3956 0 -1 54944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_96_27
timestamp 1606120353
transform 1 0 3588 0 -1 54944
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_96_32
timestamp 1606120353
transform 1 0 4048 0 -1 54944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_96_44
timestamp 1606120353
transform 1 0 5152 0 -1 54944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_96_56
timestamp 1606120353
transform 1 0 6256 0 -1 54944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_96_68
timestamp 1606120353
transform 1 0 7360 0 -1 54944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_96_80
timestamp 1606120353
transform 1 0 8464 0 -1 54944
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_715
timestamp 1606120353
transform 1 0 9568 0 -1 54944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_96_93
timestamp 1606120353
transform 1 0 9660 0 -1 54944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_96_105
timestamp 1606120353
transform 1 0 10764 0 -1 54944
box 0 -48 1104 592
use sky130_fd_sc_hd__buf_1  _0962_
timestamp 1606120353
transform 1 0 12144 0 -1 54944
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0970_
timestamp 1606120353
transform 1 0 13156 0 -1 54944
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__C
timestamp 1606120353
transform 1 0 12972 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__A
timestamp 1606120353
transform 1 0 12604 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__D
timestamp 1606120353
transform 1 0 11960 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_96_117
timestamp 1606120353
transform 1 0 11868 0 -1 54944
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_96_123
timestamp 1606120353
transform 1 0 12420 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_96_127
timestamp 1606120353
transform 1 0 12788 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_96_134
timestamp 1606120353
transform 1 0 13432 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_96_138
timestamp 1606120353
transform 1 0 13800 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__A
timestamp 1606120353
transform 1 0 13616 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__D
timestamp 1606120353
transform 1 0 13984 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0972_
timestamp 1606120353
transform 1 0 14168 0 -1 54944
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_96_145
timestamp 1606120353
transform 1 0 14444 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__B
timestamp 1606120353
transform 1 0 14628 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_96_149
timestamp 1606120353
transform 1 0 14812 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__C
timestamp 1606120353
transform 1 0 14996 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_716
timestamp 1606120353
transform 1 0 15180 0 -1 54944
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_96_154
timestamp 1606120353
transform 1 0 15272 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _1031_
timestamp 1606120353
transform 1 0 15640 0 -1 54944
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__D
timestamp 1606120353
transform 1 0 16652 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__A
timestamp 1606120353
transform 1 0 15456 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__C
timestamp 1606120353
transform 1 0 17020 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_96_167
timestamp 1606120353
transform 1 0 16468 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_96_171
timestamp 1606120353
transform 1 0 16836 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_96_175
timestamp 1606120353
transform 1 0 17204 0 -1 54944
box 0 -48 368 592
use sky130_fd_sc_hd__and4_4  _0955_
timestamp 1606120353
transform 1 0 17848 0 -1 54944
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__B
timestamp 1606120353
transform 1 0 17664 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__B
timestamp 1606120353
transform 1 0 18860 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A2
timestamp 1606120353
transform 1 0 19228 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_96_179
timestamp 1606120353
transform 1 0 17572 0 -1 54944
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_96_191
timestamp 1606120353
transform 1 0 18676 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_96_195
timestamp 1606120353
transform 1 0 19044 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0911_
timestamp 1606120353
transform 1 0 20884 0 -1 54944
box 0 -48 1196 592
use sky130_fd_sc_hd__buf_1  _0979_
timestamp 1606120353
transform 1 0 19412 0 -1 54944
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_717
timestamp 1606120353
transform 1 0 20792 0 -1 54944
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A
timestamp 1606120353
transform 1 0 19872 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A1
timestamp 1606120353
transform 1 0 20240 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__B1
timestamp 1606120353
transform 1 0 20608 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_96_202
timestamp 1606120353
transform 1 0 19688 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_96_206
timestamp 1606120353
transform 1 0 20056 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_96_210
timestamp 1606120353
transform 1 0 20424 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0906_
timestamp 1606120353
transform 1 0 22816 0 -1 54944
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__B
timestamp 1606120353
transform 1 0 22264 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__A1
timestamp 1606120353
transform 1 0 22632 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_96_228
timestamp 1606120353
transform 1 0 22080 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_96_232
timestamp 1606120353
transform 1 0 22448 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__B1_N
timestamp 1606120353
transform 1 0 24196 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__A1
timestamp 1606120353
transform 1 0 24564 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_96_249
timestamp 1606120353
transform 1 0 24012 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_96_253
timestamp 1606120353
transform 1 0 24380 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_96_257
timestamp 1606120353
transform 1 0 24748 0 -1 54944
box 0 -48 1104 592
use sky130_fd_sc_hd__a21bo_4  _0937_
timestamp 1606120353
transform 1 0 26496 0 -1 54944
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_718
timestamp 1606120353
transform 1 0 26404 0 -1 54944
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__CLK
timestamp 1606120353
transform 1 0 26128 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_96_269
timestamp 1606120353
transform 1 0 25852 0 -1 54944
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_96_274
timestamp 1606120353
transform 1 0 26312 0 -1 54944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1606120353
transform -1 0 28888 0 -1 54944
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_96_289
timestamp 1606120353
transform 1 0 27692 0 -1 54944
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_96_297
timestamp 1606120353
transform 1 0 28428 0 -1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1606120353
transform 1 0 1104 0 1 54944
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_97_3
timestamp 1606120353
transform 1 0 1380 0 1 54944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_97_15
timestamp 1606120353
transform 1 0 2484 0 1 54944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_97_27
timestamp 1606120353
transform 1 0 3588 0 1 54944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_97_39
timestamp 1606120353
transform 1 0 4692 0 1 54944
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_719
timestamp 1606120353
transform 1 0 6716 0 1 54944
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_97_51
timestamp 1606120353
transform 1 0 5796 0 1 54944
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_97_59
timestamp 1606120353
transform 1 0 6532 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_97_62
timestamp 1606120353
transform 1 0 6808 0 1 54944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_97_74
timestamp 1606120353
transform 1 0 7912 0 1 54944
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_97_86
timestamp 1606120353
transform 1 0 9016 0 1 54944
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__D
timestamp 1606120353
transform 1 0 10488 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__CLK
timestamp 1606120353
transform 1 0 10856 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_97_98
timestamp 1606120353
transform 1 0 10120 0 1 54944
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_97_104
timestamp 1606120353
transform 1 0 10672 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_97_108
timestamp 1606120353
transform 1 0 11040 0 1 54944
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_720
timestamp 1606120353
transform 1 0 12328 0 1 54944
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__A
timestamp 1606120353
transform 1 0 13248 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__A
timestamp 1606120353
transform 1 0 12880 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_120
timestamp 1606120353
transform 1 0 12144 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_97_123
timestamp 1606120353
transform 1 0 12420 0 1 54944
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_97_127
timestamp 1606120353
transform 1 0 12788 0 1 54944
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_97_130
timestamp 1606120353
transform 1 0 13064 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1004_
timestamp 1606120353
transform 1 0 13432 0 1 54944
box 0 -48 276 592
use sky130_fd_sc_hd__or4_4  _1024_
timestamp 1606120353
transform 1 0 14444 0 1 54944
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__A
timestamp 1606120353
transform 1 0 14168 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_97_137
timestamp 1606120353
transform 1 0 13708 0 1 54944
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_97_141
timestamp 1606120353
transform 1 0 14076 0 1 54944
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_97_144
timestamp 1606120353
transform 1 0 14352 0 1 54944
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_97_154
timestamp 1606120353
transform 1 0 15272 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _1014_
timestamp 1606120353
transform 1 0 16008 0 1 54944
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__B
timestamp 1606120353
transform 1 0 17020 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__B
timestamp 1606120353
transform 1 0 15824 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__A
timestamp 1606120353
transform 1 0 15456 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_158
timestamp 1606120353
transform 1 0 15640 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_171
timestamp 1606120353
transform 1 0 16836 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_175
timestamp 1606120353
transform 1 0 17204 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0978_
timestamp 1606120353
transform 1 0 18032 0 1 54944
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_721
timestamp 1606120353
transform 1 0 17940 0 1 54944
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__B
timestamp 1606120353
transform 1 0 17756 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__A
timestamp 1606120353
transform 1 0 17388 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__D
timestamp 1606120353
transform 1 0 19044 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_179
timestamp 1606120353
transform 1 0 17572 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_193
timestamp 1606120353
transform 1 0 18860 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_197
timestamp 1606120353
transform 1 0 19228 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0966_
timestamp 1606120353
transform 1 0 20056 0 1 54944
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__B1
timestamp 1606120353
transform 1 0 21160 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__A
timestamp 1606120353
transform 1 0 19872 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__C
timestamp 1606120353
transform 1 0 19412 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_97_201
timestamp 1606120353
transform 1 0 19596 0 1 54944
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_97_215
timestamp 1606120353
transform 1 0 20884 0 1 54944
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_97_220
timestamp 1606120353
transform 1 0 21344 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__a21o_4  _0909_
timestamp 1606120353
transform 1 0 21712 0 1 54944
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__A
timestamp 1606120353
transform 1 0 21528 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__A2
timestamp 1606120353
transform 1 0 23368 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A1
timestamp 1606120353
transform 1 0 23000 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_236
timestamp 1606120353
transform 1 0 22816 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_240
timestamp 1606120353
transform 1 0 23184 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0925_
timestamp 1606120353
transform 1 0 24196 0 1 54944
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_722
timestamp 1606120353
transform 1 0 23552 0 1 54944
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__D
timestamp 1606120353
transform 1 0 23828 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_245
timestamp 1606120353
transform 1 0 23644 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_97_249
timestamp 1606120353
transform 1 0 24012 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_97_264
timestamp 1606120353
transform 1 0 25392 0 1 54944
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1185_
timestamp 1606120353
transform 1 0 26128 0 1 54944
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__D
timestamp 1606120353
transform 1 0 25944 0 1 54944
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1606120353
transform -1 0 28888 0 1 54944
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_97_291
timestamp 1606120353
transform 1 0 27876 0 1 54944
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1606120353
transform 1 0 1104 0 -1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_98_3
timestamp 1606120353
transform 1 0 1380 0 -1 56032
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_98_15
timestamp 1606120353
transform 1 0 2484 0 -1 56032
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_723
timestamp 1606120353
transform 1 0 3956 0 -1 56032
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_98_27
timestamp 1606120353
transform 1 0 3588 0 -1 56032
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_98_32
timestamp 1606120353
transform 1 0 4048 0 -1 56032
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_98_44
timestamp 1606120353
transform 1 0 5152 0 -1 56032
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_98_56
timestamp 1606120353
transform 1 0 6256 0 -1 56032
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_98_68
timestamp 1606120353
transform 1 0 7360 0 -1 56032
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_98_80
timestamp 1606120353
transform 1 0 8464 0 -1 56032
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1150_
timestamp 1606120353
transform 1 0 10488 0 -1 56032
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_724
timestamp 1606120353
transform 1 0 9568 0 -1 56032
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_98_93
timestamp 1606120353
transform 1 0 9660 0 -1 56032
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_98_101
timestamp 1606120353
transform 1 0 10396 0 -1 56032
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _1025_
timestamp 1606120353
transform 1 0 13156 0 -1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_98_121
timestamp 1606120353
transform 1 0 12236 0 -1 56032
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_98_129
timestamp 1606120353
transform 1 0 12972 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_134
timestamp 1606120353
transform 1 0 13432 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_138
timestamp 1606120353
transform 1 0 13800 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__A
timestamp 1606120353
transform 1 0 13616 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__A2
timestamp 1606120353
transform 1 0 13984 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0969_
timestamp 1606120353
transform 1 0 14168 0 -1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_98_145
timestamp 1606120353
transform 1 0 14444 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__C
timestamp 1606120353
transform 1 0 14628 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_149
timestamp 1606120353
transform 1 0 14812 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__A1
timestamp 1606120353
transform 1 0 14996 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_725
timestamp 1606120353
transform 1 0 15180 0 -1 56032
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_98_154
timestamp 1606120353
transform 1 0 15272 0 -1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__buf_1  _0977_
timestamp 1606120353
transform 1 0 15548 0 -1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__or4_4  _1000_
timestamp 1606120353
transform 1 0 16560 0 -1 56032
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__C
timestamp 1606120353
transform 1 0 16376 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__C
timestamp 1606120353
transform 1 0 16008 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_160
timestamp 1606120353
transform 1 0 15824 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_164
timestamp 1606120353
transform 1 0 16192 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _1052_
timestamp 1606120353
transform 1 0 18768 0 -1 56032
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A
timestamp 1606120353
transform 1 0 18032 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__B
timestamp 1606120353
transform 1 0 17572 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__B
timestamp 1606120353
transform 1 0 18400 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_177
timestamp 1606120353
transform 1 0 17388 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_98_181
timestamp 1606120353
transform 1 0 17756 0 -1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_98_186
timestamp 1606120353
transform 1 0 18216 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_190
timestamp 1606120353
transform 1 0 18584 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1001_
timestamp 1606120353
transform 1 0 20884 0 -1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_726
timestamp 1606120353
transform 1 0 20792 0 -1 56032
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__A1
timestamp 1606120353
transform 1 0 20056 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__A
timestamp 1606120353
transform 1 0 21344 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__B1
timestamp 1606120353
transform 1 0 20424 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_204
timestamp 1606120353
transform 1 0 19872 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_208
timestamp 1606120353
transform 1 0 20240 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_212
timestamp 1606120353
transform 1 0 20608 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_218
timestamp 1606120353
transform 1 0 21160 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__nor2_4  _0910_
timestamp 1606120353
transform 1 0 21896 0 -1 56032
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A2
timestamp 1606120353
transform 1 0 21712 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_clk_A
timestamp 1606120353
transform 1 0 22908 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__CLK
timestamp 1606120353
transform 1 0 23276 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_222
timestamp 1606120353
transform 1 0 21528 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_235
timestamp 1606120353
transform 1 0 22724 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_239
timestamp 1606120353
transform 1 0 23092 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1178_
timestamp 1606120353
transform 1 0 23460 0 -1 56032
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_8  FILLER_98_262
timestamp 1606120353
transform 1 0 25208 0 -1 56032
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_727
timestamp 1606120353
transform 1 0 26404 0 -1 56032
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__CLK
timestamp 1606120353
transform 1 0 26128 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_98_270
timestamp 1606120353
transform 1 0 25944 0 -1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_98_274
timestamp 1606120353
transform 1 0 26312 0 -1 56032
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_98_276
timestamp 1606120353
transform 1 0 26496 0 -1 56032
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1606120353
transform -1 0 28888 0 -1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_98_288
timestamp 1606120353
transform 1 0 27600 0 -1 56032
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_98_296
timestamp 1606120353
transform 1 0 28336 0 -1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1193_
timestamp 1606120353
transform 1 0 1380 0 -1 57120
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1606120353
transform 1 0 1104 0 1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1606120353
transform 1 0 1104 0 -1 57120
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__D
timestamp 1606120353
transform 1 0 1564 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__CLK
timestamp 1606120353
transform 1 0 1932 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_99_3
timestamp 1606120353
transform 1 0 1380 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_99_7
timestamp 1606120353
transform 1 0 1748 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_99_11
timestamp 1606120353
transform 1 0 2116 0 1 56032
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_100_22
timestamp 1606120353
transform 1 0 3128 0 -1 57120
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_732
timestamp 1606120353
transform 1 0 3956 0 -1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_99_23
timestamp 1606120353
transform 1 0 3220 0 1 56032
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_99_35
timestamp 1606120353
transform 1 0 4324 0 1 56032
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_100_30
timestamp 1606120353
transform 1 0 3864 0 -1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_100_32
timestamp 1606120353
transform 1 0 4048 0 -1 57120
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_100_44
timestamp 1606120353
transform 1 0 5152 0 -1 57120
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_728
timestamp 1606120353
transform 1 0 6716 0 1 56032
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1158__CLK
timestamp 1606120353
transform 1 0 6992 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_99_47
timestamp 1606120353
transform 1 0 5428 0 1 56032
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_99_59
timestamp 1606120353
transform 1 0 6532 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_99_62
timestamp 1606120353
transform 1 0 6808 0 1 56032
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_100_56
timestamp 1606120353
transform 1 0 6256 0 -1 57120
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_100_66
timestamp 1606120353
transform 1 0 7176 0 -1 57120
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_99_74
timestamp 1606120353
transform 1 0 7912 0 1 56032
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_99_86
timestamp 1606120353
transform 1 0 9016 0 1 56032
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_100_78
timestamp 1606120353
transform 1 0 8280 0 -1 57120
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_733
timestamp 1606120353
transform 1 0 9568 0 -1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_99_98
timestamp 1606120353
transform 1 0 10120 0 1 56032
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_99_110
timestamp 1606120353
transform 1 0 11224 0 1 56032
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_100_90
timestamp 1606120353
transform 1 0 9384 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_100_93
timestamp 1606120353
transform 1 0 9660 0 -1 57120
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_100_105
timestamp 1606120353
transform 1 0 10764 0 -1 57120
box 0 -48 1104 592
use sky130_fd_sc_hd__buf_1  _1015_
timestamp 1606120353
transform 1 0 13156 0 -1 57120
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_729
timestamp 1606120353
transform 1 0 12328 0 1 56032
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__A
timestamp 1606120353
transform 1 0 13156 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_99_123
timestamp 1606120353
transform 1 0 12420 0 1 56032
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_100_117
timestamp 1606120353
transform 1 0 11868 0 -1 57120
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_100_129
timestamp 1606120353
transform 1 0 12972 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_99_133
timestamp 1606120353
transform 1 0 13340 0 1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_100_134
timestamp 1606120353
transform 1 0 13432 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__A
timestamp 1606120353
transform 1 0 13616 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__B1
timestamp 1606120353
transform 1 0 13616 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_99_138
timestamp 1606120353
transform 1 0 13800 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_100_138
timestamp 1606120353
transform 1 0 13800 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__A
timestamp 1606120353
transform 1 0 13984 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__B1
timestamp 1606120353
transform 1 0 13984 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1006_
timestamp 1606120353
transform 1 0 14168 0 -1 57120
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_99_142
timestamp 1606120353
transform 1 0 14168 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_100_149
timestamp 1606120353
transform 1 0 14812 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_100_145
timestamp 1606120353
transform 1 0 14444 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__D
timestamp 1606120353
transform 1 0 14996 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__D
timestamp 1606120353
transform 1 0 14628 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__B
timestamp 1606120353
transform 1 0 14352 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_734
timestamp 1606120353
transform 1 0 15180 0 -1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__or4_4  _1021_
timestamp 1606120353
transform 1 0 14536 0 1 56032
box 0 -48 828 592
use sky130_fd_sc_hd__o21ai_4  _1063_
timestamp 1606120353
transform 1 0 15272 0 -1 57120
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_99_159
timestamp 1606120353
transform 1 0 15732 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_99_155
timestamp 1606120353
transform 1 0 15364 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__C
timestamp 1606120353
transform 1 0 15548 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__B
timestamp 1606120353
transform 1 0 15916 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _1005_
timestamp 1606120353
transform 1 0 16100 0 1 56032
box 0 -48 828 592
use sky130_fd_sc_hd__fill_1  FILLER_100_171
timestamp 1606120353
transform 1 0 16836 0 -1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_100_167
timestamp 1606120353
transform 1 0 16468 0 -1 57120
box 0 -48 368 592
use sky130_fd_sc_hd__decap_3  FILLER_99_172
timestamp 1606120353
transform 1 0 16928 0 1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A
timestamp 1606120353
transform 1 0 16928 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_100_174
timestamp 1606120353
transform 1 0 17112 0 -1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__A
timestamp 1606120353
transform 1 0 17204 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _1017_
timestamp 1606120353
transform 1 0 17204 0 -1 57120
box 0 -48 828 592
use sky130_fd_sc_hd__fill_2  FILLER_100_184
timestamp 1606120353
transform 1 0 18032 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_99_177
timestamp 1606120353
transform 1 0 17388 0 1 56032
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__A
timestamp 1606120353
transform 1 0 17756 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__C
timestamp 1606120353
transform 1 0 18216 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_730
timestamp 1606120353
transform 1 0 17940 0 1 56032
box 0 -48 92 592
use sky130_fd_sc_hd__or4_4  _0973_
timestamp 1606120353
transform 1 0 18032 0 1 56032
box 0 -48 828 592
use sky130_fd_sc_hd__fill_1  FILLER_100_192
timestamp 1606120353
transform 1 0 18768 0 -1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_100_188
timestamp 1606120353
transform 1 0 18400 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_99_197
timestamp 1606120353
transform 1 0 19228 0 1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_99_193
timestamp 1606120353
transform 1 0 18860 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__D
timestamp 1606120353
transform 1 0 18584 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__C
timestamp 1606120353
transform 1 0 19044 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1016_
timestamp 1606120353
transform 1 0 18860 0 -1 57120
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_100_206
timestamp 1606120353
transform 1 0 20056 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__A1
timestamp 1606120353
transform 1 0 20240 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__A1
timestamp 1606120353
transform 1 0 19504 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_clk
timestamp 1606120353
transform 1 0 19688 0 1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_100_218
timestamp 1606120353
transform 1 0 21160 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_100_210
timestamp 1606120353
transform 1 0 20424 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_99_218
timestamp 1606120353
transform 1 0 21160 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__A2
timestamp 1606120353
transform 1 0 21344 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__B1
timestamp 1606120353
transform 1 0 21344 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__A2
timestamp 1606120353
transform 1 0 20608 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_735
timestamp 1606120353
transform 1 0 20792 0 -1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__buf_1  _1043_
timestamp 1606120353
transform 1 0 20884 0 -1 57120
box 0 -48 276 592
use sky130_fd_sc_hd__o21ai_4  _1054_
timestamp 1606120353
transform 1 0 19964 0 1 56032
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_2  FILLER_100_226
timestamp 1606120353
transform 1 0 21896 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_100_222
timestamp 1606120353
transform 1 0 21528 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_99_229
timestamp 1606120353
transform 1 0 22172 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_99_222
timestamp 1606120353
transform 1 0 21528 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__A2
timestamp 1606120353
transform 1 0 22080 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__A2
timestamp 1606120353
transform 1 0 21712 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__A
timestamp 1606120353
transform 1 0 21712 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0965_
timestamp 1606120353
transform 1 0 21896 0 1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_100_234
timestamp 1606120353
transform 1 0 22632 0 -1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_100_230
timestamp 1606120353
transform 1 0 22264 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_99_237
timestamp 1606120353
transform 1 0 22908 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_99_233
timestamp 1606120353
transform 1 0 22540 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__B1
timestamp 1606120353
transform 1 0 22448 0 -1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A
timestamp 1606120353
transform 1 0 22356 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__A
timestamp 1606120353
transform 1 0 22724 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__inv_8  _0866_
timestamp 1606120353
transform 1 0 22724 0 -1 57120
box 0 -48 828 592
use sky130_fd_sc_hd__decap_3  FILLER_99_241
timestamp 1606120353
transform 1 0 23276 0 1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__B1
timestamp 1606120353
transform 1 0 23092 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_731
timestamp 1606120353
transform 1 0 23552 0 1 56032
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_99_245
timestamp 1606120353
transform 1 0 23644 0 1 56032
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_99_257
timestamp 1606120353
transform 1 0 24748 0 1 56032
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_100_244
timestamp 1606120353
transform 1 0 23552 0 -1 57120
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_100_256
timestamp 1606120353
transform 1 0 24656 0 -1 57120
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1195_
timestamp 1606120353
transform 1 0 26128 0 1 56032
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_736
timestamp 1606120353
transform 1 0 26404 0 -1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__D
timestamp 1606120353
transform 1 0 25944 0 1 56032
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_99_269
timestamp 1606120353
transform 1 0 25852 0 1 56032
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_100_268
timestamp 1606120353
transform 1 0 25760 0 -1 57120
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_100_274
timestamp 1606120353
transform 1 0 26312 0 -1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_100_276
timestamp 1606120353
transform 1 0 26496 0 -1 57120
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1606120353
transform -1 0 28888 0 1 56032
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1606120353
transform -1 0 28888 0 -1 57120
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_99_291
timestamp 1606120353
transform 1 0 27876 0 1 56032
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_100_288
timestamp 1606120353
transform 1 0 27600 0 -1 57120
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_100_296
timestamp 1606120353
transform 1 0 28336 0 -1 57120
box 0 -48 276 592
use sky130_fd_sc_hd__a21bo_4  _0935_
timestamp 1606120353
transform 1 0 2576 0 1 57120
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1606120353
transform 1 0 1104 0 1 57120
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__B1_N
timestamp 1606120353
transform 1 0 2392 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__A1
timestamp 1606120353
transform 1 0 2024 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_101_3
timestamp 1606120353
transform 1 0 1380 0 1 57120
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_101_9
timestamp 1606120353
transform 1 0 1932 0 1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_101_12
timestamp 1606120353
transform 1 0 2208 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_101_29
timestamp 1606120353
transform 1 0 3772 0 1 57120
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_101_41
timestamp 1606120353
transform 1 0 4876 0 1 57120
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1158_
timestamp 1606120353
transform 1 0 6992 0 1 57120
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_737
timestamp 1606120353
transform 1 0 6716 0 1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1158__D
timestamp 1606120353
transform 1 0 6532 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_101_53
timestamp 1606120353
transform 1 0 5980 0 1 57120
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_101_62
timestamp 1606120353
transform 1 0 6808 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_101_83
timestamp 1606120353
transform 1 0 8740 0 1 57120
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_101_95
timestamp 1606120353
transform 1 0 9844 0 1 57120
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_101_107
timestamp 1606120353
transform 1 0 10948 0 1 57120
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_738
timestamp 1606120353
transform 1 0 12328 0 1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_clk_A
timestamp 1606120353
transform 1 0 11960 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_101_115
timestamp 1606120353
transform 1 0 11684 0 1 57120
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_101_120
timestamp 1606120353
transform 1 0 12144 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_101_123
timestamp 1606120353
transform 1 0 12420 0 1 57120
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_101_131
timestamp 1606120353
transform 1 0 13156 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1059_
timestamp 1606120353
transform 1 0 13524 0 1 57120
box 0 -48 276 592
use sky130_fd_sc_hd__o21ai_4  _1069_
timestamp 1606120353
transform 1 0 14536 0 1 57120
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__A1
timestamp 1606120353
transform 1 0 14352 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__A1
timestamp 1606120353
transform 1 0 13984 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__A
timestamp 1606120353
transform 1 0 13340 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_101_138
timestamp 1606120353
transform 1 0 13800 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_101_142
timestamp 1606120353
transform 1 0 14168 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0974_
timestamp 1606120353
transform 1 0 16928 0 1 57120
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__D
timestamp 1606120353
transform 1 0 16744 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__A
timestamp 1606120353
transform 1 0 16100 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_101_159
timestamp 1606120353
transform 1 0 15732 0 1 57120
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_101_165
timestamp 1606120353
transform 1 0 16284 0 1 57120
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_101_169
timestamp 1606120353
transform 1 0 16652 0 1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_101_175
timestamp 1606120353
transform 1 0 17204 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__or4_4  _0982_
timestamp 1606120353
transform 1 0 18032 0 1 57120
box 0 -48 828 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_739
timestamp 1606120353
transform 1 0 17940 0 1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__B
timestamp 1606120353
transform 1 0 17388 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__C
timestamp 1606120353
transform 1 0 17756 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__D
timestamp 1606120353
transform 1 0 19044 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_101_179
timestamp 1606120353
transform 1 0 17572 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_101_193
timestamp 1606120353
transform 1 0 18860 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_101_197
timestamp 1606120353
transform 1 0 19228 0 1 57120
box 0 -48 276 592
use sky130_fd_sc_hd__o21ai_4  _1053_
timestamp 1606120353
transform 1 0 19688 0 1 57120
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__A1
timestamp 1606120353
transform 1 0 19504 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__A2
timestamp 1606120353
transform 1 0 21068 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_101_215
timestamp 1606120353
transform 1 0 20884 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_101_219
timestamp 1606120353
transform 1 0 21252 0 1 57120
box 0 -48 276 592
use sky130_fd_sc_hd__inv_8  _0861_
timestamp 1606120353
transform 1 0 21712 0 1 57120
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__A
timestamp 1606120353
transform 1 0 21528 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__B1
timestamp 1606120353
transform 1 0 23368 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__A1
timestamp 1606120353
transform 1 0 22724 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_101_233
timestamp 1606120353
transform 1 0 22540 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_101_237
timestamp 1606120353
transform 1 0 22908 0 1 57120
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_101_241
timestamp 1606120353
transform 1 0 23276 0 1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_740
timestamp 1606120353
transform 1 0 23552 0 1 57120
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A2
timestamp 1606120353
transform 1 0 23828 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A1
timestamp 1606120353
transform 1 0 24196 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_101_245
timestamp 1606120353
transform 1 0 23644 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_101_249
timestamp 1606120353
transform 1 0 24012 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_101_253
timestamp 1606120353
transform 1 0 24380 0 1 57120
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_101_265
timestamp 1606120353
transform 1 0 25484 0 1 57120
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_101_277
timestamp 1606120353
transform 1 0 26588 0 1 57120
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1606120353
transform -1 0 28888 0 1 57120
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_101_289
timestamp 1606120353
transform 1 0 27692 0 1 57120
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_101_297
timestamp 1606120353
transform 1 0 28428 0 1 57120
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1606120353
transform 1 0 1104 0 -1 58208
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__A2
timestamp 1606120353
transform 1 0 2576 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__CLK
timestamp 1606120353
transform 1 0 3128 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_102_3
timestamp 1606120353
transform 1 0 1380 0 -1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_102_15
timestamp 1606120353
transform 1 0 2484 0 -1 58208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_102_18
timestamp 1606120353
transform 1 0 2760 0 -1 58208
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_741
timestamp 1606120353
transform 1 0 3956 0 -1 58208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_102_24
timestamp 1606120353
transform 1 0 3312 0 -1 58208
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_102_30
timestamp 1606120353
transform 1 0 3864 0 -1 58208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_102_32
timestamp 1606120353
transform 1 0 4048 0 -1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_102_44
timestamp 1606120353
transform 1 0 5152 0 -1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_102_56
timestamp 1606120353
transform 1 0 6256 0 -1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_102_68
timestamp 1606120353
transform 1 0 7360 0 -1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_102_80
timestamp 1606120353
transform 1 0 8464 0 -1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_742
timestamp 1606120353
transform 1 0 9568 0 -1 58208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_102_93
timestamp 1606120353
transform 1 0 9660 0 -1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_102_105
timestamp 1606120353
transform 1 0 10764 0 -1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_clk
timestamp 1606120353
transform 1 0 11960 0 -1 58208
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_102_117
timestamp 1606120353
transform 1 0 11868 0 -1 58208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_102_121
timestamp 1606120353
transform 1 0 12236 0 -1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_102_137
timestamp 1606120353
transform 1 0 13708 0 -1 58208
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_102_133
timestamp 1606120353
transform 1 0 13340 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__B1
timestamp 1606120353
transform 1 0 13984 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__A
timestamp 1606120353
transform 1 0 13524 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _1022_
timestamp 1606120353
transform 1 0 14168 0 -1 58208
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_102_149
timestamp 1606120353
transform 1 0 14812 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_102_145
timestamp 1606120353
transform 1 0 14444 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__A2
timestamp 1606120353
transform 1 0 14996 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__A2
timestamp 1606120353
transform 1 0 14628 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_743
timestamp 1606120353
transform 1 0 15180 0 -1 58208
box 0 -48 92 592
use sky130_fd_sc_hd__o21ai_4  _1068_
timestamp 1606120353
transform 1 0 15272 0 -1 58208
box 0 -48 1196 592
use sky130_fd_sc_hd__or4_4  _0991_
timestamp 1606120353
transform 1 0 17204 0 -1 58208
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__A
timestamp 1606120353
transform 1 0 17020 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__B1
timestamp 1606120353
transform 1 0 16652 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_102_167
timestamp 1606120353
transform 1 0 16468 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_102_171
timestamp 1606120353
transform 1 0 16836 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _1013_
timestamp 1606120353
transform 1 0 18860 0 -1 58208
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__B
timestamp 1606120353
transform 1 0 18216 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A
timestamp 1606120353
transform 1 0 18584 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_102_184
timestamp 1606120353
transform 1 0 18032 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_102_188
timestamp 1606120353
transform 1 0 18400 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_102_192
timestamp 1606120353
transform 1 0 18768 0 -1 58208
box 0 -48 92 592
use sky130_fd_sc_hd__o21a_4  _1049_
timestamp 1606120353
transform 1 0 20884 0 -1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_744
timestamp 1606120353
transform 1 0 20792 0 -1 58208
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__A1
timestamp 1606120353
transform 1 0 20424 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_102_206
timestamp 1606120353
transform 1 0 20056 0 -1 58208
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_102_212
timestamp 1606120353
transform 1 0 20608 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__B1
timestamp 1606120353
transform 1 0 22172 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__A
timestamp 1606120353
transform 1 0 22540 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__B1
timestamp 1606120353
transform 1 0 22908 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__A
timestamp 1606120353
transform 1 0 23276 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_102_227
timestamp 1606120353
transform 1 0 21988 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_102_231
timestamp 1606120353
transform 1 0 22356 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_102_235
timestamp 1606120353
transform 1 0 22724 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_102_239
timestamp 1606120353
transform 1 0 23092 0 -1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _0868_
timestamp 1606120353
transform 1 0 23552 0 -1 58208
box 0 -48 1196 592
use sky130_fd_sc_hd__fill_1  FILLER_102_243
timestamp 1606120353
transform 1 0 23460 0 -1 58208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_102_257
timestamp 1606120353
transform 1 0 24748 0 -1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_745
timestamp 1606120353
transform 1 0 26404 0 -1 58208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_102_269
timestamp 1606120353
transform 1 0 25852 0 -1 58208
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_102_276
timestamp 1606120353
transform 1 0 26496 0 -1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1606120353
transform -1 0 28888 0 -1 58208
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_102_288
timestamp 1606120353
transform 1 0 27600 0 -1 58208
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_102_296
timestamp 1606120353
transform 1 0 28336 0 -1 58208
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1221_
timestamp 1606120353
transform 1 0 3128 0 1 58208
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1606120353
transform 1 0 1104 0 1 58208
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__D
timestamp 1606120353
transform 1 0 2944 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_103_3
timestamp 1606120353
transform 1 0 1380 0 1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_103_15
timestamp 1606120353
transform 1 0 2484 0 1 58208
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_103_19
timestamp 1606120353
transform 1 0 2852 0 1 58208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_103_41
timestamp 1606120353
transform 1 0 4876 0 1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_746
timestamp 1606120353
transform 1 0 6716 0 1 58208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_103_53
timestamp 1606120353
transform 1 0 5980 0 1 58208
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_103_62
timestamp 1606120353
transform 1 0 6808 0 1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_103_74
timestamp 1606120353
transform 1 0 7912 0 1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_103_86
timestamp 1606120353
transform 1 0 9016 0 1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_103_98
timestamp 1606120353
transform 1 0 10120 0 1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_103_110
timestamp 1606120353
transform 1 0 11224 0 1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_747
timestamp 1606120353
transform 1 0 12328 0 1 58208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_103_123
timestamp 1606120353
transform 1 0 12420 0 1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__buf_1  _1018_
timestamp 1606120353
transform 1 0 14260 0 1 58208
box 0 -48 276 592
use sky130_fd_sc_hd__o21ai_4  _1062_
timestamp 1606120353
transform 1 0 15272 0 1 58208
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__A1
timestamp 1606120353
transform 1 0 15088 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__A
timestamp 1606120353
transform 1 0 14720 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__A2
timestamp 1606120353
transform 1 0 14076 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_103_135
timestamp 1606120353
transform 1 0 13524 0 1 58208
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_103_146
timestamp 1606120353
transform 1 0 14536 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_103_150
timestamp 1606120353
transform 1 0 14904 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__A1
timestamp 1606120353
transform 1 0 16652 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__D
timestamp 1606120353
transform 1 0 17204 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_103_167
timestamp 1606120353
transform 1 0 16468 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_103_171
timestamp 1606120353
transform 1 0 16836 0 1 58208
box 0 -48 368 592
use sky130_fd_sc_hd__o21a_4  _0989_
timestamp 1606120353
transform 1 0 18584 0 1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_748
timestamp 1606120353
transform 1 0 17940 0 1 58208
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__A2
timestamp 1606120353
transform 1 0 18400 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__A1
timestamp 1606120353
transform 1 0 17756 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_103_177
timestamp 1606120353
transform 1 0 17388 0 1 58208
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_103_184
timestamp 1606120353
transform 1 0 18032 0 1 58208
box 0 -48 368 592
use sky130_fd_sc_hd__o21a_4  _1012_
timestamp 1606120353
transform 1 0 20424 0 1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__A2
timestamp 1606120353
transform 1 0 20240 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__B1
timestamp 1606120353
transform 1 0 19872 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_103_202
timestamp 1606120353
transform 1 0 19688 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_103_206
timestamp 1606120353
transform 1 0 20056 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_103_222
timestamp 1606120353
transform 1 0 21528 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__A2
timestamp 1606120353
transform 1 0 21712 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_103_226
timestamp 1606120353
transform 1 0 21896 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__A1
timestamp 1606120353
transform 1 0 22080 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0983_
timestamp 1606120353
transform 1 0 22264 0 1 58208
box 0 -48 276 592
use sky130_fd_sc_hd__decap_4  FILLER_103_233
timestamp 1606120353
transform 1 0 22540 0 1 58208
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_103_240
timestamp 1606120353
transform 1 0 23184 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_103_237
timestamp 1606120353
transform 1 0 22908 0 1 58208
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__A1
timestamp 1606120353
transform 1 0 23000 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__A2
timestamp 1606120353
transform 1 0 23368 0 1 58208
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0867_
timestamp 1606120353
transform 1 0 23644 0 1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_749
timestamp 1606120353
transform 1 0 23552 0 1 58208
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_103_257
timestamp 1606120353
transform 1 0 24748 0 1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_103_269
timestamp 1606120353
transform 1 0 25852 0 1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_103_281
timestamp 1606120353
transform 1 0 26956 0 1 58208
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1606120353
transform -1 0 28888 0 1 58208
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_103_293
timestamp 1606120353
transform 1 0 28060 0 1 58208
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1606120353
transform 1 0 1104 0 -1 59296
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_104_3
timestamp 1606120353
transform 1 0 1380 0 -1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_104_15
timestamp 1606120353
transform 1 0 2484 0 -1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_750
timestamp 1606120353
transform 1 0 3956 0 -1 59296
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_104_27
timestamp 1606120353
transform 1 0 3588 0 -1 59296
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_104_32
timestamp 1606120353
transform 1 0 4048 0 -1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_104_44
timestamp 1606120353
transform 1 0 5152 0 -1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_104_56
timestamp 1606120353
transform 1 0 6256 0 -1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_104_68
timestamp 1606120353
transform 1 0 7360 0 -1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_104_80
timestamp 1606120353
transform 1 0 8464 0 -1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_751
timestamp 1606120353
transform 1 0 9568 0 -1 59296
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_104_93
timestamp 1606120353
transform 1 0 9660 0 -1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_104_105
timestamp 1606120353
transform 1 0 10764 0 -1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_104_117
timestamp 1606120353
transform 1 0 11868 0 -1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_104_129
timestamp 1606120353
transform 1 0 12972 0 -1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_752
timestamp 1606120353
transform 1 0 15180 0 -1 59296
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__A2
timestamp 1606120353
transform 1 0 14996 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__B1
timestamp 1606120353
transform 1 0 14628 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_104_141
timestamp 1606120353
transform 1 0 14076 0 -1 59296
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_104_149
timestamp 1606120353
transform 1 0 14812 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_104_154
timestamp 1606120353
transform 1 0 15272 0 -1 59296
box 0 -48 368 592
use sky130_fd_sc_hd__o21ai_4  _1060_
timestamp 1606120353
transform 1 0 15824 0 -1 59296
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__A1
timestamp 1606120353
transform 1 0 17204 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__B1
timestamp 1606120353
transform 1 0 15640 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_104_173
timestamp 1606120353
transform 1 0 17020 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _1061_
timestamp 1606120353
transform 1 0 17756 0 -1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__A1
timestamp 1606120353
transform 1 0 19044 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__A2
timestamp 1606120353
transform 1 0 17572 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_104_177
timestamp 1606120353
transform 1 0 17388 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_104_193
timestamp 1606120353
transform 1 0 18860 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_104_197
timestamp 1606120353
transform 1 0 19228 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__A2
timestamp 1606120353
transform 1 0 19412 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__buf_1  _0992_
timestamp 1606120353
transform 1 0 19596 0 -1 59296
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_104_204
timestamp 1606120353
transform 1 0 19872 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__A
timestamp 1606120353
transform 1 0 20056 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_104_208
timestamp 1606120353
transform 1 0 20240 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__B1
timestamp 1606120353
transform 1 0 20424 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_104_212
timestamp 1606120353
transform 1 0 20608 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_104_215
timestamp 1606120353
transform 1 0 20884 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_753
timestamp 1606120353
transform 1 0 20792 0 -1 59296
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_104_219
timestamp 1606120353
transform 1 0 21252 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__B1
timestamp 1606120353
transform 1 0 21068 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _0862_
timestamp 1606120353
transform 1 0 21436 0 -1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__inv_8  _0864_
timestamp 1606120353
transform 1 0 23276 0 -1 59296
box 0 -48 828 592
use sky130_fd_sc_hd__decap_8  FILLER_104_233
timestamp 1606120353
transform 1 0 22540 0 -1 59296
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__B1
timestamp 1606120353
transform 1 0 24288 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_104_250
timestamp 1606120353
transform 1 0 24104 0 -1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_104_254
timestamp 1606120353
transform 1 0 24472 0 -1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_754
timestamp 1606120353
transform 1 0 26404 0 -1 59296
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_104_266
timestamp 1606120353
transform 1 0 25576 0 -1 59296
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_104_274
timestamp 1606120353
transform 1 0 26312 0 -1 59296
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_104_276
timestamp 1606120353
transform 1 0 26496 0 -1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1606120353
transform -1 0 28888 0 -1 59296
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_104_288
timestamp 1606120353
transform 1 0 27600 0 -1 59296
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_104_296
timestamp 1606120353
transform 1 0 28336 0 -1 59296
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1606120353
transform 1 0 1104 0 1 59296
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1606120353
transform 1 0 1104 0 -1 60384
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__D
timestamp 1606120353
transform 1 0 1564 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_105_3
timestamp 1606120353
transform 1 0 1380 0 1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_105_15
timestamp 1606120353
transform 1 0 2484 0 1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_106_3
timestamp 1606120353
transform 1 0 1380 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_106_7
timestamp 1606120353
transform 1 0 1748 0 -1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_106_19
timestamp 1606120353
transform 1 0 2852 0 -1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_759
timestamp 1606120353
transform 1 0 3956 0 -1 60384
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_105_27
timestamp 1606120353
transform 1 0 3588 0 1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_105_39
timestamp 1606120353
transform 1 0 4692 0 1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_106_32
timestamp 1606120353
transform 1 0 4048 0 -1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_106_44
timestamp 1606120353
transform 1 0 5152 0 -1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_755
timestamp 1606120353
transform 1 0 6716 0 1 59296
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_105_51
timestamp 1606120353
transform 1 0 5796 0 1 59296
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_105_59
timestamp 1606120353
transform 1 0 6532 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_105_62
timestamp 1606120353
transform 1 0 6808 0 1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_106_56
timestamp 1606120353
transform 1 0 6256 0 -1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_105_74
timestamp 1606120353
transform 1 0 7912 0 1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_105_86
timestamp 1606120353
transform 1 0 9016 0 1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_106_68
timestamp 1606120353
transform 1 0 7360 0 -1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_106_80
timestamp 1606120353
transform 1 0 8464 0 -1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_760
timestamp 1606120353
transform 1 0 9568 0 -1 60384
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_105_98
timestamp 1606120353
transform 1 0 10120 0 1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_105_110
timestamp 1606120353
transform 1 0 11224 0 1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_106_93
timestamp 1606120353
transform 1 0 9660 0 -1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_106_105
timestamp 1606120353
transform 1 0 10764 0 -1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_756
timestamp 1606120353
transform 1 0 12328 0 1 59296
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_105_123
timestamp 1606120353
transform 1 0 12420 0 1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_106_117
timestamp 1606120353
transform 1 0 11868 0 -1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_106_129
timestamp 1606120353
transform 1 0 12972 0 -1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_761
timestamp 1606120353
transform 1 0 15180 0 -1 60384
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__B1
timestamp 1606120353
transform 1 0 15180 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__B1
timestamp 1606120353
transform 1 0 14812 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_105_135
timestamp 1606120353
transform 1 0 13524 0 1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_105_147
timestamp 1606120353
transform 1 0 14628 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_105_151
timestamp 1606120353
transform 1 0 14996 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_106_141
timestamp 1606120353
transform 1 0 14076 0 -1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_106_154
timestamp 1606120353
transform 1 0 15272 0 -1 60384
box 0 -48 368 592
use sky130_fd_sc_hd__decap_4  FILLER_106_165
timestamp 1606120353
transform 1 0 16284 0 -1 60384
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_106_161
timestamp 1606120353
transform 1 0 15916 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_106_158
timestamp 1606120353
transform 1 0 15640 0 -1 60384
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_105_155
timestamp 1606120353
transform 1 0 15364 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__A1
timestamp 1606120353
transform 1 0 15732 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__A2
timestamp 1606120353
transform 1 0 15548 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__A2
timestamp 1606120353
transform 1 0 16100 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_105_175
timestamp 1606120353
transform 1 0 17204 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_105_171
timestamp 1606120353
transform 1 0 16836 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__A1
timestamp 1606120353
transform 1 0 16652 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__A2
timestamp 1606120353
transform 1 0 17020 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__o21a_4  _1067_
timestamp 1606120353
transform 1 0 15732 0 1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__o21a_4  _1057_
timestamp 1606120353
transform 1 0 16836 0 -1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_106_187
timestamp 1606120353
transform 1 0 18308 0 -1 60384
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_106_183
timestamp 1606120353
transform 1 0 17940 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_105_184
timestamp 1606120353
transform 1 0 18032 0 1 59296
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_105_179
timestamp 1606120353
transform 1 0 17572 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__B1
timestamp 1606120353
transform 1 0 17388 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__B1
timestamp 1606120353
transform 1 0 18124 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A2
timestamp 1606120353
transform 1 0 17756 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_757
timestamp 1606120353
transform 1 0 17940 0 1 59296
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_105_188
timestamp 1606120353
transform 1 0 18400 0 1 59296
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__B1
timestamp 1606120353
transform 1 0 18676 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A1
timestamp 1606120353
transform 1 0 18492 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _0990_
timestamp 1606120353
transform 1 0 18676 0 1 59296
box 0 -48 1196 592
use sky130_fd_sc_hd__o21ai_4  _0976_
timestamp 1606120353
transform 1 0 18860 0 -1 60384
box 0 -48 1196 592
use sky130_fd_sc_hd__o21ai_4  _0863_
timestamp 1606120353
transform 1 0 20700 0 1 59296
box 0 -48 1196 592
use sky130_fd_sc_hd__o21ai_4  _1051_
timestamp 1606120353
transform 1 0 20884 0 -1 60384
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_762
timestamp 1606120353
transform 1 0 20792 0 -1 60384
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A2
timestamp 1606120353
transform 1 0 20516 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A1
timestamp 1606120353
transform 1 0 20148 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__B1
timestamp 1606120353
transform 1 0 20608 0 -1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_105_204
timestamp 1606120353
transform 1 0 19872 0 1 59296
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_105_209
timestamp 1606120353
transform 1 0 20332 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_106_206
timestamp 1606120353
transform 1 0 20056 0 -1 60384
box 0 -48 552 592
use sky130_fd_sc_hd__inv_8  _0857_
timestamp 1606120353
transform 1 0 22816 0 -1 60384
box 0 -48 828 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__A1
timestamp 1606120353
transform 1 0 22080 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__A2
timestamp 1606120353
transform 1 0 22448 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__A
timestamp 1606120353
transform 1 0 22816 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_105_226
timestamp 1606120353
transform 1 0 21896 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_105_230
timestamp 1606120353
transform 1 0 22264 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_105_234
timestamp 1606120353
transform 1 0 22632 0 1 59296
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_105_238
timestamp 1606120353
transform 1 0 23000 0 1 59296
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILLER_106_228
timestamp 1606120353
transform 1 0 22080 0 -1 60384
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_758
timestamp 1606120353
transform 1 0 23552 0 1 59296
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_105_245
timestamp 1606120353
transform 1 0 23644 0 1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_105_257
timestamp 1606120353
transform 1 0 24748 0 1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_106_245
timestamp 1606120353
transform 1 0 23644 0 -1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_106_257
timestamp 1606120353
transform 1 0 24748 0 -1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_763
timestamp 1606120353
transform 1 0 26404 0 -1 60384
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_105_269
timestamp 1606120353
transform 1 0 25852 0 1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_105_281
timestamp 1606120353
transform 1 0 26956 0 1 59296
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_106_269
timestamp 1606120353
transform 1 0 25852 0 -1 60384
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_106_276
timestamp 1606120353
transform 1 0 26496 0 -1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1606120353
transform -1 0 28888 0 1 59296
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1606120353
transform -1 0 28888 0 -1 60384
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_105_293
timestamp 1606120353
transform 1 0 28060 0 1 59296
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILLER_106_288
timestamp 1606120353
transform 1 0 27600 0 -1 60384
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_106_296
timestamp 1606120353
transform 1 0 28336 0 -1 60384
box 0 -48 276 592
use sky130_fd_sc_hd__dfxtp_4  _1219_
timestamp 1606120353
transform 1 0 1380 0 1 60384
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1606120353
transform 1 0 1104 0 1 60384
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_107_22
timestamp 1606120353
transform 1 0 3128 0 1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_107_34
timestamp 1606120353
transform 1 0 4232 0 1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_764
timestamp 1606120353
transform 1 0 6716 0 1 60384
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_107_46
timestamp 1606120353
transform 1 0 5336 0 1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_107_58
timestamp 1606120353
transform 1 0 6440 0 1 60384
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_107_62
timestamp 1606120353
transform 1 0 6808 0 1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_107_74
timestamp 1606120353
transform 1 0 7912 0 1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_107_86
timestamp 1606120353
transform 1 0 9016 0 1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_107_98
timestamp 1606120353
transform 1 0 10120 0 1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_107_110
timestamp 1606120353
transform 1 0 11224 0 1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_765
timestamp 1606120353
transform 1 0 12328 0 1 60384
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_107_123
timestamp 1606120353
transform 1 0 12420 0 1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_107_135
timestamp 1606120353
transform 1 0 13524 0 1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_107_147
timestamp 1606120353
transform 1 0 14628 0 1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__o21a_4  _1019_
timestamp 1606120353
transform 1 0 16100 0 1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__A1
timestamp 1606120353
transform 1 0 15916 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_107_159
timestamp 1606120353
transform 1 0 15732 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_107_175
timestamp 1606120353
transform 1 0 17204 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__o21ai_4  _0993_
timestamp 1606120353
transform 1 0 18032 0 1 60384
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_766
timestamp 1606120353
transform 1 0 17940 0 1 60384
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__A1
timestamp 1606120353
transform 1 0 17756 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__A1
timestamp 1606120353
transform 1 0 17388 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_107_179
timestamp 1606120353
transform 1 0 17572 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_107_197
timestamp 1606120353
transform 1 0 19228 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__dfxtp_4  _1186_
timestamp 1606120353
transform 1 0 20608 0 1 60384
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__D
timestamp 1606120353
transform 1 0 20424 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__A
timestamp 1606120353
transform 1 0 19412 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_107_201
timestamp 1606120353
transform 1 0 19596 0 1 60384
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_107_209
timestamp 1606120353
transform 1 0 20332 0 1 60384
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__B1_N
timestamp 1606120353
transform 1 0 22540 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__A2
timestamp 1606120353
transform 1 0 22908 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_107_231
timestamp 1606120353
transform 1 0 22356 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_107_235
timestamp 1606120353
transform 1 0 22724 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_107_239
timestamp 1606120353
transform 1 0 23092 0 1 60384
box 0 -48 368 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_767
timestamp 1606120353
transform 1 0 23552 0 1 60384
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_107_243
timestamp 1606120353
transform 1 0 23460 0 1 60384
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_107_245
timestamp 1606120353
transform 1 0 23644 0 1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_107_257
timestamp 1606120353
transform 1 0 24748 0 1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__B1_N
timestamp 1606120353
transform 1 0 26496 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__A2
timestamp 1606120353
transform 1 0 26864 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__A1
timestamp 1606120353
transform 1 0 27232 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_107_269
timestamp 1606120353
transform 1 0 25852 0 1 60384
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_107_275
timestamp 1606120353
transform 1 0 26404 0 1 60384
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_107_278
timestamp 1606120353
transform 1 0 26680 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_107_282
timestamp 1606120353
transform 1 0 27048 0 1 60384
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_107_286
timestamp 1606120353
transform 1 0 27416 0 1 60384
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1606120353
transform -1 0 28888 0 1 60384
box 0 -48 276 592
use sky130_fd_sc_hd__fill_1  FILLER_107_298
timestamp 1606120353
transform 1 0 28520 0 1 60384
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1606120353
transform 1 0 1104 0 -1 61472
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__CLK
timestamp 1606120353
transform 1 0 1564 0 -1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_108_3
timestamp 1606120353
transform 1 0 1380 0 -1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_108_7
timestamp 1606120353
transform 1 0 1748 0 -1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_108_19
timestamp 1606120353
transform 1 0 2852 0 -1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_768
timestamp 1606120353
transform 1 0 3956 0 -1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_108_32
timestamp 1606120353
transform 1 0 4048 0 -1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_108_44
timestamp 1606120353
transform 1 0 5152 0 -1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_108_56
timestamp 1606120353
transform 1 0 6256 0 -1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_108_68
timestamp 1606120353
transform 1 0 7360 0 -1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_108_80
timestamp 1606120353
transform 1 0 8464 0 -1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_769
timestamp 1606120353
transform 1 0 9568 0 -1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_108_93
timestamp 1606120353
transform 1 0 9660 0 -1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_108_105
timestamp 1606120353
transform 1 0 10764 0 -1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__CLK
timestamp 1606120353
transform 1 0 12420 0 -1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_108_117
timestamp 1606120353
transform 1 0 11868 0 -1 61472
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_108_125
timestamp 1606120353
transform 1 0 12604 0 -1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_770
timestamp 1606120353
transform 1 0 15180 0 -1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_108_137
timestamp 1606120353
transform 1 0 13708 0 -1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_108_149
timestamp 1606120353
transform 1 0 14812 0 -1 61472
box 0 -48 368 592
use sky130_fd_sc_hd__decap_8  FILLER_108_154
timestamp 1606120353
transform 1 0 15272 0 -1 61472
box 0 -48 736 592
use sky130_fd_sc_hd__o21ai_4  _1058_
timestamp 1606120353
transform 1 0 17204 0 -1 61472
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__B1
timestamp 1606120353
transform 1 0 16100 0 -1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__A2
timestamp 1606120353
transform 1 0 17020 0 -1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_108_162
timestamp 1606120353
transform 1 0 16008 0 -1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_108_165
timestamp 1606120353
transform 1 0 16284 0 -1 61472
box 0 -48 736 592
use sky130_fd_sc_hd__buf_1  _0985_
timestamp 1606120353
transform 1 0 19136 0 -1 61472
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__A2
timestamp 1606120353
transform 1 0 18584 0 -1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__A2
timestamp 1606120353
transform 1 0 18952 0 -1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_108_188
timestamp 1606120353
transform 1 0 18400 0 -1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_108_192
timestamp 1606120353
transform 1 0 18768 0 -1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__a21bo_4  _0927_
timestamp 1606120353
transform 1 0 21252 0 -1 61472
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_771
timestamp 1606120353
transform 1 0 20792 0 -1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__A1
timestamp 1606120353
transform 1 0 21068 0 -1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__CLK
timestamp 1606120353
transform 1 0 20608 0 -1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_108_199
timestamp 1606120353
transform 1 0 19412 0 -1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_108_211
timestamp 1606120353
transform 1 0 20516 0 -1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_108_215
timestamp 1606120353
transform 1 0 20884 0 -1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_108_232
timestamp 1606120353
transform 1 0 22448 0 -1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_108_244
timestamp 1606120353
transform 1 0 23552 0 -1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_108_256
timestamp 1606120353
transform 1 0 24656 0 -1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__a21bo_4  _0928_
timestamp 1606120353
transform 1 0 26496 0 -1 61472
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_772
timestamp 1606120353
transform 1 0 26404 0 -1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__CLK
timestamp 1606120353
transform 1 0 26128 0 -1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_108_268
timestamp 1606120353
transform 1 0 25760 0 -1 61472
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_108_274
timestamp 1606120353
transform 1 0 26312 0 -1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1606120353
transform -1 0 28888 0 -1 61472
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_108_289
timestamp 1606120353
transform 1 0 27692 0 -1 61472
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_108_297
timestamp 1606120353
transform 1 0 28428 0 -1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1606120353
transform 1 0 1104 0 1 61472
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_109_3
timestamp 1606120353
transform 1 0 1380 0 1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_109_15
timestamp 1606120353
transform 1 0 2484 0 1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_109_27
timestamp 1606120353
transform 1 0 3588 0 1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_109_39
timestamp 1606120353
transform 1 0 4692 0 1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_773
timestamp 1606120353
transform 1 0 6716 0 1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_109_51
timestamp 1606120353
transform 1 0 5796 0 1 61472
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_109_59
timestamp 1606120353
transform 1 0 6532 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_109_62
timestamp 1606120353
transform 1 0 6808 0 1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_109_74
timestamp 1606120353
transform 1 0 7912 0 1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_109_86
timestamp 1606120353
transform 1 0 9016 0 1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_109_98
timestamp 1606120353
transform 1 0 10120 0 1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_109_110
timestamp 1606120353
transform 1 0 11224 0 1 61472
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1213_
timestamp 1606120353
transform 1 0 12420 0 1 61472
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_774
timestamp 1606120353
transform 1 0 12328 0 1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__D
timestamp 1606120353
transform 1 0 12144 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_109_118
timestamp 1606120353
transform 1 0 11960 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_109_142
timestamp 1606120353
transform 1 0 14168 0 1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_109_154
timestamp 1606120353
transform 1 0 15272 0 1 61472
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__A1
timestamp 1606120353
transform 1 0 15916 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__A2
timestamp 1606120353
transform 1 0 16284 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__B1
timestamp 1606120353
transform 1 0 17204 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__B1
timestamp 1606120353
transform 1 0 16652 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_109_160
timestamp 1606120353
transform 1 0 15824 0 1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_109_163
timestamp 1606120353
transform 1 0 16100 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_109_167
timestamp 1606120353
transform 1 0 16468 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_109_171
timestamp 1606120353
transform 1 0 16836 0 1 61472
box 0 -48 368 592
use sky130_fd_sc_hd__o21ai_4  _1050_
timestamp 1606120353
transform 1 0 18952 0 1 61472
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_775
timestamp 1606120353
transform 1 0 17940 0 1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__A1
timestamp 1606120353
transform 1 0 18768 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_109_177
timestamp 1606120353
transform 1 0 17388 0 1 61472
box 0 -48 552 592
use sky130_fd_sc_hd__decap_8  FILLER_109_184
timestamp 1606120353
transform 1 0 18032 0 1 61472
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_109_207
timestamp 1606120353
transform 1 0 20148 0 1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_109_219
timestamp 1606120353
transform 1 0 21252 0 1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_109_231
timestamp 1606120353
transform 1 0 22356 0 1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_776
timestamp 1606120353
transform 1 0 23552 0 1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_109_243
timestamp 1606120353
transform 1 0 23460 0 1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_109_245
timestamp 1606120353
transform 1 0 23644 0 1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_109_257
timestamp 1606120353
transform 1 0 24748 0 1 61472
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1225_
timestamp 1606120353
transform 1 0 26128 0 1 61472
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__D
timestamp 1606120353
transform 1 0 25944 0 1 61472
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_109_269
timestamp 1606120353
transform 1 0 25852 0 1 61472
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1606120353
transform -1 0 28888 0 1 61472
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_109_291
timestamp 1606120353
transform 1 0 27876 0 1 61472
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1606120353
transform 1 0 1104 0 -1 62560
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_110_3
timestamp 1606120353
transform 1 0 1380 0 -1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_110_15
timestamp 1606120353
transform 1 0 2484 0 -1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_777
timestamp 1606120353
transform 1 0 3956 0 -1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_110_27
timestamp 1606120353
transform 1 0 3588 0 -1 62560
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_110_32
timestamp 1606120353
transform 1 0 4048 0 -1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_110_44
timestamp 1606120353
transform 1 0 5152 0 -1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_110_56
timestamp 1606120353
transform 1 0 6256 0 -1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_110_68
timestamp 1606120353
transform 1 0 7360 0 -1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_110_80
timestamp 1606120353
transform 1 0 8464 0 -1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_778
timestamp 1606120353
transform 1 0 9568 0 -1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_110_93
timestamp 1606120353
transform 1 0 9660 0 -1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_110_105
timestamp 1606120353
transform 1 0 10764 0 -1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_110_117
timestamp 1606120353
transform 1 0 11868 0 -1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_110_129
timestamp 1606120353
transform 1 0 12972 0 -1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_779
timestamp 1606120353
transform 1 0 15180 0 -1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_110_141
timestamp 1606120353
transform 1 0 14076 0 -1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_110_154
timestamp 1606120353
transform 1 0 15272 0 -1 62560
box 0 -48 552 592
use sky130_fd_sc_hd__o21a_4  _1071_
timestamp 1606120353
transform 1 0 15916 0 -1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_110_160
timestamp 1606120353
transform 1 0 15824 0 -1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_110_173
timestamp 1606120353
transform 1 0 17020 0 -1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__B1
timestamp 1606120353
transform 1 0 18952 0 -1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_110_185
timestamp 1606120353
transform 1 0 18124 0 -1 62560
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_110_193
timestamp 1606120353
transform 1 0 18860 0 -1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_110_196
timestamp 1606120353
transform 1 0 19136 0 -1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_780
timestamp 1606120353
transform 1 0 20792 0 -1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_110_208
timestamp 1606120353
transform 1 0 20240 0 -1 62560
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_110_215
timestamp 1606120353
transform 1 0 20884 0 -1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_110_227
timestamp 1606120353
transform 1 0 21988 0 -1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_110_239
timestamp 1606120353
transform 1 0 23092 0 -1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_110_251
timestamp 1606120353
transform 1 0 24196 0 -1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_110_263
timestamp 1606120353
transform 1 0 25300 0 -1 62560
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_781
timestamp 1606120353
transform 1 0 26404 0 -1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__CLK
timestamp 1606120353
transform 1 0 26128 0 -1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_110_271
timestamp 1606120353
transform 1 0 26036 0 -1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_110_274
timestamp 1606120353
transform 1 0 26312 0 -1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_110_276
timestamp 1606120353
transform 1 0 26496 0 -1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1606120353
transform -1 0 28888 0 -1 62560
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_110_288
timestamp 1606120353
transform 1 0 27600 0 -1 62560
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_110_296
timestamp 1606120353
transform 1 0 28336 0 -1 62560
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1606120353
transform 1 0 1104 0 1 62560
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_111_3
timestamp 1606120353
transform 1 0 1380 0 1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_111_15
timestamp 1606120353
transform 1 0 2484 0 1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_111_27
timestamp 1606120353
transform 1 0 3588 0 1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_111_39
timestamp 1606120353
transform 1 0 4692 0 1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_782
timestamp 1606120353
transform 1 0 6716 0 1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_111_51
timestamp 1606120353
transform 1 0 5796 0 1 62560
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_111_59
timestamp 1606120353
transform 1 0 6532 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_111_62
timestamp 1606120353
transform 1 0 6808 0 1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_111_74
timestamp 1606120353
transform 1 0 7912 0 1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_111_86
timestamp 1606120353
transform 1 0 9016 0 1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_111_98
timestamp 1606120353
transform 1 0 10120 0 1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_111_110
timestamp 1606120353
transform 1 0 11224 0 1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_783
timestamp 1606120353
transform 1 0 12328 0 1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_111_123
timestamp 1606120353
transform 1 0 12420 0 1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__A1
timestamp 1606120353
transform 1 0 15272 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_111_135
timestamp 1606120353
transform 1 0 13524 0 1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_111_147
timestamp 1606120353
transform 1 0 14628 0 1 62560
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_111_153
timestamp 1606120353
transform 1 0 15180 0 1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__A2
timestamp 1606120353
transform 1 0 15640 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__B1
timestamp 1606120353
transform 1 0 16008 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_111_156
timestamp 1606120353
transform 1 0 15456 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_111_160
timestamp 1606120353
transform 1 0 15824 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_111_164
timestamp 1606120353
transform 1 0 16192 0 1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_111_176
timestamp 1606120353
transform 1 0 17296 0 1 62560
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_784
timestamp 1606120353
transform 1 0 17940 0 1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_111_182
timestamp 1606120353
transform 1 0 17848 0 1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_111_184
timestamp 1606120353
transform 1 0 18032 0 1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_111_196
timestamp 1606120353
transform 1 0 19136 0 1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_111_208
timestamp 1606120353
transform 1 0 20240 0 1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_111_220
timestamp 1606120353
transform 1 0 21344 0 1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A1
timestamp 1606120353
transform 1 0 23368 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_111_232
timestamp 1606120353
transform 1 0 22448 0 1 62560
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_111_240
timestamp 1606120353
transform 1 0 23184 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_785
timestamp 1606120353
transform 1 0 23552 0 1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__B1_N
timestamp 1606120353
transform 1 0 23828 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A2
timestamp 1606120353
transform 1 0 24196 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_111_245
timestamp 1606120353
transform 1 0 23644 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_111_249
timestamp 1606120353
transform 1 0 24012 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_111_253
timestamp 1606120353
transform 1 0 24380 0 1 62560
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1187_
timestamp 1606120353
transform 1 0 26128 0 1 62560
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__D
timestamp 1606120353
transform 1 0 25944 0 1 62560
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_111_265
timestamp 1606120353
transform 1 0 25484 0 1 62560
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_111_269
timestamp 1606120353
transform 1 0 25852 0 1 62560
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1606120353
transform -1 0 28888 0 1 62560
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_111_291
timestamp 1606120353
transform 1 0 27876 0 1 62560
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1606120353
transform 1 0 1104 0 -1 63648
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1606120353
transform 1 0 1104 0 1 63648
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_112_3
timestamp 1606120353
transform 1 0 1380 0 -1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_112_15
timestamp 1606120353
transform 1 0 2484 0 -1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_113_3
timestamp 1606120353
transform 1 0 1380 0 1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_113_15
timestamp 1606120353
transform 1 0 2484 0 1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_786
timestamp 1606120353
transform 1 0 3956 0 -1 63648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_112_27
timestamp 1606120353
transform 1 0 3588 0 -1 63648
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_112_32
timestamp 1606120353
transform 1 0 4048 0 -1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_112_44
timestamp 1606120353
transform 1 0 5152 0 -1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_113_27
timestamp 1606120353
transform 1 0 3588 0 1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_113_39
timestamp 1606120353
transform 1 0 4692 0 1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_791
timestamp 1606120353
transform 1 0 6716 0 1 63648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_112_56
timestamp 1606120353
transform 1 0 6256 0 -1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_113_51
timestamp 1606120353
transform 1 0 5796 0 1 63648
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_113_59
timestamp 1606120353
transform 1 0 6532 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_113_62
timestamp 1606120353
transform 1 0 6808 0 1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_112_68
timestamp 1606120353
transform 1 0 7360 0 -1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_112_80
timestamp 1606120353
transform 1 0 8464 0 -1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_113_74
timestamp 1606120353
transform 1 0 7912 0 1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_113_86
timestamp 1606120353
transform 1 0 9016 0 1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_787
timestamp 1606120353
transform 1 0 9568 0 -1 63648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_112_93
timestamp 1606120353
transform 1 0 9660 0 -1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_112_105
timestamp 1606120353
transform 1 0 10764 0 -1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_113_98
timestamp 1606120353
transform 1 0 10120 0 1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_113_110
timestamp 1606120353
transform 1 0 11224 0 1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_792
timestamp 1606120353
transform 1 0 12328 0 1 63648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_112_117
timestamp 1606120353
transform 1 0 11868 0 -1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_112_129
timestamp 1606120353
transform 1 0 12972 0 -1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_113_123
timestamp 1606120353
transform 1 0 12420 0 1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__o21ai_4  _1077_
timestamp 1606120353
transform 1 0 15272 0 -1 63648
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_788
timestamp 1606120353
transform 1 0 15180 0 -1 63648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_112_141
timestamp 1606120353
transform 1 0 14076 0 -1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_113_135
timestamp 1606120353
transform 1 0 13524 0 1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_113_147
timestamp 1606120353
transform 1 0 14628 0 1 63648
box 0 -48 736 592
use sky130_fd_sc_hd__o21ai_4  _1078_
timestamp 1606120353
transform 1 0 15916 0 1 63648
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__A1
timestamp 1606120353
transform 1 0 15732 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__B1
timestamp 1606120353
transform 1 0 15364 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_112_167
timestamp 1606120353
transform 1 0 16468 0 -1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_113_157
timestamp 1606120353
transform 1 0 15548 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_113_174
timestamp 1606120353
transform 1 0 17112 0 1 63648
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1181_
timestamp 1606120353
transform 1 0 18768 0 1 63648
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_793
timestamp 1606120353
transform 1 0 17940 0 1 63648
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1181__D
timestamp 1606120353
transform 1 0 18584 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1181__CLK
timestamp 1606120353
transform 1 0 18768 0 -1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_112_179
timestamp 1606120353
transform 1 0 17572 0 -1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_112_191
timestamp 1606120353
transform 1 0 18676 0 -1 63648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_112_194
timestamp 1606120353
transform 1 0 18952 0 -1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_113_182
timestamp 1606120353
transform 1 0 17848 0 1 63648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_113_184
timestamp 1606120353
transform 1 0 18032 0 1 63648
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_789
timestamp 1606120353
transform 1 0 20792 0 -1 63648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_112_206
timestamp 1606120353
transform 1 0 20056 0 -1 63648
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_112_215
timestamp 1606120353
transform 1 0 20884 0 -1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_113_211
timestamp 1606120353
transform 1 0 20516 0 1 63648
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_113_219
timestamp 1606120353
transform 1 0 21252 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__D
timestamp 1606120353
transform 1 0 21436 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__CLK
timestamp 1606120353
transform 1 0 21804 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_112_227
timestamp 1606120353
transform 1 0 21988 0 -1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_112_239
timestamp 1606120353
transform 1 0 23092 0 -1 63648
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_113_223
timestamp 1606120353
transform 1 0 21620 0 1 63648
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_113_227
timestamp 1606120353
transform 1 0 21988 0 1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_113_239
timestamp 1606120353
transform 1 0 23092 0 1 63648
box 0 -48 368 592
use sky130_fd_sc_hd__a21bo_4  _0933_
timestamp 1606120353
transform 1 0 23460 0 -1 63648
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_794
timestamp 1606120353
transform 1 0 23552 0 1 63648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_112_256
timestamp 1606120353
transform 1 0 24656 0 -1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_113_243
timestamp 1606120353
transform 1 0 23460 0 1 63648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_113_245
timestamp 1606120353
transform 1 0 23644 0 1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_113_257
timestamp 1606120353
transform 1 0 24748 0 1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_790
timestamp 1606120353
transform 1 0 26404 0 -1 63648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_112_268
timestamp 1606120353
transform 1 0 25760 0 -1 63648
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_112_274
timestamp 1606120353
transform 1 0 26312 0 -1 63648
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_112_276
timestamp 1606120353
transform 1 0 26496 0 -1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_113_269
timestamp 1606120353
transform 1 0 25852 0 1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_113_281
timestamp 1606120353
transform 1 0 26956 0 1 63648
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1606120353
transform -1 0 28888 0 -1 63648
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1606120353
transform -1 0 28888 0 1 63648
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_112_288
timestamp 1606120353
transform 1 0 27600 0 -1 63648
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_112_296
timestamp 1606120353
transform 1 0 28336 0 -1 63648
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_113_293
timestamp 1606120353
transform 1 0 28060 0 1 63648
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1606120353
transform 1 0 1104 0 -1 64736
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_114_3
timestamp 1606120353
transform 1 0 1380 0 -1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_114_15
timestamp 1606120353
transform 1 0 2484 0 -1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_795
timestamp 1606120353
transform 1 0 3956 0 -1 64736
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_114_27
timestamp 1606120353
transform 1 0 3588 0 -1 64736
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_114_32
timestamp 1606120353
transform 1 0 4048 0 -1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_114_44
timestamp 1606120353
transform 1 0 5152 0 -1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_114_56
timestamp 1606120353
transform 1 0 6256 0 -1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_114_68
timestamp 1606120353
transform 1 0 7360 0 -1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_114_80
timestamp 1606120353
transform 1 0 8464 0 -1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_796
timestamp 1606120353
transform 1 0 9568 0 -1 64736
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_114_93
timestamp 1606120353
transform 1 0 9660 0 -1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_114_105
timestamp 1606120353
transform 1 0 10764 0 -1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_114_117
timestamp 1606120353
transform 1 0 11868 0 -1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_114_129
timestamp 1606120353
transform 1 0 12972 0 -1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_797
timestamp 1606120353
transform 1 0 15180 0 -1 64736
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__B1
timestamp 1606120353
transform 1 0 14996 0 -1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_114_141
timestamp 1606120353
transform 1 0 14076 0 -1 64736
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_114_149
timestamp 1606120353
transform 1 0 14812 0 -1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_114_154
timestamp 1606120353
transform 1 0 15272 0 -1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__A2
timestamp 1606120353
transform 1 0 15916 0 -1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__A2
timestamp 1606120353
transform 1 0 15456 0 -1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_114_158
timestamp 1606120353
transform 1 0 15640 0 -1 64736
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_114_163
timestamp 1606120353
transform 1 0 16100 0 -1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_114_175
timestamp 1606120353
transform 1 0 17204 0 -1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_114_187
timestamp 1606120353
transform 1 0 18308 0 -1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_798
timestamp 1606120353
transform 1 0 20792 0 -1 64736
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_114_199
timestamp 1606120353
transform 1 0 19412 0 -1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_114_211
timestamp 1606120353
transform 1 0 20516 0 -1 64736
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_114_215
timestamp 1606120353
transform 1 0 20884 0 -1 64736
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1191_
timestamp 1606120353
transform 1 0 21436 0 -1 64736
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_12  FILLER_114_240
timestamp 1606120353
transform 1 0 23184 0 -1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_114_252
timestamp 1606120353
transform 1 0 24288 0 -1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_114_264
timestamp 1606120353
transform 1 0 25392 0 -1 64736
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_799
timestamp 1606120353
transform 1 0 26404 0 -1 64736
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_114_272
timestamp 1606120353
transform 1 0 26128 0 -1 64736
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_114_276
timestamp 1606120353
transform 1 0 26496 0 -1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1606120353
transform -1 0 28888 0 -1 64736
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_114_288
timestamp 1606120353
transform 1 0 27600 0 -1 64736
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_114_296
timestamp 1606120353
transform 1 0 28336 0 -1 64736
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_230
timestamp 1606120353
transform 1 0 1104 0 1 64736
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_115_3
timestamp 1606120353
transform 1 0 1380 0 1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_115_15
timestamp 1606120353
transform 1 0 2484 0 1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_115_27
timestamp 1606120353
transform 1 0 3588 0 1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_115_39
timestamp 1606120353
transform 1 0 4692 0 1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_800
timestamp 1606120353
transform 1 0 6716 0 1 64736
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_115_51
timestamp 1606120353
transform 1 0 5796 0 1 64736
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_115_59
timestamp 1606120353
transform 1 0 6532 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_115_62
timestamp 1606120353
transform 1 0 6808 0 1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_115_74
timestamp 1606120353
transform 1 0 7912 0 1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_115_86
timestamp 1606120353
transform 1 0 9016 0 1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_115_98
timestamp 1606120353
transform 1 0 10120 0 1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_115_110
timestamp 1606120353
transform 1 0 11224 0 1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_801
timestamp 1606120353
transform 1 0 12328 0 1 64736
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_115_123
timestamp 1606120353
transform 1 0 12420 0 1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__o21ai_4  _1072_
timestamp 1606120353
transform 1 0 15180 0 1 64736
box 0 -48 1196 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__A1
timestamp 1606120353
transform 1 0 14996 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__A1
timestamp 1606120353
transform 1 0 14628 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__A2
timestamp 1606120353
transform 1 0 14260 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_115_135
timestamp 1606120353
transform 1 0 13524 0 1 64736
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_115_145
timestamp 1606120353
transform 1 0 14444 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_115_149
timestamp 1606120353
transform 1 0 14812 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__A2
timestamp 1606120353
transform 1 0 17112 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__B1
timestamp 1606120353
transform 1 0 16560 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_115_166
timestamp 1606120353
transform 1 0 16376 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_115_170
timestamp 1606120353
transform 1 0 16744 0 1 64736
box 0 -48 368 592
use sky130_fd_sc_hd__fill_2  FILLER_115_176
timestamp 1606120353
transform 1 0 17296 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_802
timestamp 1606120353
transform 1 0 17940 0 1 64736
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__A1
timestamp 1606120353
transform 1 0 17480 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__B1
timestamp 1606120353
transform 1 0 18216 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_115_180
timestamp 1606120353
transform 1 0 17664 0 1 64736
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_115_184
timestamp 1606120353
transform 1 0 18032 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_115_188
timestamp 1606120353
transform 1 0 18400 0 1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_115_200
timestamp 1606120353
transform 1 0 19504 0 1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_115_212
timestamp 1606120353
transform 1 0 20608 0 1 64736
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_115_220
timestamp 1606120353
transform 1 0 21344 0 1 64736
box 0 -48 276 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_clk
timestamp 1606120353
transform 1 0 21620 0 1 64736
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_clk_A
timestamp 1606120353
transform 1 0 22080 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_115_226
timestamp 1606120353
transform 1 0 21896 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_115_230
timestamp 1606120353
transform 1 0 22264 0 1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_115_242
timestamp 1606120353
transform 1 0 23368 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_803
timestamp 1606120353
transform 1 0 23552 0 1 64736
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_clk
timestamp 1606120353
transform 1 0 24380 0 1 64736
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_clk_A
timestamp 1606120353
transform 1 0 24840 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_115_245
timestamp 1606120353
transform 1 0 23644 0 1 64736
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_115_256
timestamp 1606120353
transform 1 0 24656 0 1 64736
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_115_260
timestamp 1606120353
transform 1 0 25024 0 1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_115_272
timestamp 1606120353
transform 1 0 26128 0 1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_115_284
timestamp 1606120353
transform 1 0 27232 0 1 64736
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_231
timestamp 1606120353
transform -1 0 28888 0 1 64736
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_115_296
timestamp 1606120353
transform 1 0 28336 0 1 64736
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_232
timestamp 1606120353
transform 1 0 1104 0 -1 65824
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_116_3
timestamp 1606120353
transform 1 0 1380 0 -1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_116_15
timestamp 1606120353
transform 1 0 2484 0 -1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_804
timestamp 1606120353
transform 1 0 3956 0 -1 65824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_116_27
timestamp 1606120353
transform 1 0 3588 0 -1 65824
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_116_32
timestamp 1606120353
transform 1 0 4048 0 -1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_116_44
timestamp 1606120353
transform 1 0 5152 0 -1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_116_56
timestamp 1606120353
transform 1 0 6256 0 -1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_116_68
timestamp 1606120353
transform 1 0 7360 0 -1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_116_80
timestamp 1606120353
transform 1 0 8464 0 -1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_805
timestamp 1606120353
transform 1 0 9568 0 -1 65824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_116_93
timestamp 1606120353
transform 1 0 9660 0 -1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_116_105
timestamp 1606120353
transform 1 0 10764 0 -1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_116_117
timestamp 1606120353
transform 1 0 11868 0 -1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_116_129
timestamp 1606120353
transform 1 0 12972 0 -1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__o21ai_4  _1073_
timestamp 1606120353
transform 1 0 15272 0 -1 65824
box 0 -48 1196 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_806
timestamp 1606120353
transform 1 0 15180 0 -1 65824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_116_141
timestamp 1606120353
transform 1 0 14076 0 -1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_116_167
timestamp 1606120353
transform 1 0 16468 0 -1 65824
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_116_175
timestamp 1606120353
transform 1 0 17204 0 -1 65824
box 0 -48 276 592
use sky130_fd_sc_hd__o21ai_4  _1023_
timestamp 1606120353
transform 1 0 17480 0 -1 65824
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_12  FILLER_116_191
timestamp 1606120353
transform 1 0 18676 0 -1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_807
timestamp 1606120353
transform 1 0 20792 0 -1 65824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_116_203
timestamp 1606120353
transform 1 0 19780 0 -1 65824
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_116_211
timestamp 1606120353
transform 1 0 20516 0 -1 65824
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_116_215
timestamp 1606120353
transform 1 0 20884 0 -1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_116_227
timestamp 1606120353
transform 1 0 21988 0 -1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_116_239
timestamp 1606120353
transform 1 0 23092 0 -1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_116_251
timestamp 1606120353
transform 1 0 24196 0 -1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_116_263
timestamp 1606120353
transform 1 0 25300 0 -1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_808
timestamp 1606120353
transform 1 0 26404 0 -1 65824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_116_276
timestamp 1606120353
transform 1 0 26496 0 -1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_233
timestamp 1606120353
transform -1 0 28888 0 -1 65824
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_116_288
timestamp 1606120353
transform 1 0 27600 0 -1 65824
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_116_296
timestamp 1606120353
transform 1 0 28336 0 -1 65824
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_234
timestamp 1606120353
transform 1 0 1104 0 1 65824
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_117_3
timestamp 1606120353
transform 1 0 1380 0 1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_117_15
timestamp 1606120353
transform 1 0 2484 0 1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_117_27
timestamp 1606120353
transform 1 0 3588 0 1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_117_39
timestamp 1606120353
transform 1 0 4692 0 1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_809
timestamp 1606120353
transform 1 0 6716 0 1 65824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_117_51
timestamp 1606120353
transform 1 0 5796 0 1 65824
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_117_59
timestamp 1606120353
transform 1 0 6532 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_117_62
timestamp 1606120353
transform 1 0 6808 0 1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_117_74
timestamp 1606120353
transform 1 0 7912 0 1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_117_86
timestamp 1606120353
transform 1 0 9016 0 1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_117_98
timestamp 1606120353
transform 1 0 10120 0 1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_117_110
timestamp 1606120353
transform 1 0 11224 0 1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_810
timestamp 1606120353
transform 1 0 12328 0 1 65824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_117_123
timestamp 1606120353
transform 1 0 12420 0 1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_117_135
timestamp 1606120353
transform 1 0 13524 0 1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_117_147
timestamp 1606120353
transform 1 0 14628 0 1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__A1
timestamp 1606120353
transform 1 0 16744 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__A2
timestamp 1606120353
transform 1 0 17112 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__B1
timestamp 1606120353
transform 1 0 16376 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_117_159
timestamp 1606120353
transform 1 0 15732 0 1 65824
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_117_165
timestamp 1606120353
transform 1 0 16284 0 1 65824
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_117_168
timestamp 1606120353
transform 1 0 16560 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_117_172
timestamp 1606120353
transform 1 0 16928 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_117_176
timestamp 1606120353
transform 1 0 17296 0 1 65824
box 0 -48 368 592
use sky130_fd_sc_hd__dfxtp_4  _1217_
timestamp 1606120353
transform 1 0 18032 0 1 65824
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_811
timestamp 1606120353
transform 1 0 17940 0 1 65824
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__D
timestamp 1606120353
transform 1 0 17756 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_117_180
timestamp 1606120353
transform 1 0 17664 0 1 65824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_117_203
timestamp 1606120353
transform 1 0 19780 0 1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_117_215
timestamp 1606120353
transform 1 0 20884 0 1 65824
box 0 -48 736 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_clk_A
timestamp 1606120353
transform 1 0 21620 0 1 65824
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_117_225
timestamp 1606120353
transform 1 0 21804 0 1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_117_237
timestamp 1606120353
transform 1 0 22908 0 1 65824
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_812
timestamp 1606120353
transform 1 0 23552 0 1 65824
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_117_243
timestamp 1606120353
transform 1 0 23460 0 1 65824
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_117_245
timestamp 1606120353
transform 1 0 23644 0 1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_117_257
timestamp 1606120353
transform 1 0 24748 0 1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_117_269
timestamp 1606120353
transform 1 0 25852 0 1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_117_281
timestamp 1606120353
transform 1 0 26956 0 1 65824
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_235
timestamp 1606120353
transform -1 0 28888 0 1 65824
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_117_293
timestamp 1606120353
transform 1 0 28060 0 1 65824
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_236
timestamp 1606120353
transform 1 0 1104 0 -1 66912
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_238
timestamp 1606120353
transform 1 0 1104 0 1 66912
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_118_3
timestamp 1606120353
transform 1 0 1380 0 -1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_118_15
timestamp 1606120353
transform 1 0 2484 0 -1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_119_3
timestamp 1606120353
transform 1 0 1380 0 1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_119_15
timestamp 1606120353
transform 1 0 2484 0 1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_813
timestamp 1606120353
transform 1 0 3956 0 -1 66912
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_118_27
timestamp 1606120353
transform 1 0 3588 0 -1 66912
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_118_32
timestamp 1606120353
transform 1 0 4048 0 -1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_118_44
timestamp 1606120353
transform 1 0 5152 0 -1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_119_27
timestamp 1606120353
transform 1 0 3588 0 1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_119_39
timestamp 1606120353
transform 1 0 4692 0 1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_818
timestamp 1606120353
transform 1 0 6716 0 1 66912
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_118_56
timestamp 1606120353
transform 1 0 6256 0 -1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_119_51
timestamp 1606120353
transform 1 0 5796 0 1 66912
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_119_59
timestamp 1606120353
transform 1 0 6532 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_119_62
timestamp 1606120353
transform 1 0 6808 0 1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_118_68
timestamp 1606120353
transform 1 0 7360 0 -1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_118_80
timestamp 1606120353
transform 1 0 8464 0 -1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_119_74
timestamp 1606120353
transform 1 0 7912 0 1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_119_86
timestamp 1606120353
transform 1 0 9016 0 1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_814
timestamp 1606120353
transform 1 0 9568 0 -1 66912
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_clk
timestamp 1606120353
transform 1 0 10672 0 1 66912
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_clk_A
timestamp 1606120353
transform 1 0 11132 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_118_93
timestamp 1606120353
transform 1 0 9660 0 -1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_118_105
timestamp 1606120353
transform 1 0 10764 0 -1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_119_98
timestamp 1606120353
transform 1 0 10120 0 1 66912
box 0 -48 552 592
use sky130_fd_sc_hd__fill_2  FILLER_119_107
timestamp 1606120353
transform 1 0 10948 0 1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_819
timestamp 1606120353
transform 1 0 12328 0 1 66912
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_118_117
timestamp 1606120353
transform 1 0 11868 0 -1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_118_129
timestamp 1606120353
transform 1 0 12972 0 -1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_119_111
timestamp 1606120353
transform 1 0 11316 0 1 66912
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_119_119
timestamp 1606120353
transform 1 0 12052 0 1 66912
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_119_123
timestamp 1606120353
transform 1 0 12420 0 1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_815
timestamp 1606120353
transform 1 0 15180 0 -1 66912
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_118_141
timestamp 1606120353
transform 1 0 14076 0 -1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_118_154
timestamp 1606120353
transform 1 0 15272 0 -1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_119_135
timestamp 1606120353
transform 1 0 13524 0 1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_119_147
timestamp 1606120353
transform 1 0 14628 0 1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__o21ai_4  _1020_
timestamp 1606120353
transform 1 0 16744 0 -1 66912
box 0 -48 1196 592
use sky130_fd_sc_hd__decap_4  FILLER_118_166
timestamp 1606120353
transform 1 0 16376 0 -1 66912
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_119_159
timestamp 1606120353
transform 1 0 15732 0 1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_119_171
timestamp 1606120353
transform 1 0 16836 0 1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_820
timestamp 1606120353
transform 1 0 17940 0 1 66912
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__CLK
timestamp 1606120353
transform 1 0 18124 0 -1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_118_183
timestamp 1606120353
transform 1 0 17940 0 -1 66912
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_118_187
timestamp 1606120353
transform 1 0 18308 0 -1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_119_184
timestamp 1606120353
transform 1 0 18032 0 1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_119_196
timestamp 1606120353
transform 1 0 19136 0 1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_816
timestamp 1606120353
transform 1 0 20792 0 -1 66912
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_118_199
timestamp 1606120353
transform 1 0 19412 0 -1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_118_211
timestamp 1606120353
transform 1 0 20516 0 -1 66912
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_118_215
timestamp 1606120353
transform 1 0 20884 0 -1 66912
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_119_208
timestamp 1606120353
transform 1 0 20240 0 1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_119_220
timestamp 1606120353
transform 1 0 21344 0 1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_clk
timestamp 1606120353
transform 1 0 21620 0 -1 66912
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_118_226
timestamp 1606120353
transform 1 0 21896 0 -1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_118_238
timestamp 1606120353
transform 1 0 23000 0 -1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_119_232
timestamp 1606120353
transform 1 0 22448 0 1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_821
timestamp 1606120353
transform 1 0 23552 0 1 66912
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_118_250
timestamp 1606120353
transform 1 0 24104 0 -1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_118_262
timestamp 1606120353
transform 1 0 25208 0 -1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_119_245
timestamp 1606120353
transform 1 0 23644 0 1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_119_257
timestamp 1606120353
transform 1 0 24748 0 1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_817
timestamp 1606120353
transform 1 0 26404 0 -1 66912
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_118_274
timestamp 1606120353
transform 1 0 26312 0 -1 66912
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_118_276
timestamp 1606120353
transform 1 0 26496 0 -1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_119_269
timestamp 1606120353
transform 1 0 25852 0 1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_119_281
timestamp 1606120353
transform 1 0 26956 0 1 66912
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_237
timestamp 1606120353
transform -1 0 28888 0 -1 66912
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_239
timestamp 1606120353
transform -1 0 28888 0 1 66912
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_118_288
timestamp 1606120353
transform 1 0 27600 0 -1 66912
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_118_296
timestamp 1606120353
transform 1 0 28336 0 -1 66912
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_119_293
timestamp 1606120353
transform 1 0 28060 0 1 66912
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_240
timestamp 1606120353
transform 1 0 1104 0 -1 68000
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_120_3
timestamp 1606120353
transform 1 0 1380 0 -1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_120_15
timestamp 1606120353
transform 1 0 2484 0 -1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_822
timestamp 1606120353
transform 1 0 3956 0 -1 68000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_120_27
timestamp 1606120353
transform 1 0 3588 0 -1 68000
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_120_32
timestamp 1606120353
transform 1 0 4048 0 -1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_120_44
timestamp 1606120353
transform 1 0 5152 0 -1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_120_56
timestamp 1606120353
transform 1 0 6256 0 -1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_120_68
timestamp 1606120353
transform 1 0 7360 0 -1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_120_80
timestamp 1606120353
transform 1 0 8464 0 -1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_823
timestamp 1606120353
transform 1 0 9568 0 -1 68000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_120_93
timestamp 1606120353
transform 1 0 9660 0 -1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_120_105
timestamp 1606120353
transform 1 0 10764 0 -1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_120_117
timestamp 1606120353
transform 1 0 11868 0 -1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_120_129
timestamp 1606120353
transform 1 0 12972 0 -1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_824
timestamp 1606120353
transform 1 0 15180 0 -1 68000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_120_141
timestamp 1606120353
transform 1 0 14076 0 -1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_120_154
timestamp 1606120353
transform 1 0 15272 0 -1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_120_166
timestamp 1606120353
transform 1 0 16376 0 -1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_120_178
timestamp 1606120353
transform 1 0 17480 0 -1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_120_190
timestamp 1606120353
transform 1 0 18584 0 -1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_825
timestamp 1606120353
transform 1 0 20792 0 -1 68000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_120_202
timestamp 1606120353
transform 1 0 19688 0 -1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_120_215
timestamp 1606120353
transform 1 0 20884 0 -1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_120_227
timestamp 1606120353
transform 1 0 21988 0 -1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_120_239
timestamp 1606120353
transform 1 0 23092 0 -1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_120_251
timestamp 1606120353
transform 1 0 24196 0 -1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_120_263
timestamp 1606120353
transform 1 0 25300 0 -1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_826
timestamp 1606120353
transform 1 0 26404 0 -1 68000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_120_276
timestamp 1606120353
transform 1 0 26496 0 -1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_241
timestamp 1606120353
transform -1 0 28888 0 -1 68000
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_120_288
timestamp 1606120353
transform 1 0 27600 0 -1 68000
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_120_296
timestamp 1606120353
transform 1 0 28336 0 -1 68000
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_242
timestamp 1606120353
transform 1 0 1104 0 1 68000
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_121_3
timestamp 1606120353
transform 1 0 1380 0 1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_121_15
timestamp 1606120353
transform 1 0 2484 0 1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_121_27
timestamp 1606120353
transform 1 0 3588 0 1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_121_39
timestamp 1606120353
transform 1 0 4692 0 1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_827
timestamp 1606120353
transform 1 0 6716 0 1 68000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_121_51
timestamp 1606120353
transform 1 0 5796 0 1 68000
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_121_59
timestamp 1606120353
transform 1 0 6532 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_121_62
timestamp 1606120353
transform 1 0 6808 0 1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_clk
timestamp 1606120353
transform 1 0 9108 0 1 68000
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_121_74
timestamp 1606120353
transform 1 0 7912 0 1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_121_86
timestamp 1606120353
transform 1 0 9016 0 1 68000
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_clk_A
timestamp 1606120353
transform 1 0 9568 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_121_90
timestamp 1606120353
transform 1 0 9384 0 1 68000
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_121_94
timestamp 1606120353
transform 1 0 9752 0 1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_121_106
timestamp 1606120353
transform 1 0 10856 0 1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_828
timestamp 1606120353
transform 1 0 12328 0 1 68000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_121_118
timestamp 1606120353
transform 1 0 11960 0 1 68000
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_121_123
timestamp 1606120353
transform 1 0 12420 0 1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_121_135
timestamp 1606120353
transform 1 0 13524 0 1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_121_147
timestamp 1606120353
transform 1 0 14628 0 1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_121_159
timestamp 1606120353
transform 1 0 15732 0 1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_121_171
timestamp 1606120353
transform 1 0 16836 0 1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_829
timestamp 1606120353
transform 1 0 17940 0 1 68000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_121_184
timestamp 1606120353
transform 1 0 18032 0 1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_121_196
timestamp 1606120353
transform 1 0 19136 0 1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_121_208
timestamp 1606120353
transform 1 0 20240 0 1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_121_220
timestamp 1606120353
transform 1 0 21344 0 1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_121_232
timestamp 1606120353
transform 1 0 22448 0 1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_830
timestamp 1606120353
transform 1 0 23552 0 1 68000
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_121_245
timestamp 1606120353
transform 1 0 23644 0 1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_121_257
timestamp 1606120353
transform 1 0 24748 0 1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_121_269
timestamp 1606120353
transform 1 0 25852 0 1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_121_281
timestamp 1606120353
transform 1 0 26956 0 1 68000
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_243
timestamp 1606120353
transform -1 0 28888 0 1 68000
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_121_293
timestamp 1606120353
transform 1 0 28060 0 1 68000
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_244
timestamp 1606120353
transform 1 0 1104 0 -1 69088
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_122_3
timestamp 1606120353
transform 1 0 1380 0 -1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_122_15
timestamp 1606120353
transform 1 0 2484 0 -1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_831
timestamp 1606120353
transform 1 0 3956 0 -1 69088
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_122_27
timestamp 1606120353
transform 1 0 3588 0 -1 69088
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_122_32
timestamp 1606120353
transform 1 0 4048 0 -1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_122_44
timestamp 1606120353
transform 1 0 5152 0 -1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_122_56
timestamp 1606120353
transform 1 0 6256 0 -1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_122_68
timestamp 1606120353
transform 1 0 7360 0 -1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_122_80
timestamp 1606120353
transform 1 0 8464 0 -1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_832
timestamp 1606120353
transform 1 0 9568 0 -1 69088
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_122_93
timestamp 1606120353
transform 1 0 9660 0 -1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_122_105
timestamp 1606120353
transform 1 0 10764 0 -1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_122_117
timestamp 1606120353
transform 1 0 11868 0 -1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_122_129
timestamp 1606120353
transform 1 0 12972 0 -1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_833
timestamp 1606120353
transform 1 0 15180 0 -1 69088
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_122_141
timestamp 1606120353
transform 1 0 14076 0 -1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_122_154
timestamp 1606120353
transform 1 0 15272 0 -1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_122_166
timestamp 1606120353
transform 1 0 16376 0 -1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_122_178
timestamp 1606120353
transform 1 0 17480 0 -1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_122_190
timestamp 1606120353
transform 1 0 18584 0 -1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_834
timestamp 1606120353
transform 1 0 20792 0 -1 69088
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_122_202
timestamp 1606120353
transform 1 0 19688 0 -1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_122_215
timestamp 1606120353
transform 1 0 20884 0 -1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_122_227
timestamp 1606120353
transform 1 0 21988 0 -1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_122_239
timestamp 1606120353
transform 1 0 23092 0 -1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_122_251
timestamp 1606120353
transform 1 0 24196 0 -1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_122_263
timestamp 1606120353
transform 1 0 25300 0 -1 69088
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_835
timestamp 1606120353
transform 1 0 26404 0 -1 69088
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__CLK
timestamp 1606120353
transform 1 0 26128 0 -1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_122_271
timestamp 1606120353
transform 1 0 26036 0 -1 69088
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_122_274
timestamp 1606120353
transform 1 0 26312 0 -1 69088
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_122_276
timestamp 1606120353
transform 1 0 26496 0 -1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_245
timestamp 1606120353
transform -1 0 28888 0 -1 69088
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_122_288
timestamp 1606120353
transform 1 0 27600 0 -1 69088
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_122_296
timestamp 1606120353
transform 1 0 28336 0 -1 69088
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_246
timestamp 1606120353
transform 1 0 1104 0 1 69088
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__D
timestamp 1606120353
transform 1 0 1564 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__CLK
timestamp 1606120353
transform 1 0 1932 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_123_3
timestamp 1606120353
transform 1 0 1380 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_123_7
timestamp 1606120353
transform 1 0 1748 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_123_11
timestamp 1606120353
transform 1 0 2116 0 1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_123_23
timestamp 1606120353
transform 1 0 3220 0 1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_123_35
timestamp 1606120353
transform 1 0 4324 0 1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_836
timestamp 1606120353
transform 1 0 6716 0 1 69088
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_123_47
timestamp 1606120353
transform 1 0 5428 0 1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_123_59
timestamp 1606120353
transform 1 0 6532 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_123_62
timestamp 1606120353
transform 1 0 6808 0 1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_123_74
timestamp 1606120353
transform 1 0 7912 0 1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_123_86
timestamp 1606120353
transform 1 0 9016 0 1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_123_98
timestamp 1606120353
transform 1 0 10120 0 1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_1  FILLER_123_110
timestamp 1606120353
transform 1 0 11224 0 1 69088
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_837
timestamp 1606120353
transform 1 0 12328 0 1 69088
box 0 -48 92 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_clk
timestamp 1606120353
transform 1 0 11316 0 1 69088
box 0 -48 276 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_clk_A
timestamp 1606120353
transform 1 0 11776 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_123_114
timestamp 1606120353
transform 1 0 11592 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__decap_4  FILLER_123_118
timestamp 1606120353
transform 1 0 11960 0 1 69088
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_123_123
timestamp 1606120353
transform 1 0 12420 0 1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_123_135
timestamp 1606120353
transform 1 0 13524 0 1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_123_147
timestamp 1606120353
transform 1 0 14628 0 1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_123_159
timestamp 1606120353
transform 1 0 15732 0 1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_123_171
timestamp 1606120353
transform 1 0 16836 0 1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_838
timestamp 1606120353
transform 1 0 17940 0 1 69088
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_123_184
timestamp 1606120353
transform 1 0 18032 0 1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_123_196
timestamp 1606120353
transform 1 0 19136 0 1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_123_208
timestamp 1606120353
transform 1 0 20240 0 1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_123_220
timestamp 1606120353
transform 1 0 21344 0 1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_123_232
timestamp 1606120353
transform 1 0 22448 0 1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_839
timestamp 1606120353
transform 1 0 23552 0 1 69088
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_123_245
timestamp 1606120353
transform 1 0 23644 0 1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_123_257
timestamp 1606120353
transform 1 0 24748 0 1 69088
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1159_
timestamp 1606120353
transform 1 0 26128 0 1 69088
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__D
timestamp 1606120353
transform 1 0 25944 0 1 69088
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_123_269
timestamp 1606120353
transform 1 0 25852 0 1 69088
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  PHY_247
timestamp 1606120353
transform -1 0 28888 0 1 69088
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_123_291
timestamp 1606120353
transform 1 0 27876 0 1 69088
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1201_
timestamp 1606120353
transform 1 0 1380 0 -1 70176
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_3  PHY_248
timestamp 1606120353
transform 1 0 1104 0 -1 70176
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_124_22
timestamp 1606120353
transform 1 0 3128 0 -1 70176
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_840
timestamp 1606120353
transform 1 0 3956 0 -1 70176
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_124_30
timestamp 1606120353
transform 1 0 3864 0 -1 70176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_124_32
timestamp 1606120353
transform 1 0 4048 0 -1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_124_44
timestamp 1606120353
transform 1 0 5152 0 -1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_124_56
timestamp 1606120353
transform 1 0 6256 0 -1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_124_68
timestamp 1606120353
transform 1 0 7360 0 -1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_124_80
timestamp 1606120353
transform 1 0 8464 0 -1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_841
timestamp 1606120353
transform 1 0 9568 0 -1 70176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_124_93
timestamp 1606120353
transform 1 0 9660 0 -1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_124_105
timestamp 1606120353
transform 1 0 10764 0 -1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_124_117
timestamp 1606120353
transform 1 0 11868 0 -1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_124_129
timestamp 1606120353
transform 1 0 12972 0 -1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_842
timestamp 1606120353
transform 1 0 15180 0 -1 70176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_124_141
timestamp 1606120353
transform 1 0 14076 0 -1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_124_154
timestamp 1606120353
transform 1 0 15272 0 -1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_124_166
timestamp 1606120353
transform 1 0 16376 0 -1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_124_178
timestamp 1606120353
transform 1 0 17480 0 -1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_124_190
timestamp 1606120353
transform 1 0 18584 0 -1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_843
timestamp 1606120353
transform 1 0 20792 0 -1 70176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_124_202
timestamp 1606120353
transform 1 0 19688 0 -1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_124_215
timestamp 1606120353
transform 1 0 20884 0 -1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_124_227
timestamp 1606120353
transform 1 0 21988 0 -1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_124_239
timestamp 1606120353
transform 1 0 23092 0 -1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_124_251
timestamp 1606120353
transform 1 0 24196 0 -1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_124_263
timestamp 1606120353
transform 1 0 25300 0 -1 70176
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_844
timestamp 1606120353
transform 1 0 26404 0 -1 70176
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__CLK
timestamp 1606120353
transform 1 0 26128 0 -1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_124_271
timestamp 1606120353
transform 1 0 26036 0 -1 70176
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_124_274
timestamp 1606120353
transform 1 0 26312 0 -1 70176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_124_276
timestamp 1606120353
transform 1 0 26496 0 -1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_249
timestamp 1606120353
transform -1 0 28888 0 -1 70176
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_124_288
timestamp 1606120353
transform 1 0 27600 0 -1 70176
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_124_296
timestamp 1606120353
transform 1 0 28336 0 -1 70176
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_250
timestamp 1606120353
transform 1 0 1104 0 1 70176
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_252
timestamp 1606120353
transform 1 0 1104 0 -1 71264
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_125_3
timestamp 1606120353
transform 1 0 1380 0 1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_125_15
timestamp 1606120353
transform 1 0 2484 0 1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_126_3
timestamp 1606120353
transform 1 0 1380 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_126_15
timestamp 1606120353
transform 1 0 2484 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_849
timestamp 1606120353
transform 1 0 3956 0 -1 71264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_125_27
timestamp 1606120353
transform 1 0 3588 0 1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_125_39
timestamp 1606120353
transform 1 0 4692 0 1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_126_27
timestamp 1606120353
transform 1 0 3588 0 -1 71264
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_126_32
timestamp 1606120353
transform 1 0 4048 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_126_44
timestamp 1606120353
transform 1 0 5152 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_845
timestamp 1606120353
transform 1 0 6716 0 1 70176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_125_51
timestamp 1606120353
transform 1 0 5796 0 1 70176
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_125_59
timestamp 1606120353
transform 1 0 6532 0 1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_125_62
timestamp 1606120353
transform 1 0 6808 0 1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_126_56
timestamp 1606120353
transform 1 0 6256 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_125_74
timestamp 1606120353
transform 1 0 7912 0 1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_125_86
timestamp 1606120353
transform 1 0 9016 0 1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_126_68
timestamp 1606120353
transform 1 0 7360 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_126_80
timestamp 1606120353
transform 1 0 8464 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_850
timestamp 1606120353
transform 1 0 9568 0 -1 71264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_125_98
timestamp 1606120353
transform 1 0 10120 0 1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_125_110
timestamp 1606120353
transform 1 0 11224 0 1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_126_93
timestamp 1606120353
transform 1 0 9660 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_126_105
timestamp 1606120353
transform 1 0 10764 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_846
timestamp 1606120353
transform 1 0 12328 0 1 70176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_125_123
timestamp 1606120353
transform 1 0 12420 0 1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_126_117
timestamp 1606120353
transform 1 0 11868 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_126_129
timestamp 1606120353
transform 1 0 12972 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_851
timestamp 1606120353
transform 1 0 15180 0 -1 71264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_125_135
timestamp 1606120353
transform 1 0 13524 0 1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_125_147
timestamp 1606120353
transform 1 0 14628 0 1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_126_141
timestamp 1606120353
transform 1 0 14076 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_126_154
timestamp 1606120353
transform 1 0 15272 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_125_159
timestamp 1606120353
transform 1 0 15732 0 1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_125_171
timestamp 1606120353
transform 1 0 16836 0 1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_126_166
timestamp 1606120353
transform 1 0 16376 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_847
timestamp 1606120353
transform 1 0 17940 0 1 70176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_125_184
timestamp 1606120353
transform 1 0 18032 0 1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_125_196
timestamp 1606120353
transform 1 0 19136 0 1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_126_178
timestamp 1606120353
transform 1 0 17480 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_126_190
timestamp 1606120353
transform 1 0 18584 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1203_
timestamp 1606120353
transform 1 0 20884 0 -1 71264
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_852
timestamp 1606120353
transform 1 0 20792 0 -1 71264
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__D
timestamp 1606120353
transform 1 0 20884 0 1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__CLK
timestamp 1606120353
transform 1 0 21252 0 1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_125_208
timestamp 1606120353
transform 1 0 20240 0 1 70176
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_125_214
timestamp 1606120353
transform 1 0 20792 0 1 70176
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_125_217
timestamp 1606120353
transform 1 0 21068 0 1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_126_202
timestamp 1606120353
transform 1 0 19688 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_125_221
timestamp 1606120353
transform 1 0 21436 0 1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_125_233
timestamp 1606120353
transform 1 0 22540 0 1 70176
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_125_241
timestamp 1606120353
transform 1 0 23276 0 1 70176
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_126_234
timestamp 1606120353
transform 1 0 22632 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_848
timestamp 1606120353
transform 1 0 23552 0 1 70176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_125_245
timestamp 1606120353
transform 1 0 23644 0 1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_125_257
timestamp 1606120353
transform 1 0 24748 0 1 70176
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_126_246
timestamp 1606120353
transform 1 0 23736 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_126_258
timestamp 1606120353
transform 1 0 24840 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1222_
timestamp 1606120353
transform 1 0 26128 0 1 70176
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_853
timestamp 1606120353
transform 1 0 26404 0 -1 71264
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__D
timestamp 1606120353
transform 1 0 25944 0 1 70176
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_125_269
timestamp 1606120353
transform 1 0 25852 0 1 70176
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_126_270
timestamp 1606120353
transform 1 0 25944 0 -1 71264
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_126_274
timestamp 1606120353
transform 1 0 26312 0 -1 71264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_126_276
timestamp 1606120353
transform 1 0 26496 0 -1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_251
timestamp 1606120353
transform -1 0 28888 0 1 70176
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_253
timestamp 1606120353
transform -1 0 28888 0 -1 71264
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_125_291
timestamp 1606120353
transform 1 0 27876 0 1 70176
box 0 -48 736 592
use sky130_fd_sc_hd__decap_8  FILLER_126_288
timestamp 1606120353
transform 1 0 27600 0 -1 71264
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_126_296
timestamp 1606120353
transform 1 0 28336 0 -1 71264
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_254
timestamp 1606120353
transform 1 0 1104 0 1 71264
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_127_3
timestamp 1606120353
transform 1 0 1380 0 1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_127_15
timestamp 1606120353
transform 1 0 2484 0 1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_127_27
timestamp 1606120353
transform 1 0 3588 0 1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_127_39
timestamp 1606120353
transform 1 0 4692 0 1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_854
timestamp 1606120353
transform 1 0 6716 0 1 71264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_127_51
timestamp 1606120353
transform 1 0 5796 0 1 71264
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_127_59
timestamp 1606120353
transform 1 0 6532 0 1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_127_62
timestamp 1606120353
transform 1 0 6808 0 1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_127_74
timestamp 1606120353
transform 1 0 7912 0 1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_127_86
timestamp 1606120353
transform 1 0 9016 0 1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_127_98
timestamp 1606120353
transform 1 0 10120 0 1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_127_110
timestamp 1606120353
transform 1 0 11224 0 1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_855
timestamp 1606120353
transform 1 0 12328 0 1 71264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_127_123
timestamp 1606120353
transform 1 0 12420 0 1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_127_135
timestamp 1606120353
transform 1 0 13524 0 1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_127_147
timestamp 1606120353
transform 1 0 14628 0 1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_127_159
timestamp 1606120353
transform 1 0 15732 0 1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_127_171
timestamp 1606120353
transform 1 0 16836 0 1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_856
timestamp 1606120353
transform 1 0 17940 0 1 71264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_127_184
timestamp 1606120353
transform 1 0 18032 0 1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_127_196
timestamp 1606120353
transform 1 0 19136 0 1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__D
timestamp 1606120353
transform 1 0 20884 0 1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__CLK
timestamp 1606120353
transform 1 0 21252 0 1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_127_208
timestamp 1606120353
transform 1 0 20240 0 1 71264
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_127_214
timestamp 1606120353
transform 1 0 20792 0 1 71264
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_127_217
timestamp 1606120353
transform 1 0 21068 0 1 71264
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_127_221
timestamp 1606120353
transform 1 0 21436 0 1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_127_233
timestamp 1606120353
transform 1 0 22540 0 1 71264
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_127_241
timestamp 1606120353
transform 1 0 23276 0 1 71264
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_857
timestamp 1606120353
transform 1 0 23552 0 1 71264
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_127_245
timestamp 1606120353
transform 1 0 23644 0 1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_127_257
timestamp 1606120353
transform 1 0 24748 0 1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_127_269
timestamp 1606120353
transform 1 0 25852 0 1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_127_281
timestamp 1606120353
transform 1 0 26956 0 1 71264
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_255
timestamp 1606120353
transform -1 0 28888 0 1 71264
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_127_293
timestamp 1606120353
transform 1 0 28060 0 1 71264
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_256
timestamp 1606120353
transform 1 0 1104 0 -1 72352
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_128_3
timestamp 1606120353
transform 1 0 1380 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_128_15
timestamp 1606120353
transform 1 0 2484 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_858
timestamp 1606120353
transform 1 0 3956 0 -1 72352
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_128_27
timestamp 1606120353
transform 1 0 3588 0 -1 72352
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_128_32
timestamp 1606120353
transform 1 0 4048 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_128_44
timestamp 1606120353
transform 1 0 5152 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_128_56
timestamp 1606120353
transform 1 0 6256 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_128_68
timestamp 1606120353
transform 1 0 7360 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_128_80
timestamp 1606120353
transform 1 0 8464 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_859
timestamp 1606120353
transform 1 0 9568 0 -1 72352
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_128_93
timestamp 1606120353
transform 1 0 9660 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_128_105
timestamp 1606120353
transform 1 0 10764 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_128_117
timestamp 1606120353
transform 1 0 11868 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_128_129
timestamp 1606120353
transform 1 0 12972 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_860
timestamp 1606120353
transform 1 0 15180 0 -1 72352
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_128_141
timestamp 1606120353
transform 1 0 14076 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_128_154
timestamp 1606120353
transform 1 0 15272 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_128_166
timestamp 1606120353
transform 1 0 16376 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_128_178
timestamp 1606120353
transform 1 0 17480 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_128_190
timestamp 1606120353
transform 1 0 18584 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1199_
timestamp 1606120353
transform 1 0 20884 0 -1 72352
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_861
timestamp 1606120353
transform 1 0 20792 0 -1 72352
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_128_202
timestamp 1606120353
transform 1 0 19688 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_128_234
timestamp 1606120353
transform 1 0 22632 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_128_246
timestamp 1606120353
transform 1 0 23736 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_128_258
timestamp 1606120353
transform 1 0 24840 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_862
timestamp 1606120353
transform 1 0 26404 0 -1 72352
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_128_270
timestamp 1606120353
transform 1 0 25944 0 -1 72352
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_128_274
timestamp 1606120353
transform 1 0 26312 0 -1 72352
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_128_276
timestamp 1606120353
transform 1 0 26496 0 -1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_257
timestamp 1606120353
transform -1 0 28888 0 -1 72352
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_128_288
timestamp 1606120353
transform 1 0 27600 0 -1 72352
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_128_296
timestamp 1606120353
transform 1 0 28336 0 -1 72352
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_258
timestamp 1606120353
transform 1 0 1104 0 1 72352
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_129_3
timestamp 1606120353
transform 1 0 1380 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_129_15
timestamp 1606120353
transform 1 0 2484 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_129_27
timestamp 1606120353
transform 1 0 3588 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_129_39
timestamp 1606120353
transform 1 0 4692 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_863
timestamp 1606120353
transform 1 0 6716 0 1 72352
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_129_51
timestamp 1606120353
transform 1 0 5796 0 1 72352
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_129_59
timestamp 1606120353
transform 1 0 6532 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_129_62
timestamp 1606120353
transform 1 0 6808 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_129_74
timestamp 1606120353
transform 1 0 7912 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_129_86
timestamp 1606120353
transform 1 0 9016 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_129_98
timestamp 1606120353
transform 1 0 10120 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_129_110
timestamp 1606120353
transform 1 0 11224 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_864
timestamp 1606120353
transform 1 0 12328 0 1 72352
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__D
timestamp 1606120353
transform 1 0 12696 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__CLK
timestamp 1606120353
transform 1 0 13064 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  FILLER_129_123
timestamp 1606120353
transform 1 0 12420 0 1 72352
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_129_128
timestamp 1606120353
transform 1 0 12880 0 1 72352
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_129_132
timestamp 1606120353
transform 1 0 13248 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_129_144
timestamp 1606120353
transform 1 0 14352 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_129_156
timestamp 1606120353
transform 1 0 15456 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_129_168
timestamp 1606120353
transform 1 0 16560 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_865
timestamp 1606120353
transform 1 0 17940 0 1 72352
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_129_180
timestamp 1606120353
transform 1 0 17664 0 1 72352
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_129_184
timestamp 1606120353
transform 1 0 18032 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_129_196
timestamp 1606120353
transform 1 0 19136 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_129_208
timestamp 1606120353
transform 1 0 20240 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_129_220
timestamp 1606120353
transform 1 0 21344 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_129_232
timestamp 1606120353
transform 1 0 22448 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_866
timestamp 1606120353
transform 1 0 23552 0 1 72352
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_129_245
timestamp 1606120353
transform 1 0 23644 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_129_257
timestamp 1606120353
transform 1 0 24748 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_129_269
timestamp 1606120353
transform 1 0 25852 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_129_281
timestamp 1606120353
transform 1 0 26956 0 1 72352
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_259
timestamp 1606120353
transform -1 0 28888 0 1 72352
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_129_293
timestamp 1606120353
transform 1 0 28060 0 1 72352
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_260
timestamp 1606120353
transform 1 0 1104 0 -1 73440
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_130_3
timestamp 1606120353
transform 1 0 1380 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_130_15
timestamp 1606120353
transform 1 0 2484 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_867
timestamp 1606120353
transform 1 0 3956 0 -1 73440
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_130_27
timestamp 1606120353
transform 1 0 3588 0 -1 73440
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_130_32
timestamp 1606120353
transform 1 0 4048 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_130_44
timestamp 1606120353
transform 1 0 5152 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_130_56
timestamp 1606120353
transform 1 0 6256 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_130_68
timestamp 1606120353
transform 1 0 7360 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_130_80
timestamp 1606120353
transform 1 0 8464 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_868
timestamp 1606120353
transform 1 0 9568 0 -1 73440
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_130_93
timestamp 1606120353
transform 1 0 9660 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_130_105
timestamp 1606120353
transform 1 0 10764 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1153_
timestamp 1606120353
transform 1 0 12696 0 -1 73440
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_8  FILLER_130_117
timestamp 1606120353
transform 1 0 11868 0 -1 73440
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_130_125
timestamp 1606120353
transform 1 0 12604 0 -1 73440
box 0 -48 92 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_869
timestamp 1606120353
transform 1 0 15180 0 -1 73440
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_130_145
timestamp 1606120353
transform 1 0 14444 0 -1 73440
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_130_154
timestamp 1606120353
transform 1 0 15272 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_130_166
timestamp 1606120353
transform 1 0 16376 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_130_178
timestamp 1606120353
transform 1 0 17480 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_130_190
timestamp 1606120353
transform 1 0 18584 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_870
timestamp 1606120353
transform 1 0 20792 0 -1 73440
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_130_202
timestamp 1606120353
transform 1 0 19688 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_130_215
timestamp 1606120353
transform 1 0 20884 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_130_227
timestamp 1606120353
transform 1 0 21988 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_130_239
timestamp 1606120353
transform 1 0 23092 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_130_251
timestamp 1606120353
transform 1 0 24196 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_130_263
timestamp 1606120353
transform 1 0 25300 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_871
timestamp 1606120353
transform 1 0 26404 0 -1 73440
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_130_276
timestamp 1606120353
transform 1 0 26496 0 -1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_261
timestamp 1606120353
transform -1 0 28888 0 -1 73440
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_130_288
timestamp 1606120353
transform 1 0 27600 0 -1 73440
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_130_296
timestamp 1606120353
transform 1 0 28336 0 -1 73440
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_262
timestamp 1606120353
transform 1 0 1104 0 1 73440
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_131_3
timestamp 1606120353
transform 1 0 1380 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_131_15
timestamp 1606120353
transform 1 0 2484 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_131_27
timestamp 1606120353
transform 1 0 3588 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_131_39
timestamp 1606120353
transform 1 0 4692 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_872
timestamp 1606120353
transform 1 0 6716 0 1 73440
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_131_51
timestamp 1606120353
transform 1 0 5796 0 1 73440
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_131_59
timestamp 1606120353
transform 1 0 6532 0 1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_131_62
timestamp 1606120353
transform 1 0 6808 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_131_74
timestamp 1606120353
transform 1 0 7912 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_131_86
timestamp 1606120353
transform 1 0 9016 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_131_98
timestamp 1606120353
transform 1 0 10120 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_131_110
timestamp 1606120353
transform 1 0 11224 0 1 73440
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_873
timestamp 1606120353
transform 1 0 12328 0 1 73440
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__D
timestamp 1606120353
transform 1 0 12144 0 1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__CLK
timestamp 1606120353
transform 1 0 12604 0 1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_131_118
timestamp 1606120353
transform 1 0 11960 0 1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_131_123
timestamp 1606120353
transform 1 0 12420 0 1 73440
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_131_127
timestamp 1606120353
transform 1 0 12788 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_131_139
timestamp 1606120353
transform 1 0 13892 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_131_151
timestamp 1606120353
transform 1 0 14996 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_131_163
timestamp 1606120353
transform 1 0 16100 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_131_175
timestamp 1606120353
transform 1 0 17204 0 1 73440
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_874
timestamp 1606120353
transform 1 0 17940 0 1 73440
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_131_184
timestamp 1606120353
transform 1 0 18032 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_131_196
timestamp 1606120353
transform 1 0 19136 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_131_208
timestamp 1606120353
transform 1 0 20240 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_131_220
timestamp 1606120353
transform 1 0 21344 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_131_232
timestamp 1606120353
transform 1 0 22448 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_875
timestamp 1606120353
transform 1 0 23552 0 1 73440
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_131_245
timestamp 1606120353
transform 1 0 23644 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_131_257
timestamp 1606120353
transform 1 0 24748 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_131_269
timestamp 1606120353
transform 1 0 25852 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_131_281
timestamp 1606120353
transform 1 0 26956 0 1 73440
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_263
timestamp 1606120353
transform -1 0 28888 0 1 73440
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_131_293
timestamp 1606120353
transform 1 0 28060 0 1 73440
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_264
timestamp 1606120353
transform 1 0 1104 0 -1 74528
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_266
timestamp 1606120353
transform 1 0 1104 0 1 74528
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_132_3
timestamp 1606120353
transform 1 0 1380 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_132_15
timestamp 1606120353
transform 1 0 2484 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_133_3
timestamp 1606120353
transform 1 0 1380 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_133_15
timestamp 1606120353
transform 1 0 2484 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_876
timestamp 1606120353
transform 1 0 3956 0 -1 74528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_132_27
timestamp 1606120353
transform 1 0 3588 0 -1 74528
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_132_32
timestamp 1606120353
transform 1 0 4048 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_132_44
timestamp 1606120353
transform 1 0 5152 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_133_27
timestamp 1606120353
transform 1 0 3588 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_133_39
timestamp 1606120353
transform 1 0 4692 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_881
timestamp 1606120353
transform 1 0 6716 0 1 74528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_132_56
timestamp 1606120353
transform 1 0 6256 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_133_51
timestamp 1606120353
transform 1 0 5796 0 1 74528
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_133_59
timestamp 1606120353
transform 1 0 6532 0 1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_133_62
timestamp 1606120353
transform 1 0 6808 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_132_68
timestamp 1606120353
transform 1 0 7360 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_132_80
timestamp 1606120353
transform 1 0 8464 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_133_74
timestamp 1606120353
transform 1 0 7912 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_133_86
timestamp 1606120353
transform 1 0 9016 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_877
timestamp 1606120353
transform 1 0 9568 0 -1 74528
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__D
timestamp 1606120353
transform 1 0 10396 0 1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__CLK
timestamp 1606120353
transform 1 0 10764 0 1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_132_93
timestamp 1606120353
transform 1 0 9660 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_132_105
timestamp 1606120353
transform 1 0 10764 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_133_98
timestamp 1606120353
transform 1 0 10120 0 1 74528
box 0 -48 276 592
use sky130_fd_sc_hd__fill_2  FILLER_133_103
timestamp 1606120353
transform 1 0 10580 0 1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_133_107
timestamp 1606120353
transform 1 0 10948 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1161_
timestamp 1606120353
transform 1 0 12144 0 -1 74528
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_882
timestamp 1606120353
transform 1 0 12328 0 1 74528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_132_117
timestamp 1606120353
transform 1 0 11868 0 -1 74528
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  FILLER_133_119
timestamp 1606120353
transform 1 0 12052 0 1 74528
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_133_123
timestamp 1606120353
transform 1 0 12420 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_878
timestamp 1606120353
transform 1 0 15180 0 -1 74528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_132_139
timestamp 1606120353
transform 1 0 13892 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_132_151
timestamp 1606120353
transform 1 0 14996 0 -1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_132_154
timestamp 1606120353
transform 1 0 15272 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_133_135
timestamp 1606120353
transform 1 0 13524 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_133_147
timestamp 1606120353
transform 1 0 14628 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_132_166
timestamp 1606120353
transform 1 0 16376 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_133_159
timestamp 1606120353
transform 1 0 15732 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_133_171
timestamp 1606120353
transform 1 0 16836 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_133_184
timestamp 1606120353
transform 1 0 18032 0 1 74528
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_883
timestamp 1606120353
transform 1 0 17940 0 1 74528
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_133_192
timestamp 1606120353
transform 1 0 18768 0 1 74528
box 0 -48 92 592
use sky130_fd_sc_hd__fill_1  FILLER_132_194
timestamp 1606120353
transform 1 0 18952 0 -1 74528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_132_190
timestamp 1606120353
transform 1 0 18584 0 -1 74528
box 0 -48 368 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__CLK
timestamp 1606120353
transform 1 0 19044 0 -1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__D
timestamp 1606120353
transform 1 0 18860 0 1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_132_197
timestamp 1606120353
transform 1 0 19228 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_132_178
timestamp 1606120353
transform 1 0 17480 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1170_
timestamp 1606120353
transform 1 0 19044 0 1 74528
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_879
timestamp 1606120353
transform 1 0 20792 0 -1 74528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_132_209
timestamp 1606120353
transform 1 0 20332 0 -1 74528
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_132_213
timestamp 1606120353
transform 1 0 20700 0 -1 74528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_132_215
timestamp 1606120353
transform 1 0 20884 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_133_214
timestamp 1606120353
transform 1 0 20792 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_132_227
timestamp 1606120353
transform 1 0 21988 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_132_239
timestamp 1606120353
transform 1 0 23092 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_133_226
timestamp 1606120353
transform 1 0 21896 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_133_238
timestamp 1606120353
transform 1 0 23000 0 1 74528
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_884
timestamp 1606120353
transform 1 0 23552 0 1 74528
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__D
timestamp 1606120353
transform 1 0 23828 0 1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__CLK
timestamp 1606120353
transform 1 0 24196 0 1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_132_251
timestamp 1606120353
transform 1 0 24196 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_132_263
timestamp 1606120353
transform 1 0 25300 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_133_245
timestamp 1606120353
transform 1 0 23644 0 1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_133_249
timestamp 1606120353
transform 1 0 24012 0 1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_133_253
timestamp 1606120353
transform 1 0 24380 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_880
timestamp 1606120353
transform 1 0 26404 0 -1 74528
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_132_276
timestamp 1606120353
transform 1 0 26496 0 -1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_133_265
timestamp 1606120353
transform 1 0 25484 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_133_277
timestamp 1606120353
transform 1 0 26588 0 1 74528
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_265
timestamp 1606120353
transform -1 0 28888 0 -1 74528
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_267
timestamp 1606120353
transform -1 0 28888 0 1 74528
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_132_288
timestamp 1606120353
transform 1 0 27600 0 -1 74528
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_132_296
timestamp 1606120353
transform 1 0 28336 0 -1 74528
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_133_289
timestamp 1606120353
transform 1 0 27692 0 1 74528
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_133_297
timestamp 1606120353
transform 1 0 28428 0 1 74528
box 0 -48 184 592
use sky130_fd_sc_hd__decap_3  PHY_268
timestamp 1606120353
transform 1 0 1104 0 -1 75616
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_134_3
timestamp 1606120353
transform 1 0 1380 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_134_15
timestamp 1606120353
transform 1 0 2484 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_885
timestamp 1606120353
transform 1 0 3956 0 -1 75616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_134_27
timestamp 1606120353
transform 1 0 3588 0 -1 75616
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_134_32
timestamp 1606120353
transform 1 0 4048 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_134_44
timestamp 1606120353
transform 1 0 5152 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_134_56
timestamp 1606120353
transform 1 0 6256 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_134_68
timestamp 1606120353
transform 1 0 7360 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_134_80
timestamp 1606120353
transform 1 0 8464 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1224_
timestamp 1606120353
transform 1 0 10396 0 -1 75616
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_886
timestamp 1606120353
transform 1 0 9568 0 -1 75616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_134_93
timestamp 1606120353
transform 1 0 9660 0 -1 75616
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_134_120
timestamp 1606120353
transform 1 0 12144 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_134_132
timestamp 1606120353
transform 1 0 13248 0 -1 75616
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_887
timestamp 1606120353
transform 1 0 15180 0 -1 75616
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__CLK
timestamp 1606120353
transform 1 0 13524 0 -1 75616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_134_137
timestamp 1606120353
transform 1 0 13708 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_4  FILLER_134_149
timestamp 1606120353
transform 1 0 14812 0 -1 75616
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_134_154
timestamp 1606120353
transform 1 0 15272 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_134_166
timestamp 1606120353
transform 1 0 16376 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_134_178
timestamp 1606120353
transform 1 0 17480 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_134_190
timestamp 1606120353
transform 1 0 18584 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_888
timestamp 1606120353
transform 1 0 20792 0 -1 75616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_134_202
timestamp 1606120353
transform 1 0 19688 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_134_215
timestamp 1606120353
transform 1 0 20884 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_134_227
timestamp 1606120353
transform 1 0 21988 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_134_239
timestamp 1606120353
transform 1 0 23092 0 -1 75616
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1198_
timestamp 1606120353
transform 1 0 23644 0 -1 75616
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_8  FILLER_134_264
timestamp 1606120353
transform 1 0 25392 0 -1 75616
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_889
timestamp 1606120353
transform 1 0 26404 0 -1 75616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_3  FILLER_134_272
timestamp 1606120353
transform 1 0 26128 0 -1 75616
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_134_276
timestamp 1606120353
transform 1 0 26496 0 -1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_269
timestamp 1606120353
transform -1 0 28888 0 -1 75616
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_134_288
timestamp 1606120353
transform 1 0 27600 0 -1 75616
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_134_296
timestamp 1606120353
transform 1 0 28336 0 -1 75616
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_270
timestamp 1606120353
transform 1 0 1104 0 1 75616
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_135_3
timestamp 1606120353
transform 1 0 1380 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_135_15
timestamp 1606120353
transform 1 0 2484 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_135_27
timestamp 1606120353
transform 1 0 3588 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_135_39
timestamp 1606120353
transform 1 0 4692 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_890
timestamp 1606120353
transform 1 0 6716 0 1 75616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_135_51
timestamp 1606120353
transform 1 0 5796 0 1 75616
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_135_59
timestamp 1606120353
transform 1 0 6532 0 1 75616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_135_62
timestamp 1606120353
transform 1 0 6808 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_135_74
timestamp 1606120353
transform 1 0 7912 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_135_86
timestamp 1606120353
transform 1 0 9016 0 1 75616
box 0 -48 552 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__D
timestamp 1606120353
transform 1 0 9660 0 1 75616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__CLK
timestamp 1606120353
transform 1 0 10028 0 1 75616
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_135_92
timestamp 1606120353
transform 1 0 9568 0 1 75616
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_135_95
timestamp 1606120353
transform 1 0 9844 0 1 75616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_135_99
timestamp 1606120353
transform 1 0 10212 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_891
timestamp 1606120353
transform 1 0 12328 0 1 75616
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__D
timestamp 1606120353
transform 1 0 12144 0 1 75616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__CLK
timestamp 1606120353
transform 1 0 12604 0 1 75616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_8  FILLER_135_111
timestamp 1606120353
transform 1 0 11316 0 1 75616
box 0 -48 736 592
use sky130_fd_sc_hd__fill_1  FILLER_135_119
timestamp 1606120353
transform 1 0 12052 0 1 75616
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_135_123
timestamp 1606120353
transform 1 0 12420 0 1 75616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_135_127
timestamp 1606120353
transform 1 0 12788 0 1 75616
box 0 -48 552 592
use sky130_fd_sc_hd__dfxtp_4  _1220_
timestamp 1606120353
transform 1 0 13524 0 1 75616
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__D
timestamp 1606120353
transform 1 0 13340 0 1 75616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_135_154
timestamp 1606120353
transform 1 0 15272 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_135_166
timestamp 1606120353
transform 1 0 16376 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_892
timestamp 1606120353
transform 1 0 17940 0 1 75616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_135_178
timestamp 1606120353
transform 1 0 17480 0 1 75616
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_135_182
timestamp 1606120353
transform 1 0 17848 0 1 75616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_135_184
timestamp 1606120353
transform 1 0 18032 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_135_196
timestamp 1606120353
transform 1 0 19136 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__D
timestamp 1606120353
transform 1 0 20884 0 1 75616
box 0 -48 184 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__CLK
timestamp 1606120353
transform 1 0 21252 0 1 75616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_6  FILLER_135_208
timestamp 1606120353
transform 1 0 20240 0 1 75616
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_135_214
timestamp 1606120353
transform 1 0 20792 0 1 75616
box 0 -48 92 592
use sky130_fd_sc_hd__fill_2  FILLER_135_217
timestamp 1606120353
transform 1 0 21068 0 1 75616
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_135_221
timestamp 1606120353
transform 1 0 21436 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_135_233
timestamp 1606120353
transform 1 0 22540 0 1 75616
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_135_241
timestamp 1606120353
transform 1 0 23276 0 1 75616
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_893
timestamp 1606120353
transform 1 0 23552 0 1 75616
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_135_245
timestamp 1606120353
transform 1 0 23644 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_135_257
timestamp 1606120353
transform 1 0 24748 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_135_269
timestamp 1606120353
transform 1 0 25852 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_135_281
timestamp 1606120353
transform 1 0 26956 0 1 75616
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_271
timestamp 1606120353
transform -1 0 28888 0 1 75616
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_135_293
timestamp 1606120353
transform 1 0 28060 0 1 75616
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_272
timestamp 1606120353
transform 1 0 1104 0 -1 76704
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_136_3
timestamp 1606120353
transform 1 0 1380 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_136_15
timestamp 1606120353
transform 1 0 2484 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_894
timestamp 1606120353
transform 1 0 3956 0 -1 76704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_136_27
timestamp 1606120353
transform 1 0 3588 0 -1 76704
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_136_32
timestamp 1606120353
transform 1 0 4048 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_136_44
timestamp 1606120353
transform 1 0 5152 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_136_56
timestamp 1606120353
transform 1 0 6256 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_136_68
timestamp 1606120353
transform 1 0 7360 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_136_80
timestamp 1606120353
transform 1 0 8464 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1128_
timestamp 1606120353
transform 1 0 9660 0 -1 76704
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_895
timestamp 1606120353
transform 1 0 9568 0 -1 76704
box 0 -48 92 592
use sky130_fd_sc_hd__dfxtp_4  _1177_
timestamp 1606120353
transform 1 0 12144 0 -1 76704
box 0 -48 1748 592
use sky130_fd_sc_hd__decap_8  FILLER_136_112
timestamp 1606120353
transform 1 0 11408 0 -1 76704
box 0 -48 736 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_896
timestamp 1606120353
transform 1 0 15180 0 -1 76704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_136_139
timestamp 1606120353
transform 1 0 13892 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_136_151
timestamp 1606120353
transform 1 0 14996 0 -1 76704
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_136_154
timestamp 1606120353
transform 1 0 15272 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_136_166
timestamp 1606120353
transform 1 0 16376 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__CLK
timestamp 1606120353
transform 1 0 19320 0 -1 76704
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_136_178
timestamp 1606120353
transform 1 0 17480 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_8  FILLER_136_190
timestamp 1606120353
transform 1 0 18584 0 -1 76704
box 0 -48 736 592
use sky130_fd_sc_hd__dfxtp_4  _1171_
timestamp 1606120353
transform 1 0 20884 0 -1 76704
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_897
timestamp 1606120353
transform 1 0 20792 0 -1 76704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_136_200
timestamp 1606120353
transform 1 0 19504 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__fill_2  FILLER_136_212
timestamp 1606120353
transform 1 0 20608 0 -1 76704
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_136_234
timestamp 1606120353
transform 1 0 22632 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_136_246
timestamp 1606120353
transform 1 0 23736 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_136_258
timestamp 1606120353
transform 1 0 24840 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_898
timestamp 1606120353
transform 1 0 26404 0 -1 76704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_136_270
timestamp 1606120353
transform 1 0 25944 0 -1 76704
box 0 -48 368 592
use sky130_fd_sc_hd__fill_1  FILLER_136_274
timestamp 1606120353
transform 1 0 26312 0 -1 76704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_136_276
timestamp 1606120353
transform 1 0 26496 0 -1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_273
timestamp 1606120353
transform -1 0 28888 0 -1 76704
box 0 -48 276 592
use sky130_fd_sc_hd__decap_8  FILLER_136_288
timestamp 1606120353
transform 1 0 27600 0 -1 76704
box 0 -48 736 592
use sky130_fd_sc_hd__decap_3  FILLER_136_296
timestamp 1606120353
transform 1 0 28336 0 -1 76704
box 0 -48 276 592
use sky130_fd_sc_hd__decap_3  PHY_274
timestamp 1606120353
transform 1 0 1104 0 1 76704
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_137_3
timestamp 1606120353
transform 1 0 1380 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_137_15
timestamp 1606120353
transform 1 0 2484 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_137_27
timestamp 1606120353
transform 1 0 3588 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_137_39
timestamp 1606120353
transform 1 0 4692 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_899
timestamp 1606120353
transform 1 0 6716 0 1 76704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_8  FILLER_137_51
timestamp 1606120353
transform 1 0 5796 0 1 76704
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_137_59
timestamp 1606120353
transform 1 0 6532 0 1 76704
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_137_62
timestamp 1606120353
transform 1 0 6808 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_137_74
timestamp 1606120353
transform 1 0 7912 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_137_86
timestamp 1606120353
transform 1 0 9016 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_137_98
timestamp 1606120353
transform 1 0 10120 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_137_110
timestamp 1606120353
transform 1 0 11224 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_900
timestamp 1606120353
transform 1 0 12328 0 1 76704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_137_123
timestamp 1606120353
transform 1 0 12420 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1226_
timestamp 1606120353
transform 1 0 13800 0 1 76704
box 0 -48 1748 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__D
timestamp 1606120353
transform 1 0 13616 0 1 76704
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_137_135
timestamp 1606120353
transform 1 0 13524 0 1 76704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_137_157
timestamp 1606120353
transform 1 0 15548 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_137_169
timestamp 1606120353
transform 1 0 16652 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__dfxtp_4  _1182_
timestamp 1606120353
transform 1 0 19320 0 1 76704
box 0 -48 1748 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_901
timestamp 1606120353
transform 1 0 17940 0 1 76704
box 0 -48 92 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__D
timestamp 1606120353
transform 1 0 19136 0 1 76704
box 0 -48 184 592
use sky130_fd_sc_hd__fill_2  FILLER_137_181
timestamp 1606120353
transform 1 0 17756 0 1 76704
box 0 -48 184 592
use sky130_fd_sc_hd__decap_12  FILLER_137_184
timestamp 1606120353
transform 1 0 18032 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_137_217
timestamp 1606120353
transform 1 0 21068 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_137_229
timestamp 1606120353
transform 1 0 22172 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_137_241
timestamp 1606120353
transform 1 0 23276 0 1 76704
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_902
timestamp 1606120353
transform 1 0 23552 0 1 76704
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_137_245
timestamp 1606120353
transform 1 0 23644 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_137_257
timestamp 1606120353
transform 1 0 24748 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_137_269
timestamp 1606120353
transform 1 0 25852 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_137_281
timestamp 1606120353
transform 1 0 26956 0 1 76704
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_275
timestamp 1606120353
transform -1 0 28888 0 1 76704
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_137_293
timestamp 1606120353
transform 1 0 28060 0 1 76704
box 0 -48 552 592
use sky130_fd_sc_hd__decap_3  PHY_276
timestamp 1606120353
transform 1 0 1104 0 -1 77792
box 0 -48 276 592
use sky130_fd_sc_hd__decap_12  FILLER_138_3
timestamp 1606120353
transform 1 0 1380 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_138_15
timestamp 1606120353
transform 1 0 2484 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_903
timestamp 1606120353
transform 1 0 3956 0 -1 77792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_4  FILLER_138_27
timestamp 1606120353
transform 1 0 3588 0 -1 77792
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_138_32
timestamp 1606120353
transform 1 0 4048 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_138_44
timestamp 1606120353
transform 1 0 5152 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_904
timestamp 1606120353
transform 1 0 6808 0 -1 77792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_138_56
timestamp 1606120353
transform 1 0 6256 0 -1 77792
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_138_63
timestamp 1606120353
transform 1 0 6900 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_138_75
timestamp 1606120353
transform 1 0 8004 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_138_87
timestamp 1606120353
transform 1 0 9108 0 -1 77792
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_905
timestamp 1606120353
transform 1 0 9660 0 -1 77792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_138_94
timestamp 1606120353
transform 1 0 9752 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_138_106
timestamp 1606120353
transform 1 0 10856 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_906
timestamp 1606120353
transform 1 0 12512 0 -1 77792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_138_118
timestamp 1606120353
transform 1 0 11960 0 -1 77792
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_138_125
timestamp 1606120353
transform 1 0 12604 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__CLK
timestamp 1606120353
transform 1 0 13800 0 -1 77792
box 0 -48 184 592
use sky130_fd_sc_hd__fill_1  FILLER_138_137
timestamp 1606120353
transform 1 0 13708 0 -1 77792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_138_140
timestamp 1606120353
transform 1 0 13984 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  FILLER_138_152
timestamp 1606120353
transform 1 0 15088 0 -1 77792
box 0 -48 276 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_907
timestamp 1606120353
transform 1 0 15364 0 -1 77792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_138_156
timestamp 1606120353
transform 1 0 15456 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_138_168
timestamp 1606120353
transform 1 0 16560 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_908
timestamp 1606120353
transform 1 0 18216 0 -1 77792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_138_180
timestamp 1606120353
transform 1 0 17664 0 -1 77792
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_138_187
timestamp 1606120353
transform 1 0 18308 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_909
timestamp 1606120353
transform 1 0 21068 0 -1 77792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_138_199
timestamp 1606120353
transform 1 0 19412 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_138_211
timestamp 1606120353
transform 1 0 20516 0 -1 77792
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_138_218
timestamp 1606120353
transform 1 0 21160 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_138_230
timestamp 1606120353
transform 1 0 22264 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_6  FILLER_138_242
timestamp 1606120353
transform 1 0 23368 0 -1 77792
box 0 -48 552 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_910
timestamp 1606120353
transform 1 0 23920 0 -1 77792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_12  FILLER_138_249
timestamp 1606120353
transform 1 0 24012 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_138_261
timestamp 1606120353
transform 1 0 25116 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_911
timestamp 1606120353
transform 1 0 26772 0 -1 77792
box 0 -48 92 592
use sky130_fd_sc_hd__decap_6  FILLER_138_273
timestamp 1606120353
transform 1 0 26220 0 -1 77792
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_138_280
timestamp 1606120353
transform 1 0 26864 0 -1 77792
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_3  PHY_277
timestamp 1606120353
transform -1 0 28888 0 -1 77792
box 0 -48 276 592
use sky130_fd_sc_hd__decap_6  FILLER_138_292
timestamp 1606120353
transform 1 0 27968 0 -1 77792
box 0 -48 552 592
use sky130_fd_sc_hd__fill_1  FILLER_138_298
timestamp 1606120353
transform 1 0 28520 0 -1 77792
box 0 -48 92 592
<< labels >>
rlabel metal3 s 29200 11568 30000 11688 6 addr_r[0]
port 0 nsew default input
rlabel metal3 s 29200 72088 30000 72208 6 addr_r[10]
port 1 nsew default input
rlabel metal3 s 29200 40128 30000 40248 6 addr_r[11]
port 2 nsew default input
rlabel metal2 s 11058 79200 11114 80000 6 addr_r[12]
port 3 nsew default input
rlabel metal3 s 29200 63248 30000 63368 6 addr_r[13]
port 4 nsew default input
rlabel metal3 s 0 43528 800 43648 6 addr_r[1]
port 5 nsew default input
rlabel metal2 s 9678 79200 9734 80000 6 addr_r[2]
port 6 nsew default input
rlabel metal2 s 28078 0 28134 800 6 addr_r[3]
port 7 nsew default input
rlabel metal3 s 0 26528 800 26648 6 addr_r[4]
port 8 nsew default input
rlabel metal3 s 0 66648 800 66768 6 addr_r[5]
port 9 nsew default input
rlabel metal3 s 0 7488 800 7608 6 addr_r[6]
port 10 nsew default input
rlabel metal3 s 0 13608 800 13728 6 addr_r[7]
port 11 nsew default input
rlabel metal2 s 9218 0 9274 800 6 addr_r[8]
port 12 nsew default input
rlabel metal3 s 0 59848 800 59968 6 addr_r[9]
port 13 nsew default input
rlabel metal2 s 25318 0 25374 800 6 addr_w[0]
port 14 nsew default input
rlabel metal3 s 0 10208 800 10328 6 addr_w[10]
port 15 nsew default input
rlabel metal3 s 0 50328 800 50448 6 addr_w[11]
port 16 nsew default input
rlabel metal3 s 29200 8848 30000 8968 6 addr_w[12]
port 17 nsew default input
rlabel metal2 s 14738 0 14794 800 6 addr_w[13]
port 18 nsew default input
rlabel metal2 s 19338 0 19394 800 6 addr_w[1]
port 19 nsew default input
rlabel metal3 s 29200 34688 30000 34808 6 addr_w[2]
port 20 nsew default input
rlabel metal3 s 29200 8 30000 128 6 addr_w[3]
port 21 nsew default input
rlabel metal3 s 29200 15648 30000 15768 6 addr_w[4]
port 22 nsew default input
rlabel metal3 s 0 70048 800 70168 6 addr_w[5]
port 23 nsew default input
rlabel metal3 s 0 2048 800 2168 6 addr_w[6]
port 24 nsew default input
rlabel metal2 s 3698 0 3754 800 6 addr_w[7]
port 25 nsew default input
rlabel metal3 s 0 53728 800 53848 6 addr_w[8]
port 26 nsew default input
rlabel metal3 s 0 51688 800 51808 6 addr_w[9]
port 27 nsew default input
rlabel metal3 s 29200 49648 30000 49768 6 baseaddr_r_sync[0]
port 28 nsew default tristate
rlabel metal2 s 14738 79200 14794 80000 6 baseaddr_r_sync[1]
port 29 nsew default tristate
rlabel metal3 s 29200 21768 30000 21888 6 baseaddr_r_sync[2]
port 30 nsew default tristate
rlabel metal2 s 17958 0 18014 800 6 baseaddr_r_sync[3]
port 31 nsew default tristate
rlabel metal3 s 29200 30608 30000 30728 6 baseaddr_r_sync[4]
port 32 nsew default tristate
rlabel metal2 s 20258 0 20314 800 6 baseaddr_r_sync[5]
port 33 nsew default tristate
rlabel metal3 s 29200 26528 30000 26648 6 baseaddr_r_sync[6]
port 34 nsew default tristate
rlabel metal3 s 0 61888 800 62008 6 baseaddr_r_sync[7]
port 35 nsew default tristate
rlabel metal2 s 16578 79200 16634 80000 6 baseaddr_r_sync[8]
port 36 nsew default tristate
rlabel metal3 s 0 76848 800 76968 6 baseaddr_w_sync[0]
port 37 nsew default tristate
rlabel metal3 s 29200 73448 30000 73568 6 baseaddr_w_sync[1]
port 38 nsew default tristate
rlabel metal2 s 5998 0 6054 800 6 baseaddr_w_sync[2]
port 39 nsew default tristate
rlabel metal3 s 0 71408 800 71528 6 baseaddr_w_sync[3]
port 40 nsew default tristate
rlabel metal2 s 938 79200 994 80000 6 baseaddr_w_sync[4]
port 41 nsew default tristate
rlabel metal2 s 23478 79200 23534 80000 6 baseaddr_w_sync[5]
port 42 nsew default tristate
rlabel metal2 s 24858 0 24914 800 6 baseaddr_w_sync[6]
port 43 nsew default tristate
rlabel metal3 s 0 33328 800 33448 6 baseaddr_w_sync[7]
port 44 nsew default tristate
rlabel metal3 s 29200 12248 30000 12368 6 baseaddr_w_sync[8]
port 45 nsew default tristate
rlabel metal3 s 0 22448 800 22568 6 clk
port 46 nsew default input
rlabel metal2 s 14278 79200 14334 80000 6 conf[0]
port 47 nsew default input
rlabel metal2 s 18418 0 18474 800 6 conf[1]
port 48 nsew default input
rlabel metal3 s 29200 45568 30000 45688 6 conf[2]
port 49 nsew default input
rlabel metal3 s 29200 19048 30000 19168 6 csb
port 50 nsew default input
rlabel metal2 s 27618 79200 27674 80000 6 csb0_sync
port 51 nsew default tristate
rlabel metal3 s 0 58488 800 58608 6 csb1_sync
port 52 nsew default tristate
rlabel metal3 s 29200 13608 30000 13728 6 d_fabric_in[0]
port 53 nsew default input
rlabel metal3 s 29200 2048 30000 2168 6 d_fabric_in[10]
port 54 nsew default input
rlabel metal2 s 10138 79200 10194 80000 6 d_fabric_in[11]
port 55 nsew default input
rlabel metal3 s 29200 78208 30000 78328 6 d_fabric_in[12]
port 56 nsew default input
rlabel metal3 s 0 30608 800 30728 6 d_fabric_in[13]
port 57 nsew default input
rlabel metal3 s 0 688 800 808 6 d_fabric_in[14]
port 58 nsew default input
rlabel metal3 s 0 63928 800 64048 6 d_fabric_in[15]
port 59 nsew default input
rlabel metal2 s 17498 79200 17554 80000 6 d_fabric_in[16]
port 60 nsew default input
rlabel metal3 s 29200 76848 30000 76968 6 d_fabric_in[17]
port 61 nsew default input
rlabel metal3 s 29200 66648 30000 66768 6 d_fabric_in[18]
port 62 nsew default input
rlabel metal2 s 28078 79200 28134 80000 6 d_fabric_in[19]
port 63 nsew default input
rlabel metal3 s 0 6808 800 6928 6 d_fabric_in[1]
port 64 nsew default input
rlabel metal2 s 20718 0 20774 800 6 d_fabric_in[20]
port 65 nsew default input
rlabel metal3 s 29200 64608 30000 64728 6 d_fabric_in[21]
port 66 nsew default input
rlabel metal3 s 29200 14968 30000 15088 6 d_fabric_in[22]
port 67 nsew default input
rlabel metal3 s 29200 56448 30000 56568 6 d_fabric_in[23]
port 68 nsew default input
rlabel metal3 s 0 37408 800 37528 6 d_fabric_in[24]
port 69 nsew default input
rlabel metal2 s 20258 79200 20314 80000 6 d_fabric_in[25]
port 70 nsew default input
rlabel metal3 s 0 72088 800 72208 6 d_fabric_in[26]
port 71 nsew default input
rlabel metal3 s 0 57128 800 57248 6 d_fabric_in[27]
port 72 nsew default input
rlabel metal3 s 29200 53048 30000 53168 6 d_fabric_in[28]
port 73 nsew default input
rlabel metal3 s 29200 59848 30000 59968 6 d_fabric_in[29]
port 74 nsew default input
rlabel metal2 s 27158 0 27214 800 6 d_fabric_in[2]
port 75 nsew default input
rlabel metal3 s 29200 20408 30000 20528 6 d_fabric_in[30]
port 76 nsew default input
rlabel metal3 s 0 41488 800 41608 6 d_fabric_in[31]
port 77 nsew default input
rlabel metal3 s 29200 5448 30000 5568 6 d_fabric_in[3]
port 78 nsew default input
rlabel metal2 s 17958 79200 18014 80000 6 d_fabric_in[4]
port 79 nsew default input
rlabel metal2 s 13358 79200 13414 80000 6 d_fabric_in[5]
port 80 nsew default input
rlabel metal3 s 0 44888 800 45008 6 d_fabric_in[6]
port 81 nsew default input
rlabel metal3 s 29200 79568 30000 79688 6 d_fabric_in[7]
port 82 nsew default input
rlabel metal3 s 0 45568 800 45688 6 d_fabric_in[8]
port 83 nsew default input
rlabel metal2 s 1398 0 1454 800 6 d_fabric_in[9]
port 84 nsew default input
rlabel metal2 s 12898 0 12954 800 6 d_fabric_out[0]
port 85 nsew default tristate
rlabel metal3 s 0 3408 800 3528 6 d_fabric_out[10]
port 86 nsew default tristate
rlabel metal3 s 29200 688 30000 808 6 d_fabric_out[11]
port 87 nsew default tristate
rlabel metal3 s 29200 70048 30000 70168 6 d_fabric_out[12]
port 88 nsew default tristate
rlabel metal2 s 15198 0 15254 800 6 d_fabric_out[13]
port 89 nsew default tristate
rlabel metal3 s 29200 3408 30000 3528 6 d_fabric_out[14]
port 90 nsew default tristate
rlabel metal2 s 1858 79200 1914 80000 6 d_fabric_out[15]
port 91 nsew default tristate
rlabel metal3 s 29200 58488 30000 58608 6 d_fabric_out[16]
port 92 nsew default tristate
rlabel metal2 s 12438 79200 12494 80000 6 d_fabric_out[17]
port 93 nsew default tristate
rlabel metal2 s 26238 0 26294 800 6 d_fabric_out[18]
port 94 nsew default tristate
rlabel metal3 s 29200 31968 30000 32088 6 d_fabric_out[19]
port 95 nsew default tristate
rlabel metal2 s 29458 0 29514 800 6 d_fabric_out[1]
port 96 nsew default tristate
rlabel metal2 s 13818 0 13874 800 6 d_fabric_out[20]
port 97 nsew default tristate
rlabel metal3 s 0 28568 800 28688 6 d_fabric_out[21]
port 98 nsew default tristate
rlabel metal3 s 0 27208 800 27328 6 d_fabric_out[22]
port 99 nsew default tristate
rlabel metal3 s 0 21768 800 21888 6 d_fabric_out[23]
port 100 nsew default tristate
rlabel metal3 s 29200 46928 30000 47048 6 d_fabric_out[24]
port 101 nsew default tristate
rlabel metal3 s 0 4088 800 4208 6 d_fabric_out[25]
port 102 nsew default tristate
rlabel metal3 s 0 8848 800 8968 6 d_fabric_out[26]
port 103 nsew default tristate
rlabel metal3 s 0 14968 800 15088 6 d_fabric_out[27]
port 104 nsew default tristate
rlabel metal2 s 2318 79200 2374 80000 6 d_fabric_out[28]
port 105 nsew default tristate
rlabel metal3 s 0 48288 800 48408 6 d_fabric_out[29]
port 106 nsew default tristate
rlabel metal3 s 0 78208 800 78328 6 d_fabric_out[2]
port 107 nsew default tristate
rlabel metal2 s 5538 79200 5594 80000 6 d_fabric_out[30]
port 108 nsew default tristate
rlabel metal2 s 29918 79200 29974 80000 6 d_fabric_out[31]
port 109 nsew default tristate
rlabel metal2 s 21178 79200 21234 80000 6 d_fabric_out[3]
port 110 nsew default tristate
rlabel metal3 s 29200 6808 30000 6928 6 d_fabric_out[4]
port 111 nsew default tristate
rlabel metal3 s 29200 68688 30000 68808 6 d_fabric_out[5]
port 112 nsew default tristate
rlabel metal3 s 29200 65288 30000 65408 6 d_fabric_out[6]
port 113 nsew default tristate
rlabel metal3 s 29200 53728 30000 53848 6 d_fabric_out[7]
port 114 nsew default tristate
rlabel metal3 s 0 25168 800 25288 6 d_fabric_out[8]
port 115 nsew default tristate
rlabel metal3 s 0 46928 800 47048 6 d_fabric_out[9]
port 116 nsew default tristate
rlabel metal2 s 478 0 534 800 6 d_sram_in[0]
port 117 nsew default tristate
rlabel metal3 s 29200 43528 30000 43648 6 d_sram_in[10]
port 118 nsew default tristate
rlabel metal3 s 29200 42168 30000 42288 6 d_sram_in[11]
port 119 nsew default tristate
rlabel metal2 s 6458 79200 6514 80000 6 d_sram_in[12]
port 120 nsew default tristate
rlabel metal3 s 0 55088 800 55208 6 d_sram_in[13]
port 121 nsew default tristate
rlabel metal3 s 0 5448 800 5568 6 d_sram_in[14]
port 122 nsew default tristate
rlabel metal3 s 0 31968 800 32088 6 d_sram_in[15]
port 123 nsew default tristate
rlabel metal3 s 29200 38088 30000 38208 6 d_sram_in[16]
port 124 nsew default tristate
rlabel metal3 s 29200 28568 30000 28688 6 d_sram_in[17]
port 125 nsew default tristate
rlabel metal2 s 2318 0 2374 800 6 d_sram_in[18]
port 126 nsew default tristate
rlabel metal3 s 29200 74808 30000 74928 6 d_sram_in[19]
port 127 nsew default tristate
rlabel metal3 s 0 79568 800 79688 6 d_sram_in[1]
port 128 nsew default tristate
rlabel metal3 s 0 68008 800 68128 6 d_sram_in[20]
port 129 nsew default tristate
rlabel metal3 s 29200 61888 30000 62008 6 d_sram_in[21]
port 130 nsew default tristate
rlabel metal2 s 17038 0 17094 800 6 d_sram_in[22]
port 131 nsew default tristate
rlabel metal2 s 21638 0 21694 800 6 d_sram_in[23]
port 132 nsew default tristate
rlabel metal3 s 29200 23128 30000 23248 6 d_sram_in[24]
port 133 nsew default tristate
rlabel metal2 s 25778 79200 25834 80000 6 d_sram_in[25]
port 134 nsew default tristate
rlabel metal2 s 8298 0 8354 800 6 d_sram_in[26]
port 135 nsew default tristate
rlabel metal3 s 0 75488 800 75608 6 d_sram_in[27]
port 136 nsew default tristate
rlabel metal3 s 0 38768 800 38888 6 d_sram_in[28]
port 137 nsew default tristate
rlabel metal3 s 29200 23808 30000 23928 6 d_sram_in[29]
port 138 nsew default tristate
rlabel metal2 s 6918 0 6974 800 6 d_sram_in[2]
port 139 nsew default tristate
rlabel metal2 s 6918 79200 6974 80000 6 d_sram_in[30]
port 140 nsew default tristate
rlabel metal3 s 29200 35368 30000 35488 6 d_sram_in[31]
port 141 nsew default tristate
rlabel metal3 s 0 53048 800 53168 6 d_sram_in[3]
port 142 nsew default tristate
rlabel metal2 s 3238 79200 3294 80000 6 d_sram_in[4]
port 143 nsew default tristate
rlabel metal3 s 29200 41488 30000 41608 6 d_sram_in[5]
port 144 nsew default tristate
rlabel metal3 s 0 65288 800 65408 6 d_sram_in[6]
port 145 nsew default tristate
rlabel metal3 s 29200 8168 30000 8288 6 d_sram_in[7]
port 146 nsew default tristate
rlabel metal3 s 29200 4088 30000 4208 6 d_sram_in[8]
port 147 nsew default tristate
rlabel metal3 s 29200 44888 30000 45008 6 d_sram_in[9]
port 148 nsew default tristate
rlabel metal3 s 0 35368 800 35488 6 d_sram_out[0]
port 149 nsew default input
rlabel metal2 s 10138 0 10194 800 6 d_sram_out[10]
port 150 nsew default input
rlabel metal3 s 0 36728 800 36848 6 d_sram_out[11]
port 151 nsew default input
rlabel metal3 s 0 63248 800 63368 6 d_sram_out[12]
port 152 nsew default input
rlabel metal2 s 8758 79200 8814 80000 6 d_sram_out[13]
port 153 nsew default input
rlabel metal3 s 0 15648 800 15768 6 d_sram_out[14]
port 154 nsew default input
rlabel metal2 s 24398 79200 24454 80000 6 d_sram_out[15]
port 155 nsew default input
rlabel metal2 s 11518 0 11574 800 6 d_sram_out[16]
port 156 nsew default input
rlabel metal3 s 29200 76168 30000 76288 6 d_sram_out[17]
port 157 nsew default input
rlabel metal2 s 23938 0 23994 800 6 d_sram_out[18]
port 158 nsew default input
rlabel metal2 s 22098 79200 22154 80000 6 d_sram_out[19]
port 159 nsew default input
rlabel metal3 s 29200 61208 30000 61328 6 d_sram_out[1]
port 160 nsew default input
rlabel metal3 s 29200 27208 30000 27328 6 d_sram_out[20]
port 161 nsew default input
rlabel metal3 s 0 17008 800 17128 6 d_sram_out[21]
port 162 nsew default input
rlabel metal2 s 2778 0 2834 800 6 d_sram_out[22]
port 163 nsew default input
rlabel metal2 s 22558 79200 22614 80000 6 d_sram_out[23]
port 164 nsew default input
rlabel metal3 s 29200 17008 30000 17128 6 d_sram_out[24]
port 165 nsew default input
rlabel metal3 s 0 12248 800 12368 6 d_sram_out[25]
port 166 nsew default input
rlabel metal2 s 24858 79200 24914 80000 6 d_sram_out[26]
port 167 nsew default input
rlabel metal3 s 29200 25168 30000 25288 6 d_sram_out[27]
port 168 nsew default input
rlabel metal2 s 12438 0 12494 800 6 d_sram_out[28]
port 169 nsew default input
rlabel metal2 s 28538 0 28594 800 6 d_sram_out[29]
port 170 nsew default input
rlabel metal3 s 29200 71408 30000 71528 6 d_sram_out[2]
port 171 nsew default input
rlabel metal3 s 0 40128 800 40248 6 d_sram_out[30]
port 172 nsew default input
rlabel metal3 s 0 48968 800 49088 6 d_sram_out[31]
port 173 nsew default input
rlabel metal3 s 29200 38768 30000 38888 6 d_sram_out[3]
port 174 nsew default input
rlabel metal2 s 10598 0 10654 800 6 d_sram_out[4]
port 175 nsew default input
rlabel metal2 s 4618 0 4674 800 6 d_sram_out[5]
port 176 nsew default input
rlabel metal3 s 29200 55088 30000 55208 6 d_sram_out[6]
port 177 nsew default input
rlabel metal3 s 0 60528 800 60648 6 d_sram_out[7]
port 178 nsew default input
rlabel metal3 s 0 29928 800 30048 6 d_sram_out[8]
port 179 nsew default input
rlabel metal3 s 0 20408 800 20528 6 d_sram_out[9]
port 180 nsew default input
rlabel metal2 s 18878 79200 18934 80000 6 out_reg
port 181 nsew default input
rlabel metal3 s 0 23808 800 23928 6 reb
port 182 nsew default input
rlabel metal3 s 29200 18368 30000 18488 6 w_mask[0]
port 183 nsew default tristate
rlabel metal2 s 4618 79200 4674 80000 6 w_mask[10]
port 184 nsew default tristate
rlabel metal3 s 29200 68008 30000 68128 6 w_mask[11]
port 185 nsew default tristate
rlabel metal2 s 18 0 74 800 6 w_mask[12]
port 186 nsew default tristate
rlabel metal3 s 0 19048 800 19168 6 w_mask[13]
port 187 nsew default tristate
rlabel metal2 s 16118 0 16174 800 6 w_mask[14]
port 188 nsew default tristate
rlabel metal2 s 7378 0 7434 800 6 w_mask[15]
port 189 nsew default tristate
rlabel metal2 s 19798 79200 19854 80000 6 w_mask[16]
port 190 nsew default tristate
rlabel metal2 s 28998 79200 29054 80000 6 w_mask[17]
port 191 nsew default tristate
rlabel metal3 s 29200 57128 30000 57248 6 w_mask[18]
port 192 nsew default tristate
rlabel metal2 s 23018 0 23074 800 6 w_mask[19]
port 193 nsew default tristate
rlabel metal3 s 29200 10208 30000 10328 6 w_mask[1]
port 194 nsew default tristate
rlabel metal3 s 0 74808 800 74928 6 w_mask[20]
port 195 nsew default tristate
rlabel metal3 s 0 56448 800 56568 6 w_mask[21]
port 196 nsew default tristate
rlabel metal2 s 15658 79200 15714 80000 6 w_mask[22]
port 197 nsew default tristate
rlabel metal3 s 0 10888 800 11008 6 w_mask[23]
port 198 nsew default tristate
rlabel metal2 s 5078 0 5134 800 6 w_mask[24]
port 199 nsew default tristate
rlabel metal3 s 0 42168 800 42288 6 w_mask[25]
port 200 nsew default tristate
rlabel metal2 s 11978 79200 12034 80000 6 w_mask[26]
port 201 nsew default tristate
rlabel metal3 s 0 73448 800 73568 6 w_mask[27]
port 202 nsew default tristate
rlabel metal2 s 7838 79200 7894 80000 6 w_mask[28]
port 203 nsew default tristate
rlabel metal2 s 26698 79200 26754 80000 6 w_mask[29]
port 204 nsew default tristate
rlabel metal2 s 18 79200 74 80000 6 w_mask[2]
port 205 nsew default tristate
rlabel metal2 s 22558 0 22614 800 6 w_mask[30]
port 206 nsew default tristate
rlabel metal3 s 0 18368 800 18488 6 w_mask[31]
port 207 nsew default tristate
rlabel metal3 s 29200 51688 30000 51808 6 w_mask[3]
port 208 nsew default tristate
rlabel metal3 s 29200 48288 30000 48408 6 w_mask[4]
port 209 nsew default tristate
rlabel metal2 s 4158 79200 4214 80000 6 w_mask[5]
port 210 nsew default tristate
rlabel metal3 s 29200 36728 30000 36848 6 w_mask[6]
port 211 nsew default tristate
rlabel metal3 s 29200 29928 30000 30048 6 w_mask[7]
port 212 nsew default tristate
rlabel metal3 s 29200 50328 30000 50448 6 w_mask[8]
port 213 nsew default tristate
rlabel metal3 s 29200 33328 30000 33448 6 w_mask[9]
port 214 nsew default tristate
rlabel metal3 s 0 68688 800 68808 6 web
port 215 nsew default input
rlabel metal3 s 0 34008 800 34128 6 web0_sync
port 216 nsew default tristate
rlabel metal5 s 1104 15301 28888 15621 6 VPWR
port 217 nsew default input
rlabel metal5 s 1104 28635 28888 28955 6 VGND
port 218 nsew default input
<< end >>
