magic
tech sky130A
magscale 1 2
timestamp 1607333050
<< locali >>
rect 22661 56899 22695 57001
rect 14105 55131 14139 55369
rect 17049 54655 17083 54825
rect 29561 48059 29595 48161
rect 12541 37179 12575 37417
rect 17877 35683 17911 35785
rect 12449 34935 12483 35173
rect 19349 33303 19383 33609
rect 20821 33371 20855 33473
rect 13277 31671 13311 31977
rect 14473 30039 14507 30141
rect 11437 29563 11471 29801
rect 20177 29495 20211 29801
rect 21833 29495 21867 29801
rect 21741 28475 21775 28645
rect 11621 27999 11655 28101
rect 21281 27999 21315 28169
rect 22109 27319 22143 27625
rect 22201 27387 22235 27625
rect 22385 26775 22419 27013
rect 20177 25687 20211 25925
rect 13093 24055 13127 24157
rect 21833 22967 21867 23205
<< viali >>
rect 24317 77537 24351 77571
rect 24041 77469 24075 77503
rect 18061 77333 18095 77367
rect 25605 77333 25639 77367
rect 29469 77333 29503 77367
rect 22661 77129 22695 77163
rect 24409 77129 24443 77163
rect 29101 77129 29135 77163
rect 31033 77129 31067 77163
rect 24133 77061 24167 77095
rect 15393 76993 15427 77027
rect 15761 76993 15795 77027
rect 17877 76993 17911 77027
rect 18337 76993 18371 77027
rect 24869 76993 24903 77027
rect 29745 76993 29779 77027
rect 15485 76925 15519 76959
rect 18061 76925 18095 76959
rect 21097 76925 21131 76959
rect 21373 76925 21407 76959
rect 24593 76925 24627 76959
rect 29469 76925 29503 76959
rect 17141 76857 17175 76891
rect 19441 76789 19475 76823
rect 20913 76789 20947 76823
rect 26157 76789 26191 76823
rect 21557 76449 21591 76483
rect 15577 76381 15611 76415
rect 17601 76381 17635 76415
rect 17877 76381 17911 76415
rect 21833 76381 21867 76415
rect 28825 76381 28859 76415
rect 29101 76381 29135 76415
rect 21189 76313 21223 76347
rect 18981 76245 19015 76279
rect 22937 76245 22971 76279
rect 24133 76245 24167 76279
rect 24685 76245 24719 76279
rect 30389 76245 30423 76279
rect 21649 76041 21683 76075
rect 28917 76041 28951 76075
rect 29469 75973 29503 76007
rect 18337 75905 18371 75939
rect 18889 75905 18923 75939
rect 19165 75837 19199 75871
rect 25697 75837 25731 75871
rect 25881 75837 25915 75871
rect 26157 75837 26191 75871
rect 18797 75769 18831 75803
rect 27537 75769 27571 75803
rect 17693 75701 17727 75735
rect 20269 75701 20303 75735
rect 22017 75701 22051 75735
rect 29837 75429 29871 75463
rect 30573 75361 30607 75395
rect 29745 75293 29779 75327
rect 30665 75293 30699 75327
rect 18981 75157 19015 75191
rect 25973 75157 26007 75191
rect 30389 74953 30423 74987
rect 19717 74817 19751 74851
rect 20085 74817 20119 74851
rect 19809 74749 19843 74783
rect 21189 74613 21223 74647
rect 29653 74613 29687 74647
rect 30113 74613 30147 74647
rect 19901 74341 19935 74375
rect 19533 72573 19567 72607
rect 19809 72573 19843 72607
rect 19349 72505 19383 72539
rect 21097 72437 21131 72471
rect 19533 71893 19567 71927
rect 22661 71009 22695 71043
rect 22937 71009 22971 71043
rect 24317 70941 24351 70975
rect 23029 70601 23063 70635
rect 22753 70465 22787 70499
rect 23949 69853 23983 69887
rect 24225 69853 24259 69887
rect 25329 69717 25363 69751
rect 24317 69513 24351 69547
rect 25973 69513 26007 69547
rect 24041 69445 24075 69479
rect 26157 69309 26191 69343
rect 26433 69241 26467 69275
rect 22845 68833 22879 68867
rect 25237 68833 25271 68867
rect 22569 68765 22603 68799
rect 23949 68629 23983 68663
rect 25053 68629 25087 68663
rect 22661 68425 22695 68459
rect 23949 68289 23983 68323
rect 24317 68289 24351 68323
rect 23029 68221 23063 68255
rect 24041 68221 24075 68255
rect 25697 68153 25731 68187
rect 24133 67609 24167 67643
rect 25145 67609 25179 67643
rect 26433 67337 26467 67371
rect 26617 67133 26651 67167
rect 26985 66997 27019 67031
rect 1777 65365 1811 65399
rect 1593 65161 1627 65195
rect 1777 65025 1811 65059
rect 2053 64957 2087 64991
rect 3433 64889 3467 64923
rect 1593 64277 1627 64311
rect 1869 63937 1903 63971
rect 4261 63937 4295 63971
rect 1593 63869 1627 63903
rect 3985 63869 4019 63903
rect 4169 63869 4203 63903
rect 4997 63869 5031 63903
rect 5089 63869 5123 63903
rect 3249 63801 3283 63835
rect 3617 63733 3651 63767
rect 1685 63529 1719 63563
rect 4261 63529 4295 63563
rect 4997 63393 5031 63427
rect 14105 63393 14139 63427
rect 21281 63393 21315 63427
rect 21741 63393 21775 63427
rect 4721 63325 4755 63359
rect 21097 63325 21131 63359
rect 13921 63257 13955 63291
rect 21741 63257 21775 63291
rect 6285 63189 6319 63223
rect 18705 63189 18739 63223
rect 19073 63189 19107 63223
rect 4721 62985 4755 63019
rect 20361 62985 20395 63019
rect 18613 62849 18647 62883
rect 18797 62849 18831 62883
rect 19809 62849 19843 62883
rect 22293 62849 22327 62883
rect 19073 62781 19107 62815
rect 19533 62781 19567 62815
rect 20729 62781 20763 62815
rect 21097 62781 21131 62815
rect 21373 62781 21407 62815
rect 21557 62781 21591 62815
rect 22017 62781 22051 62815
rect 5181 62645 5215 62679
rect 13921 62645 13955 62679
rect 18613 62305 18647 62339
rect 19073 62305 19107 62339
rect 26525 62305 26559 62339
rect 26801 62305 26835 62339
rect 18429 62237 18463 62271
rect 19073 62169 19107 62203
rect 21189 62101 21223 62135
rect 21557 62101 21591 62135
rect 22017 62101 22051 62135
rect 27905 62101 27939 62135
rect 18337 61897 18371 61931
rect 26617 61897 26651 61931
rect 26893 61829 26927 61863
rect 13369 61693 13403 61727
rect 13185 61557 13219 61591
rect 13737 61557 13771 61591
rect 18613 61557 18647 61591
rect 18981 61557 19015 61591
rect 21097 61557 21131 61591
rect 19901 61353 19935 61387
rect 10977 61217 11011 61251
rect 19717 61217 19751 61251
rect 20729 61217 20763 61251
rect 21649 61217 21683 61251
rect 21925 61217 21959 61251
rect 21281 61149 21315 61183
rect 19625 61081 19659 61115
rect 21925 61081 21959 61115
rect 10793 61013 10827 61047
rect 20177 61013 20211 61047
rect 22569 61013 22603 61047
rect 25329 61013 25363 61047
rect 10885 60809 10919 60843
rect 18981 60809 19015 60843
rect 21281 60809 21315 60843
rect 20637 60741 20671 60775
rect 25421 60673 25455 60707
rect 30849 60673 30883 60707
rect 31217 60673 31251 60707
rect 35725 60673 35759 60707
rect 36093 60673 36127 60707
rect 18797 60605 18831 60639
rect 19717 60605 19751 60639
rect 19993 60605 20027 60639
rect 20269 60605 20303 60639
rect 20637 60605 20671 60639
rect 22293 60605 22327 60639
rect 22431 60605 22465 60639
rect 22569 60605 22603 60639
rect 25145 60605 25179 60639
rect 25329 60605 25363 60639
rect 26157 60605 26191 60639
rect 26249 60605 26283 60639
rect 30941 60605 30975 60639
rect 35817 60605 35851 60639
rect 18705 60537 18739 60571
rect 21741 60537 21775 60571
rect 23397 60537 23431 60571
rect 19349 60469 19383 60503
rect 21649 60469 21683 60503
rect 23029 60469 23063 60503
rect 32321 60469 32355 60503
rect 37381 60469 37415 60503
rect 20361 60265 20395 60299
rect 24501 60265 24535 60299
rect 25329 60265 25363 60299
rect 29561 60265 29595 60299
rect 30941 60265 30975 60299
rect 23305 60197 23339 60231
rect 19257 60129 19291 60163
rect 19404 60129 19438 60163
rect 21281 60129 21315 60163
rect 21741 60129 21775 60163
rect 22845 60129 22879 60163
rect 27261 60129 27295 60163
rect 29745 60129 29779 60163
rect 19165 60061 19199 60095
rect 19625 60061 19659 60095
rect 20729 60061 20763 60095
rect 21097 60061 21131 60095
rect 21833 60061 21867 60095
rect 26617 60061 26651 60095
rect 18337 59993 18371 60027
rect 22661 59993 22695 60027
rect 23029 59993 23063 60027
rect 18613 59925 18647 59959
rect 19533 59925 19567 59959
rect 19901 59925 19935 59959
rect 22293 59925 22327 59959
rect 23857 59925 23891 59959
rect 24225 59925 24259 59959
rect 30205 59925 30239 59959
rect 35817 59925 35851 59959
rect 17877 59721 17911 59755
rect 22845 59721 22879 59755
rect 25513 59721 25547 59755
rect 18797 59653 18831 59687
rect 22293 59653 22327 59687
rect 27261 59653 27295 59687
rect 19625 59585 19659 59619
rect 20637 59585 20671 59619
rect 21373 59585 21407 59619
rect 21649 59585 21683 59619
rect 23949 59585 23983 59619
rect 25973 59585 26007 59619
rect 26617 59585 26651 59619
rect 30389 59585 30423 59619
rect 18613 59517 18647 59551
rect 20177 59517 20211 59551
rect 20453 59517 20487 59551
rect 21833 59517 21867 59551
rect 22385 59517 22419 59551
rect 24225 59517 24259 59551
rect 26341 59517 26375 59551
rect 26801 59517 26835 59551
rect 27261 59517 27295 59551
rect 27813 59517 27847 59551
rect 30021 59517 30055 59551
rect 30297 59517 30331 59551
rect 31125 59517 31159 59551
rect 31217 59517 31251 59551
rect 29745 59449 29779 59483
rect 18429 59381 18463 59415
rect 19349 59381 19383 59415
rect 20913 59381 20947 59415
rect 23305 59381 23339 59415
rect 28181 59381 28215 59415
rect 29101 59381 29135 59415
rect 1593 59177 1627 59211
rect 21557 59177 21591 59211
rect 22385 59177 22419 59211
rect 19257 59109 19291 59143
rect 20361 59109 20395 59143
rect 26525 59109 26559 59143
rect 29101 59109 29135 59143
rect 16681 59041 16715 59075
rect 17693 59041 17727 59075
rect 20913 59041 20947 59075
rect 23029 59041 23063 59075
rect 23305 59041 23339 59075
rect 24777 59041 24811 59075
rect 25237 59041 25271 59075
rect 27353 59041 27387 59075
rect 27537 59041 27571 59075
rect 29837 59041 29871 59075
rect 35173 59041 35207 59075
rect 35449 59041 35483 59075
rect 18061 58973 18095 59007
rect 19625 58973 19659 59007
rect 20729 58973 20763 59007
rect 21281 58973 21315 59007
rect 22661 58973 22695 59007
rect 24593 58973 24627 59007
rect 27077 58973 27111 59007
rect 29009 58973 29043 59007
rect 29929 58973 29963 59007
rect 19533 58905 19567 58939
rect 21189 58905 21223 58939
rect 23397 58905 23431 58939
rect 25237 58905 25271 58939
rect 26341 58905 26375 58939
rect 16865 58837 16899 58871
rect 17233 58837 17267 58871
rect 17601 58837 17635 58871
rect 17831 58837 17865 58871
rect 17969 58837 18003 58871
rect 18337 58837 18371 58871
rect 18981 58837 19015 58871
rect 19395 58837 19429 58871
rect 19901 58837 19935 58871
rect 21051 58837 21085 58871
rect 21925 58837 21959 58871
rect 24041 58837 24075 58871
rect 36553 58837 36587 58871
rect 16865 58633 16899 58667
rect 17141 58633 17175 58667
rect 19054 58633 19088 58667
rect 19349 58633 19383 58667
rect 22937 58633 22971 58667
rect 25145 58633 25179 58667
rect 35265 58633 35299 58667
rect 18797 58565 18831 58599
rect 19165 58565 19199 58599
rect 25881 58565 25915 58599
rect 26433 58565 26467 58599
rect 27721 58565 27755 58599
rect 1593 58497 1627 58531
rect 1869 58497 1903 58531
rect 19257 58497 19291 58531
rect 21189 58497 21223 58531
rect 23489 58497 23523 58531
rect 23949 58497 23983 58531
rect 24777 58497 24811 58531
rect 16957 58429 16991 58463
rect 17417 58429 17451 58463
rect 18429 58429 18463 58463
rect 21741 58429 21775 58463
rect 22017 58429 22051 58463
rect 22201 58429 22235 58463
rect 24225 58429 24259 58463
rect 24593 58429 24627 58463
rect 25697 58429 25731 58463
rect 26893 58429 26927 58463
rect 27445 58429 27479 58463
rect 27721 58429 27755 58463
rect 28273 58429 28307 58463
rect 28917 58429 28951 58463
rect 18889 58361 18923 58395
rect 20913 58361 20947 58395
rect 2973 58293 3007 58327
rect 16497 58293 16531 58327
rect 17877 58293 17911 58327
rect 19993 58293 20027 58327
rect 20545 58293 20579 58327
rect 22569 58293 22603 58327
rect 25513 58293 25547 58327
rect 26801 58293 26835 58327
rect 29561 58293 29595 58327
rect 35541 58293 35575 58327
rect 1685 58089 1719 58123
rect 15669 58089 15703 58123
rect 19717 58089 19751 58123
rect 25789 58089 25823 58123
rect 26341 58089 26375 58123
rect 29009 58089 29043 58123
rect 17509 58021 17543 58055
rect 20729 58021 20763 58055
rect 20913 58021 20947 58055
rect 15485 57953 15519 57987
rect 16489 57953 16523 57987
rect 17877 57953 17911 57987
rect 19073 57953 19107 57987
rect 23121 57953 23155 57987
rect 23535 57953 23569 57987
rect 24501 57953 24535 57987
rect 25329 57953 25363 57987
rect 28457 57953 28491 57987
rect 19441 57885 19475 57919
rect 20177 57885 20211 57919
rect 21281 57885 21315 57919
rect 22753 57885 22787 57919
rect 25053 57885 25087 57919
rect 25513 57885 25547 57919
rect 27629 57885 27663 57919
rect 28181 57885 28215 57919
rect 28641 57885 28675 57919
rect 18613 57817 18647 57851
rect 19211 57817 19245 57851
rect 23397 57817 23431 57851
rect 24317 57817 24351 57851
rect 16405 57749 16439 57783
rect 16681 57749 16715 57783
rect 17049 57749 17083 57783
rect 17417 57749 17451 57783
rect 18981 57749 19015 57783
rect 19349 57749 19383 57783
rect 21051 57749 21085 57783
rect 21189 57749 21223 57783
rect 21373 57749 21407 57783
rect 22017 57749 22051 57783
rect 22385 57749 22419 57783
rect 23949 57749 23983 57783
rect 26985 57749 27019 57783
rect 27445 57749 27479 57783
rect 14289 57545 14323 57579
rect 14749 57545 14783 57579
rect 17877 57545 17911 57579
rect 19303 57545 19337 57579
rect 19625 57545 19659 57579
rect 20269 57545 20303 57579
rect 21557 57545 21591 57579
rect 24133 57545 24167 57579
rect 25605 57545 25639 57579
rect 29009 57545 29043 57579
rect 18337 57477 18371 57511
rect 18705 57477 18739 57511
rect 19441 57477 19475 57511
rect 20913 57477 20947 57511
rect 25237 57477 25271 57511
rect 27261 57477 27295 57511
rect 15209 57409 15243 57443
rect 19533 57409 19567 57443
rect 21741 57409 21775 57443
rect 27353 57409 27387 57443
rect 29285 57409 29319 57443
rect 35173 57409 35207 57443
rect 15485 57341 15519 57375
rect 16865 57341 16899 57375
rect 18153 57341 18187 57375
rect 20729 57341 20763 57375
rect 22293 57341 22327 57375
rect 22431 57341 22465 57375
rect 22569 57341 22603 57375
rect 23121 57341 23155 57375
rect 24317 57341 24351 57375
rect 25881 57341 25915 57375
rect 27905 57341 27939 57375
rect 28181 57341 28215 57375
rect 28365 57341 28399 57375
rect 29377 57341 29411 57375
rect 35265 57341 35299 57375
rect 35541 57341 35575 57375
rect 15025 57273 15059 57307
rect 17509 57273 17543 57307
rect 19165 57273 19199 57307
rect 25789 57273 25823 57307
rect 26893 57273 26927 57307
rect 18981 57205 19015 57239
rect 20545 57205 20579 57239
rect 21189 57205 21223 57239
rect 23397 57205 23431 57239
rect 24501 57205 24535 57239
rect 28641 57205 28675 57239
rect 36645 57205 36679 57239
rect 18245 57001 18279 57035
rect 18613 57001 18647 57035
rect 18981 57001 19015 57035
rect 20177 57001 20211 57035
rect 20729 57001 20763 57035
rect 22661 57001 22695 57035
rect 22845 57001 22879 57035
rect 26709 57001 26743 57035
rect 21097 56933 21131 56967
rect 21465 56933 21499 56967
rect 14197 56865 14231 56899
rect 15669 56865 15703 56899
rect 17049 56865 17083 56899
rect 18061 56865 18095 56899
rect 19073 56865 19107 56899
rect 22017 56865 22051 56899
rect 22293 56865 22327 56899
rect 22661 56865 22695 56899
rect 23121 56865 23155 56899
rect 23305 56865 23339 56899
rect 23673 56865 23707 56899
rect 24225 56865 24259 56899
rect 25237 56865 25271 56899
rect 26525 56865 26559 56899
rect 28365 56865 28399 56899
rect 28825 56865 28859 56899
rect 15393 56797 15427 56831
rect 17877 56797 17911 56831
rect 19441 56797 19475 56831
rect 22477 56797 22511 56831
rect 24409 56797 24443 56831
rect 27813 56797 27847 56831
rect 28181 56797 28215 56831
rect 17601 56729 17635 56763
rect 19349 56729 19383 56763
rect 25421 56729 25455 56763
rect 27445 56729 27479 56763
rect 28917 56729 28951 56763
rect 13737 56661 13771 56695
rect 14013 56661 14047 56695
rect 14381 56661 14415 56695
rect 14749 56661 14783 56695
rect 15117 56661 15151 56695
rect 19211 56661 19245 56695
rect 19533 56661 19567 56695
rect 24685 56661 24719 56695
rect 25145 56661 25179 56695
rect 25697 56661 25731 56695
rect 26065 56661 26099 56695
rect 35265 56661 35299 56695
rect 13277 56457 13311 56491
rect 15761 56457 15795 56491
rect 16865 56457 16899 56491
rect 17877 56457 17911 56491
rect 18429 56457 18463 56491
rect 19809 56457 19843 56491
rect 21373 56457 21407 56491
rect 21557 56457 21591 56491
rect 23305 56457 23339 56491
rect 27169 56457 27203 56491
rect 27537 56457 27571 56491
rect 17141 56389 17175 56423
rect 18705 56389 18739 56423
rect 19073 56389 19107 56423
rect 19671 56389 19705 56423
rect 21262 56389 21296 56423
rect 24869 56389 24903 56423
rect 14197 56321 14231 56355
rect 14657 56321 14691 56355
rect 19901 56321 19935 56355
rect 20545 56321 20579 56355
rect 21465 56321 21499 56355
rect 25237 56321 25271 56355
rect 26065 56321 26099 56355
rect 28365 56321 28399 56355
rect 13369 56253 13403 56287
rect 14381 56253 14415 56287
rect 16957 56253 16991 56287
rect 18521 56253 18555 56287
rect 19533 56253 19567 56287
rect 22109 56253 22143 56287
rect 23673 56253 23707 56287
rect 24133 56253 24167 56287
rect 25145 56253 25179 56287
rect 25973 56253 26007 56287
rect 27813 56253 27847 56287
rect 13921 56185 13955 56219
rect 20913 56185 20947 56219
rect 21097 56185 21131 56219
rect 13553 56117 13587 56151
rect 16497 56117 16531 56151
rect 17509 56117 17543 56151
rect 19349 56117 19383 56151
rect 20177 56117 20211 56151
rect 22569 56117 22603 56151
rect 23029 56117 23063 56151
rect 23857 56117 23891 56151
rect 24501 56117 24535 56151
rect 26525 56117 26559 56151
rect 28641 56117 28675 56151
rect 14381 55913 14415 55947
rect 17509 55913 17543 55947
rect 18705 55913 18739 55947
rect 19073 55913 19107 55947
rect 20269 55913 20303 55947
rect 24317 55913 24351 55947
rect 26985 55913 27019 55947
rect 28549 55913 28583 55947
rect 13737 55845 13771 55879
rect 16129 55845 16163 55879
rect 19993 55845 20027 55879
rect 12173 55777 12207 55811
rect 13185 55777 13219 55811
rect 14197 55777 14231 55811
rect 16865 55777 16899 55811
rect 18337 55777 18371 55811
rect 19257 55777 19291 55811
rect 20913 55777 20947 55811
rect 21097 55777 21131 55811
rect 22937 55777 22971 55811
rect 23213 55777 23247 55811
rect 24225 55777 24259 55811
rect 24961 55777 24995 55811
rect 25237 55777 25271 55811
rect 26617 55777 26651 55811
rect 28273 55777 28307 55811
rect 33149 55777 33183 55811
rect 15485 55709 15519 55743
rect 16497 55709 16531 55743
rect 17233 55709 17267 55743
rect 18429 55709 18463 55743
rect 19625 55709 19659 55743
rect 21741 55709 21775 55743
rect 22385 55709 22419 55743
rect 23397 55709 23431 55743
rect 24133 55709 24167 55743
rect 32873 55709 32907 55743
rect 14105 55641 14139 55675
rect 16037 55641 16071 55675
rect 16405 55641 16439 55675
rect 12357 55573 12391 55607
rect 13369 55573 13403 55607
rect 14933 55573 14967 55607
rect 16294 55573 16328 55607
rect 19422 55573 19456 55607
rect 19533 55573 19567 55607
rect 20729 55573 20763 55607
rect 21189 55573 21223 55607
rect 22293 55573 22327 55607
rect 23673 55573 23707 55607
rect 25605 55573 25639 55607
rect 25973 55573 26007 55607
rect 27721 55573 27755 55607
rect 31861 55573 31895 55607
rect 34253 55573 34287 55607
rect 12265 55369 12299 55403
rect 12725 55369 12759 55403
rect 14013 55369 14047 55403
rect 14105 55369 14139 55403
rect 14381 55369 14415 55403
rect 15117 55369 15151 55403
rect 17785 55369 17819 55403
rect 19809 55369 19843 55403
rect 23029 55369 23063 55403
rect 25053 55369 25087 55403
rect 33241 55369 33275 55403
rect 13369 55301 13403 55335
rect 13737 55233 13771 55267
rect 12817 55165 12851 55199
rect 13829 55165 13863 55199
rect 15006 55301 15040 55335
rect 24501 55301 24535 55335
rect 26341 55301 26375 55335
rect 14749 55233 14783 55267
rect 15209 55233 15243 55267
rect 17141 55233 17175 55267
rect 20177 55233 20211 55267
rect 21649 55233 21683 55267
rect 22385 55233 22419 55267
rect 22661 55233 22695 55267
rect 25605 55233 25639 55267
rect 28457 55233 28491 55267
rect 31585 55233 31619 55267
rect 31861 55233 31895 55267
rect 32781 55233 32815 55267
rect 33609 55233 33643 55267
rect 16221 55165 16255 55199
rect 16757 55165 16791 55199
rect 18705 55165 18739 55199
rect 19625 55165 19659 55199
rect 21189 55165 21223 55199
rect 21741 55165 21775 55199
rect 23673 55165 23707 55199
rect 24041 55165 24075 55199
rect 24501 55165 24535 55199
rect 26433 55165 26467 55199
rect 26893 55165 26927 55199
rect 27997 55165 28031 55199
rect 28825 55165 28859 55199
rect 32689 55165 32723 55199
rect 14105 55097 14139 55131
rect 14841 55097 14875 55131
rect 15577 55097 15611 55131
rect 16405 55097 16439 55131
rect 18061 55097 18095 55131
rect 25973 55097 26007 55131
rect 31953 55097 31987 55131
rect 13001 55029 13035 55063
rect 15853 55029 15887 55063
rect 16589 55029 16623 55063
rect 16681 55029 16715 55063
rect 17509 55029 17543 55063
rect 19349 55029 19383 55063
rect 20453 55029 20487 55063
rect 21833 55029 21867 55063
rect 23489 55029 23523 55063
rect 26525 55029 26559 55063
rect 28181 55029 28215 55063
rect 13645 54825 13679 54859
rect 14933 54825 14967 54859
rect 16773 54825 16807 54859
rect 17049 54825 17083 54859
rect 17601 54825 17635 54859
rect 22017 54825 22051 54859
rect 23581 54825 23615 54859
rect 23949 54825 23983 54859
rect 27905 54825 27939 54859
rect 14105 54757 14139 54791
rect 15577 54757 15611 54791
rect 15761 54757 15795 54791
rect 13185 54689 13219 54723
rect 14197 54689 14231 54723
rect 19441 54757 19475 54791
rect 19993 54757 20027 54791
rect 26525 54757 26559 54791
rect 17417 54689 17451 54723
rect 19349 54689 19383 54723
rect 19533 54689 19567 54723
rect 21557 54689 21591 54723
rect 21741 54689 21775 54723
rect 22569 54689 22603 54723
rect 22753 54689 22787 54723
rect 25053 54689 25087 54723
rect 25421 54689 25455 54723
rect 26985 54689 27019 54723
rect 27353 54689 27387 54723
rect 28641 54689 28675 54723
rect 16129 54621 16163 54655
rect 17049 54621 17083 54655
rect 18613 54621 18647 54655
rect 19165 54621 19199 54655
rect 23121 54621 23155 54655
rect 25145 54621 25179 54655
rect 25513 54621 25547 54655
rect 27445 54621 27479 54655
rect 28917 54621 28951 54655
rect 14381 54553 14415 54587
rect 16037 54553 16071 54587
rect 17233 54553 17267 54587
rect 20637 54553 20671 54587
rect 24317 54553 24351 54587
rect 13369 54485 13403 54519
rect 15899 54485 15933 54519
rect 16405 54485 16439 54519
rect 20361 54485 20395 54519
rect 21097 54485 21131 54519
rect 24501 54485 24535 54519
rect 25881 54485 25915 54519
rect 26341 54485 26375 54519
rect 30021 54485 30055 54519
rect 31769 54485 31803 54519
rect 13185 54281 13219 54315
rect 14289 54281 14323 54315
rect 16865 54281 16899 54315
rect 17601 54281 17635 54315
rect 19993 54281 20027 54315
rect 23121 54281 23155 54315
rect 24317 54281 24351 54315
rect 27905 54281 27939 54315
rect 28733 54281 28767 54315
rect 29101 54281 29135 54315
rect 17141 54213 17175 54247
rect 19625 54213 19659 54247
rect 23489 54213 23523 54247
rect 14841 54145 14875 54179
rect 16497 54145 16531 54179
rect 20177 54145 20211 54179
rect 20913 54145 20947 54179
rect 22431 54145 22465 54179
rect 25237 54145 25271 54179
rect 25605 54145 25639 54179
rect 27261 54145 27295 54179
rect 13737 54077 13771 54111
rect 13829 54077 13863 54111
rect 15117 54077 15151 54111
rect 18613 54077 18647 54111
rect 18797 54077 18831 54111
rect 18889 54077 18923 54111
rect 19349 54077 19383 54111
rect 21557 54077 21591 54111
rect 22293 54077 22327 54111
rect 22569 54077 22603 54111
rect 24041 54077 24075 54111
rect 25145 54077 25179 54111
rect 25513 54077 25547 54111
rect 26525 54077 26559 54111
rect 26801 54077 26835 54111
rect 27537 54077 27571 54111
rect 28089 54077 28123 54111
rect 20545 54009 20579 54043
rect 21281 54009 21315 54043
rect 21741 54009 21775 54043
rect 24501 54009 24535 54043
rect 26893 54009 26927 54043
rect 14013 53941 14047 53975
rect 14749 53941 14783 53975
rect 18521 53941 18555 53975
rect 20361 53941 20395 53975
rect 20453 53941 20487 53975
rect 25973 53941 26007 53975
rect 26341 53941 26375 53975
rect 26709 53941 26743 53975
rect 28273 53941 28307 53975
rect 14105 53737 14139 53771
rect 15853 53737 15887 53771
rect 17049 53737 17083 53771
rect 19441 53737 19475 53771
rect 19533 53737 19567 53771
rect 20361 53737 20395 53771
rect 20637 53737 20671 53771
rect 21189 53737 21223 53771
rect 22753 53737 22787 53771
rect 15117 53669 15151 53703
rect 15761 53669 15795 53703
rect 15945 53669 15979 53703
rect 16313 53669 16347 53703
rect 16589 53669 16623 53703
rect 19257 53669 19291 53703
rect 19625 53669 19659 53703
rect 21557 53669 21591 53703
rect 23489 53669 23523 53703
rect 14197 53601 14231 53635
rect 15577 53601 15611 53635
rect 17141 53601 17175 53635
rect 17509 53601 17543 53635
rect 17969 53601 18003 53635
rect 19993 53601 20027 53635
rect 21649 53601 21683 53635
rect 22477 53601 22511 53635
rect 23765 53601 23799 53635
rect 24133 53601 24167 53635
rect 24501 53601 24535 53635
rect 27353 53601 27387 53635
rect 27537 53601 27571 53635
rect 27721 53601 27755 53635
rect 28181 53601 28215 53635
rect 22569 53533 22603 53567
rect 14381 53465 14415 53499
rect 17969 53465 18003 53499
rect 19073 53465 19107 53499
rect 24409 53465 24443 53499
rect 25697 53465 25731 53499
rect 27169 53465 27203 53499
rect 14749 53397 14783 53431
rect 18613 53397 18647 53431
rect 23121 53397 23155 53431
rect 24961 53397 24995 53431
rect 25421 53397 25455 53431
rect 26249 53397 26283 53431
rect 26709 53397 26743 53431
rect 15117 53193 15151 53227
rect 16681 53193 16715 53227
rect 17785 53193 17819 53227
rect 19533 53193 19567 53227
rect 22661 53193 22695 53227
rect 23489 53193 23523 53227
rect 24777 53193 24811 53227
rect 29561 53193 29595 53227
rect 14289 53125 14323 53159
rect 14933 53125 14967 53159
rect 18981 53125 19015 53159
rect 19993 53125 20027 53159
rect 20913 53125 20947 53159
rect 22017 53125 22051 53159
rect 23765 53125 23799 53159
rect 14565 53057 14599 53091
rect 16773 53057 16807 53091
rect 17141 53057 17175 53091
rect 20637 53057 20671 53091
rect 24133 53057 24167 53091
rect 25973 53057 26007 53091
rect 13921 52989 13955 53023
rect 15301 52989 15335 53023
rect 15393 52989 15427 53023
rect 16405 52989 16439 53023
rect 16552 52989 16586 53023
rect 17509 52989 17543 53023
rect 18153 52989 18187 53023
rect 18521 52989 18555 53023
rect 18981 52989 19015 53023
rect 20085 52989 20119 53023
rect 21373 52989 21407 53023
rect 22109 52989 22143 53023
rect 22293 52989 22327 53023
rect 23673 52989 23707 53023
rect 23949 52989 23983 53023
rect 25237 52989 25271 53023
rect 26893 52989 26927 53023
rect 27077 52989 27111 53023
rect 27537 52989 27571 53023
rect 28457 52989 28491 53023
rect 25605 52921 25639 52955
rect 15577 52853 15611 52887
rect 15945 52853 15979 52887
rect 16313 52853 16347 52887
rect 20269 52853 20303 52887
rect 23029 52853 23063 52887
rect 25053 52853 25087 52887
rect 25421 52853 25455 52887
rect 25513 52853 25547 52887
rect 26525 52853 26559 52887
rect 27169 52853 27203 52887
rect 28089 52853 28123 52887
rect 14749 52649 14783 52683
rect 16865 52649 16899 52683
rect 18337 52649 18371 52683
rect 21097 52649 21131 52683
rect 21649 52649 21683 52683
rect 23765 52649 23799 52683
rect 24041 52649 24075 52683
rect 25697 52649 25731 52683
rect 28733 52649 28767 52683
rect 29101 52649 29135 52683
rect 15853 52581 15887 52615
rect 16221 52581 16255 52615
rect 17049 52581 17083 52615
rect 20361 52581 20395 52615
rect 24961 52581 24995 52615
rect 27445 52581 27479 52615
rect 10517 52513 10551 52547
rect 15669 52513 15703 52547
rect 15761 52513 15795 52547
rect 16589 52513 16623 52547
rect 17923 52513 17957 52547
rect 18889 52513 18923 52547
rect 19441 52513 19475 52547
rect 19809 52513 19843 52547
rect 20637 52513 20671 52547
rect 20913 52513 20947 52547
rect 22661 52513 22695 52547
rect 23121 52513 23155 52547
rect 24685 52513 24719 52547
rect 25973 52513 26007 52547
rect 28181 52513 28215 52547
rect 29469 52513 29503 52547
rect 10241 52445 10275 52479
rect 11897 52445 11931 52479
rect 15485 52445 15519 52479
rect 17601 52445 17635 52479
rect 17739 52445 17773 52479
rect 22477 52445 22511 52479
rect 27353 52445 27387 52479
rect 28273 52445 28307 52479
rect 29193 52445 29227 52479
rect 30757 52445 30791 52479
rect 15117 52377 15151 52411
rect 19717 52377 19751 52411
rect 23121 52377 23155 52411
rect 18705 52309 18739 52343
rect 22109 52309 22143 52343
rect 25237 52309 25271 52343
rect 26801 52309 26835 52343
rect 27077 52309 27111 52343
rect 10241 52105 10275 52139
rect 10701 52105 10735 52139
rect 15485 52105 15519 52139
rect 15853 52105 15887 52139
rect 19073 52105 19107 52139
rect 21005 52105 21039 52139
rect 23029 52105 23063 52139
rect 24133 52105 24167 52139
rect 25145 52105 25179 52139
rect 25513 52105 25547 52139
rect 27721 52105 27755 52139
rect 29745 52105 29779 52139
rect 14473 52037 14507 52071
rect 22293 52037 22327 52071
rect 23673 52037 23707 52071
rect 28365 52037 28399 52071
rect 16129 51969 16163 52003
rect 16681 51969 16715 52003
rect 18061 51969 18095 52003
rect 18797 51969 18831 52003
rect 27353 51969 27387 52003
rect 30205 51969 30239 52003
rect 30573 51969 30607 52003
rect 14841 51901 14875 51935
rect 16957 51901 16991 51935
rect 17141 51901 17175 51935
rect 18245 51901 18279 51935
rect 19533 51901 19567 51935
rect 19901 51901 19935 51935
rect 20269 51901 20303 51935
rect 20453 51901 20487 51935
rect 21557 51901 21591 51935
rect 22385 51901 22419 51935
rect 22569 51901 22603 51935
rect 23489 51901 23523 51935
rect 23949 51901 23983 51935
rect 25237 51901 25271 51935
rect 25329 51901 25363 51935
rect 26801 51901 26835 51935
rect 26893 51901 26927 51935
rect 28181 51901 28215 51935
rect 28641 51901 28675 51935
rect 29101 51901 29135 51935
rect 29285 51901 29319 51935
rect 30297 51901 30331 51935
rect 17877 51833 17911 51867
rect 18429 51833 18463 51867
rect 23857 51833 23891 51867
rect 26065 51833 26099 51867
rect 26617 51833 26651 51867
rect 26985 51833 27019 51867
rect 15209 51765 15243 51799
rect 17509 51765 17543 51799
rect 18337 51765 18371 51799
rect 19717 51765 19751 51799
rect 21465 51765 21499 51799
rect 24685 51765 24719 51799
rect 26433 51765 26467 51799
rect 28089 51765 28123 51799
rect 29469 51765 29503 51799
rect 31861 51765 31895 51799
rect 15117 51561 15151 51595
rect 15485 51561 15519 51595
rect 18521 51561 18555 51595
rect 18797 51561 18831 51595
rect 20269 51561 20303 51595
rect 21373 51561 21407 51595
rect 21833 51561 21867 51595
rect 23305 51561 23339 51595
rect 25881 51561 25915 51595
rect 27905 51561 27939 51595
rect 30665 51561 30699 51595
rect 15853 51493 15887 51527
rect 16589 51493 16623 51527
rect 16957 51493 16991 51527
rect 24593 51493 24627 51527
rect 26249 51493 26283 51527
rect 27261 51493 27295 51527
rect 16037 51425 16071 51459
rect 17417 51425 17451 51459
rect 17877 51425 17911 51459
rect 19809 51425 19843 51459
rect 20913 51425 20947 51459
rect 21925 51425 21959 51459
rect 22293 51425 22327 51459
rect 22753 51425 22787 51459
rect 23949 51425 23983 51459
rect 24041 51425 24075 51459
rect 24133 51425 24167 51459
rect 24961 51425 24995 51459
rect 25237 51425 25271 51459
rect 25421 51425 25455 51459
rect 26801 51425 26835 51459
rect 26985 51425 27019 51459
rect 29193 51425 29227 51459
rect 29285 51425 29319 51459
rect 30205 51425 30239 51459
rect 31401 51425 31435 51459
rect 33885 51425 33919 51459
rect 17233 51357 17267 51391
rect 18981 51357 19015 51391
rect 19533 51357 19567 51391
rect 19993 51357 20027 51391
rect 20729 51357 20763 51391
rect 23029 51357 23063 51391
rect 28365 51357 28399 51391
rect 28457 51357 28491 51391
rect 17969 51289 18003 51323
rect 21097 51289 21131 51323
rect 29745 51289 29779 51323
rect 14749 51221 14783 51255
rect 16221 51221 16255 51255
rect 23673 51221 23707 51255
rect 25605 51221 25639 51255
rect 27537 51221 27571 51255
rect 30113 51221 30147 51255
rect 30389 51221 30423 51255
rect 31217 51221 31251 51255
rect 33701 51221 33735 51255
rect 15301 51017 15335 51051
rect 16037 51017 16071 51051
rect 19809 51017 19843 51051
rect 20361 51017 20395 51051
rect 22017 51017 22051 51051
rect 22293 51017 22327 51051
rect 22661 51017 22695 51051
rect 24869 51017 24903 51051
rect 28457 51017 28491 51051
rect 30389 51017 30423 51051
rect 31769 51017 31803 51051
rect 15669 50949 15703 50983
rect 18889 50949 18923 50983
rect 24133 50949 24167 50983
rect 17141 50881 17175 50915
rect 25237 50881 25271 50915
rect 26617 50881 26651 50915
rect 29285 50881 29319 50915
rect 14657 50813 14691 50847
rect 15117 50813 15151 50847
rect 16681 50813 16715 50847
rect 16957 50813 16991 50847
rect 18061 50813 18095 50847
rect 18613 50813 18647 50847
rect 18981 50813 19015 50847
rect 20821 50813 20855 50847
rect 21005 50813 21039 50847
rect 21373 50813 21407 50847
rect 22477 50813 22511 50847
rect 22937 50813 22971 50847
rect 23397 50813 23431 50847
rect 23949 50813 23983 50847
rect 24961 50813 24995 50847
rect 27797 50813 27831 50847
rect 29377 50813 29411 50847
rect 30849 50813 30883 50847
rect 31309 50813 31343 50847
rect 33701 50813 33735 50847
rect 15025 50745 15059 50779
rect 16129 50745 16163 50779
rect 17509 50745 17543 50779
rect 17877 50745 17911 50779
rect 27261 50745 27295 50779
rect 27445 50745 27479 50779
rect 27721 50745 27755 50779
rect 28181 50745 28215 50779
rect 19533 50677 19567 50711
rect 20821 50677 20855 50711
rect 24409 50677 24443 50711
rect 26893 50677 26927 50711
rect 27629 50677 27663 50711
rect 29009 50677 29043 50711
rect 30757 50677 30791 50711
rect 31033 50677 31067 50711
rect 17693 50473 17727 50507
rect 18061 50473 18095 50507
rect 20637 50473 20671 50507
rect 23581 50473 23615 50507
rect 26801 50473 26835 50507
rect 27169 50473 27203 50507
rect 30941 50473 30975 50507
rect 21189 50405 21223 50439
rect 22845 50405 22879 50439
rect 26341 50405 26375 50439
rect 15577 50337 15611 50371
rect 18797 50337 18831 50371
rect 19257 50337 19291 50371
rect 19993 50337 20027 50371
rect 21741 50337 21775 50371
rect 22293 50337 22327 50371
rect 22661 50337 22695 50371
rect 24225 50337 24259 50371
rect 24501 50337 24535 50371
rect 24961 50337 24995 50371
rect 27537 50337 27571 50371
rect 28365 50337 28399 50371
rect 28457 50337 28491 50371
rect 31493 50337 31527 50371
rect 15301 50269 15335 50303
rect 17325 50269 17359 50303
rect 18521 50269 18555 50303
rect 19533 50269 19567 50303
rect 23673 50269 23707 50303
rect 24685 50269 24719 50303
rect 25789 50269 25823 50303
rect 27629 50269 27663 50303
rect 29561 50269 29595 50303
rect 29837 50269 29871 50303
rect 21649 50201 21683 50235
rect 15025 50133 15059 50167
rect 16681 50133 16715 50167
rect 23121 50133 23155 50167
rect 25513 50133 25547 50167
rect 28917 50133 28951 50167
rect 29285 50133 29319 50167
rect 17141 49929 17175 49963
rect 17417 49929 17451 49963
rect 17877 49929 17911 49963
rect 19441 49929 19475 49963
rect 21465 49929 21499 49963
rect 26433 49929 26467 49963
rect 28365 49929 28399 49963
rect 28917 49929 28951 49963
rect 32229 49929 32263 49963
rect 14473 49861 14507 49895
rect 18889 49861 18923 49895
rect 24869 49861 24903 49895
rect 26893 49861 26927 49895
rect 15393 49793 15427 49827
rect 15761 49793 15795 49827
rect 16221 49793 16255 49827
rect 23489 49793 23523 49827
rect 25237 49793 25271 49827
rect 25421 49793 25455 49827
rect 26157 49793 26191 49827
rect 27077 49793 27111 49827
rect 29469 49793 29503 49827
rect 30297 49793 30331 49827
rect 30665 49793 30699 49827
rect 31217 49793 31251 49827
rect 14749 49725 14783 49759
rect 15209 49725 15243 49759
rect 15945 49725 15979 49759
rect 16313 49725 16347 49759
rect 18245 49725 18279 49759
rect 18613 49725 18647 49759
rect 18889 49725 18923 49759
rect 19901 49725 19935 49759
rect 20085 49725 20119 49759
rect 20361 49725 20395 49759
rect 20821 49725 20855 49759
rect 21097 49725 21131 49759
rect 22201 49725 22235 49759
rect 22385 49725 22419 49759
rect 23121 49725 23155 49759
rect 23857 49725 23891 49759
rect 23949 49725 23983 49759
rect 24133 49725 24167 49759
rect 27537 49725 27571 49759
rect 27721 49725 27755 49759
rect 27905 49725 27939 49759
rect 28733 49725 28767 49759
rect 29101 49725 29135 49759
rect 29377 49725 29411 49759
rect 30205 49725 30239 49759
rect 31033 49725 31067 49759
rect 31309 49725 31343 49759
rect 21833 49657 21867 49691
rect 25789 49657 25823 49691
rect 22201 49589 22235 49623
rect 24317 49589 24351 49623
rect 25605 49589 25639 49623
rect 25697 49589 25731 49623
rect 17417 49385 17451 49419
rect 19349 49385 19383 49419
rect 19625 49385 19659 49419
rect 20269 49385 20303 49419
rect 20729 49385 20763 49419
rect 21281 49385 21315 49419
rect 23213 49385 23247 49419
rect 23581 49385 23615 49419
rect 25145 49385 25179 49419
rect 25513 49385 25547 49419
rect 27813 49385 27847 49419
rect 29653 49385 29687 49419
rect 30941 49385 30975 49419
rect 13277 49317 13311 49351
rect 21649 49317 21683 49351
rect 26525 49317 26559 49351
rect 27537 49317 27571 49351
rect 27997 49317 28031 49351
rect 13737 49249 13771 49283
rect 13921 49249 13955 49283
rect 14105 49249 14139 49283
rect 14749 49249 14783 49283
rect 15393 49249 15427 49283
rect 15669 49249 15703 49283
rect 18245 49249 18279 49283
rect 18797 49249 18831 49283
rect 19809 49249 19843 49283
rect 21741 49249 21775 49283
rect 22293 49249 22327 49283
rect 22661 49249 22695 49283
rect 23673 49249 23707 49283
rect 24041 49249 24075 49283
rect 24501 49249 24535 49283
rect 26709 49249 26743 49283
rect 28549 49249 28583 49283
rect 28825 49249 28859 49283
rect 29929 49249 29963 49283
rect 17785 49181 17819 49215
rect 18061 49181 18095 49215
rect 24777 49181 24811 49215
rect 27077 49181 27111 49215
rect 29009 49181 29043 49215
rect 29837 49181 29871 49215
rect 13185 49113 13219 49147
rect 18705 49113 18739 49147
rect 22569 49113 22603 49147
rect 15025 49045 15059 49079
rect 16957 49045 16991 49079
rect 19993 49045 20027 49079
rect 25881 49045 25915 49079
rect 26249 49045 26283 49079
rect 31217 49045 31251 49079
rect 13185 48841 13219 48875
rect 15761 48841 15795 48875
rect 17417 48841 17451 48875
rect 17877 48841 17911 48875
rect 18245 48841 18279 48875
rect 18613 48841 18647 48875
rect 20545 48841 20579 48875
rect 21005 48841 21039 48875
rect 25789 48841 25823 48875
rect 28733 48841 28767 48875
rect 31033 48841 31067 48875
rect 31401 48841 31435 48875
rect 15393 48773 15427 48807
rect 23121 48773 23155 48807
rect 26617 48773 26651 48807
rect 12817 48705 12851 48739
rect 18981 48705 19015 48739
rect 19257 48705 19291 48739
rect 19901 48705 19935 48739
rect 23489 48705 23523 48739
rect 25513 48705 25547 48739
rect 27721 48705 27755 48739
rect 29469 48705 29503 48739
rect 30297 48705 30331 48739
rect 13277 48637 13311 48671
rect 13553 48637 13587 48671
rect 18061 48637 18095 48671
rect 19441 48637 19475 48671
rect 19993 48637 20027 48671
rect 21189 48637 21223 48671
rect 21649 48637 21683 48671
rect 22201 48637 22235 48671
rect 22569 48637 22603 48671
rect 22753 48637 22787 48671
rect 23765 48637 23799 48671
rect 24961 48637 24995 48671
rect 26801 48637 26835 48671
rect 26985 48637 27019 48671
rect 27169 48637 27203 48671
rect 28181 48637 28215 48671
rect 29653 48637 29687 48671
rect 30113 48637 30147 48671
rect 31217 48637 31251 48671
rect 31677 48637 31711 48671
rect 24777 48569 24811 48603
rect 25145 48569 25179 48603
rect 14657 48501 14691 48535
rect 17141 48501 17175 48535
rect 20913 48501 20947 48535
rect 21557 48501 21591 48535
rect 23949 48501 23983 48535
rect 24317 48501 24351 48535
rect 24685 48501 24719 48535
rect 25053 48501 25087 48535
rect 26249 48501 26283 48535
rect 27997 48501 28031 48535
rect 28365 48501 28399 48535
rect 29101 48501 29135 48535
rect 30665 48501 30699 48535
rect 13737 48297 13771 48331
rect 17969 48297 18003 48331
rect 22017 48297 22051 48331
rect 25605 48297 25639 48331
rect 28181 48297 28215 48331
rect 28641 48297 28675 48331
rect 29469 48297 29503 48331
rect 29837 48297 29871 48331
rect 11621 48229 11655 48263
rect 15117 48229 15151 48263
rect 18429 48229 18463 48263
rect 18797 48229 18831 48263
rect 20545 48229 20579 48263
rect 22385 48229 22419 48263
rect 23029 48229 23063 48263
rect 26525 48229 26559 48263
rect 30757 48229 30791 48263
rect 12265 48161 12299 48195
rect 12633 48161 12667 48195
rect 12817 48161 12851 48195
rect 13921 48161 13955 48195
rect 15761 48161 15795 48195
rect 15945 48161 15979 48195
rect 16129 48161 16163 48195
rect 19073 48161 19107 48195
rect 19441 48161 19475 48195
rect 19809 48161 19843 48195
rect 21189 48161 21223 48195
rect 21465 48161 21499 48195
rect 22569 48161 22603 48195
rect 23305 48161 23339 48195
rect 23857 48161 23891 48195
rect 24225 48161 24259 48195
rect 24593 48161 24627 48195
rect 25145 48161 25179 48195
rect 26985 48161 27019 48195
rect 27169 48161 27203 48195
rect 27353 48161 27387 48195
rect 27813 48161 27847 48195
rect 28549 48161 28583 48195
rect 28825 48161 28859 48195
rect 29561 48161 29595 48195
rect 29929 48161 29963 48195
rect 30021 48161 30055 48195
rect 12173 48093 12207 48127
rect 13829 48093 13863 48127
rect 19993 48093 20027 48127
rect 21373 48093 21407 48127
rect 22477 48093 22511 48127
rect 24685 48093 24719 48127
rect 31125 48093 31159 48127
rect 13369 48025 13403 48059
rect 15577 48025 15611 48059
rect 29561 48025 29595 48059
rect 11437 47957 11471 47991
rect 14105 47957 14139 47991
rect 14657 47957 14691 47991
rect 23765 47957 23799 47991
rect 26249 47957 26283 47991
rect 30205 47957 30239 47991
rect 31493 47957 31527 47991
rect 10977 47753 11011 47787
rect 11345 47753 11379 47787
rect 14289 47753 14323 47787
rect 16681 47753 16715 47787
rect 18613 47753 18647 47787
rect 18981 47753 19015 47787
rect 19349 47753 19383 47787
rect 19625 47753 19659 47787
rect 21465 47753 21499 47787
rect 23489 47753 23523 47787
rect 26985 47753 27019 47787
rect 29101 47753 29135 47787
rect 31125 47753 31159 47787
rect 11713 47685 11747 47719
rect 12173 47685 12207 47719
rect 23121 47685 23155 47719
rect 27537 47685 27571 47719
rect 32413 47685 32447 47719
rect 12541 47617 12575 47651
rect 14381 47617 14415 47651
rect 21189 47617 21223 47651
rect 22753 47617 22787 47651
rect 25421 47617 25455 47651
rect 25513 47617 25547 47651
rect 13001 47549 13035 47583
rect 13369 47549 13403 47583
rect 13461 47549 13495 47583
rect 14657 47549 14691 47583
rect 16313 47549 16347 47583
rect 16865 47549 16899 47583
rect 17325 47549 17359 47583
rect 19441 47549 19475 47583
rect 20361 47549 20395 47583
rect 21097 47549 21131 47583
rect 21925 47549 21959 47583
rect 22661 47549 22695 47583
rect 24225 47549 24259 47583
rect 24501 47549 24535 47583
rect 24685 47549 24719 47583
rect 25697 47549 25731 47583
rect 27721 47549 27755 47583
rect 27905 47549 27939 47583
rect 28089 47549 28123 47583
rect 29285 47549 29319 47583
rect 29745 47549 29779 47583
rect 30849 47549 30883 47583
rect 30941 47549 30975 47583
rect 31677 47549 31711 47583
rect 32229 47549 32263 47583
rect 32689 47549 32723 47583
rect 23673 47481 23707 47515
rect 24961 47481 24995 47515
rect 25881 47481 25915 47515
rect 26249 47481 26283 47515
rect 30389 47481 30423 47515
rect 13921 47413 13955 47447
rect 15761 47413 15795 47447
rect 17049 47413 17083 47447
rect 19993 47413 20027 47447
rect 25789 47413 25823 47447
rect 26617 47413 26651 47447
rect 28549 47413 28583 47447
rect 29377 47413 29411 47447
rect 30665 47413 30699 47447
rect 12725 47209 12759 47243
rect 13645 47209 13679 47243
rect 19993 47209 20027 47243
rect 21189 47209 21223 47243
rect 21465 47209 21499 47243
rect 22477 47209 22511 47243
rect 23121 47209 23155 47243
rect 24593 47209 24627 47243
rect 25421 47209 25455 47243
rect 25789 47209 25823 47243
rect 26249 47209 26283 47243
rect 28457 47209 28491 47243
rect 29837 47209 29871 47243
rect 30205 47209 30239 47243
rect 30665 47209 30699 47243
rect 31401 47209 31435 47243
rect 31769 47209 31803 47243
rect 13369 47141 13403 47175
rect 14381 47141 14415 47175
rect 15853 47141 15887 47175
rect 16129 47141 16163 47175
rect 23581 47141 23615 47175
rect 24317 47141 24351 47175
rect 25053 47141 25087 47175
rect 26525 47141 26559 47175
rect 30757 47141 30791 47175
rect 11621 47073 11655 47107
rect 13921 47073 13955 47107
rect 15393 47073 15427 47107
rect 16681 47073 16715 47107
rect 19809 47073 19843 47107
rect 21005 47073 21039 47107
rect 22017 47073 22051 47107
rect 22293 47073 22327 47107
rect 23489 47073 23523 47107
rect 25237 47073 25271 47107
rect 27169 47073 27203 47107
rect 27537 47073 27571 47107
rect 29009 47073 29043 47107
rect 29377 47073 29411 47107
rect 29469 47073 29503 47107
rect 30573 47073 30607 47107
rect 32137 47073 32171 47107
rect 11345 47005 11379 47039
rect 13829 47005 13863 47039
rect 15301 47005 15335 47039
rect 16957 47005 16991 47039
rect 18337 47005 18371 47039
rect 20729 47005 20763 47039
rect 23949 47005 23983 47039
rect 27077 47005 27111 47039
rect 27629 47005 27663 47039
rect 28089 47005 28123 47039
rect 30389 47005 30423 47039
rect 31125 47005 31159 47039
rect 20361 46937 20395 46971
rect 21925 46937 21959 46971
rect 22109 46937 22143 46971
rect 28825 46937 28859 46971
rect 1593 46869 1627 46903
rect 14933 46869 14967 46903
rect 23746 46869 23780 46903
rect 23857 46869 23891 46903
rect 32321 46869 32355 46903
rect 11713 46665 11747 46699
rect 13829 46665 13863 46699
rect 19901 46665 19935 46699
rect 21189 46665 21223 46699
rect 21557 46665 21591 46699
rect 25237 46665 25271 46699
rect 27445 46665 27479 46699
rect 29101 46665 29135 46699
rect 29653 46665 29687 46699
rect 32137 46665 32171 46699
rect 21925 46597 21959 46631
rect 32505 46597 32539 46631
rect 1685 46529 1719 46563
rect 12725 46529 12759 46563
rect 14933 46529 14967 46563
rect 20913 46529 20947 46563
rect 22477 46529 22511 46563
rect 24685 46529 24719 46563
rect 26157 46529 26191 46563
rect 26709 46529 26743 46563
rect 30113 46529 30147 46563
rect 32873 46529 32907 46563
rect 1409 46461 1443 46495
rect 12449 46461 12483 46495
rect 15393 46461 15427 46495
rect 15577 46461 15611 46495
rect 15761 46461 15795 46495
rect 20545 46461 20579 46495
rect 21005 46461 21039 46495
rect 22017 46461 22051 46495
rect 22109 46461 22143 46495
rect 22293 46461 22327 46495
rect 23121 46461 23155 46495
rect 23489 46461 23523 46495
rect 24593 46461 24627 46495
rect 26065 46461 26099 46495
rect 26985 46461 27019 46495
rect 27169 46461 27203 46495
rect 28089 46461 28123 46495
rect 28181 46461 28215 46495
rect 29837 46461 29871 46495
rect 3065 46393 3099 46427
rect 16221 46393 16255 46427
rect 16773 46393 16807 46427
rect 11437 46325 11471 46359
rect 12265 46325 12299 46359
rect 14381 46325 14415 46359
rect 14749 46325 14783 46359
rect 17141 46325 17175 46359
rect 25697 46325 25731 46359
rect 28365 46325 28399 46359
rect 28733 46325 28767 46359
rect 31217 46325 31251 46359
rect 31769 46325 31803 46359
rect 1685 46121 1719 46155
rect 8861 46121 8895 46155
rect 12541 46121 12575 46155
rect 13369 46121 13403 46155
rect 13737 46121 13771 46155
rect 15577 46121 15611 46155
rect 21373 46121 21407 46155
rect 23673 46121 23707 46155
rect 25789 46121 25823 46155
rect 27169 46121 27203 46155
rect 28365 46121 28399 46155
rect 28641 46121 28675 46155
rect 29101 46121 29135 46155
rect 30389 46121 30423 46155
rect 31217 46121 31251 46155
rect 14381 46053 14415 46087
rect 26801 46053 26835 46087
rect 12817 45985 12851 46019
rect 13921 45985 13955 46019
rect 21465 45985 21499 46019
rect 22109 45985 22143 46019
rect 22477 45985 22511 46019
rect 22753 45985 22787 46019
rect 24869 45985 24903 46019
rect 27537 45985 27571 46019
rect 28089 45985 28123 46019
rect 28273 45985 28307 46019
rect 29285 45985 29319 46019
rect 29929 45985 29963 46019
rect 30757 45985 30791 46019
rect 32137 45985 32171 46019
rect 32229 45985 32263 46019
rect 13829 45917 13863 45951
rect 22937 45917 22971 45951
rect 24041 45917 24075 45951
rect 24593 45917 24627 45951
rect 25053 45917 25087 45951
rect 21649 45849 21683 45883
rect 22569 45849 22603 45883
rect 13001 45781 13035 45815
rect 14933 45781 14967 45815
rect 25421 45781 25455 45815
rect 26249 45781 26283 45815
rect 30941 45781 30975 45815
rect 31585 45781 31619 45815
rect 32413 45781 32447 45815
rect 14749 45577 14783 45611
rect 22477 45577 22511 45611
rect 23121 45577 23155 45611
rect 27629 45577 27663 45611
rect 28733 45577 28767 45611
rect 30757 45577 30791 45611
rect 32137 45577 32171 45611
rect 32505 45577 32539 45611
rect 22753 45509 22787 45543
rect 24041 45509 24075 45543
rect 28089 45509 28123 45543
rect 29101 45509 29135 45543
rect 9873 45441 9907 45475
rect 13369 45441 13403 45475
rect 25237 45441 25271 45475
rect 26065 45441 26099 45475
rect 30021 45441 30055 45475
rect 8769 45373 8803 45407
rect 8953 45373 8987 45407
rect 9781 45373 9815 45407
rect 13645 45373 13679 45407
rect 22569 45373 22603 45407
rect 24777 45373 24811 45407
rect 25145 45373 25179 45407
rect 26157 45373 26191 45407
rect 26801 45373 26835 45407
rect 26893 45373 26927 45407
rect 27169 45373 27203 45407
rect 27353 45373 27387 45407
rect 28181 45373 28215 45407
rect 29561 45373 29595 45407
rect 31125 45373 31159 45407
rect 9045 45305 9079 45339
rect 24317 45305 24351 45339
rect 25697 45305 25731 45339
rect 29285 45305 29319 45339
rect 29653 45305 29687 45339
rect 30849 45305 30883 45339
rect 31033 45305 31067 45339
rect 31217 45305 31251 45339
rect 31585 45305 31619 45339
rect 12817 45237 12851 45271
rect 13277 45237 13311 45271
rect 21465 45237 21499 45271
rect 22017 45237 22051 45271
rect 23489 45237 23523 45271
rect 28365 45237 28399 45271
rect 29469 45237 29503 45271
rect 30297 45237 30331 45271
rect 8861 45033 8895 45067
rect 13553 45033 13587 45067
rect 14381 45033 14415 45067
rect 22477 45033 22511 45067
rect 22753 45033 22787 45067
rect 23121 45033 23155 45067
rect 23765 45033 23799 45067
rect 24685 45033 24719 45067
rect 26709 45033 26743 45067
rect 27445 45033 27479 45067
rect 29377 45033 29411 45067
rect 30941 45033 30975 45067
rect 31493 45033 31527 45067
rect 24317 44965 24351 44999
rect 1777 44897 1811 44931
rect 13737 44897 13771 44931
rect 13829 44897 13863 44931
rect 22293 44897 22327 44931
rect 23857 44897 23891 44931
rect 24869 44897 24903 44931
rect 25053 44897 25087 44931
rect 25145 44897 25179 44931
rect 26525 44897 26559 44931
rect 28181 44897 28215 44931
rect 28549 44897 28583 44931
rect 28733 44897 28767 44931
rect 29561 44897 29595 44931
rect 1501 44829 1535 44863
rect 28273 44829 28307 44863
rect 29837 44829 29871 44863
rect 12541 44761 12575 44795
rect 13461 44761 13495 44795
rect 26341 44761 26375 44795
rect 3065 44693 3099 44727
rect 12909 44693 12943 44727
rect 14013 44693 14047 44727
rect 22201 44693 22235 44727
rect 25329 44693 25363 44727
rect 25973 44693 26007 44727
rect 27077 44693 27111 44727
rect 27629 44693 27663 44727
rect 31861 44693 31895 44727
rect 1685 44489 1719 44523
rect 8125 44489 8159 44523
rect 14289 44489 14323 44523
rect 15485 44489 15519 44523
rect 15945 44489 15979 44523
rect 24869 44489 24903 44523
rect 26801 44489 26835 44523
rect 27261 44489 27295 44523
rect 28733 44489 28767 44523
rect 31125 44489 31159 44523
rect 37657 44489 37691 44523
rect 14013 44421 14047 44455
rect 25329 44421 25363 44455
rect 8585 44353 8619 44387
rect 12541 44353 12575 44387
rect 12909 44353 12943 44387
rect 24593 44353 24627 44387
rect 25513 44353 25547 44387
rect 28273 44353 28307 44387
rect 30849 44353 30883 44387
rect 31677 44353 31711 44387
rect 36001 44353 36035 44387
rect 2053 44285 2087 44319
rect 8309 44285 8343 44319
rect 13093 44285 13127 44319
rect 13461 44285 13495 44319
rect 13553 44285 13587 44319
rect 15669 44285 15703 44319
rect 23397 44285 23431 44319
rect 23949 44285 23983 44319
rect 24041 44285 24075 44319
rect 24225 44285 24259 44319
rect 25605 44285 25639 44319
rect 26341 44285 26375 44319
rect 26433 44285 26467 44319
rect 27813 44285 27847 44319
rect 28181 44285 28215 44319
rect 29101 44285 29135 44319
rect 29285 44285 29319 44319
rect 29745 44285 29779 44319
rect 30757 44285 30791 44319
rect 30941 44285 30975 44319
rect 36093 44285 36127 44319
rect 36369 44285 36403 44319
rect 9965 44217 9999 44251
rect 11897 44217 11931 44251
rect 27353 44217 27387 44251
rect 30389 44217 30423 44251
rect 12173 44149 12207 44183
rect 22385 44149 22419 44183
rect 29377 44149 29411 44183
rect 8309 43945 8343 43979
rect 12541 43945 12575 43979
rect 13185 43945 13219 43979
rect 17785 43945 17819 43979
rect 23857 43945 23891 43979
rect 24777 43945 24811 43979
rect 25973 43945 26007 43979
rect 26341 43945 26375 43979
rect 26617 43945 26651 43979
rect 27997 43945 28031 43979
rect 29653 43945 29687 43979
rect 36093 43945 36127 43979
rect 30021 43877 30055 43911
rect 10977 43809 11011 43843
rect 15393 43809 15427 43843
rect 17969 43809 18003 43843
rect 20913 43809 20947 43843
rect 23673 43809 23707 43843
rect 24225 43809 24259 43843
rect 24869 43809 24903 43843
rect 25237 43809 25271 43843
rect 26525 43809 26559 43843
rect 27077 43809 27111 43843
rect 28365 43809 28399 43843
rect 29193 43809 29227 43843
rect 30205 43809 30239 43843
rect 11253 43741 11287 43775
rect 15301 43741 15335 43775
rect 21189 43741 21223 43775
rect 28457 43741 28491 43775
rect 29285 43741 29319 43775
rect 30665 43741 30699 43775
rect 23581 43673 23615 43707
rect 27629 43673 27663 43707
rect 15577 43605 15611 43639
rect 22293 43605 22327 43639
rect 30389 43605 30423 43639
rect 11069 43401 11103 43435
rect 11345 43401 11379 43435
rect 15301 43401 15335 43435
rect 17785 43401 17819 43435
rect 21005 43401 21039 43435
rect 27905 43401 27939 43435
rect 28273 43401 28307 43435
rect 28641 43401 28675 43435
rect 30665 43401 30699 43435
rect 21281 43333 21315 43367
rect 24409 43333 24443 43367
rect 29009 43333 29043 43367
rect 13093 43265 13127 43299
rect 14749 43265 14783 43299
rect 15669 43265 15703 43299
rect 24593 43265 24627 43299
rect 25513 43265 25547 43299
rect 25973 43265 26007 43299
rect 27445 43265 27479 43299
rect 29377 43265 29411 43299
rect 30297 43265 30331 43299
rect 13369 43197 13403 43231
rect 25421 43197 25455 43231
rect 26525 43197 26559 43231
rect 27353 43197 27387 43231
rect 30205 43197 30239 43231
rect 24685 43129 24719 43163
rect 26617 43129 26651 43163
rect 29469 43129 29503 43163
rect 12909 43061 12943 43095
rect 23857 43061 23891 43095
rect 26341 43061 26375 43095
rect 14105 42857 14139 42891
rect 24501 42857 24535 42891
rect 24961 42857 24995 42891
rect 26341 42857 26375 42891
rect 28365 42857 28399 42891
rect 29929 42857 29963 42891
rect 12909 42721 12943 42755
rect 13093 42721 13127 42755
rect 13277 42721 13311 42755
rect 20913 42721 20947 42755
rect 21189 42721 21223 42755
rect 24133 42721 24167 42755
rect 26801 42721 26835 42755
rect 27261 42721 27295 42755
rect 27629 42721 27663 42755
rect 28641 42721 28675 42755
rect 29469 42721 29503 42755
rect 33793 42721 33827 42755
rect 26709 42653 26743 42687
rect 27997 42653 28031 42687
rect 28733 42653 28767 42687
rect 29561 42653 29595 42687
rect 34069 42653 34103 42687
rect 35173 42653 35207 42687
rect 12725 42585 12759 42619
rect 19625 42517 19659 42551
rect 22293 42517 22327 42551
rect 25237 42517 25271 42551
rect 25697 42517 25731 42551
rect 12633 42313 12667 42347
rect 21005 42313 21039 42347
rect 25513 42313 25547 42347
rect 26985 42313 27019 42347
rect 27445 42313 27479 42347
rect 28089 42313 28123 42347
rect 29009 42313 29043 42347
rect 29469 42313 29503 42347
rect 34161 42313 34195 42347
rect 13277 42245 13311 42279
rect 14381 42245 14415 42279
rect 21281 42245 21315 42279
rect 27721 42245 27755 42279
rect 28641 42245 28675 42279
rect 13001 42177 13035 42211
rect 25789 42177 25823 42211
rect 26617 42177 26651 42211
rect 12449 42109 12483 42143
rect 14565 42109 14599 42143
rect 14749 42109 14783 42143
rect 14933 42109 14967 42143
rect 19533 42109 19567 42143
rect 19717 42109 19751 42143
rect 19809 42109 19843 42143
rect 24041 42109 24075 42143
rect 24501 42109 24535 42143
rect 25697 42109 25731 42143
rect 26525 42109 26559 42143
rect 27537 42109 27571 42143
rect 20269 42041 20303 42075
rect 23949 42041 23983 42075
rect 12265 41973 12299 42007
rect 14013 41973 14047 42007
rect 19073 41973 19107 42007
rect 19349 41973 19383 42007
rect 24317 41973 24351 42007
rect 33885 41973 33919 42007
rect 12541 41769 12575 41803
rect 14197 41769 14231 41803
rect 21097 41769 21131 41803
rect 25605 41769 25639 41803
rect 26801 41769 26835 41803
rect 5733 41701 5767 41735
rect 13645 41701 13679 41735
rect 4353 41633 4387 41667
rect 13185 41633 13219 41667
rect 19901 41633 19935 41667
rect 23489 41633 23523 41667
rect 4077 41565 4111 41599
rect 10333 41565 10367 41599
rect 10609 41565 10643 41599
rect 13093 41565 13127 41599
rect 19165 41565 19199 41599
rect 23765 41565 23799 41599
rect 27261 41565 27295 41599
rect 27537 41565 27571 41599
rect 28917 41565 28951 41599
rect 29285 41565 29319 41599
rect 11713 41429 11747 41463
rect 19533 41429 19567 41463
rect 24869 41429 24903 41463
rect 10425 41225 10459 41259
rect 23857 41225 23891 41259
rect 27353 41225 27387 41259
rect 27721 41225 27755 41259
rect 29101 41225 29135 41259
rect 19257 41157 19291 41191
rect 24225 41157 24259 41191
rect 18613 41089 18647 41123
rect 19625 41089 19659 41123
rect 21005 41089 21039 41123
rect 29377 41089 29411 41123
rect 30297 41089 30331 41123
rect 18061 41021 18095 41055
rect 19165 41021 19199 41055
rect 19441 41021 19475 41055
rect 20269 41021 20303 41055
rect 20545 41021 20579 41055
rect 21097 41021 21131 41055
rect 21373 41021 21407 41055
rect 30205 41021 30239 41055
rect 4445 40953 4479 40987
rect 13185 40953 13219 40987
rect 29469 40953 29503 40987
rect 4077 40885 4111 40919
rect 10793 40885 10827 40919
rect 13461 40885 13495 40919
rect 18245 40885 18279 40919
rect 18981 40885 19015 40919
rect 22477 40885 22511 40919
rect 21097 40681 21131 40715
rect 21741 40681 21775 40715
rect 23489 40681 23523 40715
rect 2421 40613 2455 40647
rect 2973 40613 3007 40647
rect 13001 40613 13035 40647
rect 2605 40545 2639 40579
rect 13829 40545 13863 40579
rect 15945 40545 15979 40579
rect 17693 40545 17727 40579
rect 18981 40545 19015 40579
rect 19349 40545 19383 40579
rect 19717 40545 19751 40579
rect 19993 40545 20027 40579
rect 20085 40545 20119 40579
rect 20269 40545 20303 40579
rect 20729 40545 20763 40579
rect 20913 40545 20947 40579
rect 22109 40545 22143 40579
rect 22385 40545 22419 40579
rect 35265 40545 35299 40579
rect 11345 40477 11379 40511
rect 11621 40477 11655 40511
rect 17785 40477 17819 40511
rect 34989 40477 35023 40511
rect 1685 40341 1719 40375
rect 14013 40341 14047 40375
rect 16129 40341 16163 40375
rect 18797 40341 18831 40375
rect 21373 40341 21407 40375
rect 25697 40341 25731 40375
rect 29285 40341 29319 40375
rect 36369 40341 36403 40375
rect 17141 40137 17175 40171
rect 23121 40137 23155 40171
rect 35449 40137 35483 40171
rect 11713 40069 11747 40103
rect 35173 40069 35207 40103
rect 1593 40001 1627 40035
rect 18337 40001 18371 40035
rect 20821 40001 20855 40035
rect 21373 40001 21407 40035
rect 26157 40001 26191 40035
rect 1869 39933 1903 39967
rect 13093 39933 13127 39967
rect 13553 39933 13587 39967
rect 15577 39933 15611 39967
rect 15945 39933 15979 39967
rect 16497 39933 16531 39967
rect 17877 39933 17911 39967
rect 21097 39933 21131 39967
rect 23397 39933 23431 39967
rect 25145 39933 25179 39967
rect 26295 39933 26329 39967
rect 26433 39933 26467 39967
rect 3249 39865 3283 39899
rect 16037 39865 16071 39899
rect 18797 39865 18831 39899
rect 20545 39865 20579 39899
rect 25605 39865 25639 39899
rect 11437 39797 11471 39831
rect 13277 39797 13311 39831
rect 13921 39797 13955 39831
rect 15209 39797 15243 39831
rect 18613 39797 18647 39831
rect 22477 39797 22511 39831
rect 25513 39797 25547 39831
rect 2789 39593 2823 39627
rect 19073 39593 19107 39627
rect 21097 39593 21131 39627
rect 22753 39593 22787 39627
rect 25145 39593 25179 39627
rect 1593 39525 1627 39559
rect 18797 39525 18831 39559
rect 19993 39525 20027 39559
rect 20269 39525 20303 39559
rect 26525 39525 26559 39559
rect 15577 39457 15611 39491
rect 17877 39457 17911 39491
rect 18245 39457 18279 39491
rect 19901 39457 19935 39491
rect 21373 39457 21407 39491
rect 25053 39457 25087 39491
rect 26617 39457 26651 39491
rect 35357 39457 35391 39491
rect 14473 39389 14507 39423
rect 15485 39389 15519 39423
rect 16037 39389 16071 39423
rect 17233 39389 17267 39423
rect 17785 39389 17819 39423
rect 18337 39389 18371 39423
rect 21649 39389 21683 39423
rect 34713 39389 34747 39423
rect 13829 39321 13863 39355
rect 17141 39321 17175 39355
rect 2421 39253 2455 39287
rect 14197 39253 14231 39287
rect 15025 39253 15059 39287
rect 16313 39253 16347 39287
rect 16681 39253 16715 39287
rect 20729 39253 20763 39287
rect 9413 39049 9447 39083
rect 16313 39049 16347 39083
rect 16773 39049 16807 39083
rect 17785 39049 17819 39083
rect 19349 39049 19383 39083
rect 21005 39049 21039 39083
rect 22385 39049 22419 39083
rect 26341 39049 26375 39083
rect 29745 39049 29779 39083
rect 35173 39049 35207 39083
rect 20039 38981 20073 39015
rect 20177 38981 20211 39015
rect 26709 38981 26743 39015
rect 1685 38913 1719 38947
rect 9873 38913 9907 38947
rect 13277 38913 13311 38947
rect 18061 38913 18095 38947
rect 18613 38913 18647 38947
rect 19073 38913 19107 38947
rect 20269 38913 20303 38947
rect 24409 38913 24443 38947
rect 25053 38913 25087 38947
rect 25973 38913 26007 38947
rect 27353 38913 27387 38947
rect 27813 38913 27847 38947
rect 30205 38913 30239 38947
rect 1409 38845 1443 38879
rect 9137 38845 9171 38879
rect 9597 38845 9631 38879
rect 13737 38845 13771 38879
rect 14105 38845 14139 38879
rect 14289 38845 14323 38879
rect 14749 38845 14783 38879
rect 15117 38845 15151 38879
rect 15669 38845 15703 38879
rect 16497 38845 16531 38879
rect 16589 38845 16623 38879
rect 17325 38845 17359 38879
rect 18889 38845 18923 38879
rect 19809 38845 19843 38879
rect 20637 38845 20671 38879
rect 21465 38845 21499 38879
rect 21925 38845 21959 38879
rect 24777 38845 24811 38879
rect 25421 38845 25455 38879
rect 25789 38845 25823 38879
rect 27629 38845 27663 38879
rect 29929 38845 29963 38879
rect 13645 38777 13679 38811
rect 19901 38777 19935 38811
rect 21373 38777 21407 38811
rect 24041 38777 24075 38811
rect 26801 38777 26835 38811
rect 2789 38709 2823 38743
rect 11161 38709 11195 38743
rect 12909 38709 12943 38743
rect 16037 38709 16071 38743
rect 21649 38709 21683 38743
rect 31309 38709 31343 38743
rect 1685 38505 1719 38539
rect 1961 38505 1995 38539
rect 15945 38505 15979 38539
rect 19993 38505 20027 38539
rect 20729 38505 20763 38539
rect 21741 38505 21775 38539
rect 25697 38505 25731 38539
rect 26893 38505 26927 38539
rect 27169 38505 27203 38539
rect 29929 38505 29963 38539
rect 13277 38437 13311 38471
rect 18153 38437 18187 38471
rect 11805 38369 11839 38403
rect 11989 38369 12023 38403
rect 12357 38369 12391 38403
rect 12541 38369 12575 38403
rect 14197 38369 14231 38403
rect 14381 38369 14415 38403
rect 16037 38369 16071 38403
rect 16405 38369 16439 38403
rect 16865 38369 16899 38403
rect 19073 38369 19107 38403
rect 19441 38369 19475 38403
rect 21005 38369 21039 38403
rect 24409 38369 24443 38403
rect 25237 38369 25271 38403
rect 27997 38369 28031 38403
rect 11345 38301 11379 38335
rect 13369 38301 13403 38335
rect 13921 38301 13955 38335
rect 18705 38301 18739 38335
rect 20913 38301 20947 38335
rect 24501 38301 24535 38335
rect 25329 38301 25363 38335
rect 27721 38301 27755 38335
rect 16865 38233 16899 38267
rect 17509 38233 17543 38267
rect 19349 38233 19383 38267
rect 11161 38165 11195 38199
rect 12817 38165 12851 38199
rect 14749 38165 14783 38199
rect 15117 38165 15151 38199
rect 15485 38165 15519 38199
rect 20269 38165 20303 38199
rect 21189 38165 21223 38199
rect 24133 38165 24167 38199
rect 27629 38165 27663 38199
rect 29101 38165 29135 38199
rect 11069 37961 11103 37995
rect 13645 37961 13679 37995
rect 14105 37961 14139 37995
rect 15853 37961 15887 37995
rect 17417 37961 17451 37995
rect 17877 37961 17911 37995
rect 19809 37961 19843 37995
rect 23489 37961 23523 37995
rect 26249 37961 26283 37995
rect 28181 37961 28215 37995
rect 28641 37961 28675 37995
rect 11437 37893 11471 37927
rect 15485 37893 15519 37927
rect 24041 37893 24075 37927
rect 12541 37825 12575 37859
rect 14841 37825 14875 37859
rect 16497 37825 16531 37859
rect 21649 37825 21683 37859
rect 24777 37825 24811 37859
rect 25053 37825 25087 37859
rect 27813 37825 27847 37859
rect 12633 37757 12667 37791
rect 13185 37757 13219 37791
rect 13369 37757 13403 37791
rect 14933 37757 14967 37791
rect 16589 37757 16623 37791
rect 16957 37757 16991 37791
rect 17141 37757 17175 37791
rect 18245 37757 18279 37791
rect 18797 37757 18831 37791
rect 18889 37757 18923 37791
rect 19533 37757 19567 37791
rect 20453 37757 20487 37791
rect 20637 37757 20671 37791
rect 20821 37757 20855 37791
rect 24409 37757 24443 37791
rect 25421 37757 25455 37791
rect 25697 37757 25731 37791
rect 26617 37757 26651 37791
rect 26893 37757 26927 37791
rect 27721 37757 27755 37791
rect 10701 37689 10735 37723
rect 15945 37689 15979 37723
rect 19993 37689 20027 37723
rect 25973 37689 26007 37723
rect 26985 37689 27019 37723
rect 11897 37621 11931 37655
rect 12173 37621 12207 37655
rect 15117 37621 15151 37655
rect 18153 37621 18187 37655
rect 21281 37621 21315 37655
rect 12173 37417 12207 37451
rect 12541 37417 12575 37451
rect 13185 37417 13219 37451
rect 15485 37417 15519 37451
rect 18153 37417 18187 37451
rect 18429 37417 18463 37451
rect 20085 37417 20119 37451
rect 20453 37417 20487 37451
rect 25145 37417 25179 37451
rect 27169 37417 27203 37451
rect 33517 37417 33551 37451
rect 10609 37281 10643 37315
rect 10793 37281 10827 37315
rect 11069 37281 11103 37315
rect 16313 37349 16347 37383
rect 13737 37281 13771 37315
rect 14197 37281 14231 37315
rect 15301 37281 15335 37315
rect 16129 37281 16163 37315
rect 16957 37281 16991 37315
rect 17325 37281 17359 37315
rect 17877 37281 17911 37315
rect 18521 37281 18555 37315
rect 18981 37281 19015 37315
rect 19165 37281 19199 37315
rect 27445 37281 27479 37315
rect 32413 37281 32447 37315
rect 13461 37213 13495 37247
rect 16865 37213 16899 37247
rect 17417 37213 17451 37247
rect 23121 37213 23155 37247
rect 23397 37213 23431 37247
rect 32137 37213 32171 37247
rect 12541 37145 12575 37179
rect 14197 37145 14231 37179
rect 12817 37077 12851 37111
rect 14749 37077 14783 37111
rect 15117 37077 15151 37111
rect 24501 37077 24535 37111
rect 9965 36873 9999 36907
rect 16221 36873 16255 36907
rect 16681 36873 16715 36907
rect 17509 36873 17543 36907
rect 20177 36873 20211 36907
rect 20545 36873 20579 36907
rect 21649 36873 21683 36907
rect 23213 36873 23247 36907
rect 26801 36873 26835 36907
rect 27445 36873 27479 36907
rect 32505 36873 32539 36907
rect 14381 36805 14415 36839
rect 11529 36737 11563 36771
rect 12265 36737 12299 36771
rect 13553 36737 13587 36771
rect 14473 36737 14507 36771
rect 15853 36737 15887 36771
rect 25329 36737 25363 36771
rect 10885 36669 10919 36703
rect 11897 36669 11931 36703
rect 12633 36669 12667 36703
rect 13461 36669 13495 36703
rect 14933 36669 14967 36703
rect 15209 36669 15243 36703
rect 15301 36669 15335 36703
rect 15669 36669 15703 36703
rect 16957 36669 16991 36703
rect 18245 36669 18279 36703
rect 18797 36669 18831 36703
rect 19073 36669 19107 36703
rect 25421 36669 25455 36703
rect 25697 36669 25731 36703
rect 12725 36601 12759 36635
rect 14013 36601 14047 36635
rect 17877 36601 17911 36635
rect 10241 36533 10275 36567
rect 10609 36533 10643 36567
rect 17141 36533 17175 36567
rect 18153 36533 18187 36567
rect 19533 36533 19567 36567
rect 19901 36533 19935 36567
rect 20913 36533 20947 36567
rect 21281 36533 21315 36567
rect 23857 36533 23891 36567
rect 32137 36533 32171 36567
rect 10977 36329 11011 36363
rect 11621 36329 11655 36363
rect 13277 36329 13311 36363
rect 14841 36329 14875 36363
rect 17509 36329 17543 36363
rect 18613 36329 18647 36363
rect 18981 36329 19015 36363
rect 24501 36329 24535 36363
rect 29561 36329 29595 36363
rect 15301 36261 15335 36295
rect 18337 36261 18371 36295
rect 21741 36261 21775 36295
rect 11069 36193 11103 36227
rect 12265 36193 12299 36227
rect 12817 36193 12851 36227
rect 13001 36193 13035 36227
rect 15761 36193 15795 36227
rect 15945 36193 15979 36227
rect 16129 36193 16163 36227
rect 16681 36193 16715 36227
rect 17601 36193 17635 36227
rect 17785 36193 17819 36227
rect 17877 36193 17911 36227
rect 19165 36193 19199 36227
rect 19349 36193 19383 36227
rect 20913 36193 20947 36227
rect 23397 36193 23431 36227
rect 28181 36193 28215 36227
rect 12081 36125 12115 36159
rect 16405 36125 16439 36159
rect 19717 36125 19751 36159
rect 21373 36125 21407 36159
rect 22569 36125 22603 36159
rect 23121 36125 23155 36159
rect 25421 36125 25455 36159
rect 28457 36125 28491 36159
rect 20361 36057 20395 36091
rect 11253 35989 11287 36023
rect 11989 35989 12023 36023
rect 14013 35989 14047 36023
rect 14565 35989 14599 36023
rect 17049 35989 17083 36023
rect 19993 35989 20027 36023
rect 21097 35989 21131 36023
rect 22109 35989 22143 36023
rect 10793 35785 10827 35819
rect 11069 35785 11103 35819
rect 11713 35785 11747 35819
rect 12081 35785 12115 35819
rect 12817 35785 12851 35819
rect 13737 35785 13771 35819
rect 16037 35785 16071 35819
rect 16359 35785 16393 35819
rect 16497 35785 16531 35819
rect 16681 35785 16715 35819
rect 17325 35785 17359 35819
rect 17693 35785 17727 35819
rect 17877 35785 17911 35819
rect 18521 35785 18555 35819
rect 23213 35785 23247 35819
rect 28549 35785 28583 35819
rect 20453 35717 20487 35751
rect 10425 35649 10459 35683
rect 15025 35649 15059 35683
rect 15301 35649 15335 35683
rect 16589 35649 16623 35683
rect 17877 35649 17911 35683
rect 18061 35649 18095 35683
rect 20913 35649 20947 35683
rect 12725 35581 12759 35615
rect 13369 35581 13403 35615
rect 14381 35581 14415 35615
rect 14565 35581 14599 35615
rect 14841 35581 14875 35615
rect 18245 35581 18279 35615
rect 18337 35581 18371 35615
rect 19625 35581 19659 35615
rect 21189 35581 21223 35615
rect 12541 35513 12575 35547
rect 13921 35513 13955 35547
rect 16221 35513 16255 35547
rect 20177 35513 20211 35547
rect 22569 35513 22603 35547
rect 28273 35513 28307 35547
rect 10057 35445 10091 35479
rect 15761 35445 15795 35479
rect 19165 35445 19199 35479
rect 19809 35445 19843 35479
rect 23949 35445 23983 35479
rect 1777 35241 1811 35275
rect 11345 35241 11379 35275
rect 11713 35241 11747 35275
rect 13093 35241 13127 35275
rect 17509 35241 17543 35275
rect 18337 35241 18371 35275
rect 19717 35241 19751 35275
rect 21189 35241 21223 35275
rect 22753 35241 22787 35275
rect 10609 35173 10643 35207
rect 12357 35173 12391 35207
rect 12449 35173 12483 35207
rect 12725 35173 12759 35207
rect 13185 35173 13219 35207
rect 15301 35173 15335 35207
rect 16773 35173 16807 35207
rect 17693 35173 17727 35207
rect 18061 35173 18095 35207
rect 19441 35173 19475 35207
rect 22477 35173 22511 35207
rect 10241 35105 10275 35139
rect 11897 35105 11931 35139
rect 11805 35037 11839 35071
rect 10977 34969 11011 35003
rect 13829 35105 13863 35139
rect 14197 35105 14231 35139
rect 15945 35105 15979 35139
rect 16037 35105 16071 35139
rect 16313 35105 16347 35139
rect 17601 35105 17635 35139
rect 18889 35105 18923 35139
rect 19073 35105 19107 35139
rect 20453 35105 20487 35139
rect 21373 35105 21407 35139
rect 21557 35105 21591 35139
rect 21925 35105 21959 35139
rect 13737 35037 13771 35071
rect 14289 35037 14323 35071
rect 16405 35037 16439 35071
rect 17325 35037 17359 35071
rect 21833 35037 21867 35071
rect 23581 35037 23615 35071
rect 20085 34969 20119 35003
rect 24225 34969 24259 35003
rect 9413 34901 9447 34935
rect 12449 34901 12483 34935
rect 14657 34901 14691 34935
rect 15025 34901 15059 34935
rect 17141 34901 17175 34935
rect 18705 34901 18739 34935
rect 23121 34901 23155 34935
rect 23857 34901 23891 34935
rect 3065 34697 3099 34731
rect 8953 34697 8987 34731
rect 9229 34697 9263 34731
rect 11529 34697 11563 34731
rect 13369 34697 13403 34731
rect 13737 34697 13771 34731
rect 15577 34697 15611 34731
rect 16294 34697 16328 34731
rect 16773 34697 16807 34731
rect 19901 34697 19935 34731
rect 21465 34697 21499 34731
rect 23213 34697 23247 34731
rect 24685 34697 24719 34731
rect 27813 34697 27847 34731
rect 16405 34629 16439 34663
rect 19441 34629 19475 34663
rect 20821 34629 20855 34663
rect 21189 34629 21223 34663
rect 1685 34561 1719 34595
rect 9689 34561 9723 34595
rect 11897 34561 11931 34595
rect 12449 34561 12483 34595
rect 13829 34561 13863 34595
rect 16497 34561 16531 34595
rect 18797 34561 18831 34595
rect 26157 34561 26191 34595
rect 26525 34561 26559 34595
rect 29101 34561 29135 34595
rect 30665 34561 30699 34595
rect 1961 34493 1995 34527
rect 9413 34493 9447 34527
rect 12541 34493 12575 34527
rect 13001 34493 13035 34527
rect 14289 34493 14323 34527
rect 14473 34493 14507 34527
rect 14657 34493 14691 34527
rect 14933 34493 14967 34527
rect 15209 34493 15243 34527
rect 16037 34493 16071 34527
rect 17417 34493 17451 34527
rect 17877 34493 17911 34527
rect 18153 34493 18187 34527
rect 19073 34493 19107 34527
rect 19625 34493 19659 34527
rect 19717 34493 19751 34527
rect 21005 34493 21039 34527
rect 21833 34493 21867 34527
rect 22017 34493 22051 34527
rect 22569 34493 22603 34527
rect 23949 34493 23983 34527
rect 26249 34493 26283 34527
rect 29285 34493 29319 34527
rect 29561 34493 29595 34527
rect 12173 34425 12207 34459
rect 16129 34425 16163 34459
rect 22937 34425 22971 34459
rect 10977 34357 11011 34391
rect 20453 34357 20487 34391
rect 22201 34357 22235 34391
rect 24225 34357 24259 34391
rect 10609 34153 10643 34187
rect 12449 34153 12483 34187
rect 16313 34153 16347 34187
rect 17877 34153 17911 34187
rect 18797 34153 18831 34187
rect 19441 34153 19475 34187
rect 21189 34153 21223 34187
rect 24133 34153 24167 34187
rect 25053 34153 25087 34187
rect 29285 34153 29319 34187
rect 10333 34085 10367 34119
rect 11529 34085 11563 34119
rect 16405 34085 16439 34119
rect 17969 34085 18003 34119
rect 18337 34085 18371 34119
rect 19625 34085 19659 34119
rect 8861 34017 8895 34051
rect 11161 34017 11195 34051
rect 13001 34017 13035 34051
rect 13369 34017 13403 34051
rect 13553 34017 13587 34051
rect 16221 34017 16255 34051
rect 17785 34017 17819 34051
rect 19533 34017 19567 34051
rect 20913 34017 20947 34051
rect 21097 34017 21131 34051
rect 22753 34017 22787 34051
rect 27629 34017 27663 34051
rect 32413 34017 32447 34051
rect 11897 33949 11931 33983
rect 12817 33949 12851 33983
rect 15025 33949 15059 33983
rect 16037 33949 16071 33983
rect 16773 33949 16807 33983
rect 17601 33949 17635 33983
rect 19257 33949 19291 33983
rect 19993 33949 20027 33983
rect 23029 33949 23063 33983
rect 27353 33949 27387 33983
rect 32137 33949 32171 33983
rect 22109 33881 22143 33915
rect 25421 33881 25455 33915
rect 1777 33813 1811 33847
rect 8125 33813 8159 33847
rect 8493 33813 8527 33847
rect 8677 33813 8711 33847
rect 9505 33813 9539 33847
rect 9965 33813 9999 33847
rect 12265 33813 12299 33847
rect 13921 33813 13955 33847
rect 14289 33813 14323 33847
rect 14657 33813 14691 33847
rect 15577 33813 15611 33847
rect 15945 33813 15979 33847
rect 17417 33813 17451 33847
rect 19165 33813 19199 33847
rect 20269 33813 20303 33847
rect 20729 33813 20763 33847
rect 21741 33813 21775 33847
rect 22477 33813 22511 33847
rect 24685 33813 24719 33847
rect 26249 33813 26283 33847
rect 28733 33813 28767 33847
rect 33517 33813 33551 33847
rect 6469 33609 6503 33643
rect 7573 33609 7607 33643
rect 9413 33609 9447 33643
rect 10057 33609 10091 33643
rect 16865 33609 16899 33643
rect 17509 33609 17543 33643
rect 17877 33609 17911 33643
rect 19349 33609 19383 33643
rect 22201 33609 22235 33643
rect 23949 33609 23983 33643
rect 25605 33609 25639 33643
rect 27445 33609 27479 33643
rect 27813 33609 27847 33643
rect 32229 33609 32263 33643
rect 32505 33609 32539 33643
rect 10425 33541 10459 33575
rect 9045 33473 9079 33507
rect 11529 33473 11563 33507
rect 12449 33473 12483 33507
rect 14289 33473 14323 33507
rect 15669 33473 15703 33507
rect 6653 33405 6687 33439
rect 9505 33405 9539 33439
rect 10517 33405 10551 33439
rect 11069 33405 11103 33439
rect 11345 33405 11379 33439
rect 12265 33405 12299 33439
rect 13001 33405 13035 33439
rect 13277 33405 13311 33439
rect 13461 33405 13495 33439
rect 14841 33405 14875 33439
rect 15025 33405 15059 33439
rect 15117 33405 15151 33439
rect 15577 33405 15611 33439
rect 16589 33405 16623 33439
rect 16681 33405 16715 33439
rect 18337 33405 18371 33439
rect 7113 33337 7147 33371
rect 18061 33337 18095 33371
rect 18429 33337 18463 33371
rect 18797 33337 18831 33371
rect 19625 33473 19659 33507
rect 20361 33473 20395 33507
rect 20821 33473 20855 33507
rect 21189 33473 21223 33507
rect 19533 33405 19567 33439
rect 19809 33405 19843 33439
rect 20913 33405 20947 33439
rect 21925 33405 21959 33439
rect 23489 33405 23523 33439
rect 24133 33405 24167 33439
rect 24317 33405 24351 33439
rect 24685 33405 24719 33439
rect 24869 33405 24903 33439
rect 25237 33405 25271 33439
rect 19993 33337 20027 33371
rect 20821 33337 20855 33371
rect 21557 33337 21591 33371
rect 22845 33337 22879 33371
rect 25881 33337 25915 33371
rect 7849 33269 7883 33303
rect 8309 33269 8343 33303
rect 8585 33269 8619 33303
rect 9689 33269 9723 33303
rect 11897 33269 11931 33303
rect 13829 33269 13863 33303
rect 14197 33269 14231 33303
rect 16037 33269 16071 33303
rect 16405 33269 16439 33303
rect 18245 33269 18279 33303
rect 19073 33269 19107 33303
rect 19349 33269 19383 33303
rect 19901 33269 19935 33303
rect 21373 33269 21407 33303
rect 21465 33269 21499 33303
rect 23121 33269 23155 33303
rect 23305 33269 23339 33303
rect 26249 33269 26283 33303
rect 8125 33065 8159 33099
rect 8769 33065 8803 33099
rect 9505 33065 9539 33099
rect 11069 33065 11103 33099
rect 15485 33065 15519 33099
rect 17601 33065 17635 33099
rect 18613 33065 18647 33099
rect 20085 33065 20119 33099
rect 21925 33065 21959 33099
rect 25881 33065 25915 33099
rect 26709 33065 26743 33099
rect 8493 32997 8527 33031
rect 13185 32997 13219 33031
rect 16589 32997 16623 33031
rect 16773 32997 16807 33031
rect 21281 32997 21315 33031
rect 8585 32929 8619 32963
rect 9137 32929 9171 32963
rect 12173 32929 12207 32963
rect 13829 32929 13863 32963
rect 14197 32929 14231 32963
rect 14289 32929 14323 32963
rect 15301 32929 15335 32963
rect 16405 32929 16439 32963
rect 16681 32929 16715 32963
rect 17969 32929 18003 32963
rect 19533 32929 19567 32963
rect 21097 32929 21131 32963
rect 21189 32929 21223 32963
rect 22569 32929 22603 32963
rect 24225 32929 24259 32963
rect 27169 32929 27203 32963
rect 28641 32929 28675 32963
rect 28917 32929 28951 32963
rect 9689 32861 9723 32895
rect 9965 32861 9999 32895
rect 13093 32861 13127 32895
rect 13737 32861 13771 32895
rect 17141 32861 17175 32895
rect 18337 32861 18371 32895
rect 19349 32861 19383 32895
rect 20913 32861 20947 32895
rect 21649 32861 21683 32895
rect 22477 32861 22511 32895
rect 23673 32861 23707 32895
rect 23949 32861 23983 32895
rect 25329 32861 25363 32895
rect 12633 32793 12667 32827
rect 18245 32793 18279 32827
rect 22385 32793 22419 32827
rect 26341 32793 26375 32827
rect 11713 32725 11747 32759
rect 12081 32725 12115 32759
rect 12357 32725 12391 32759
rect 14657 32725 14691 32759
rect 15025 32725 15059 32759
rect 15945 32725 15979 32759
rect 18134 32725 18168 32759
rect 18981 32725 19015 32759
rect 19717 32725 19751 32759
rect 20729 32725 20763 32759
rect 22753 32725 22787 32759
rect 23305 32725 23339 32759
rect 30021 32725 30055 32759
rect 4905 32521 4939 32555
rect 5457 32521 5491 32555
rect 7757 32521 7791 32555
rect 9137 32521 9171 32555
rect 10425 32521 10459 32555
rect 11897 32521 11931 32555
rect 12173 32521 12207 32555
rect 12725 32521 12759 32555
rect 15393 32521 15427 32555
rect 16083 32521 16117 32555
rect 16957 32521 16991 32555
rect 17417 32521 17451 32555
rect 20545 32521 20579 32555
rect 22477 32521 22511 32555
rect 25053 32521 25087 32555
rect 25605 32521 25639 32555
rect 27169 32521 27203 32555
rect 28273 32521 28307 32555
rect 28457 32521 28491 32555
rect 28917 32521 28951 32555
rect 13093 32453 13127 32487
rect 16221 32453 16255 32487
rect 20802 32453 20836 32487
rect 20913 32453 20947 32487
rect 29469 32453 29503 32487
rect 8769 32385 8803 32419
rect 9505 32385 9539 32419
rect 10987 32385 11021 32419
rect 11529 32385 11563 32419
rect 13461 32385 13495 32419
rect 16313 32385 16347 32419
rect 19625 32385 19659 32419
rect 21005 32385 21039 32419
rect 22201 32385 22235 32419
rect 25973 32385 26007 32419
rect 5089 32317 5123 32351
rect 8217 32317 8251 32351
rect 8309 32317 8343 32351
rect 9597 32317 9631 32351
rect 9689 32317 9723 32351
rect 11069 32317 11103 32351
rect 12541 32317 12575 32351
rect 14013 32317 14047 32351
rect 14289 32317 14323 32351
rect 14381 32317 14415 32351
rect 14657 32317 14691 32351
rect 14933 32317 14967 32351
rect 15761 32317 15795 32351
rect 17693 32317 17727 32351
rect 18337 32317 18371 32351
rect 18797 32317 18831 32351
rect 18981 32317 19015 32351
rect 19165 32317 19199 32351
rect 19809 32317 19843 32351
rect 22293 32317 22327 32351
rect 23397 32317 23431 32351
rect 23673 32317 23707 32351
rect 23949 32317 23983 32351
rect 26157 32317 26191 32351
rect 27353 32317 27387 32351
rect 27629 32317 27663 32351
rect 28641 32317 28675 32351
rect 10149 32249 10183 32283
rect 10885 32249 10919 32283
rect 13553 32249 13587 32283
rect 15945 32249 15979 32283
rect 20637 32249 20671 32283
rect 21649 32249 21683 32283
rect 22109 32249 22143 32283
rect 26985 32249 27019 32283
rect 7389 32181 7423 32215
rect 8125 32181 8159 32215
rect 16589 32181 16623 32215
rect 17509 32181 17543 32215
rect 20177 32181 20211 32215
rect 21281 32181 21315 32215
rect 23029 32181 23063 32215
rect 26341 32181 26375 32215
rect 26617 32181 26651 32215
rect 7389 31977 7423 32011
rect 8493 31977 8527 32011
rect 10333 31977 10367 32011
rect 12817 31977 12851 32011
rect 13277 31977 13311 32011
rect 14657 31977 14691 32011
rect 16497 31977 16531 32011
rect 18981 31977 19015 32011
rect 21189 31977 21223 32011
rect 23305 31977 23339 32011
rect 24869 31977 24903 32011
rect 25145 31977 25179 32011
rect 8033 31909 8067 31943
rect 13093 31909 13127 31943
rect 7573 31841 7607 31875
rect 8585 31841 8619 31875
rect 10057 31841 10091 31875
rect 9137 31773 9171 31807
rect 10517 31773 10551 31807
rect 10793 31773 10827 31807
rect 7757 31705 7791 31739
rect 8769 31705 8803 31739
rect 9505 31705 9539 31739
rect 13461 31909 13495 31943
rect 13829 31909 13863 31943
rect 14013 31909 14047 31943
rect 19993 31909 20027 31943
rect 22845 31909 22879 31943
rect 23765 31909 23799 31943
rect 24409 31909 24443 31943
rect 26157 31909 26191 31943
rect 13921 31841 13955 31875
rect 14381 31841 14415 31875
rect 15577 31841 15611 31875
rect 15761 31841 15795 31875
rect 16129 31841 16163 31875
rect 16681 31841 16715 31875
rect 17601 31841 17635 31875
rect 18337 31841 18371 31875
rect 18429 31841 18463 31875
rect 18797 31841 18831 31875
rect 21373 31841 21407 31875
rect 21557 31841 21591 31875
rect 21925 31841 21959 31875
rect 22477 31841 22511 31875
rect 23581 31841 23615 31875
rect 23673 31841 23707 31875
rect 24961 31841 24995 31875
rect 26985 31841 27019 31875
rect 29193 31841 29227 31875
rect 29469 31841 29503 31875
rect 13645 31773 13679 31807
rect 15117 31773 15151 31807
rect 17509 31773 17543 31807
rect 23397 31773 23431 31807
rect 24133 31773 24167 31807
rect 25421 31773 25455 31807
rect 26709 31773 26743 31807
rect 28089 31773 28123 31807
rect 30573 31773 30607 31807
rect 25789 31705 25823 31739
rect 7113 31637 7147 31671
rect 11897 31637 11931 31671
rect 13277 31637 13311 31671
rect 17049 31637 17083 31671
rect 19625 31637 19659 31671
rect 20729 31637 20763 31671
rect 11897 31433 11931 31467
rect 13829 31433 13863 31467
rect 15853 31433 15887 31467
rect 22569 31433 22603 31467
rect 23121 31433 23155 31467
rect 26065 31433 26099 31467
rect 26801 31433 26835 31467
rect 27077 31433 27111 31467
rect 27445 31433 27479 31467
rect 28089 31433 28123 31467
rect 29469 31433 29503 31467
rect 14105 31365 14139 31399
rect 16221 31365 16255 31399
rect 19533 31365 19567 31399
rect 23489 31365 23523 31399
rect 6653 31297 6687 31331
rect 7573 31297 7607 31331
rect 7849 31297 7883 31331
rect 10701 31297 10735 31331
rect 10793 31297 10827 31331
rect 14749 31297 14783 31331
rect 15485 31297 15519 31331
rect 16405 31297 16439 31331
rect 17141 31297 17175 31331
rect 18797 31297 18831 31331
rect 19625 31297 19659 31331
rect 21189 31297 21223 31331
rect 21925 31297 21959 31331
rect 23673 31297 23707 31331
rect 25697 31297 25731 31331
rect 28457 31297 28491 31331
rect 12449 31229 12483 31263
rect 12909 31229 12943 31263
rect 13277 31229 13311 31263
rect 13369 31229 13403 31263
rect 14933 31229 14967 31263
rect 18337 31229 18371 31263
rect 19809 31229 19843 31263
rect 21097 31229 21131 31263
rect 21373 31229 21407 31263
rect 25237 31229 25271 31263
rect 26249 31229 26283 31263
rect 27261 31229 27295 31263
rect 27721 31229 27755 31263
rect 10333 31161 10367 31195
rect 11069 31161 11103 31195
rect 11161 31161 11195 31195
rect 11529 31161 11563 31195
rect 15117 31161 15151 31195
rect 16681 31161 16715 31195
rect 16773 31161 16807 31195
rect 17877 31161 17911 31195
rect 18061 31161 18095 31195
rect 18429 31161 18463 31195
rect 19073 31161 19107 31195
rect 19901 31161 19935 31195
rect 19993 31161 20027 31195
rect 20361 31161 20395 31195
rect 21557 31161 21591 31195
rect 23857 31161 23891 31195
rect 24041 31161 24075 31195
rect 24409 31161 24443 31195
rect 25145 31161 25179 31195
rect 7021 31093 7055 31127
rect 7481 31093 7515 31127
rect 8953 31093 8987 31127
rect 9597 31093 9631 31127
rect 9965 31093 9999 31127
rect 10977 31093 11011 31127
rect 12265 31093 12299 31127
rect 14565 31093 14599 31127
rect 15025 31093 15059 31127
rect 16589 31093 16623 31127
rect 17509 31093 17543 31127
rect 18245 31093 18279 31127
rect 20637 31093 20671 31127
rect 21465 31093 21499 31127
rect 22201 31093 22235 31127
rect 23949 31093 23983 31127
rect 24685 31093 24719 31127
rect 25421 31093 25455 31127
rect 26433 31093 26467 31127
rect 28825 31093 28859 31127
rect 29837 31093 29871 31127
rect 6745 30889 6779 30923
rect 7757 30889 7791 30923
rect 8769 30889 8803 30923
rect 10333 30889 10367 30923
rect 11253 30889 11287 30923
rect 13553 30889 13587 30923
rect 15485 30889 15519 30923
rect 18061 30889 18095 30923
rect 18797 30889 18831 30923
rect 19257 30889 19291 30923
rect 20729 30889 20763 30923
rect 21189 30889 21223 30923
rect 21925 30889 21959 30923
rect 22937 30889 22971 30923
rect 23765 30889 23799 30923
rect 24685 30889 24719 30923
rect 25973 30889 26007 30923
rect 13829 30821 13863 30855
rect 14013 30821 14047 30855
rect 14381 30821 14415 30855
rect 16313 30821 16347 30855
rect 16681 30821 16715 30855
rect 17049 30821 17083 30855
rect 18153 30821 18187 30855
rect 21281 30821 21315 30855
rect 21649 30821 21683 30855
rect 22385 30821 22419 30855
rect 7573 30753 7607 30787
rect 8585 30753 8619 30787
rect 10149 30753 10183 30787
rect 11805 30753 11839 30787
rect 12173 30753 12207 30787
rect 13921 30753 13955 30787
rect 15025 30753 15059 30787
rect 15301 30753 15335 30787
rect 16497 30753 16531 30787
rect 16589 30753 16623 30787
rect 17325 30753 17359 30787
rect 19625 30753 19659 30787
rect 19809 30753 19843 30787
rect 21097 30753 21131 30787
rect 22477 30753 22511 30787
rect 22753 30753 22787 30787
rect 24041 30753 24075 30787
rect 7481 30685 7515 30719
rect 9045 30685 9079 30719
rect 10057 30685 10091 30719
rect 11621 30685 11655 30719
rect 12081 30685 12115 30719
rect 12725 30685 12759 30719
rect 13185 30685 13219 30719
rect 13645 30685 13679 30719
rect 14749 30685 14783 30719
rect 18521 30685 18555 30719
rect 20913 30685 20947 30719
rect 24409 30685 24443 30719
rect 27169 30685 27203 30719
rect 27445 30685 27479 30719
rect 7113 30617 7147 30651
rect 18429 30617 18463 30651
rect 20361 30617 20395 30651
rect 22569 30617 22603 30651
rect 24317 30617 24351 30651
rect 25605 30617 25639 30651
rect 8125 30549 8159 30583
rect 8493 30549 8527 30583
rect 9413 30549 9447 30583
rect 10885 30549 10919 30583
rect 15761 30549 15795 30583
rect 16221 30549 16255 30583
rect 18318 30549 18352 30583
rect 19993 30549 20027 30583
rect 24179 30549 24213 30583
rect 25329 30549 25363 30583
rect 26709 30549 26743 30583
rect 28549 30549 28583 30583
rect 7573 30345 7607 30379
rect 9137 30345 9171 30379
rect 9965 30345 9999 30379
rect 11805 30345 11839 30379
rect 14197 30345 14231 30379
rect 16313 30345 16347 30379
rect 23305 30345 23339 30379
rect 24133 30345 24167 30379
rect 6285 30277 6319 30311
rect 12173 30277 12207 30311
rect 12725 30277 12759 30311
rect 17877 30277 17911 30311
rect 19073 30277 19107 30311
rect 22017 30277 22051 30311
rect 22293 30277 22327 30311
rect 26617 30277 26651 30311
rect 28733 30277 28767 30311
rect 7665 30209 7699 30243
rect 8125 30209 8159 30243
rect 13185 30209 13219 30243
rect 13921 30209 13955 30243
rect 14749 30209 14783 30243
rect 15485 30209 15519 30243
rect 17141 30209 17175 30243
rect 18061 30209 18095 30243
rect 19993 30209 20027 30243
rect 23673 30209 23707 30243
rect 8309 30141 8343 30175
rect 8677 30141 8711 30175
rect 8769 30141 8803 30175
rect 9781 30141 9815 30175
rect 11069 30141 11103 30175
rect 13093 30141 13127 30175
rect 13369 30141 13403 30175
rect 14473 30141 14507 30175
rect 14933 30141 14967 30175
rect 17509 30141 17543 30175
rect 18245 30141 18279 30175
rect 19901 30141 19935 30175
rect 20177 30141 20211 30175
rect 20545 30141 20579 30175
rect 21189 30141 21223 30175
rect 21649 30141 21683 30175
rect 22477 30141 22511 30175
rect 23949 30141 23983 30175
rect 25973 30141 26007 30175
rect 26801 30141 26835 30175
rect 26893 30141 26927 30175
rect 7205 30073 7239 30107
rect 10793 30073 10827 30107
rect 11161 30073 11195 30107
rect 11529 30073 11563 30107
rect 13553 30073 13587 30107
rect 14565 30073 14599 30107
rect 15117 30073 15151 30107
rect 16405 30073 16439 30107
rect 16773 30073 16807 30107
rect 18429 30073 18463 30107
rect 18797 30073 18831 30107
rect 22937 30073 22971 30107
rect 23857 30073 23891 30107
rect 25237 30073 25271 30107
rect 25421 30073 25455 30107
rect 25605 30073 25639 30107
rect 27353 30073 27387 30107
rect 28089 30073 28123 30107
rect 6653 30005 6687 30039
rect 9689 30005 9723 30039
rect 10333 30005 10367 30039
rect 10701 30005 10735 30039
rect 10977 30005 11011 30039
rect 13461 30005 13495 30039
rect 14473 30005 14507 30039
rect 15025 30005 15059 30039
rect 15853 30005 15887 30039
rect 16589 30005 16623 30039
rect 16681 30005 16715 30039
rect 18337 30005 18371 30039
rect 19533 30005 19567 30039
rect 22661 30005 22695 30039
rect 24685 30005 24719 30039
rect 25053 30005 25087 30039
rect 25513 30005 25547 30039
rect 26249 30005 26283 30039
rect 27629 30005 27663 30039
rect 28457 30005 28491 30039
rect 29469 30005 29503 30039
rect 2973 29801 3007 29835
rect 6745 29801 6779 29835
rect 9505 29801 9539 29835
rect 10333 29801 10367 29835
rect 11437 29801 11471 29835
rect 13277 29801 13311 29835
rect 14841 29801 14875 29835
rect 15485 29801 15519 29835
rect 16037 29801 16071 29835
rect 17233 29801 17267 29835
rect 17693 29801 17727 29835
rect 17969 29801 18003 29835
rect 18981 29801 19015 29835
rect 20177 29801 20211 29835
rect 20361 29801 20395 29835
rect 21189 29801 21223 29835
rect 21833 29801 21867 29835
rect 21925 29801 21959 29835
rect 22293 29801 22327 29835
rect 23581 29801 23615 29835
rect 23949 29801 23983 29835
rect 25605 29801 25639 29835
rect 25973 29801 26007 29835
rect 26709 29801 26743 29835
rect 27629 29801 27663 29835
rect 28273 29801 28307 29835
rect 8493 29733 8527 29767
rect 1409 29665 1443 29699
rect 7113 29665 7147 29699
rect 9137 29665 9171 29699
rect 9781 29665 9815 29699
rect 10793 29665 10827 29699
rect 1685 29597 1719 29631
rect 6837 29597 6871 29631
rect 12173 29733 12207 29767
rect 12541 29733 12575 29767
rect 16221 29733 16255 29767
rect 16589 29733 16623 29767
rect 18153 29733 18187 29767
rect 19349 29733 19383 29767
rect 11989 29665 12023 29699
rect 12081 29665 12115 29699
rect 14197 29665 14231 29699
rect 16405 29665 16439 29699
rect 16497 29665 16531 29699
rect 18061 29665 18095 29699
rect 19533 29665 19567 29699
rect 11805 29597 11839 29631
rect 13369 29597 13403 29631
rect 13921 29597 13955 29631
rect 14381 29597 14415 29631
rect 16957 29597 16991 29631
rect 17785 29597 17819 29631
rect 18521 29597 18555 29631
rect 19441 29597 19475 29631
rect 19993 29597 20027 29631
rect 9965 29529 9999 29563
rect 10977 29529 11011 29563
rect 11345 29529 11379 29563
rect 11437 29529 11471 29563
rect 21281 29733 21315 29767
rect 21097 29665 21131 29699
rect 20913 29597 20947 29631
rect 21649 29597 21683 29631
rect 24777 29733 24811 29767
rect 25329 29733 25363 29767
rect 26893 29733 26927 29767
rect 27261 29733 27295 29767
rect 23029 29665 23063 29699
rect 24041 29665 24075 29699
rect 24317 29665 24351 29699
rect 26525 29665 26559 29699
rect 26801 29665 26835 29699
rect 24133 29529 24167 29563
rect 10701 29461 10735 29495
rect 11713 29461 11747 29495
rect 12817 29461 12851 29495
rect 20177 29461 20211 29495
rect 20637 29461 20671 29495
rect 21833 29461 21867 29495
rect 22937 29461 22971 29495
rect 27905 29461 27939 29495
rect 28733 29461 28767 29495
rect 1961 29257 1995 29291
rect 6653 29257 6687 29291
rect 7113 29257 7147 29291
rect 9413 29257 9447 29291
rect 9781 29257 9815 29291
rect 10241 29257 10275 29291
rect 10517 29257 10551 29291
rect 11897 29257 11931 29291
rect 12265 29257 12299 29291
rect 12725 29257 12759 29291
rect 15577 29257 15611 29291
rect 16221 29257 16255 29291
rect 16405 29257 16439 29291
rect 17509 29257 17543 29291
rect 19717 29257 19751 29291
rect 20177 29257 20211 29291
rect 23121 29257 23155 29291
rect 23489 29257 23523 29291
rect 25605 29257 25639 29291
rect 26065 29257 26099 29291
rect 27997 29257 28031 29291
rect 29469 29257 29503 29291
rect 11529 29189 11563 29223
rect 13277 29189 13311 29223
rect 14933 29189 14967 29223
rect 21373 29189 21407 29223
rect 21833 29189 21867 29223
rect 27629 29189 27663 29223
rect 28273 29189 28307 29223
rect 7573 29121 7607 29155
rect 14289 29121 14323 29155
rect 17785 29121 17819 29155
rect 20361 29121 20395 29155
rect 21925 29121 21959 29155
rect 23949 29121 23983 29155
rect 26249 29121 26283 29155
rect 27169 29121 27203 29155
rect 7297 29053 7331 29087
rect 10333 29053 10367 29087
rect 10885 29053 10919 29087
rect 11345 29053 11379 29087
rect 13829 29053 13863 29087
rect 14013 29053 14047 29087
rect 14381 29053 14415 29087
rect 15393 29053 15427 29087
rect 15853 29053 15887 29087
rect 16681 29053 16715 29087
rect 20545 29053 20579 29087
rect 22201 29053 22235 29087
rect 23673 29053 23707 29087
rect 27077 29053 27111 29087
rect 28089 29053 28123 29087
rect 28549 29053 28583 29087
rect 11253 28985 11287 29019
rect 13369 28985 13403 29019
rect 15301 28985 15335 29019
rect 16589 28985 16623 29019
rect 17141 28985 17175 29019
rect 18429 28985 18463 29019
rect 18613 28985 18647 29019
rect 18981 28985 19015 29019
rect 19349 28985 19383 29019
rect 20729 28985 20763 29019
rect 21097 28985 21131 29019
rect 22293 28985 22327 29019
rect 22661 28985 22695 29019
rect 25329 28985 25363 29019
rect 26341 28985 26375 29019
rect 29009 28985 29043 29019
rect 1685 28917 1719 28951
rect 8677 28917 8711 28951
rect 18797 28917 18831 28951
rect 18889 28917 18923 28951
rect 20637 28917 20671 28951
rect 22109 28917 22143 28951
rect 9413 28713 9447 28747
rect 10609 28713 10643 28747
rect 11805 28713 11839 28747
rect 12357 28713 12391 28747
rect 13829 28713 13863 28747
rect 14749 28713 14783 28747
rect 16957 28713 16991 28747
rect 18613 28713 18647 28747
rect 20361 28713 20395 28747
rect 21925 28713 21959 28747
rect 22661 28713 22695 28747
rect 23581 28713 23615 28747
rect 23949 28713 23983 28747
rect 25145 28713 25179 28747
rect 25881 28713 25915 28747
rect 26249 28713 26283 28747
rect 27629 28713 27663 28747
rect 27997 28713 28031 28747
rect 29009 28713 29043 28747
rect 7573 28645 7607 28679
rect 9137 28645 9171 28679
rect 18797 28645 18831 28679
rect 19993 28645 20027 28679
rect 20729 28645 20763 28679
rect 21097 28645 21131 28679
rect 21281 28645 21315 28679
rect 21741 28645 21775 28679
rect 22845 28645 22879 28679
rect 26525 28645 26559 28679
rect 8217 28577 8251 28611
rect 8585 28577 8619 28611
rect 8769 28577 8803 28611
rect 10793 28577 10827 28611
rect 12909 28577 12943 28611
rect 13277 28577 13311 28611
rect 16129 28577 16163 28611
rect 17417 28577 17451 28611
rect 18705 28577 18739 28611
rect 21189 28577 21223 28611
rect 8309 28509 8343 28543
rect 12817 28509 12851 28543
rect 13185 28509 13219 28543
rect 15301 28509 15335 28543
rect 15853 28509 15887 28543
rect 16313 28509 16347 28543
rect 18429 28509 18463 28543
rect 19165 28509 19199 28543
rect 20913 28509 20947 28543
rect 21649 28509 21683 28543
rect 22753 28577 22787 28611
rect 24225 28577 24259 28611
rect 28089 28577 28123 28611
rect 32689 28577 32723 28611
rect 22477 28509 22511 28543
rect 23213 28509 23247 28543
rect 26893 28509 26927 28543
rect 32413 28509 32447 28543
rect 10241 28441 10275 28475
rect 18337 28441 18371 28475
rect 21741 28441 21775 28475
rect 22293 28441 22327 28475
rect 26690 28441 26724 28475
rect 28273 28441 28307 28475
rect 6929 28373 6963 28407
rect 7297 28373 7331 28407
rect 11161 28373 11195 28407
rect 14289 28373 14323 28407
rect 15117 28373 15151 28407
rect 16681 28373 16715 28407
rect 17601 28373 17635 28407
rect 17969 28373 18003 28407
rect 19441 28373 19475 28407
rect 24317 28373 24351 28407
rect 25513 28373 25547 28407
rect 26801 28373 26835 28407
rect 27169 28373 27203 28407
rect 28549 28373 28583 28407
rect 33793 28373 33827 28407
rect 1685 28169 1719 28203
rect 2237 28169 2271 28203
rect 8401 28169 8435 28203
rect 9505 28169 9539 28203
rect 10241 28169 10275 28203
rect 10517 28169 10551 28203
rect 10793 28169 10827 28203
rect 12909 28169 12943 28203
rect 14013 28169 14047 28203
rect 17785 28169 17819 28203
rect 18521 28169 18555 28203
rect 18889 28169 18923 28203
rect 21281 28169 21315 28203
rect 22661 28169 22695 28203
rect 23949 28169 23983 28203
rect 25881 28169 25915 28203
rect 26249 28169 26283 28203
rect 28089 28169 28123 28203
rect 28641 28169 28675 28203
rect 29101 28169 29135 28203
rect 32505 28169 32539 28203
rect 32781 28169 32815 28203
rect 8769 28101 8803 28135
rect 11621 28101 11655 28135
rect 11897 28101 11931 28135
rect 20729 28101 20763 28135
rect 9137 28033 9171 28067
rect 13645 28033 13679 28067
rect 15761 28033 15795 28067
rect 16313 28033 16347 28067
rect 17417 28033 17451 28067
rect 19257 28033 19291 28067
rect 23121 28101 23155 28135
rect 25513 28101 25547 28135
rect 21557 28033 21591 28067
rect 21649 28033 21683 28067
rect 24133 28033 24167 28067
rect 25145 28033 25179 28067
rect 26709 28033 26743 28067
rect 1409 27965 1443 27999
rect 1593 27965 1627 27999
rect 7665 27965 7699 27999
rect 9321 27965 9355 27999
rect 10333 27965 10367 27999
rect 11345 27965 11379 27999
rect 11621 27965 11655 27999
rect 12725 27965 12759 27999
rect 14197 27965 14231 27999
rect 14381 27965 14415 27999
rect 14749 27965 14783 27999
rect 14933 27965 14967 27999
rect 16589 27965 16623 27999
rect 16773 27965 16807 27999
rect 18337 27965 18371 27999
rect 19625 27965 19659 27999
rect 19809 27965 19843 27999
rect 20361 27965 20395 27999
rect 20637 27965 20671 27999
rect 21281 27965 21315 27999
rect 22001 27965 22035 27999
rect 24317 27965 24351 27999
rect 24685 27965 24719 27999
rect 24869 27965 24903 27999
rect 25697 27965 25731 27999
rect 26985 27965 27019 27999
rect 29285 27965 29319 27999
rect 29745 27965 29779 27999
rect 7297 27897 7331 27931
rect 21833 27897 21867 27931
rect 22385 27897 22419 27931
rect 8033 27829 8067 27863
rect 9873 27829 9907 27863
rect 11253 27829 11287 27863
rect 11529 27829 11563 27863
rect 12265 27829 12299 27863
rect 13277 27829 13311 27863
rect 15301 27829 15335 27863
rect 17049 27829 17083 27863
rect 21097 27829 21131 27863
rect 21925 27829 21959 27863
rect 23489 27829 23523 27863
rect 26525 27829 26559 27863
rect 29469 27829 29503 27863
rect 8677 27625 8711 27659
rect 10793 27625 10827 27659
rect 12449 27625 12483 27659
rect 12909 27625 12943 27659
rect 18429 27625 18463 27659
rect 18889 27625 18923 27659
rect 20729 27625 20763 27659
rect 22109 27625 22143 27659
rect 10517 27557 10551 27591
rect 11161 27557 11195 27591
rect 13001 27557 13035 27591
rect 14841 27557 14875 27591
rect 16221 27557 16255 27591
rect 17417 27557 17451 27591
rect 17785 27557 17819 27591
rect 19993 27557 20027 27591
rect 20913 27557 20947 27591
rect 6745 27489 6779 27523
rect 10609 27489 10643 27523
rect 11713 27489 11747 27523
rect 13829 27489 13863 27523
rect 14013 27489 14047 27523
rect 15853 27489 15887 27523
rect 16037 27489 16071 27523
rect 16129 27489 16163 27523
rect 17325 27489 17359 27523
rect 17601 27489 17635 27523
rect 17693 27489 17727 27523
rect 18981 27489 19015 27523
rect 21060 27489 21094 27523
rect 21925 27489 21959 27523
rect 7021 27421 7055 27455
rect 9045 27421 9079 27455
rect 10149 27421 10183 27455
rect 11621 27421 11655 27455
rect 13553 27421 13587 27455
rect 14473 27421 14507 27455
rect 16589 27421 16623 27455
rect 18153 27421 18187 27455
rect 19349 27421 19383 27455
rect 21281 27421 21315 27455
rect 15761 27353 15795 27387
rect 19146 27353 19180 27387
rect 21189 27353 21223 27387
rect 22201 27625 22235 27659
rect 26249 27625 26283 27659
rect 26709 27625 26743 27659
rect 26985 27625 27019 27659
rect 23489 27557 23523 27591
rect 24041 27557 24075 27591
rect 24409 27557 24443 27591
rect 25789 27557 25823 27591
rect 27353 27557 27387 27591
rect 28825 27557 28859 27591
rect 22477 27489 22511 27523
rect 23213 27489 23247 27523
rect 24225 27489 24259 27523
rect 24317 27489 24351 27523
rect 26525 27489 26559 27523
rect 27537 27489 27571 27523
rect 28365 27489 28399 27523
rect 22845 27421 22879 27455
rect 24777 27421 24811 27455
rect 22201 27353 22235 27387
rect 25421 27353 25455 27387
rect 1593 27285 1627 27319
rect 8309 27285 8343 27319
rect 9413 27285 9447 27319
rect 11529 27285 11563 27319
rect 11897 27285 11931 27319
rect 16865 27285 16899 27319
rect 19257 27285 19291 27319
rect 19625 27285 19659 27319
rect 21557 27285 21591 27319
rect 22109 27285 22143 27319
rect 22293 27285 22327 27319
rect 22615 27285 22649 27319
rect 22753 27285 22787 27319
rect 23857 27285 23891 27319
rect 25053 27285 25087 27319
rect 27721 27285 27755 27319
rect 27997 27285 28031 27319
rect 7389 27081 7423 27115
rect 9505 27081 9539 27115
rect 14657 27081 14691 27115
rect 16037 27081 16071 27115
rect 16405 27081 16439 27115
rect 16865 27081 16899 27115
rect 17785 27081 17819 27115
rect 18797 27081 18831 27115
rect 22937 27081 22971 27115
rect 25421 27081 25455 27115
rect 25789 27081 25823 27115
rect 26065 27081 26099 27115
rect 27077 27081 27111 27115
rect 28457 27081 28491 27115
rect 9229 27013 9263 27047
rect 11805 27013 11839 27047
rect 12265 27013 12299 27047
rect 18429 27013 18463 27047
rect 22385 27013 22419 27047
rect 23489 27013 23523 27047
rect 23949 27013 23983 27047
rect 1869 26945 1903 26979
rect 10425 26945 10459 26979
rect 10885 26945 10919 26979
rect 13599 26945 13633 26979
rect 16589 26945 16623 26979
rect 20269 26945 20303 26979
rect 1593 26877 1627 26911
rect 8309 26877 8343 26911
rect 9321 26877 9355 26911
rect 10977 26877 11011 26911
rect 11345 26877 11379 26911
rect 11437 26877 11471 26911
rect 12909 26877 12943 26911
rect 13461 26877 13495 26911
rect 13737 26877 13771 26911
rect 14749 26877 14783 26911
rect 15209 26877 15243 26911
rect 15577 26877 15611 26911
rect 15669 26877 15703 26911
rect 16681 26877 16715 26911
rect 17417 26877 17451 26911
rect 18245 26877 18279 26911
rect 19441 26877 19475 26911
rect 19625 26877 19659 26911
rect 19993 26877 20027 26911
rect 20545 26877 20579 26911
rect 21005 26877 21039 26911
rect 3249 26809 3283 26843
rect 8861 26809 8895 26843
rect 21557 26809 21591 26843
rect 21833 26809 21867 26843
rect 21925 26809 21959 26843
rect 22293 26809 22327 26843
rect 24041 26945 24075 26979
rect 23673 26877 23707 26911
rect 23820 26877 23854 26911
rect 25237 26877 25271 26911
rect 26249 26877 26283 26911
rect 27261 26877 27295 26911
rect 27721 26877 27755 26911
rect 28089 26877 28123 26911
rect 22661 26809 22695 26843
rect 25053 26809 25087 26843
rect 7113 26741 7147 26775
rect 8493 26741 8527 26775
rect 9873 26741 9907 26775
rect 10241 26741 10275 26775
rect 12817 26741 12851 26775
rect 14289 26741 14323 26775
rect 19073 26741 19107 26775
rect 21373 26741 21407 26775
rect 21741 26741 21775 26775
rect 22385 26741 22419 26775
rect 24317 26741 24351 26775
rect 24777 26741 24811 26775
rect 26433 26741 26467 26775
rect 26709 26741 26743 26775
rect 27445 26741 27479 26775
rect 1685 26537 1719 26571
rect 7481 26537 7515 26571
rect 10057 26537 10091 26571
rect 11897 26537 11931 26571
rect 13093 26537 13127 26571
rect 14657 26537 14691 26571
rect 16405 26537 16439 26571
rect 20361 26537 20395 26571
rect 20729 26537 20763 26571
rect 22385 26537 22419 26571
rect 25789 26537 25823 26571
rect 28089 26537 28123 26571
rect 13369 26469 13403 26503
rect 15117 26469 15151 26503
rect 19165 26469 19199 26503
rect 19257 26469 19291 26503
rect 21649 26469 21683 26503
rect 22477 26469 22511 26503
rect 23765 26469 23799 26503
rect 26157 26469 26191 26503
rect 1961 26401 1995 26435
rect 6101 26401 6135 26435
rect 6377 26401 6411 26435
rect 8585 26401 8619 26435
rect 9137 26401 9171 26435
rect 9505 26401 9539 26435
rect 10793 26401 10827 26435
rect 12541 26401 12575 26435
rect 14197 26401 14231 26435
rect 15577 26401 15611 26435
rect 16681 26401 16715 26435
rect 17417 26401 17451 26435
rect 17601 26401 17635 26435
rect 18889 26401 18923 26435
rect 19073 26401 19107 26435
rect 19993 26401 20027 26435
rect 20913 26401 20947 26435
rect 22624 26401 22658 26435
rect 24409 26401 24443 26435
rect 26525 26401 26559 26435
rect 27537 26401 27571 26435
rect 10517 26333 10551 26367
rect 13921 26333 13955 26367
rect 14381 26333 14415 26367
rect 18705 26333 18739 26367
rect 19625 26333 19659 26367
rect 21060 26333 21094 26367
rect 21281 26333 21315 26367
rect 22017 26333 22051 26367
rect 22845 26333 22879 26367
rect 24041 26333 24075 26367
rect 27077 26333 27111 26367
rect 27445 26333 27479 26367
rect 8769 26265 8803 26299
rect 10333 26265 10367 26299
rect 15761 26265 15795 26299
rect 17417 26265 17451 26299
rect 18061 26265 18095 26299
rect 21189 26265 21223 26299
rect 22937 26265 22971 26299
rect 25053 26265 25087 26299
rect 25513 26265 25547 26299
rect 27721 26265 27755 26299
rect 16129 26197 16163 26231
rect 18337 26197 18371 26231
rect 22753 26197 22787 26231
rect 26709 26197 26743 26231
rect 6469 25993 6503 26027
rect 8677 25993 8711 26027
rect 13461 25993 13495 26027
rect 14933 25993 14967 26027
rect 15301 25993 15335 26027
rect 16681 25993 16715 26027
rect 17877 25993 17911 26027
rect 21097 25993 21131 26027
rect 21465 25993 21499 26027
rect 23213 25993 23247 26027
rect 25329 25993 25363 26027
rect 27077 25993 27111 26027
rect 27629 25993 27663 26027
rect 11529 25925 11563 25959
rect 20177 25925 20211 25959
rect 20729 25925 20763 25959
rect 22293 25925 22327 25959
rect 25697 25925 25731 25959
rect 9321 25857 9355 25891
rect 16405 25857 16439 25891
rect 18337 25857 18371 25891
rect 8309 25789 8343 25823
rect 9045 25789 9079 25823
rect 12265 25789 12299 25823
rect 12449 25789 12483 25823
rect 12633 25789 12667 25823
rect 13829 25789 13863 25823
rect 14013 25789 14047 25823
rect 15393 25789 15427 25823
rect 15945 25789 15979 25823
rect 16221 25789 16255 25823
rect 18153 25789 18187 25823
rect 18705 25789 18739 25823
rect 18889 25789 18923 25823
rect 19257 25789 19291 25823
rect 19625 25789 19659 25823
rect 11897 25721 11931 25755
rect 14197 25721 14231 25755
rect 14565 25721 14599 25755
rect 17509 25721 17543 25755
rect 21189 25857 21223 25891
rect 24317 25857 24351 25891
rect 24777 25857 24811 25891
rect 26709 25857 26743 25891
rect 20968 25789 21002 25823
rect 21925 25789 21959 25823
rect 22385 25789 22419 25823
rect 24501 25789 24535 25823
rect 24869 25789 24903 25823
rect 25881 25789 25915 25823
rect 26065 25789 26099 25823
rect 20821 25721 20855 25755
rect 26433 25721 26467 25755
rect 6101 25653 6135 25687
rect 10609 25653 10643 25687
rect 11161 25653 11195 25687
rect 12725 25653 12759 25687
rect 14105 25653 14139 25687
rect 17141 25653 17175 25687
rect 20177 25653 20211 25687
rect 20269 25653 20303 25687
rect 22569 25653 22603 25687
rect 22845 25653 22879 25687
rect 24133 25653 24167 25687
rect 9137 25449 9171 25483
rect 9505 25449 9539 25483
rect 11345 25449 11379 25483
rect 12173 25449 12207 25483
rect 12449 25449 12483 25483
rect 12909 25449 12943 25483
rect 13277 25449 13311 25483
rect 14749 25449 14783 25483
rect 15577 25449 15611 25483
rect 16497 25449 16531 25483
rect 20085 25449 20119 25483
rect 21097 25449 21131 25483
rect 22753 25449 22787 25483
rect 25329 25449 25363 25483
rect 26709 25449 26743 25483
rect 22477 25381 22511 25415
rect 26985 25381 27019 25415
rect 10149 25313 10183 25347
rect 10333 25313 10367 25347
rect 10701 25313 10735 25347
rect 10793 25313 10827 25347
rect 12265 25313 12299 25347
rect 13829 25313 13863 25347
rect 14197 25313 14231 25347
rect 15393 25313 15427 25347
rect 16957 25313 16991 25347
rect 17049 25313 17083 25347
rect 17233 25313 17267 25347
rect 17509 25313 17543 25347
rect 17877 25313 17911 25347
rect 18981 25313 19015 25347
rect 19533 25313 19567 25347
rect 19717 25313 19751 25347
rect 22293 25313 22327 25347
rect 23121 25313 23155 25347
rect 23397 25313 23431 25347
rect 25697 25313 25731 25347
rect 26525 25313 26559 25347
rect 9689 25245 9723 25279
rect 14289 25245 14323 25279
rect 16313 25245 16347 25279
rect 23673 25245 23707 25279
rect 26065 25245 26099 25279
rect 11805 25177 11839 25211
rect 13645 25177 13679 25211
rect 18521 25177 18555 25211
rect 19533 25177 19567 25211
rect 15117 25109 15151 25143
rect 15945 25109 15979 25143
rect 18245 25109 18279 25143
rect 20453 25109 20487 25143
rect 21465 25109 21499 25143
rect 24961 25109 24995 25143
rect 11897 24905 11931 24939
rect 14749 24905 14783 24939
rect 15393 24905 15427 24939
rect 19625 24905 19659 24939
rect 23029 24905 23063 24939
rect 23489 24905 23523 24939
rect 26617 24905 26651 24939
rect 14105 24837 14139 24871
rect 20361 24837 20395 24871
rect 8953 24769 8987 24803
rect 9413 24769 9447 24803
rect 10517 24769 10551 24803
rect 11069 24769 11103 24803
rect 14473 24769 14507 24803
rect 18061 24769 18095 24803
rect 18797 24769 18831 24803
rect 20453 24769 20487 24803
rect 22661 24769 22695 24803
rect 23673 24769 23707 24803
rect 24593 24769 24627 24803
rect 24961 24769 24995 24803
rect 25881 24769 25915 24803
rect 9137 24701 9171 24735
rect 13001 24701 13035 24735
rect 13185 24701 13219 24735
rect 13553 24701 13587 24735
rect 13737 24701 13771 24735
rect 14565 24701 14599 24735
rect 16129 24701 16163 24735
rect 16681 24701 16715 24735
rect 16865 24701 16899 24735
rect 18705 24701 18739 24735
rect 19073 24701 19107 24735
rect 19165 24701 19199 24735
rect 19901 24701 19935 24735
rect 20232 24701 20266 24735
rect 20821 24701 20855 24735
rect 21097 24701 21131 24735
rect 21649 24701 21683 24735
rect 21741 24701 21775 24735
rect 23765 24701 23799 24735
rect 25053 24701 25087 24735
rect 25513 24701 25547 24735
rect 20085 24633 20119 24667
rect 24225 24633 24259 24667
rect 8677 24565 8711 24599
rect 11437 24565 11471 24599
rect 12265 24565 12299 24599
rect 12817 24565 12851 24599
rect 15025 24565 15059 24599
rect 16129 24565 16163 24599
rect 17509 24565 17543 24599
rect 17785 24565 17819 24599
rect 21465 24565 21499 24599
rect 25237 24565 25271 24599
rect 7941 24361 7975 24395
rect 9413 24361 9447 24395
rect 10241 24361 10275 24395
rect 10609 24361 10643 24395
rect 10977 24361 11011 24395
rect 11989 24361 12023 24395
rect 13369 24361 13403 24395
rect 14749 24361 14783 24395
rect 15761 24361 15795 24395
rect 18153 24361 18187 24395
rect 19441 24361 19475 24395
rect 19901 24361 19935 24395
rect 20637 24361 20671 24395
rect 21097 24361 21131 24395
rect 21925 24361 21959 24395
rect 22753 24361 22787 24395
rect 23305 24361 23339 24395
rect 23765 24361 23799 24395
rect 24777 24361 24811 24395
rect 13645 24293 13679 24327
rect 14381 24293 14415 24327
rect 21281 24293 21315 24327
rect 24409 24293 24443 24327
rect 8125 24225 8159 24259
rect 10793 24225 10827 24259
rect 11805 24225 11839 24259
rect 12817 24225 12851 24259
rect 13921 24225 13955 24259
rect 16037 24225 16071 24259
rect 16497 24225 16531 24259
rect 16589 24225 16623 24259
rect 17601 24225 17635 24259
rect 18061 24225 18095 24259
rect 18889 24225 18923 24259
rect 19073 24225 19107 24259
rect 21189 24225 21223 24259
rect 22477 24225 22511 24259
rect 22661 24225 22695 24259
rect 23949 24225 23983 24259
rect 25237 24225 25271 24259
rect 11621 24157 11655 24191
rect 13093 24157 13127 24191
rect 13829 24157 13863 24191
rect 15853 24157 15887 24191
rect 20913 24157 20947 24191
rect 21649 24157 21683 24191
rect 22293 24157 22327 24191
rect 23857 24157 23891 24191
rect 9965 24089 9999 24123
rect 12541 24089 12575 24123
rect 16957 24089 16991 24123
rect 20269 24089 20303 24123
rect 25697 24089 25731 24123
rect 11345 24021 11379 24055
rect 13001 24021 13035 24055
rect 13093 24021 13127 24055
rect 15117 24021 15151 24055
rect 17969 24021 18003 24055
rect 25053 24021 25087 24055
rect 25421 24021 25455 24055
rect 3617 23817 3651 23851
rect 8033 23817 8067 23851
rect 11805 23817 11839 23851
rect 13829 23817 13863 23851
rect 14473 23817 14507 23851
rect 16773 23817 16807 23851
rect 17877 23817 17911 23851
rect 19993 23817 20027 23851
rect 22569 23817 22603 23851
rect 22937 23817 22971 23851
rect 23857 23817 23891 23851
rect 24225 23817 24259 23851
rect 26341 23817 26375 23851
rect 12265 23749 12299 23783
rect 16037 23749 16071 23783
rect 2053 23681 2087 23715
rect 10057 23681 10091 23715
rect 12449 23681 12483 23715
rect 14841 23681 14875 23715
rect 16497 23681 16531 23715
rect 20729 23681 20763 23715
rect 24685 23681 24719 23715
rect 2329 23613 2363 23647
rect 9781 23613 9815 23647
rect 12725 23613 12759 23647
rect 14933 23613 14967 23647
rect 15577 23613 15611 23647
rect 16589 23613 16623 23647
rect 18521 23613 18555 23647
rect 18705 23613 18739 23647
rect 19165 23613 19199 23647
rect 19441 23613 19475 23647
rect 20821 23613 20855 23647
rect 21281 23613 21315 23647
rect 21557 23613 21591 23647
rect 21741 23613 21775 23647
rect 23489 23613 23523 23647
rect 23673 23613 23707 23647
rect 24777 23613 24811 23647
rect 25053 23613 25087 23647
rect 9321 23545 9355 23579
rect 17509 23545 17543 23579
rect 20453 23545 20487 23579
rect 1869 23477 1903 23511
rect 9689 23477 9723 23511
rect 11161 23477 11195 23511
rect 16405 23477 16439 23511
rect 19441 23477 19475 23511
rect 2053 23273 2087 23307
rect 12817 23273 12851 23307
rect 15025 23273 15059 23307
rect 16589 23273 16623 23307
rect 18337 23273 18371 23307
rect 22293 23273 22327 23307
rect 23673 23273 23707 23307
rect 25605 23273 25639 23307
rect 18797 23205 18831 23239
rect 21281 23205 21315 23239
rect 21649 23205 21683 23239
rect 21833 23205 21867 23239
rect 11161 23137 11195 23171
rect 11483 23137 11517 23171
rect 11621 23137 11655 23171
rect 13829 23137 13863 23171
rect 14197 23137 14231 23171
rect 15485 23137 15519 23171
rect 17233 23137 17267 23171
rect 17601 23137 17635 23171
rect 19441 23137 19475 23171
rect 19809 23137 19843 23171
rect 19901 23137 19935 23171
rect 21097 23137 21131 23171
rect 21189 23137 21223 23171
rect 10609 23069 10643 23103
rect 11253 23069 11287 23103
rect 13277 23069 13311 23103
rect 13921 23069 13955 23103
rect 14105 23069 14139 23103
rect 15393 23069 15427 23103
rect 17693 23069 17727 23103
rect 19349 23069 19383 23103
rect 20913 23069 20947 23103
rect 17049 23001 17083 23035
rect 22477 23137 22511 23171
rect 23489 23137 23523 23171
rect 23949 23137 23983 23171
rect 24685 23137 24719 23171
rect 22661 23001 22695 23035
rect 23029 23001 23063 23035
rect 24501 23001 24535 23035
rect 1593 22933 1627 22967
rect 12081 22933 12115 22967
rect 12541 22933 12575 22967
rect 14657 22933 14691 22967
rect 15669 22933 15703 22967
rect 18613 22933 18647 22967
rect 20637 22933 20671 22967
rect 21833 22933 21867 22967
rect 21925 22933 21959 22967
rect 23305 22933 23339 22967
rect 25237 22933 25271 22967
rect 3157 22729 3191 22763
rect 10241 22729 10275 22763
rect 11805 22729 11839 22763
rect 12633 22729 12667 22763
rect 13277 22729 13311 22763
rect 15577 22729 15611 22763
rect 16037 22729 16071 22763
rect 19165 22729 19199 22763
rect 21465 22729 21499 22763
rect 22753 22729 22787 22763
rect 23857 22729 23891 22763
rect 24593 22729 24627 22763
rect 10609 22661 10643 22695
rect 10977 22661 11011 22695
rect 11345 22661 11379 22695
rect 16497 22661 16531 22695
rect 19625 22661 19659 22695
rect 15025 22593 15059 22627
rect 16589 22593 16623 22627
rect 17509 22593 17543 22627
rect 18889 22593 18923 22627
rect 20453 22593 20487 22627
rect 22385 22593 22419 22627
rect 1593 22525 1627 22559
rect 1869 22525 1903 22559
rect 12449 22525 12483 22559
rect 13645 22525 13679 22559
rect 13921 22525 13955 22559
rect 16681 22525 16715 22559
rect 18429 22525 18463 22559
rect 19993 22525 20027 22559
rect 20545 22525 20579 22559
rect 21741 22525 21775 22559
rect 23121 22525 23155 22559
rect 12265 22457 12299 22491
rect 17141 22457 17175 22491
rect 18153 22457 18187 22491
rect 18337 22457 18371 22491
rect 18521 22457 18555 22491
rect 21097 22457 21131 22491
rect 17877 22389 17911 22423
rect 19993 22389 20027 22423
rect 13277 22185 13311 22219
rect 14381 22185 14415 22219
rect 18245 22185 18279 22219
rect 20177 22185 20211 22219
rect 21741 22185 21775 22219
rect 15117 22117 15151 22151
rect 16589 22117 16623 22151
rect 17969 22117 18003 22151
rect 19809 22117 19843 22151
rect 12265 22049 12299 22083
rect 12633 22049 12667 22083
rect 13645 22049 13679 22083
rect 14197 22049 14231 22083
rect 14749 22049 14783 22083
rect 16037 22049 16071 22083
rect 16129 22049 16163 22083
rect 17509 22049 17543 22083
rect 18705 22049 18739 22083
rect 18889 22049 18923 22083
rect 21005 22049 21039 22083
rect 22109 22049 22143 22083
rect 11621 21981 11655 22015
rect 12357 21981 12391 22015
rect 12541 21981 12575 22015
rect 15945 21981 15979 22015
rect 17417 21981 17451 22015
rect 18797 21981 18831 22015
rect 20913 21981 20947 22015
rect 23121 21981 23155 22015
rect 23397 21981 23431 22015
rect 16957 21913 16991 21947
rect 1685 21845 1719 21879
rect 14013 21845 14047 21879
rect 15577 21845 15611 21879
rect 17325 21845 17359 21879
rect 19073 21845 19107 21879
rect 20453 21845 20487 21879
rect 21189 21845 21223 21879
rect 22477 21845 22511 21879
rect 24501 21845 24535 21879
rect 11345 21641 11379 21675
rect 11713 21641 11747 21675
rect 13645 21641 13679 21675
rect 14197 21641 14231 21675
rect 15761 21641 15795 21675
rect 16129 21641 16163 21675
rect 17509 21641 17543 21675
rect 19165 21641 19199 21675
rect 21373 21641 21407 21675
rect 21833 21641 21867 21675
rect 23213 21641 23247 21675
rect 26433 21641 26467 21675
rect 11989 21573 12023 21607
rect 16589 21505 16623 21539
rect 17141 21505 17175 21539
rect 18153 21505 18187 21539
rect 19625 21505 19659 21539
rect 21005 21505 21039 21539
rect 16497 21437 16531 21471
rect 16681 21437 16715 21471
rect 17877 21437 17911 21471
rect 18797 21437 18831 21471
rect 19717 21437 19751 21471
rect 19901 21437 19935 21471
rect 20361 21437 20395 21471
rect 20453 21437 20487 21471
rect 24869 21437 24903 21471
rect 25145 21437 25179 21471
rect 10977 21369 11011 21403
rect 23949 21369 23983 21403
rect 22201 21301 22235 21335
rect 24685 21301 24719 21335
rect 13093 21097 13127 21131
rect 16405 21097 16439 21131
rect 16865 21097 16899 21131
rect 18061 21097 18095 21131
rect 18521 21097 18555 21131
rect 20269 21097 20303 21131
rect 21097 21097 21131 21131
rect 21373 21097 21407 21131
rect 11713 20961 11747 20995
rect 17693 20961 17727 20995
rect 18797 20961 18831 20995
rect 18889 20961 18923 20995
rect 19349 20961 19383 20995
rect 19533 20961 19567 20995
rect 20637 20961 20671 20995
rect 20913 20961 20947 20995
rect 11989 20893 12023 20927
rect 17785 20893 17819 20927
rect 19901 20893 19935 20927
rect 24961 20757 24995 20791
rect 12081 20553 12115 20587
rect 13553 20553 13587 20587
rect 15577 20553 15611 20587
rect 17509 20553 17543 20587
rect 17877 20553 17911 20587
rect 19073 20553 19107 20587
rect 19441 20553 19475 20587
rect 13921 20485 13955 20519
rect 21557 20485 21591 20519
rect 15853 20417 15887 20451
rect 16405 20417 16439 20451
rect 18061 20417 18095 20451
rect 11805 20349 11839 20383
rect 13369 20349 13403 20383
rect 15393 20349 15427 20383
rect 16313 20349 16347 20383
rect 16957 20349 16991 20383
rect 18153 20349 18187 20383
rect 20177 20349 20211 20383
rect 20637 20349 20671 20383
rect 21005 20349 21039 20383
rect 21373 20349 21407 20383
rect 19993 20213 20027 20247
rect 12449 20009 12483 20043
rect 13921 20009 13955 20043
rect 19165 20009 19199 20043
rect 19441 20009 19475 20043
rect 20269 20009 20303 20043
rect 20545 20009 20579 20043
rect 21373 20009 21407 20043
rect 6101 19941 6135 19975
rect 18705 19941 18739 19975
rect 4445 19873 4479 19907
rect 13737 19873 13771 19907
rect 16037 19873 16071 19907
rect 17601 19873 17635 19907
rect 18153 19873 18187 19907
rect 18337 19873 18371 19907
rect 20913 19873 20947 19907
rect 4721 19805 4755 19839
rect 15945 19805 15979 19839
rect 16773 19805 16807 19839
rect 17417 19805 17451 19839
rect 21097 19737 21131 19771
rect 14933 19669 14967 19703
rect 16221 19669 16255 19703
rect 17233 19669 17267 19703
rect 16037 19465 16071 19499
rect 20085 19465 20119 19499
rect 21005 19465 21039 19499
rect 31493 19465 31527 19499
rect 12449 19329 12483 19363
rect 12725 19329 12759 19363
rect 14933 19329 14967 19363
rect 12265 19261 12299 19295
rect 14749 19261 14783 19295
rect 15025 19261 15059 19295
rect 16589 19261 16623 19295
rect 17877 19261 17911 19295
rect 18797 19261 18831 19295
rect 19027 19261 19061 19295
rect 19165 19261 19199 19295
rect 19533 19261 19567 19295
rect 19625 19261 19659 19295
rect 30113 19261 30147 19295
rect 30389 19261 30423 19295
rect 14473 19193 14507 19227
rect 15485 19193 15519 19227
rect 17141 19193 17175 19227
rect 30021 19193 30055 19227
rect 4445 19125 4479 19159
rect 4905 19125 4939 19159
rect 13829 19125 13863 19159
rect 17417 19125 17451 19159
rect 18245 19125 18279 19159
rect 20545 19125 20579 19159
rect 14197 18921 14231 18955
rect 15025 18921 15059 18955
rect 16773 18921 16807 18955
rect 17785 18921 17819 18955
rect 18429 18921 18463 18955
rect 23857 18921 23891 18955
rect 19625 18853 19659 18887
rect 11805 18785 11839 18819
rect 12541 18785 12575 18819
rect 12909 18785 12943 18819
rect 14013 18785 14047 18819
rect 15945 18785 15979 18819
rect 16313 18785 16347 18819
rect 17325 18785 17359 18819
rect 18521 18785 18555 18819
rect 18889 18785 18923 18819
rect 19441 18785 19475 18819
rect 22753 18785 22787 18819
rect 11897 18717 11931 18751
rect 12633 18717 12667 18751
rect 12817 18717 12851 18751
rect 13461 18717 13495 18751
rect 16405 18717 16439 18751
rect 22477 18717 22511 18751
rect 15761 18649 15795 18683
rect 13737 18581 13771 18615
rect 17509 18581 17543 18615
rect 30113 18581 30147 18615
rect 11989 18377 12023 18411
rect 14473 18377 14507 18411
rect 14749 18377 14783 18411
rect 16957 18377 16991 18411
rect 17325 18377 17359 18411
rect 18521 18377 18555 18411
rect 18981 18377 19015 18411
rect 22569 18377 22603 18411
rect 16313 18309 16347 18343
rect 9873 18241 9907 18275
rect 12449 18241 12483 18275
rect 12725 18241 12759 18275
rect 10149 18173 10183 18207
rect 11529 18173 11563 18207
rect 15393 18173 15427 18207
rect 15577 18173 15611 18207
rect 15761 18173 15795 18207
rect 18797 18173 18831 18207
rect 14933 18105 14967 18139
rect 16589 18105 16623 18139
rect 9689 18037 9723 18071
rect 13829 18037 13863 18071
rect 17877 18037 17911 18071
rect 22845 18037 22879 18071
rect 9873 17833 9907 17867
rect 11529 17833 11563 17867
rect 14933 17833 14967 17867
rect 18521 17833 18555 17867
rect 18981 17833 19015 17867
rect 11897 17765 11931 17799
rect 19073 17765 19107 17799
rect 12633 17697 12667 17731
rect 13001 17697 13035 17731
rect 15393 17697 15427 17731
rect 17049 17697 17083 17731
rect 17601 17697 17635 17731
rect 17785 17697 17819 17731
rect 19717 17697 19751 17731
rect 11989 17629 12023 17663
rect 12725 17629 12759 17663
rect 12909 17629 12943 17663
rect 15301 17629 15335 17663
rect 16957 17629 16991 17663
rect 13461 17493 13495 17527
rect 15577 17493 15611 17527
rect 16221 17493 16255 17527
rect 18061 17493 18095 17527
rect 8401 17289 8435 17323
rect 11713 17289 11747 17323
rect 12725 17289 12759 17323
rect 14473 17289 14507 17323
rect 14933 17289 14967 17323
rect 18245 17289 18279 17323
rect 18613 17289 18647 17323
rect 19165 17289 19199 17323
rect 12081 17221 12115 17255
rect 17417 17221 17451 17255
rect 12909 17153 12943 17187
rect 13185 17153 13219 17187
rect 15301 17153 15335 17187
rect 15669 17153 15703 17187
rect 17785 17153 17819 17187
rect 8585 17085 8619 17119
rect 15761 17085 15795 17119
rect 15945 17085 15979 17119
rect 16405 17085 16439 17119
rect 16497 17085 16531 17119
rect 17049 17017 17083 17051
rect 8953 16949 8987 16983
rect 1593 16745 1627 16779
rect 12081 16745 12115 16779
rect 15853 16745 15887 16779
rect 25329 16677 25363 16711
rect 13001 16609 13035 16643
rect 13829 16609 13863 16643
rect 14013 16609 14047 16643
rect 14197 16609 14231 16643
rect 16221 16609 16255 16643
rect 16957 16609 16991 16643
rect 17509 16609 17543 16643
rect 17693 16609 17727 16643
rect 23673 16609 23707 16643
rect 16773 16541 16807 16575
rect 23949 16541 23983 16575
rect 13645 16473 13679 16507
rect 17969 16405 18003 16439
rect 2973 16201 3007 16235
rect 13829 16201 13863 16235
rect 14105 16201 14139 16235
rect 17233 16201 17267 16235
rect 17509 16201 17543 16235
rect 10057 16133 10091 16167
rect 13461 16133 13495 16167
rect 16865 16133 16899 16167
rect 1409 16065 1443 16099
rect 1685 16065 1719 16099
rect 10241 15997 10275 16031
rect 10517 15997 10551 16031
rect 15209 15997 15243 16031
rect 15669 15997 15703 16031
rect 16405 15929 16439 15963
rect 15393 15861 15427 15895
rect 23857 15861 23891 15895
rect 24317 15861 24351 15895
rect 18429 15657 18463 15691
rect 18061 15589 18095 15623
rect 21189 15521 21223 15555
rect 20913 15453 20947 15487
rect 1593 15317 1627 15351
rect 16037 15317 16071 15351
rect 22477 15317 22511 15351
rect 15853 15113 15887 15147
rect 18337 15113 18371 15147
rect 21005 15113 21039 15147
rect 16313 15045 16347 15079
rect 13553 14977 13587 15011
rect 13829 14977 13863 15011
rect 17785 14977 17819 15011
rect 13461 14909 13495 14943
rect 15485 14909 15519 14943
rect 16497 14909 16531 14943
rect 16681 14909 16715 14943
rect 16865 14909 16899 14943
rect 18521 14909 18555 14943
rect 18705 14909 18739 14943
rect 19073 14909 19107 14943
rect 19165 14909 19199 14943
rect 15209 14841 15243 14875
rect 17509 14841 17543 14875
rect 21281 14773 21315 14807
rect 11437 14569 11471 14603
rect 13553 14569 13587 14603
rect 18981 14569 19015 14603
rect 15853 14501 15887 14535
rect 11621 14433 11655 14467
rect 15393 14433 15427 14467
rect 17877 14433 17911 14467
rect 23305 14433 23339 14467
rect 15301 14365 15335 14399
rect 17601 14365 17635 14399
rect 23121 14229 23155 14263
rect 11529 14025 11563 14059
rect 15669 14025 15703 14059
rect 17693 14025 17727 14059
rect 18337 14025 18371 14059
rect 23213 14025 23247 14059
rect 15301 13957 15335 13991
rect 24961 13957 24995 13991
rect 25145 13821 25179 13855
rect 25421 13821 25455 13855
rect 13645 13481 13679 13515
rect 21833 13481 21867 13515
rect 16773 13345 16807 13379
rect 16957 13345 16991 13379
rect 17325 13345 17359 13379
rect 22017 13345 22051 13379
rect 16497 13277 16531 13311
rect 17233 13277 17267 13311
rect 16405 12937 16439 12971
rect 17049 12937 17083 12971
rect 21925 12937 21959 12971
rect 16037 12869 16071 12903
rect 13553 12801 13587 12835
rect 13921 12801 13955 12835
rect 16773 12801 16807 12835
rect 13645 12733 13679 12767
rect 15209 12597 15243 12631
rect 17509 12393 17543 12427
rect 13185 12325 13219 12359
rect 13645 12257 13679 12291
rect 13829 12257 13863 12291
rect 14197 12257 14231 12291
rect 14381 12257 14415 12291
rect 16129 12257 16163 12291
rect 19257 12257 19291 12291
rect 19625 12257 19659 12291
rect 16405 12189 16439 12223
rect 19073 12189 19107 12223
rect 19533 12189 19567 12223
rect 15485 12053 15519 12087
rect 18429 12053 18463 12087
rect 18889 12053 18923 12087
rect 13277 11849 13311 11883
rect 14013 11849 14047 11883
rect 14933 11849 14967 11883
rect 15393 11849 15427 11883
rect 17509 11849 17543 11883
rect 18337 11849 18371 11883
rect 21005 11849 21039 11883
rect 12909 11781 12943 11815
rect 15485 11713 15519 11747
rect 19349 11713 19383 11747
rect 15761 11645 15795 11679
rect 19441 11645 19475 11679
rect 19717 11645 19751 11679
rect 17877 11577 17911 11611
rect 13645 11509 13679 11543
rect 16865 11509 16899 11543
rect 18613 11509 18647 11543
rect 19257 11237 19291 11271
rect 16221 11169 16255 11203
rect 16589 11169 16623 11203
rect 16313 11101 16347 11135
rect 16497 11101 16531 11135
rect 17601 11101 17635 11135
rect 17877 11101 17911 11135
rect 15853 11033 15887 11067
rect 19533 11033 19567 11067
rect 15301 10761 15335 10795
rect 16313 10761 16347 10795
rect 17693 10761 17727 10795
rect 16037 10693 16071 10727
rect 18245 10693 18279 10727
rect 15669 10625 15703 10659
rect 8769 10149 8803 10183
rect 1777 10081 1811 10115
rect 7113 10081 7147 10115
rect 7389 10081 7423 10115
rect 1501 10013 1535 10047
rect 3157 10013 3191 10047
rect 2053 9673 2087 9707
rect 7481 9673 7515 9707
rect 1593 9333 1627 9367
rect 7205 9333 7239 9367
rect 35909 6273 35943 6307
rect 36277 6273 36311 6307
rect 36001 6205 36035 6239
rect 37381 6069 37415 6103
rect 36001 5661 36035 5695
rect 14013 4777 14047 4811
rect 12449 4641 12483 4675
rect 12725 4573 12759 4607
rect 12725 4233 12759 4267
rect 13001 4165 13035 4199
rect 13553 4165 13587 4199
rect 19441 4097 19475 4131
rect 21189 4097 21223 4131
rect 19533 4029 19567 4063
rect 19809 4029 19843 4063
rect 14289 3689 14323 3723
rect 12725 3553 12759 3587
rect 13001 3553 13035 3587
rect 19625 3349 19659 3383
rect 12265 3145 12299 3179
rect 14933 3145 14967 3179
rect 22293 3145 22327 3179
rect 13461 3009 13495 3043
rect 13829 3009 13863 3043
rect 20637 3009 20671 3043
rect 21005 3009 21039 3043
rect 13553 2941 13587 2975
rect 20729 2941 20763 2975
rect 12817 2805 12851 2839
rect 12449 2601 12483 2635
rect 14197 2601 14231 2635
rect 20821 2601 20855 2635
rect 28457 2601 28491 2635
rect 12909 2465 12943 2499
rect 17785 2465 17819 2499
rect 18613 2465 18647 2499
rect 24593 2465 24627 2499
rect 25973 2465 26007 2499
rect 12081 2397 12115 2431
rect 12633 2397 12667 2431
rect 18153 2397 18187 2431
rect 18889 2397 18923 2431
rect 24317 2397 24351 2431
rect 26249 2397 26283 2431
rect 26900 2397 26934 2431
rect 27169 2397 27203 2431
rect 23765 2329 23799 2363
rect 19993 2261 20027 2295
rect 23489 2261 23523 2295
rect 26709 2261 26743 2295
<< metal1 >>
rect 21174 77868 21180 77920
rect 21232 77908 21238 77920
rect 24302 77908 24308 77920
rect 21232 77880 24308 77908
rect 21232 77868 21238 77880
rect 24302 77868 24308 77880
rect 24360 77868 24366 77920
rect 1104 77818 38824 77840
rect 1104 77766 19606 77818
rect 19658 77766 19670 77818
rect 19722 77766 19734 77818
rect 19786 77766 19798 77818
rect 19850 77766 38824 77818
rect 1104 77744 38824 77766
rect 3970 77664 3976 77716
rect 4028 77704 4034 77716
rect 33502 77704 33508 77716
rect 4028 77676 33508 77704
rect 4028 77664 4034 77676
rect 33502 77664 33508 77676
rect 33560 77664 33566 77716
rect 4062 77528 4068 77580
rect 4120 77568 4126 77580
rect 24302 77568 24308 77580
rect 4120 77540 24164 77568
rect 24263 77540 24308 77568
rect 4120 77528 4126 77540
rect 24029 77503 24087 77509
rect 24029 77469 24041 77503
rect 24075 77469 24087 77503
rect 24136 77500 24164 77540
rect 24302 77528 24308 77540
rect 24360 77528 24366 77580
rect 29086 77500 29092 77512
rect 24136 77472 29092 77500
rect 24029 77463 24087 77469
rect 18046 77364 18052 77376
rect 18007 77336 18052 77364
rect 18046 77324 18052 77336
rect 18104 77324 18110 77376
rect 24044 77364 24072 77463
rect 29086 77460 29092 77472
rect 29144 77460 29150 77512
rect 35342 77432 35348 77444
rect 28920 77404 35348 77432
rect 28920 77376 28948 77404
rect 35342 77392 35348 77404
rect 35400 77392 35406 77444
rect 24670 77364 24676 77376
rect 24044 77336 24676 77364
rect 24670 77324 24676 77336
rect 24728 77324 24734 77376
rect 25593 77367 25651 77373
rect 25593 77333 25605 77367
rect 25639 77364 25651 77367
rect 28074 77364 28080 77376
rect 25639 77336 28080 77364
rect 25639 77333 25651 77336
rect 25593 77327 25651 77333
rect 28074 77324 28080 77336
rect 28132 77324 28138 77376
rect 28902 77324 28908 77376
rect 28960 77324 28966 77376
rect 29454 77364 29460 77376
rect 29415 77336 29460 77364
rect 29454 77324 29460 77336
rect 29512 77324 29518 77376
rect 1104 77274 38824 77296
rect 1104 77222 4246 77274
rect 4298 77222 4310 77274
rect 4362 77222 4374 77274
rect 4426 77222 4438 77274
rect 4490 77222 34966 77274
rect 35018 77222 35030 77274
rect 35082 77222 35094 77274
rect 35146 77222 35158 77274
rect 35210 77222 38824 77274
rect 1104 77200 38824 77222
rect 22649 77163 22707 77169
rect 22649 77129 22661 77163
rect 22695 77160 22707 77163
rect 24210 77160 24216 77172
rect 22695 77132 24216 77160
rect 22695 77129 22707 77132
rect 22649 77123 22707 77129
rect 24210 77120 24216 77132
rect 24268 77120 24274 77172
rect 24394 77160 24400 77172
rect 24355 77132 24400 77160
rect 24394 77120 24400 77132
rect 24452 77120 24458 77172
rect 29086 77160 29092 77172
rect 29047 77132 29092 77160
rect 29086 77120 29092 77132
rect 29144 77120 29150 77172
rect 31021 77163 31079 77169
rect 31021 77129 31033 77163
rect 31067 77160 31079 77163
rect 32214 77160 32220 77172
rect 31067 77132 32220 77160
rect 31067 77129 31079 77132
rect 31021 77123 31079 77129
rect 32214 77120 32220 77132
rect 32272 77120 32278 77172
rect 24121 77095 24179 77101
rect 24121 77061 24133 77095
rect 24167 77092 24179 77095
rect 24302 77092 24308 77104
rect 24167 77064 24308 77092
rect 24167 77061 24179 77064
rect 24121 77055 24179 77061
rect 24302 77052 24308 77064
rect 24360 77052 24366 77104
rect 15381 77027 15439 77033
rect 15381 76993 15393 77027
rect 15427 77024 15439 77027
rect 15749 77027 15807 77033
rect 15749 77024 15761 77027
rect 15427 76996 15761 77024
rect 15427 76993 15439 76996
rect 15381 76987 15439 76993
rect 15749 76993 15761 76996
rect 15795 77024 15807 77027
rect 16114 77024 16120 77036
rect 15795 76996 16120 77024
rect 15795 76993 15807 76996
rect 15749 76987 15807 76993
rect 16114 76984 16120 76996
rect 16172 76984 16178 77036
rect 17865 77027 17923 77033
rect 17865 76993 17877 77027
rect 17911 77024 17923 77027
rect 18325 77027 18383 77033
rect 18325 77024 18337 77027
rect 17911 76996 18337 77024
rect 17911 76993 17923 76996
rect 17865 76987 17923 76993
rect 18325 76993 18337 76996
rect 18371 77024 18383 77027
rect 18414 77024 18420 77036
rect 18371 76996 18420 77024
rect 18371 76993 18383 76996
rect 18325 76987 18383 76993
rect 18414 76984 18420 76996
rect 18472 76984 18478 77036
rect 24412 77024 24440 77120
rect 24857 77027 24915 77033
rect 24857 77024 24869 77027
rect 24412 76996 24869 77024
rect 24857 76993 24869 76996
rect 24903 76993 24915 77027
rect 29104 77024 29132 77120
rect 29733 77027 29791 77033
rect 29733 77024 29745 77027
rect 29104 76996 29745 77024
rect 24857 76987 24915 76993
rect 29733 76993 29745 76996
rect 29779 76993 29791 77027
rect 29733 76987 29791 76993
rect 15470 76956 15476 76968
rect 15431 76928 15476 76956
rect 15470 76916 15476 76928
rect 15528 76916 15534 76968
rect 17586 76916 17592 76968
rect 17644 76956 17650 76968
rect 18046 76956 18052 76968
rect 17644 76928 18052 76956
rect 17644 76916 17650 76928
rect 18046 76916 18052 76928
rect 18104 76916 18110 76968
rect 21082 76956 21088 76968
rect 21043 76928 21088 76956
rect 21082 76916 21088 76928
rect 21140 76916 21146 76968
rect 21361 76959 21419 76965
rect 21361 76956 21373 76959
rect 21192 76928 21373 76956
rect 17129 76891 17187 76897
rect 17129 76857 17141 76891
rect 17175 76888 17187 76891
rect 17678 76888 17684 76900
rect 17175 76860 17684 76888
rect 17175 76857 17187 76860
rect 17129 76851 17187 76857
rect 17678 76848 17684 76860
rect 17736 76848 17742 76900
rect 19334 76780 19340 76832
rect 19392 76820 19398 76832
rect 19429 76823 19487 76829
rect 19429 76820 19441 76823
rect 19392 76792 19441 76820
rect 19392 76780 19398 76792
rect 19429 76789 19441 76792
rect 19475 76789 19487 76823
rect 20898 76820 20904 76832
rect 20859 76792 20904 76820
rect 19429 76783 19487 76789
rect 20898 76780 20904 76792
rect 20956 76820 20962 76832
rect 21192 76820 21220 76928
rect 21361 76925 21373 76928
rect 21407 76925 21419 76959
rect 21361 76919 21419 76925
rect 24581 76959 24639 76965
rect 24581 76925 24593 76959
rect 24627 76956 24639 76959
rect 24670 76956 24676 76968
rect 24627 76928 24676 76956
rect 24627 76925 24639 76928
rect 24581 76919 24639 76925
rect 24670 76916 24676 76928
rect 24728 76916 24734 76968
rect 28810 76916 28816 76968
rect 28868 76956 28874 76968
rect 29454 76956 29460 76968
rect 28868 76928 29460 76956
rect 28868 76916 28874 76928
rect 29454 76916 29460 76928
rect 29512 76916 29518 76968
rect 20956 76792 21220 76820
rect 26145 76823 26203 76829
rect 20956 76780 20962 76792
rect 26145 76789 26157 76823
rect 26191 76820 26203 76823
rect 26970 76820 26976 76832
rect 26191 76792 26976 76820
rect 26191 76789 26203 76792
rect 26145 76783 26203 76789
rect 26970 76780 26976 76792
rect 27028 76780 27034 76832
rect 1104 76730 38824 76752
rect 1104 76678 19606 76730
rect 19658 76678 19670 76730
rect 19722 76678 19734 76730
rect 19786 76678 19798 76730
rect 19850 76678 38824 76730
rect 1104 76656 38824 76678
rect 21545 76483 21603 76489
rect 21545 76449 21557 76483
rect 21591 76480 21603 76483
rect 21910 76480 21916 76492
rect 21591 76452 21916 76480
rect 21591 76449 21603 76452
rect 21545 76443 21603 76449
rect 21910 76440 21916 76452
rect 21968 76440 21974 76492
rect 15470 76372 15476 76424
rect 15528 76412 15534 76424
rect 15565 76415 15623 76421
rect 15565 76412 15577 76415
rect 15528 76384 15577 76412
rect 15528 76372 15534 76384
rect 15565 76381 15577 76384
rect 15611 76412 15623 76415
rect 17586 76412 17592 76424
rect 15611 76384 17592 76412
rect 15611 76381 15623 76384
rect 15565 76375 15623 76381
rect 17586 76372 17592 76384
rect 17644 76372 17650 76424
rect 17770 76372 17776 76424
rect 17828 76412 17834 76424
rect 17865 76415 17923 76421
rect 17865 76412 17877 76415
rect 17828 76384 17877 76412
rect 17828 76372 17834 76384
rect 17865 76381 17877 76384
rect 17911 76381 17923 76415
rect 17865 76375 17923 76381
rect 21821 76415 21879 76421
rect 21821 76381 21833 76415
rect 21867 76412 21879 76415
rect 22002 76412 22008 76424
rect 21867 76384 22008 76412
rect 21867 76381 21879 76384
rect 21821 76375 21879 76381
rect 22002 76372 22008 76384
rect 22060 76372 22066 76424
rect 28810 76412 28816 76424
rect 28771 76384 28816 76412
rect 28810 76372 28816 76384
rect 28868 76372 28874 76424
rect 28994 76372 29000 76424
rect 29052 76412 29058 76424
rect 29089 76415 29147 76421
rect 29089 76412 29101 76415
rect 29052 76384 29101 76412
rect 29052 76372 29058 76384
rect 29089 76381 29101 76384
rect 29135 76381 29147 76415
rect 29089 76375 29147 76381
rect 20530 76304 20536 76356
rect 20588 76344 20594 76356
rect 21174 76344 21180 76356
rect 20588 76316 21180 76344
rect 20588 76304 20594 76316
rect 21174 76304 21180 76316
rect 21232 76304 21238 76356
rect 17862 76236 17868 76288
rect 17920 76276 17926 76288
rect 18969 76279 19027 76285
rect 18969 76276 18981 76279
rect 17920 76248 18981 76276
rect 17920 76236 17926 76248
rect 18969 76245 18981 76248
rect 19015 76245 19027 76279
rect 22922 76276 22928 76288
rect 22883 76248 22928 76276
rect 18969 76239 19027 76245
rect 22922 76236 22928 76248
rect 22980 76236 22986 76288
rect 24118 76276 24124 76288
rect 24031 76248 24124 76276
rect 24118 76236 24124 76248
rect 24176 76276 24182 76288
rect 24670 76276 24676 76288
rect 24176 76248 24676 76276
rect 24176 76236 24182 76248
rect 24670 76236 24676 76248
rect 24728 76236 24734 76288
rect 30374 76276 30380 76288
rect 30335 76248 30380 76276
rect 30374 76236 30380 76248
rect 30432 76236 30438 76288
rect 1104 76186 38824 76208
rect 1104 76134 4246 76186
rect 4298 76134 4310 76186
rect 4362 76134 4374 76186
rect 4426 76134 4438 76186
rect 4490 76134 34966 76186
rect 35018 76134 35030 76186
rect 35082 76134 35094 76186
rect 35146 76134 35158 76186
rect 35210 76134 38824 76186
rect 1104 76112 38824 76134
rect 21637 76075 21695 76081
rect 21637 76041 21649 76075
rect 21683 76072 21695 76075
rect 22002 76072 22008 76084
rect 21683 76044 22008 76072
rect 21683 76041 21695 76044
rect 21637 76035 21695 76041
rect 22002 76032 22008 76044
rect 22060 76032 22066 76084
rect 28905 76075 28963 76081
rect 28905 76041 28917 76075
rect 28951 76072 28963 76075
rect 28994 76072 29000 76084
rect 28951 76044 29000 76072
rect 28951 76041 28963 76044
rect 28905 76035 28963 76041
rect 28994 76032 29000 76044
rect 29052 76032 29058 76084
rect 17862 76004 17868 76016
rect 17512 75976 17868 76004
rect 17512 75948 17540 75976
rect 17862 75964 17868 75976
rect 17920 75964 17926 76016
rect 28810 75964 28816 76016
rect 28868 76004 28874 76016
rect 29457 76007 29515 76013
rect 29457 76004 29469 76007
rect 28868 75976 29469 76004
rect 28868 75964 28874 75976
rect 29457 75973 29469 75976
rect 29503 75973 29515 76007
rect 29457 75967 29515 75973
rect 17494 75896 17500 75948
rect 17552 75896 17558 75948
rect 17586 75896 17592 75948
rect 17644 75936 17650 75948
rect 18325 75939 18383 75945
rect 18325 75936 18337 75939
rect 17644 75908 18337 75936
rect 17644 75896 17650 75908
rect 18325 75905 18337 75908
rect 18371 75936 18383 75939
rect 18877 75939 18935 75945
rect 18877 75936 18889 75939
rect 18371 75908 18889 75936
rect 18371 75905 18383 75908
rect 18325 75899 18383 75905
rect 18877 75905 18889 75908
rect 18923 75936 18935 75939
rect 19242 75936 19248 75948
rect 18923 75908 19248 75936
rect 18923 75905 18935 75908
rect 18877 75899 18935 75905
rect 19242 75896 19248 75908
rect 19300 75896 19306 75948
rect 19334 75896 19340 75948
rect 19392 75896 19398 75948
rect 106 75828 112 75880
rect 164 75868 170 75880
rect 934 75868 940 75880
rect 164 75840 940 75868
rect 164 75828 170 75840
rect 934 75828 940 75840
rect 992 75828 998 75880
rect 19153 75871 19211 75877
rect 19153 75868 19165 75871
rect 18984 75840 19165 75868
rect 18785 75803 18843 75809
rect 18785 75769 18797 75803
rect 18831 75800 18843 75803
rect 18984 75800 19012 75840
rect 19153 75837 19165 75840
rect 19199 75868 19211 75871
rect 19352 75868 19380 75896
rect 19199 75840 19380 75868
rect 19199 75837 19211 75840
rect 19153 75831 19211 75837
rect 25314 75828 25320 75880
rect 25372 75868 25378 75880
rect 25685 75871 25743 75877
rect 25685 75868 25697 75871
rect 25372 75840 25697 75868
rect 25372 75828 25378 75840
rect 25685 75837 25697 75840
rect 25731 75837 25743 75871
rect 25866 75868 25872 75880
rect 25827 75840 25872 75868
rect 25685 75831 25743 75837
rect 18831 75772 19012 75800
rect 25700 75800 25728 75831
rect 25866 75828 25872 75840
rect 25924 75828 25930 75880
rect 26145 75871 26203 75877
rect 26145 75868 26157 75871
rect 25976 75840 26157 75868
rect 25976 75800 26004 75840
rect 26145 75837 26157 75840
rect 26191 75837 26203 75871
rect 26145 75831 26203 75837
rect 27522 75800 27528 75812
rect 25700 75772 26004 75800
rect 27483 75772 27528 75800
rect 18831 75769 18843 75772
rect 18785 75763 18843 75769
rect 27522 75760 27528 75772
rect 27580 75760 27586 75812
rect 17681 75735 17739 75741
rect 17681 75701 17693 75735
rect 17727 75732 17739 75735
rect 17770 75732 17776 75744
rect 17727 75704 17776 75732
rect 17727 75701 17739 75704
rect 17681 75695 17739 75701
rect 17770 75692 17776 75704
rect 17828 75692 17834 75744
rect 20070 75692 20076 75744
rect 20128 75732 20134 75744
rect 20257 75735 20315 75741
rect 20257 75732 20269 75735
rect 20128 75704 20269 75732
rect 20128 75692 20134 75704
rect 20257 75701 20269 75704
rect 20303 75701 20315 75735
rect 22002 75732 22008 75744
rect 21963 75704 22008 75732
rect 20257 75695 20315 75701
rect 22002 75692 22008 75704
rect 22060 75692 22066 75744
rect 1104 75642 38824 75664
rect 1104 75590 19606 75642
rect 19658 75590 19670 75642
rect 19722 75590 19734 75642
rect 19786 75590 19798 75642
rect 19850 75590 38824 75642
rect 1104 75568 38824 75590
rect 29822 75460 29828 75472
rect 29783 75432 29828 75460
rect 29822 75420 29828 75432
rect 29880 75420 29886 75472
rect 30374 75352 30380 75404
rect 30432 75392 30438 75404
rect 30561 75395 30619 75401
rect 30561 75392 30573 75395
rect 30432 75364 30573 75392
rect 30432 75352 30438 75364
rect 30561 75361 30573 75364
rect 30607 75361 30619 75395
rect 30561 75355 30619 75361
rect 29362 75284 29368 75336
rect 29420 75324 29426 75336
rect 29733 75327 29791 75333
rect 29733 75324 29745 75327
rect 29420 75296 29745 75324
rect 29420 75284 29426 75296
rect 29733 75293 29745 75296
rect 29779 75293 29791 75327
rect 30650 75324 30656 75336
rect 30611 75296 30656 75324
rect 29733 75287 29791 75293
rect 30650 75284 30656 75296
rect 30708 75284 30714 75336
rect 18969 75191 19027 75197
rect 18969 75157 18981 75191
rect 19015 75188 19027 75191
rect 19242 75188 19248 75200
rect 19015 75160 19248 75188
rect 19015 75157 19027 75160
rect 18969 75151 19027 75157
rect 19242 75148 19248 75160
rect 19300 75148 19306 75200
rect 25958 75188 25964 75200
rect 25919 75160 25964 75188
rect 25958 75148 25964 75160
rect 26016 75148 26022 75200
rect 1104 75098 38824 75120
rect 1104 75046 4246 75098
rect 4298 75046 4310 75098
rect 4362 75046 4374 75098
rect 4426 75046 4438 75098
rect 4490 75046 34966 75098
rect 35018 75046 35030 75098
rect 35082 75046 35094 75098
rect 35146 75046 35158 75098
rect 35210 75046 38824 75098
rect 1104 75024 38824 75046
rect 30374 74984 30380 74996
rect 30335 74956 30380 74984
rect 30374 74944 30380 74956
rect 30432 74944 30438 74996
rect 19705 74851 19763 74857
rect 19705 74817 19717 74851
rect 19751 74848 19763 74851
rect 20070 74848 20076 74860
rect 19751 74820 20076 74848
rect 19751 74817 19763 74820
rect 19705 74811 19763 74817
rect 20070 74808 20076 74820
rect 20128 74808 20134 74860
rect 9674 74740 9680 74792
rect 9732 74780 9738 74792
rect 10870 74780 10876 74792
rect 9732 74752 10876 74780
rect 9732 74740 9738 74752
rect 10870 74740 10876 74752
rect 10928 74740 10934 74792
rect 15194 74740 15200 74792
rect 15252 74780 15258 74792
rect 16482 74780 16488 74792
rect 15252 74752 16488 74780
rect 15252 74740 15258 74752
rect 16482 74740 16488 74752
rect 16540 74740 16546 74792
rect 19797 74783 19855 74789
rect 19797 74749 19809 74783
rect 19843 74780 19855 74783
rect 19886 74780 19892 74792
rect 19843 74752 19892 74780
rect 19843 74749 19855 74752
rect 19797 74743 19855 74749
rect 19886 74740 19892 74752
rect 19944 74780 19950 74792
rect 20530 74780 20536 74792
rect 19944 74752 20536 74780
rect 19944 74740 19950 74752
rect 20530 74740 20536 74752
rect 20588 74740 20594 74792
rect 37366 74740 37372 74792
rect 37424 74780 37430 74792
rect 38654 74780 38660 74792
rect 37424 74752 38660 74780
rect 37424 74740 37430 74752
rect 38654 74740 38660 74752
rect 38712 74740 38718 74792
rect 2774 74604 2780 74656
rect 2832 74644 2838 74656
rect 3878 74644 3884 74656
rect 2832 74616 3884 74644
rect 2832 74604 2838 74616
rect 3878 74604 3884 74616
rect 3936 74604 3942 74656
rect 19426 74604 19432 74656
rect 19484 74644 19490 74656
rect 20070 74644 20076 74656
rect 19484 74616 20076 74644
rect 19484 74604 19490 74616
rect 20070 74604 20076 74616
rect 20128 74604 20134 74656
rect 20806 74604 20812 74656
rect 20864 74644 20870 74656
rect 21177 74647 21235 74653
rect 21177 74644 21189 74647
rect 20864 74616 21189 74644
rect 20864 74604 20870 74616
rect 21177 74613 21189 74616
rect 21223 74613 21235 74647
rect 21177 74607 21235 74613
rect 29362 74604 29368 74656
rect 29420 74644 29426 74656
rect 29641 74647 29699 74653
rect 29641 74644 29653 74647
rect 29420 74616 29653 74644
rect 29420 74604 29426 74616
rect 29641 74613 29653 74616
rect 29687 74613 29699 74647
rect 29641 74607 29699 74613
rect 30101 74647 30159 74653
rect 30101 74613 30113 74647
rect 30147 74644 30159 74647
rect 30650 74644 30656 74656
rect 30147 74616 30656 74644
rect 30147 74613 30159 74616
rect 30101 74607 30159 74613
rect 30650 74604 30656 74616
rect 30708 74604 30714 74656
rect 33134 74604 33140 74656
rect 33192 74644 33198 74656
rect 34054 74644 34060 74656
rect 33192 74616 34060 74644
rect 33192 74604 33198 74616
rect 34054 74604 34060 74616
rect 34112 74604 34118 74656
rect 1104 74554 38824 74576
rect 1104 74502 19606 74554
rect 19658 74502 19670 74554
rect 19722 74502 19734 74554
rect 19786 74502 19798 74554
rect 19850 74502 38824 74554
rect 1104 74480 38824 74502
rect 19886 74372 19892 74384
rect 19847 74344 19892 74372
rect 19886 74332 19892 74344
rect 19944 74332 19950 74384
rect 1104 74010 38824 74032
rect 1104 73958 4246 74010
rect 4298 73958 4310 74010
rect 4362 73958 4374 74010
rect 4426 73958 4438 74010
rect 4490 73958 34966 74010
rect 35018 73958 35030 74010
rect 35082 73958 35094 74010
rect 35146 73958 35158 74010
rect 35210 73958 38824 74010
rect 1104 73936 38824 73958
rect 26326 73856 26332 73908
rect 26384 73896 26390 73908
rect 27154 73896 27160 73908
rect 26384 73868 27160 73896
rect 26384 73856 26390 73868
rect 27154 73856 27160 73868
rect 27212 73856 27218 73908
rect 1104 73466 38824 73488
rect 1104 73414 19606 73466
rect 19658 73414 19670 73466
rect 19722 73414 19734 73466
rect 19786 73414 19798 73466
rect 19850 73414 38824 73466
rect 1104 73392 38824 73414
rect 19334 72972 19340 73024
rect 19392 73012 19398 73024
rect 28810 73012 28816 73024
rect 19392 72984 28816 73012
rect 19392 72972 19398 72984
rect 28810 72972 28816 72984
rect 28868 72972 28874 73024
rect 1104 72922 38824 72944
rect 1104 72870 4246 72922
rect 4298 72870 4310 72922
rect 4362 72870 4374 72922
rect 4426 72870 4438 72922
rect 4490 72870 34966 72922
rect 35018 72870 35030 72922
rect 35082 72870 35094 72922
rect 35146 72870 35158 72922
rect 35210 72870 38824 72922
rect 1104 72848 38824 72870
rect 19426 72564 19432 72616
rect 19484 72604 19490 72616
rect 19521 72607 19579 72613
rect 19521 72604 19533 72607
rect 19484 72576 19533 72604
rect 19484 72564 19490 72576
rect 19521 72573 19533 72576
rect 19567 72573 19579 72607
rect 19797 72607 19855 72613
rect 19797 72604 19809 72607
rect 19521 72567 19579 72573
rect 19628 72576 19809 72604
rect 19334 72536 19340 72548
rect 19295 72508 19340 72536
rect 19334 72496 19340 72508
rect 19392 72536 19398 72548
rect 19628 72536 19656 72576
rect 19797 72573 19809 72576
rect 19843 72573 19855 72607
rect 19797 72567 19855 72573
rect 19392 72508 19656 72536
rect 19392 72496 19398 72508
rect 21082 72468 21088 72480
rect 21043 72440 21088 72468
rect 21082 72428 21088 72440
rect 21140 72428 21146 72480
rect 1104 72378 38824 72400
rect 1104 72326 19606 72378
rect 19658 72326 19670 72378
rect 19722 72326 19734 72378
rect 19786 72326 19798 72378
rect 19850 72326 38824 72378
rect 1104 72304 38824 72326
rect 19518 71924 19524 71936
rect 19479 71896 19524 71924
rect 19518 71884 19524 71896
rect 19576 71884 19582 71936
rect 1104 71834 38824 71856
rect 1104 71782 4246 71834
rect 4298 71782 4310 71834
rect 4362 71782 4374 71834
rect 4426 71782 4438 71834
rect 4490 71782 34966 71834
rect 35018 71782 35030 71834
rect 35082 71782 35094 71834
rect 35146 71782 35158 71834
rect 35210 71782 38824 71834
rect 1104 71760 38824 71782
rect 1104 71290 38824 71312
rect 1104 71238 19606 71290
rect 19658 71238 19670 71290
rect 19722 71238 19734 71290
rect 19786 71238 19798 71290
rect 19850 71238 38824 71290
rect 1104 71216 38824 71238
rect 22094 71000 22100 71052
rect 22152 71040 22158 71052
rect 22649 71043 22707 71049
rect 22649 71040 22661 71043
rect 22152 71012 22661 71040
rect 22152 71000 22158 71012
rect 22649 71009 22661 71012
rect 22695 71040 22707 71043
rect 22738 71040 22744 71052
rect 22695 71012 22744 71040
rect 22695 71009 22707 71012
rect 22649 71003 22707 71009
rect 22738 71000 22744 71012
rect 22796 71000 22802 71052
rect 22925 71043 22983 71049
rect 22925 71009 22937 71043
rect 22971 71040 22983 71043
rect 23198 71040 23204 71052
rect 22971 71012 23204 71040
rect 22971 71009 22983 71012
rect 22925 71003 22983 71009
rect 23198 71000 23204 71012
rect 23256 71000 23262 71052
rect 24302 70972 24308 70984
rect 24263 70944 24308 70972
rect 24302 70932 24308 70944
rect 24360 70932 24366 70984
rect 1104 70746 38824 70768
rect 1104 70694 4246 70746
rect 4298 70694 4310 70746
rect 4362 70694 4374 70746
rect 4426 70694 4438 70746
rect 4490 70694 34966 70746
rect 35018 70694 35030 70746
rect 35082 70694 35094 70746
rect 35146 70694 35158 70746
rect 35210 70694 38824 70746
rect 1104 70672 38824 70694
rect 22738 70592 22744 70644
rect 22796 70632 22802 70644
rect 23017 70635 23075 70641
rect 23017 70632 23029 70635
rect 22796 70604 23029 70632
rect 22796 70592 22802 70604
rect 23017 70601 23029 70604
rect 23063 70632 23075 70635
rect 23382 70632 23388 70644
rect 23063 70604 23388 70632
rect 23063 70601 23075 70604
rect 23017 70595 23075 70601
rect 23382 70592 23388 70604
rect 23440 70592 23446 70644
rect 22741 70499 22799 70505
rect 22741 70465 22753 70499
rect 22787 70496 22799 70499
rect 23198 70496 23204 70508
rect 22787 70468 23204 70496
rect 22787 70465 22799 70468
rect 22741 70459 22799 70465
rect 23198 70456 23204 70468
rect 23256 70456 23262 70508
rect 1104 70202 38824 70224
rect 1104 70150 19606 70202
rect 19658 70150 19670 70202
rect 19722 70150 19734 70202
rect 19786 70150 19798 70202
rect 19850 70150 38824 70202
rect 1104 70128 38824 70150
rect 23474 69844 23480 69896
rect 23532 69884 23538 69896
rect 23934 69884 23940 69896
rect 23532 69856 23940 69884
rect 23532 69844 23538 69856
rect 23934 69844 23940 69856
rect 23992 69844 23998 69896
rect 24210 69884 24216 69896
rect 24171 69856 24216 69884
rect 24210 69844 24216 69856
rect 24268 69844 24274 69896
rect 24670 69708 24676 69760
rect 24728 69748 24734 69760
rect 25317 69751 25375 69757
rect 25317 69748 25329 69751
rect 24728 69720 25329 69748
rect 24728 69708 24734 69720
rect 25317 69717 25329 69720
rect 25363 69717 25375 69751
rect 25317 69711 25375 69717
rect 1104 69658 38824 69680
rect 1104 69606 4246 69658
rect 4298 69606 4310 69658
rect 4362 69606 4374 69658
rect 4426 69606 4438 69658
rect 4490 69606 34966 69658
rect 35018 69606 35030 69658
rect 35082 69606 35094 69658
rect 35146 69606 35158 69658
rect 35210 69606 38824 69658
rect 1104 69584 38824 69606
rect 23934 69504 23940 69556
rect 23992 69544 23998 69556
rect 24305 69547 24363 69553
rect 24305 69544 24317 69547
rect 23992 69516 24317 69544
rect 23992 69504 23998 69516
rect 24305 69513 24317 69516
rect 24351 69513 24363 69547
rect 25958 69544 25964 69556
rect 25919 69516 25964 69544
rect 24305 69507 24363 69513
rect 25958 69504 25964 69516
rect 26016 69504 26022 69556
rect 24029 69479 24087 69485
rect 24029 69445 24041 69479
rect 24075 69476 24087 69479
rect 24210 69476 24216 69488
rect 24075 69448 24216 69476
rect 24075 69445 24087 69448
rect 24029 69439 24087 69445
rect 24210 69436 24216 69448
rect 24268 69436 24274 69488
rect 26145 69343 26203 69349
rect 26145 69309 26157 69343
rect 26191 69340 26203 69343
rect 26191 69312 26225 69340
rect 26191 69309 26203 69312
rect 26145 69303 26203 69309
rect 25222 69232 25228 69284
rect 25280 69272 25286 69284
rect 26160 69272 26188 69303
rect 26421 69275 26479 69281
rect 26421 69272 26433 69275
rect 25280 69244 26433 69272
rect 25280 69232 25286 69244
rect 26421 69241 26433 69244
rect 26467 69241 26479 69275
rect 26421 69235 26479 69241
rect 1104 69114 38824 69136
rect 1104 69062 19606 69114
rect 19658 69062 19670 69114
rect 19722 69062 19734 69114
rect 19786 69062 19798 69114
rect 19850 69062 38824 69114
rect 1104 69040 38824 69062
rect 22830 68864 22836 68876
rect 22791 68836 22836 68864
rect 22830 68824 22836 68836
rect 22888 68824 22894 68876
rect 25222 68864 25228 68876
rect 25183 68836 25228 68864
rect 25222 68824 25228 68836
rect 25280 68824 25286 68876
rect 22554 68796 22560 68808
rect 22515 68768 22560 68796
rect 22554 68756 22560 68768
rect 22612 68796 22618 68808
rect 22738 68796 22744 68808
rect 22612 68768 22744 68796
rect 22612 68756 22618 68768
rect 22738 68756 22744 68768
rect 22796 68756 22802 68808
rect 23934 68660 23940 68672
rect 23895 68632 23940 68660
rect 23934 68620 23940 68632
rect 23992 68620 23998 68672
rect 24026 68620 24032 68672
rect 24084 68660 24090 68672
rect 25041 68663 25099 68669
rect 25041 68660 25053 68663
rect 24084 68632 25053 68660
rect 24084 68620 24090 68632
rect 25041 68629 25053 68632
rect 25087 68629 25099 68663
rect 25041 68623 25099 68629
rect 1104 68570 38824 68592
rect 1104 68518 4246 68570
rect 4298 68518 4310 68570
rect 4362 68518 4374 68570
rect 4426 68518 4438 68570
rect 4490 68518 34966 68570
rect 35018 68518 35030 68570
rect 35082 68518 35094 68570
rect 35146 68518 35158 68570
rect 35210 68518 38824 68570
rect 1104 68496 38824 68518
rect 22649 68459 22707 68465
rect 22649 68425 22661 68459
rect 22695 68456 22707 68459
rect 22830 68456 22836 68468
rect 22695 68428 22836 68456
rect 22695 68425 22707 68428
rect 22649 68419 22707 68425
rect 22830 68416 22836 68428
rect 22888 68416 22894 68468
rect 23937 68323 23995 68329
rect 23937 68289 23949 68323
rect 23983 68320 23995 68323
rect 24305 68323 24363 68329
rect 24305 68320 24317 68323
rect 23983 68292 24317 68320
rect 23983 68289 23995 68292
rect 23937 68283 23995 68289
rect 24305 68289 24317 68292
rect 24351 68320 24363 68323
rect 24670 68320 24676 68332
rect 24351 68292 24676 68320
rect 24351 68289 24363 68292
rect 24305 68283 24363 68289
rect 24670 68280 24676 68292
rect 24728 68280 24734 68332
rect 22554 68212 22560 68264
rect 22612 68252 22618 68264
rect 23017 68255 23075 68261
rect 23017 68252 23029 68255
rect 22612 68224 23029 68252
rect 22612 68212 22618 68224
rect 23017 68221 23029 68224
rect 23063 68252 23075 68255
rect 24026 68252 24032 68264
rect 23063 68224 24032 68252
rect 23063 68221 23075 68224
rect 23017 68215 23075 68221
rect 24026 68212 24032 68224
rect 24084 68212 24090 68264
rect 25685 68187 25743 68193
rect 25685 68153 25697 68187
rect 25731 68184 25743 68187
rect 25866 68184 25872 68196
rect 25731 68156 25872 68184
rect 25731 68153 25743 68156
rect 25685 68147 25743 68153
rect 25866 68144 25872 68156
rect 25924 68144 25930 68196
rect 1104 68026 38824 68048
rect 1104 67974 19606 68026
rect 19658 67974 19670 68026
rect 19722 67974 19734 68026
rect 19786 67974 19798 68026
rect 19850 67974 38824 68026
rect 1104 67952 38824 67974
rect 19334 67872 19340 67924
rect 19392 67912 19398 67924
rect 20898 67912 20904 67924
rect 19392 67884 20904 67912
rect 19392 67872 19398 67884
rect 20898 67872 20904 67884
rect 20956 67872 20962 67924
rect 13998 67600 14004 67652
rect 14056 67640 14062 67652
rect 14090 67640 14096 67652
rect 14056 67612 14096 67640
rect 14056 67600 14062 67612
rect 14090 67600 14096 67612
rect 14148 67600 14154 67652
rect 24026 67600 24032 67652
rect 24084 67640 24090 67652
rect 24121 67643 24179 67649
rect 24121 67640 24133 67643
rect 24084 67612 24133 67640
rect 24084 67600 24090 67612
rect 24121 67609 24133 67612
rect 24167 67640 24179 67643
rect 24486 67640 24492 67652
rect 24167 67612 24492 67640
rect 24167 67609 24179 67612
rect 24121 67603 24179 67609
rect 24486 67600 24492 67612
rect 24544 67600 24550 67652
rect 25133 67643 25191 67649
rect 25133 67609 25145 67643
rect 25179 67640 25191 67643
rect 25222 67640 25228 67652
rect 25179 67612 25228 67640
rect 25179 67609 25191 67612
rect 25133 67603 25191 67609
rect 25222 67600 25228 67612
rect 25280 67640 25286 67652
rect 25280 67612 26188 67640
rect 25280 67600 25286 67612
rect 26160 67572 26188 67612
rect 26418 67572 26424 67584
rect 26160 67544 26424 67572
rect 26418 67532 26424 67544
rect 26476 67532 26482 67584
rect 1104 67482 38824 67504
rect 1104 67430 4246 67482
rect 4298 67430 4310 67482
rect 4362 67430 4374 67482
rect 4426 67430 4438 67482
rect 4490 67430 34966 67482
rect 35018 67430 35030 67482
rect 35082 67430 35094 67482
rect 35146 67430 35158 67482
rect 35210 67430 38824 67482
rect 1104 67408 38824 67430
rect 26418 67368 26424 67380
rect 26379 67340 26424 67368
rect 26418 67328 26424 67340
rect 26476 67328 26482 67380
rect 26605 67167 26663 67173
rect 26605 67133 26617 67167
rect 26651 67164 26663 67167
rect 26651 67136 27016 67164
rect 26651 67133 26663 67136
rect 26605 67127 26663 67133
rect 26988 67037 27016 67136
rect 26973 67031 27031 67037
rect 26973 66997 26985 67031
rect 27019 67028 27031 67031
rect 27062 67028 27068 67040
rect 27019 67000 27068 67028
rect 27019 66997 27031 67000
rect 26973 66991 27031 66997
rect 27062 66988 27068 67000
rect 27120 66988 27126 67040
rect 1104 66938 38824 66960
rect 1104 66886 19606 66938
rect 19658 66886 19670 66938
rect 19722 66886 19734 66938
rect 19786 66886 19798 66938
rect 19850 66886 38824 66938
rect 1104 66864 38824 66886
rect 1104 66394 38824 66416
rect 1104 66342 4246 66394
rect 4298 66342 4310 66394
rect 4362 66342 4374 66394
rect 4426 66342 4438 66394
rect 4490 66342 34966 66394
rect 35018 66342 35030 66394
rect 35082 66342 35094 66394
rect 35146 66342 35158 66394
rect 35210 66342 38824 66394
rect 1104 66320 38824 66342
rect 17218 66240 17224 66292
rect 17276 66280 17282 66292
rect 17494 66280 17500 66292
rect 17276 66252 17500 66280
rect 17276 66240 17282 66252
rect 17494 66240 17500 66252
rect 17552 66240 17558 66292
rect 17218 66104 17224 66156
rect 17276 66144 17282 66156
rect 17586 66144 17592 66156
rect 17276 66116 17592 66144
rect 17276 66104 17282 66116
rect 17586 66104 17592 66116
rect 17644 66104 17650 66156
rect 1104 65850 38824 65872
rect 1104 65798 19606 65850
rect 19658 65798 19670 65850
rect 19722 65798 19734 65850
rect 19786 65798 19798 65850
rect 19850 65798 38824 65850
rect 1104 65776 38824 65798
rect 1762 65396 1768 65408
rect 1723 65368 1768 65396
rect 1762 65356 1768 65368
rect 1820 65356 1826 65408
rect 1104 65306 38824 65328
rect 1104 65254 4246 65306
rect 4298 65254 4310 65306
rect 4362 65254 4374 65306
rect 4426 65254 4438 65306
rect 4490 65254 34966 65306
rect 35018 65254 35030 65306
rect 35082 65254 35094 65306
rect 35146 65254 35158 65306
rect 35210 65254 38824 65306
rect 1104 65232 38824 65254
rect 1578 65192 1584 65204
rect 1504 65164 1584 65192
rect 1504 64988 1532 65164
rect 1578 65152 1584 65164
rect 1636 65152 1642 65204
rect 1578 65016 1584 65068
rect 1636 65056 1642 65068
rect 1762 65056 1768 65068
rect 1636 65028 1768 65056
rect 1636 65016 1642 65028
rect 1762 65016 1768 65028
rect 1820 65016 1826 65068
rect 2041 64991 2099 64997
rect 2041 64988 2053 64991
rect 1504 64960 2053 64988
rect 2041 64957 2053 64960
rect 2087 64957 2099 64991
rect 2041 64951 2099 64957
rect 3421 64923 3479 64929
rect 3421 64889 3433 64923
rect 3467 64920 3479 64923
rect 4614 64920 4620 64932
rect 3467 64892 4620 64920
rect 3467 64889 3479 64892
rect 3421 64883 3479 64889
rect 4614 64880 4620 64892
rect 4672 64880 4678 64932
rect 1104 64762 38824 64784
rect 1104 64710 19606 64762
rect 19658 64710 19670 64762
rect 19722 64710 19734 64762
rect 19786 64710 19798 64762
rect 19850 64710 38824 64762
rect 1104 64688 38824 64710
rect 1578 64308 1584 64320
rect 1539 64280 1584 64308
rect 1578 64268 1584 64280
rect 1636 64268 1642 64320
rect 1104 64218 38824 64240
rect 1104 64166 4246 64218
rect 4298 64166 4310 64218
rect 4362 64166 4374 64218
rect 4426 64166 4438 64218
rect 4490 64166 34966 64218
rect 35018 64166 35030 64218
rect 35082 64166 35094 64218
rect 35146 64166 35158 64218
rect 35210 64166 38824 64218
rect 1104 64144 38824 64166
rect 1854 63968 1860 63980
rect 1815 63940 1860 63968
rect 1854 63928 1860 63940
rect 1912 63928 1918 63980
rect 3878 63928 3884 63980
rect 3936 63968 3942 63980
rect 4249 63971 4307 63977
rect 4249 63968 4261 63971
rect 3936 63940 4261 63968
rect 3936 63928 3942 63940
rect 4249 63937 4261 63940
rect 4295 63937 4307 63971
rect 4249 63931 4307 63937
rect 1578 63900 1584 63912
rect 1491 63872 1584 63900
rect 1578 63860 1584 63872
rect 1636 63900 1642 63912
rect 2682 63900 2688 63912
rect 1636 63872 2688 63900
rect 1636 63860 1642 63872
rect 2682 63860 2688 63872
rect 2740 63860 2746 63912
rect 3973 63903 4031 63909
rect 3973 63869 3985 63903
rect 4019 63900 4031 63903
rect 4154 63900 4160 63912
rect 4019 63872 4160 63900
rect 4019 63869 4031 63872
rect 3973 63863 4031 63869
rect 4154 63860 4160 63872
rect 4212 63860 4218 63912
rect 4985 63903 5043 63909
rect 4985 63869 4997 63903
rect 5031 63869 5043 63903
rect 4985 63863 5043 63869
rect 3237 63835 3295 63841
rect 3237 63801 3249 63835
rect 3283 63832 3295 63835
rect 4246 63832 4252 63844
rect 3283 63804 4252 63832
rect 3283 63801 3295 63804
rect 3237 63795 3295 63801
rect 4246 63792 4252 63804
rect 4304 63832 4310 63844
rect 5000 63832 5028 63863
rect 5074 63860 5080 63912
rect 5132 63900 5138 63912
rect 5132 63872 5177 63900
rect 5132 63860 5138 63872
rect 4304 63804 5028 63832
rect 4304 63792 4310 63804
rect 3605 63767 3663 63773
rect 3605 63733 3617 63767
rect 3651 63764 3663 63767
rect 5074 63764 5080 63776
rect 3651 63736 5080 63764
rect 3651 63733 3663 63736
rect 3605 63727 3663 63733
rect 5074 63724 5080 63736
rect 5132 63724 5138 63776
rect 1104 63674 38824 63696
rect 1104 63622 19606 63674
rect 19658 63622 19670 63674
rect 19722 63622 19734 63674
rect 19786 63622 19798 63674
rect 19850 63622 38824 63674
rect 1104 63600 38824 63622
rect 1673 63563 1731 63569
rect 1673 63529 1685 63563
rect 1719 63560 1731 63563
rect 1854 63560 1860 63572
rect 1719 63532 1860 63560
rect 1719 63529 1731 63532
rect 1673 63523 1731 63529
rect 1854 63520 1860 63532
rect 1912 63520 1918 63572
rect 4246 63560 4252 63572
rect 4207 63532 4252 63560
rect 4246 63520 4252 63532
rect 4304 63520 4310 63572
rect 4614 63384 4620 63436
rect 4672 63424 4678 63436
rect 4985 63427 5043 63433
rect 4985 63424 4997 63427
rect 4672 63396 4997 63424
rect 4672 63384 4678 63396
rect 4985 63393 4997 63396
rect 5031 63393 5043 63427
rect 4985 63387 5043 63393
rect 13814 63384 13820 63436
rect 13872 63424 13878 63436
rect 14093 63427 14151 63433
rect 14093 63424 14105 63427
rect 13872 63396 14105 63424
rect 13872 63384 13878 63396
rect 14093 63393 14105 63396
rect 14139 63393 14151 63427
rect 14093 63387 14151 63393
rect 20346 63384 20352 63436
rect 20404 63424 20410 63436
rect 21269 63427 21327 63433
rect 21269 63424 21281 63427
rect 20404 63396 21281 63424
rect 20404 63384 20410 63396
rect 21269 63393 21281 63396
rect 21315 63393 21327 63427
rect 21269 63387 21327 63393
rect 21634 63384 21640 63436
rect 21692 63424 21698 63436
rect 21729 63427 21787 63433
rect 21729 63424 21741 63427
rect 21692 63396 21741 63424
rect 21692 63384 21698 63396
rect 21729 63393 21741 63396
rect 21775 63393 21787 63427
rect 21729 63387 21787 63393
rect 2682 63316 2688 63368
rect 2740 63356 2746 63368
rect 4709 63359 4767 63365
rect 4709 63356 4721 63359
rect 2740 63328 4721 63356
rect 2740 63316 2746 63328
rect 4709 63325 4721 63328
rect 4755 63356 4767 63359
rect 5166 63356 5172 63368
rect 4755 63328 5172 63356
rect 4755 63325 4767 63328
rect 4709 63319 4767 63325
rect 5166 63316 5172 63328
rect 5224 63316 5230 63368
rect 21082 63356 21088 63368
rect 21043 63328 21088 63356
rect 21082 63316 21088 63328
rect 21140 63316 21146 63368
rect 13909 63291 13967 63297
rect 13909 63257 13921 63291
rect 13955 63288 13967 63291
rect 13998 63288 14004 63300
rect 13955 63260 14004 63288
rect 13955 63257 13967 63260
rect 13909 63251 13967 63257
rect 13998 63248 14004 63260
rect 14056 63248 14062 63300
rect 21726 63288 21732 63300
rect 21687 63260 21732 63288
rect 21726 63248 21732 63260
rect 21784 63248 21790 63300
rect 6273 63223 6331 63229
rect 6273 63189 6285 63223
rect 6319 63220 6331 63223
rect 6914 63220 6920 63232
rect 6319 63192 6920 63220
rect 6319 63189 6331 63192
rect 6273 63183 6331 63189
rect 6914 63180 6920 63192
rect 6972 63180 6978 63232
rect 18598 63180 18604 63232
rect 18656 63220 18662 63232
rect 18693 63223 18751 63229
rect 18693 63220 18705 63223
rect 18656 63192 18705 63220
rect 18656 63180 18662 63192
rect 18693 63189 18705 63192
rect 18739 63189 18751 63223
rect 18693 63183 18751 63189
rect 18874 63180 18880 63232
rect 18932 63220 18938 63232
rect 19061 63223 19119 63229
rect 19061 63220 19073 63223
rect 18932 63192 19073 63220
rect 18932 63180 18938 63192
rect 19061 63189 19073 63192
rect 19107 63189 19119 63223
rect 19061 63183 19119 63189
rect 1104 63130 38824 63152
rect 1104 63078 4246 63130
rect 4298 63078 4310 63130
rect 4362 63078 4374 63130
rect 4426 63078 4438 63130
rect 4490 63078 34966 63130
rect 35018 63078 35030 63130
rect 35082 63078 35094 63130
rect 35146 63078 35158 63130
rect 35210 63078 38824 63130
rect 1104 63056 38824 63078
rect 4614 62976 4620 63028
rect 4672 63016 4678 63028
rect 4709 63019 4767 63025
rect 4709 63016 4721 63019
rect 4672 62988 4721 63016
rect 4672 62976 4678 62988
rect 4709 62985 4721 62988
rect 4755 62985 4767 63019
rect 20346 63016 20352 63028
rect 4709 62979 4767 62985
rect 18800 62988 20352 63016
rect 18800 62889 18828 62988
rect 20346 62976 20352 62988
rect 20404 62976 20410 63028
rect 18601 62883 18659 62889
rect 18601 62849 18613 62883
rect 18647 62880 18659 62883
rect 18785 62883 18843 62889
rect 18785 62880 18797 62883
rect 18647 62852 18797 62880
rect 18647 62849 18659 62852
rect 18601 62843 18659 62849
rect 18785 62849 18797 62852
rect 18831 62849 18843 62883
rect 18785 62843 18843 62849
rect 18874 62840 18880 62892
rect 18932 62880 18938 62892
rect 19797 62883 19855 62889
rect 18932 62852 19564 62880
rect 18932 62840 18938 62852
rect 19536 62821 19564 62852
rect 19797 62849 19809 62883
rect 19843 62880 19855 62883
rect 20070 62880 20076 62892
rect 19843 62852 20076 62880
rect 19843 62849 19855 62852
rect 19797 62843 19855 62849
rect 20070 62840 20076 62852
rect 20128 62840 20134 62892
rect 22278 62880 22284 62892
rect 22239 62852 22284 62880
rect 22278 62840 22284 62852
rect 22336 62840 22342 62892
rect 19061 62815 19119 62821
rect 19061 62781 19073 62815
rect 19107 62781 19119 62815
rect 19061 62775 19119 62781
rect 19521 62815 19579 62821
rect 19521 62781 19533 62815
rect 19567 62781 19579 62815
rect 19521 62775 19579 62781
rect 20717 62815 20775 62821
rect 20717 62781 20729 62815
rect 20763 62812 20775 62815
rect 21082 62812 21088 62824
rect 20763 62784 21088 62812
rect 20763 62781 20775 62784
rect 20717 62775 20775 62781
rect 18598 62704 18604 62756
rect 18656 62744 18662 62756
rect 19076 62744 19104 62775
rect 21082 62772 21088 62784
rect 21140 62812 21146 62824
rect 21361 62815 21419 62821
rect 21361 62812 21373 62815
rect 21140 62784 21373 62812
rect 21140 62772 21146 62784
rect 21361 62781 21373 62784
rect 21407 62812 21419 62815
rect 21450 62812 21456 62824
rect 21407 62784 21456 62812
rect 21407 62781 21419 62784
rect 21361 62775 21419 62781
rect 21450 62772 21456 62784
rect 21508 62772 21514 62824
rect 21545 62815 21603 62821
rect 21545 62781 21557 62815
rect 21591 62781 21603 62815
rect 21545 62775 21603 62781
rect 18656 62716 19104 62744
rect 18656 62704 18662 62716
rect 5166 62676 5172 62688
rect 5127 62648 5172 62676
rect 5166 62636 5172 62648
rect 5224 62636 5230 62688
rect 13814 62636 13820 62688
rect 13872 62676 13878 62688
rect 13909 62679 13967 62685
rect 13909 62676 13921 62679
rect 13872 62648 13921 62676
rect 13872 62636 13878 62648
rect 13909 62645 13921 62648
rect 13955 62645 13967 62679
rect 21560 62676 21588 62775
rect 21726 62772 21732 62824
rect 21784 62812 21790 62824
rect 22005 62815 22063 62821
rect 22005 62812 22017 62815
rect 21784 62784 22017 62812
rect 21784 62772 21790 62784
rect 22005 62781 22017 62784
rect 22051 62781 22063 62815
rect 22005 62775 22063 62781
rect 28718 62772 28724 62824
rect 28776 62812 28782 62824
rect 28902 62812 28908 62824
rect 28776 62784 28908 62812
rect 28776 62772 28782 62784
rect 28902 62772 28908 62784
rect 28960 62772 28966 62824
rect 22002 62676 22008 62688
rect 21560 62648 22008 62676
rect 13909 62639 13967 62645
rect 22002 62636 22008 62648
rect 22060 62636 22066 62688
rect 1104 62586 38824 62608
rect 1104 62534 19606 62586
rect 19658 62534 19670 62586
rect 19722 62534 19734 62586
rect 19786 62534 19798 62586
rect 19850 62534 38824 62586
rect 1104 62512 38824 62534
rect 18506 62296 18512 62348
rect 18564 62336 18570 62348
rect 18601 62339 18659 62345
rect 18601 62336 18613 62339
rect 18564 62308 18613 62336
rect 18564 62296 18570 62308
rect 18601 62305 18613 62308
rect 18647 62305 18659 62339
rect 18601 62299 18659 62305
rect 18874 62296 18880 62348
rect 18932 62336 18938 62348
rect 19061 62339 19119 62345
rect 19061 62336 19073 62339
rect 18932 62308 19073 62336
rect 18932 62296 18938 62308
rect 19061 62305 19073 62308
rect 19107 62305 19119 62339
rect 19061 62299 19119 62305
rect 26050 62296 26056 62348
rect 26108 62336 26114 62348
rect 26510 62336 26516 62348
rect 26108 62308 26516 62336
rect 26108 62296 26114 62308
rect 26510 62296 26516 62308
rect 26568 62296 26574 62348
rect 26786 62336 26792 62348
rect 26747 62308 26792 62336
rect 26786 62296 26792 62308
rect 26844 62296 26850 62348
rect 18414 62268 18420 62280
rect 18375 62240 18420 62268
rect 18414 62228 18420 62240
rect 18472 62228 18478 62280
rect 25774 62228 25780 62280
rect 25832 62268 25838 62280
rect 25958 62268 25964 62280
rect 25832 62240 25964 62268
rect 25832 62228 25838 62240
rect 25958 62228 25964 62240
rect 26016 62228 26022 62280
rect 19058 62200 19064 62212
rect 19019 62172 19064 62200
rect 19058 62160 19064 62172
rect 19116 62160 19122 62212
rect 21174 62132 21180 62144
rect 21135 62104 21180 62132
rect 21174 62092 21180 62104
rect 21232 62132 21238 62144
rect 21545 62135 21603 62141
rect 21545 62132 21557 62135
rect 21232 62104 21557 62132
rect 21232 62092 21238 62104
rect 21545 62101 21557 62104
rect 21591 62132 21603 62135
rect 21726 62132 21732 62144
rect 21591 62104 21732 62132
rect 21591 62101 21603 62104
rect 21545 62095 21603 62101
rect 21726 62092 21732 62104
rect 21784 62092 21790 62144
rect 22002 62132 22008 62144
rect 21963 62104 22008 62132
rect 22002 62092 22008 62104
rect 22060 62092 22066 62144
rect 27798 62092 27804 62144
rect 27856 62132 27862 62144
rect 27893 62135 27951 62141
rect 27893 62132 27905 62135
rect 27856 62104 27905 62132
rect 27856 62092 27862 62104
rect 27893 62101 27905 62104
rect 27939 62101 27951 62135
rect 27893 62095 27951 62101
rect 1104 62042 38824 62064
rect 1104 61990 4246 62042
rect 4298 61990 4310 62042
rect 4362 61990 4374 62042
rect 4426 61990 4438 62042
rect 4490 61990 34966 62042
rect 35018 61990 35030 62042
rect 35082 61990 35094 62042
rect 35146 61990 35158 62042
rect 35210 61990 38824 62042
rect 1104 61968 38824 61990
rect 18325 61931 18383 61937
rect 18325 61897 18337 61931
rect 18371 61928 18383 61931
rect 18414 61928 18420 61940
rect 18371 61900 18420 61928
rect 18371 61897 18383 61900
rect 18325 61891 18383 61897
rect 18414 61888 18420 61900
rect 18472 61888 18478 61940
rect 26605 61931 26663 61937
rect 26605 61897 26617 61931
rect 26651 61928 26663 61931
rect 26786 61928 26792 61940
rect 26651 61900 26792 61928
rect 26651 61897 26663 61900
rect 26605 61891 26663 61897
rect 26786 61888 26792 61900
rect 26844 61888 26850 61940
rect 26510 61820 26516 61872
rect 26568 61860 26574 61872
rect 26881 61863 26939 61869
rect 26881 61860 26893 61863
rect 26568 61832 26893 61860
rect 26568 61820 26574 61832
rect 26881 61829 26893 61832
rect 26927 61829 26939 61863
rect 26881 61823 26939 61829
rect 13357 61727 13415 61733
rect 13357 61693 13369 61727
rect 13403 61724 13415 61727
rect 13403 61696 13768 61724
rect 13403 61693 13415 61696
rect 13357 61687 13415 61693
rect 13170 61588 13176 61600
rect 13131 61560 13176 61588
rect 13170 61548 13176 61560
rect 13228 61548 13234 61600
rect 13740 61597 13768 61696
rect 13725 61591 13783 61597
rect 13725 61557 13737 61591
rect 13771 61588 13783 61591
rect 13906 61588 13912 61600
rect 13771 61560 13912 61588
rect 13771 61557 13783 61560
rect 13725 61551 13783 61557
rect 13906 61548 13912 61560
rect 13964 61548 13970 61600
rect 18506 61548 18512 61600
rect 18564 61588 18570 61600
rect 18601 61591 18659 61597
rect 18601 61588 18613 61591
rect 18564 61560 18613 61588
rect 18564 61548 18570 61560
rect 18601 61557 18613 61560
rect 18647 61557 18659 61591
rect 18601 61551 18659 61557
rect 18874 61548 18880 61600
rect 18932 61588 18938 61600
rect 18969 61591 19027 61597
rect 18969 61588 18981 61591
rect 18932 61560 18981 61588
rect 18932 61548 18938 61560
rect 18969 61557 18981 61560
rect 19015 61557 19027 61591
rect 18969 61551 19027 61557
rect 20070 61548 20076 61600
rect 20128 61588 20134 61600
rect 21085 61591 21143 61597
rect 21085 61588 21097 61591
rect 20128 61560 21097 61588
rect 20128 61548 20134 61560
rect 21085 61557 21097 61560
rect 21131 61588 21143 61591
rect 21910 61588 21916 61600
rect 21131 61560 21916 61588
rect 21131 61557 21143 61560
rect 21085 61551 21143 61557
rect 21910 61548 21916 61560
rect 21968 61548 21974 61600
rect 1104 61498 38824 61520
rect 1104 61446 19606 61498
rect 19658 61446 19670 61498
rect 19722 61446 19734 61498
rect 19786 61446 19798 61498
rect 19850 61446 38824 61498
rect 1104 61424 38824 61446
rect 19889 61387 19947 61393
rect 19889 61353 19901 61387
rect 19935 61384 19947 61387
rect 20346 61384 20352 61396
rect 19935 61356 20352 61384
rect 19935 61353 19947 61356
rect 19889 61347 19947 61353
rect 20346 61344 20352 61356
rect 20404 61344 20410 61396
rect 10962 61248 10968 61260
rect 10923 61220 10968 61248
rect 10962 61208 10968 61220
rect 11020 61208 11026 61260
rect 19334 61208 19340 61260
rect 19392 61248 19398 61260
rect 19705 61251 19763 61257
rect 19705 61248 19717 61251
rect 19392 61220 19717 61248
rect 19392 61208 19398 61220
rect 19705 61217 19717 61220
rect 19751 61217 19763 61251
rect 19705 61211 19763 61217
rect 20717 61251 20775 61257
rect 20717 61217 20729 61251
rect 20763 61248 20775 61251
rect 21637 61251 21695 61257
rect 21637 61248 21649 61251
rect 20763 61220 21649 61248
rect 20763 61217 20775 61220
rect 20717 61211 20775 61217
rect 21637 61217 21649 61220
rect 21683 61217 21695 61251
rect 21910 61248 21916 61260
rect 21871 61220 21916 61248
rect 21637 61211 21695 61217
rect 21269 61183 21327 61189
rect 21269 61149 21281 61183
rect 21315 61180 21327 61183
rect 21358 61180 21364 61192
rect 21315 61152 21364 61180
rect 21315 61149 21327 61152
rect 21269 61143 21327 61149
rect 21358 61140 21364 61152
rect 21416 61140 21422 61192
rect 21652 61180 21680 61211
rect 21910 61208 21916 61220
rect 21968 61208 21974 61260
rect 22002 61180 22008 61192
rect 21652 61152 22008 61180
rect 22002 61140 22008 61152
rect 22060 61140 22066 61192
rect 19613 61115 19671 61121
rect 19613 61081 19625 61115
rect 19659 61112 19671 61115
rect 20254 61112 20260 61124
rect 19659 61084 20260 61112
rect 19659 61081 19671 61084
rect 19613 61075 19671 61081
rect 20254 61072 20260 61084
rect 20312 61072 20318 61124
rect 20714 61072 20720 61124
rect 20772 61112 20778 61124
rect 21913 61115 21971 61121
rect 21913 61112 21925 61115
rect 20772 61084 21925 61112
rect 20772 61072 20778 61084
rect 21913 61081 21925 61084
rect 21959 61081 21971 61115
rect 21913 61075 21971 61081
rect 10778 61044 10784 61056
rect 10739 61016 10784 61044
rect 10778 61004 10784 61016
rect 10836 61004 10842 61056
rect 20070 61004 20076 61056
rect 20128 61044 20134 61056
rect 20165 61047 20223 61053
rect 20165 61044 20177 61047
rect 20128 61016 20177 61044
rect 20128 61004 20134 61016
rect 20165 61013 20177 61016
rect 20211 61013 20223 61047
rect 20165 61007 20223 61013
rect 22094 61004 22100 61056
rect 22152 61044 22158 61056
rect 22554 61044 22560 61056
rect 22152 61016 22560 61044
rect 22152 61004 22158 61016
rect 22554 61004 22560 61016
rect 22612 61004 22618 61056
rect 25317 61047 25375 61053
rect 25317 61013 25329 61047
rect 25363 61044 25375 61047
rect 26050 61044 26056 61056
rect 25363 61016 26056 61044
rect 25363 61013 25375 61016
rect 25317 61007 25375 61013
rect 26050 61004 26056 61016
rect 26108 61004 26114 61056
rect 1104 60954 38824 60976
rect 1104 60902 4246 60954
rect 4298 60902 4310 60954
rect 4362 60902 4374 60954
rect 4426 60902 4438 60954
rect 4490 60902 34966 60954
rect 35018 60902 35030 60954
rect 35082 60902 35094 60954
rect 35146 60902 35158 60954
rect 35210 60902 38824 60954
rect 1104 60880 38824 60902
rect 10873 60843 10931 60849
rect 10873 60809 10885 60843
rect 10919 60840 10931 60843
rect 10962 60840 10968 60852
rect 10919 60812 10968 60840
rect 10919 60809 10931 60812
rect 10873 60803 10931 60809
rect 10962 60800 10968 60812
rect 11020 60800 11026 60852
rect 18414 60800 18420 60852
rect 18472 60840 18478 60852
rect 18969 60843 19027 60849
rect 18969 60840 18981 60843
rect 18472 60812 18981 60840
rect 18472 60800 18478 60812
rect 18969 60809 18981 60812
rect 19015 60809 19027 60843
rect 18969 60803 19027 60809
rect 21269 60843 21327 60849
rect 21269 60809 21281 60843
rect 21315 60840 21327 60843
rect 21358 60840 21364 60852
rect 21315 60812 21364 60840
rect 21315 60809 21327 60812
rect 21269 60803 21327 60809
rect 21358 60800 21364 60812
rect 21416 60840 21422 60852
rect 23014 60840 23020 60852
rect 21416 60812 23020 60840
rect 21416 60800 21422 60812
rect 23014 60800 23020 60812
rect 23072 60800 23078 60852
rect 9398 60732 9404 60784
rect 9456 60732 9462 60784
rect 20622 60772 20628 60784
rect 20583 60744 20628 60772
rect 20622 60732 20628 60744
rect 20680 60732 20686 60784
rect 9416 60636 9444 60732
rect 20070 60664 20076 60716
rect 20128 60704 20134 60716
rect 20128 60676 20576 60704
rect 20128 60664 20134 60676
rect 20548 60648 20576 60676
rect 24302 60664 24308 60716
rect 24360 60704 24366 60716
rect 25409 60707 25467 60713
rect 25409 60704 25421 60707
rect 24360 60676 25421 60704
rect 24360 60664 24366 60676
rect 25409 60673 25421 60676
rect 25455 60673 25467 60707
rect 25409 60667 25467 60673
rect 30837 60707 30895 60713
rect 30837 60673 30849 60707
rect 30883 60704 30895 60707
rect 31202 60704 31208 60716
rect 30883 60676 31208 60704
rect 30883 60673 30895 60676
rect 30837 60667 30895 60673
rect 31202 60664 31208 60676
rect 31260 60664 31266 60716
rect 35713 60707 35771 60713
rect 35713 60673 35725 60707
rect 35759 60704 35771 60707
rect 36081 60707 36139 60713
rect 36081 60704 36093 60707
rect 35759 60676 36093 60704
rect 35759 60673 35771 60676
rect 35713 60667 35771 60673
rect 36081 60673 36093 60676
rect 36127 60704 36139 60707
rect 37458 60704 37464 60716
rect 36127 60676 37464 60704
rect 36127 60673 36139 60676
rect 36081 60667 36139 60673
rect 37458 60664 37464 60676
rect 37516 60664 37522 60716
rect 9490 60636 9496 60648
rect 9416 60608 9496 60636
rect 9490 60596 9496 60608
rect 9548 60596 9554 60648
rect 18785 60639 18843 60645
rect 18785 60605 18797 60639
rect 18831 60636 18843 60639
rect 19705 60639 19763 60645
rect 18831 60608 18865 60636
rect 18831 60605 18843 60608
rect 18785 60599 18843 60605
rect 19705 60605 19717 60639
rect 19751 60636 19763 60639
rect 19978 60636 19984 60648
rect 19751 60608 19984 60636
rect 19751 60605 19763 60608
rect 19705 60599 19763 60605
rect 18693 60571 18751 60577
rect 18693 60537 18705 60571
rect 18739 60568 18751 60571
rect 18800 60568 18828 60599
rect 19978 60596 19984 60608
rect 20036 60596 20042 60648
rect 20254 60636 20260 60648
rect 20215 60608 20260 60636
rect 20254 60596 20260 60608
rect 20312 60596 20318 60648
rect 20530 60596 20536 60648
rect 20588 60636 20594 60648
rect 20625 60639 20683 60645
rect 20625 60636 20637 60639
rect 20588 60608 20637 60636
rect 20588 60596 20594 60608
rect 20625 60605 20637 60608
rect 20671 60605 20683 60639
rect 20625 60599 20683 60605
rect 22094 60596 22100 60648
rect 22152 60636 22158 60648
rect 22281 60639 22339 60645
rect 22281 60636 22293 60639
rect 22152 60608 22293 60636
rect 22152 60596 22158 60608
rect 22281 60605 22293 60608
rect 22327 60605 22339 60639
rect 22281 60599 22339 60605
rect 19426 60568 19432 60580
rect 18739 60540 19432 60568
rect 18739 60537 18751 60540
rect 18693 60531 18751 60537
rect 19426 60528 19432 60540
rect 19484 60528 19490 60580
rect 20070 60528 20076 60580
rect 20128 60568 20134 60580
rect 21542 60568 21548 60580
rect 20128 60540 21548 60568
rect 20128 60528 20134 60540
rect 21542 60528 21548 60540
rect 21600 60568 21606 60580
rect 21729 60571 21787 60577
rect 21729 60568 21741 60571
rect 21600 60540 21741 60568
rect 21600 60528 21606 60540
rect 21729 60537 21741 60540
rect 21775 60537 21787 60571
rect 22296 60568 22324 60599
rect 22370 60596 22376 60648
rect 22428 60645 22434 60648
rect 22428 60639 22477 60645
rect 22428 60605 22431 60639
rect 22465 60605 22477 60639
rect 22554 60636 22560 60648
rect 22515 60608 22560 60636
rect 22428 60599 22477 60605
rect 22428 60596 22434 60599
rect 22554 60596 22560 60608
rect 22612 60596 22618 60648
rect 25133 60639 25191 60645
rect 25133 60605 25145 60639
rect 25179 60636 25191 60639
rect 25317 60639 25375 60645
rect 25317 60636 25329 60639
rect 25179 60608 25329 60636
rect 25179 60605 25191 60608
rect 25133 60599 25191 60605
rect 25317 60605 25329 60608
rect 25363 60605 25375 60639
rect 25317 60599 25375 60605
rect 23385 60571 23443 60577
rect 23385 60568 23397 60571
rect 22296 60540 23397 60568
rect 21729 60531 21787 60537
rect 23385 60537 23397 60540
rect 23431 60537 23443 60571
rect 25332 60568 25360 60599
rect 25498 60596 25504 60648
rect 25556 60636 25562 60648
rect 26050 60636 26056 60648
rect 25556 60608 26056 60636
rect 25556 60596 25562 60608
rect 26050 60596 26056 60608
rect 26108 60636 26114 60648
rect 26145 60639 26203 60645
rect 26145 60636 26157 60639
rect 26108 60608 26157 60636
rect 26108 60596 26114 60608
rect 26145 60605 26157 60608
rect 26191 60605 26203 60639
rect 26145 60599 26203 60605
rect 26234 60596 26240 60648
rect 26292 60636 26298 60648
rect 30926 60636 30932 60648
rect 26292 60608 26337 60636
rect 30887 60608 30932 60636
rect 26292 60596 26298 60608
rect 30926 60596 30932 60608
rect 30984 60596 30990 60648
rect 35802 60636 35808 60648
rect 35763 60608 35808 60636
rect 35802 60596 35808 60608
rect 35860 60596 35866 60648
rect 26510 60568 26516 60580
rect 25332 60540 26516 60568
rect 23385 60531 23443 60537
rect 26510 60528 26516 60540
rect 26568 60528 26574 60580
rect 19334 60500 19340 60512
rect 19295 60472 19340 60500
rect 19334 60460 19340 60472
rect 19392 60460 19398 60512
rect 21634 60500 21640 60512
rect 21595 60472 21640 60500
rect 21634 60460 21640 60472
rect 21692 60460 21698 60512
rect 22370 60460 22376 60512
rect 22428 60500 22434 60512
rect 23017 60503 23075 60509
rect 23017 60500 23029 60503
rect 22428 60472 23029 60500
rect 22428 60460 22434 60472
rect 23017 60469 23029 60472
rect 23063 60469 23075 60503
rect 32306 60500 32312 60512
rect 32267 60472 32312 60500
rect 23017 60463 23075 60469
rect 32306 60460 32312 60472
rect 32364 60460 32370 60512
rect 37366 60500 37372 60512
rect 37327 60472 37372 60500
rect 37366 60460 37372 60472
rect 37424 60460 37430 60512
rect 1104 60410 38824 60432
rect 1104 60358 19606 60410
rect 19658 60358 19670 60410
rect 19722 60358 19734 60410
rect 19786 60358 19798 60410
rect 19850 60358 38824 60410
rect 1104 60336 38824 60358
rect 20346 60296 20352 60308
rect 20307 60268 20352 60296
rect 20346 60256 20352 60268
rect 20404 60256 20410 60308
rect 21542 60256 21548 60308
rect 21600 60296 21606 60308
rect 24486 60296 24492 60308
rect 21600 60268 22968 60296
rect 24447 60268 24492 60296
rect 21600 60256 21606 60268
rect 19242 60160 19248 60172
rect 19203 60132 19248 60160
rect 19242 60120 19248 60132
rect 19300 60120 19306 60172
rect 19392 60163 19450 60169
rect 19392 60129 19404 60163
rect 19438 60160 19450 60163
rect 19702 60160 19708 60172
rect 19438 60132 19708 60160
rect 19438 60129 19450 60132
rect 19392 60123 19450 60129
rect 19702 60120 19708 60132
rect 19760 60120 19766 60172
rect 20162 60120 20168 60172
rect 20220 60160 20226 60172
rect 21744 60169 21772 60268
rect 22940 60228 22968 60268
rect 24486 60256 24492 60268
rect 24544 60256 24550 60308
rect 25314 60296 25320 60308
rect 25275 60268 25320 60296
rect 25314 60256 25320 60268
rect 25372 60256 25378 60308
rect 29546 60296 29552 60308
rect 29507 60268 29552 60296
rect 29546 60256 29552 60268
rect 29604 60256 29610 60308
rect 30466 60256 30472 60308
rect 30524 60296 30530 60308
rect 30926 60296 30932 60308
rect 30524 60268 30932 60296
rect 30524 60256 30530 60268
rect 30926 60256 30932 60268
rect 30984 60256 30990 60308
rect 23293 60231 23351 60237
rect 23293 60228 23305 60231
rect 22940 60200 23305 60228
rect 23293 60197 23305 60200
rect 23339 60197 23351 60231
rect 23293 60191 23351 60197
rect 21269 60163 21327 60169
rect 21269 60160 21281 60163
rect 20220 60132 21281 60160
rect 20220 60120 20226 60132
rect 21269 60129 21281 60132
rect 21315 60129 21327 60163
rect 21269 60123 21327 60129
rect 21729 60163 21787 60169
rect 21729 60129 21741 60163
rect 21775 60129 21787 60163
rect 22830 60160 22836 60172
rect 22791 60132 22836 60160
rect 21729 60123 21787 60129
rect 18046 60052 18052 60104
rect 18104 60092 18110 60104
rect 19153 60095 19211 60101
rect 19153 60092 19165 60095
rect 18104 60064 19165 60092
rect 18104 60052 18110 60064
rect 19153 60061 19165 60064
rect 19199 60092 19211 60095
rect 19613 60095 19671 60101
rect 19613 60092 19625 60095
rect 19199 60064 19625 60092
rect 19199 60061 19211 60064
rect 19153 60055 19211 60061
rect 19613 60061 19625 60064
rect 19659 60092 19671 60095
rect 20438 60092 20444 60104
rect 19659 60064 20444 60092
rect 19659 60061 19671 60064
rect 19613 60055 19671 60061
rect 20438 60052 20444 60064
rect 20496 60052 20502 60104
rect 20717 60095 20775 60101
rect 20717 60061 20729 60095
rect 20763 60092 20775 60095
rect 21082 60092 21088 60104
rect 20763 60064 21088 60092
rect 20763 60061 20775 60064
rect 20717 60055 20775 60061
rect 21082 60052 21088 60064
rect 21140 60052 21146 60104
rect 18325 60027 18383 60033
rect 18325 59993 18337 60027
rect 18371 60024 18383 60027
rect 20162 60024 20168 60036
rect 18371 59996 20168 60024
rect 18371 59993 18383 59996
rect 18325 59987 18383 59993
rect 20162 59984 20168 59996
rect 20220 59984 20226 60036
rect 21284 60024 21312 60123
rect 22830 60120 22836 60132
rect 22888 60120 22894 60172
rect 27249 60163 27307 60169
rect 27249 60129 27261 60163
rect 27295 60160 27307 60163
rect 27798 60160 27804 60172
rect 27295 60132 27804 60160
rect 27295 60129 27307 60132
rect 27249 60123 27307 60129
rect 27798 60120 27804 60132
rect 27856 60160 27862 60172
rect 28166 60160 28172 60172
rect 27856 60132 28172 60160
rect 27856 60120 27862 60132
rect 28166 60120 28172 60132
rect 28224 60120 28230 60172
rect 29178 60120 29184 60172
rect 29236 60160 29242 60172
rect 29733 60163 29791 60169
rect 29733 60160 29745 60163
rect 29236 60132 29745 60160
rect 29236 60120 29242 60132
rect 29733 60129 29745 60132
rect 29779 60129 29791 60163
rect 29733 60123 29791 60129
rect 21818 60092 21824 60104
rect 21779 60064 21824 60092
rect 21818 60052 21824 60064
rect 21876 60052 21882 60104
rect 26602 60092 26608 60104
rect 26563 60064 26608 60092
rect 26602 60052 26608 60064
rect 26660 60052 26666 60104
rect 22649 60027 22707 60033
rect 22649 60024 22661 60027
rect 21284 59996 22661 60024
rect 22649 59993 22661 59996
rect 22695 59993 22707 60027
rect 23014 60024 23020 60036
rect 22975 59996 23020 60024
rect 22649 59987 22707 59993
rect 23014 59984 23020 59996
rect 23072 59984 23078 60036
rect 18598 59956 18604 59968
rect 18559 59928 18604 59956
rect 18598 59916 18604 59928
rect 18656 59916 18662 59968
rect 19518 59956 19524 59968
rect 19479 59928 19524 59956
rect 19518 59916 19524 59928
rect 19576 59916 19582 59968
rect 19886 59956 19892 59968
rect 19847 59928 19892 59956
rect 19886 59916 19892 59928
rect 19944 59916 19950 59968
rect 21818 59916 21824 59968
rect 21876 59956 21882 59968
rect 22281 59959 22339 59965
rect 22281 59956 22293 59959
rect 21876 59928 22293 59956
rect 21876 59916 21882 59928
rect 22281 59925 22293 59928
rect 22327 59925 22339 59959
rect 23842 59956 23848 59968
rect 23803 59928 23848 59956
rect 22281 59919 22339 59925
rect 23842 59916 23848 59928
rect 23900 59916 23906 59968
rect 24213 59959 24271 59965
rect 24213 59925 24225 59959
rect 24259 59956 24271 59959
rect 24302 59956 24308 59968
rect 24259 59928 24308 59956
rect 24259 59925 24271 59928
rect 24213 59919 24271 59925
rect 24302 59916 24308 59928
rect 24360 59916 24366 59968
rect 29914 59916 29920 59968
rect 29972 59956 29978 59968
rect 30193 59959 30251 59965
rect 30193 59956 30205 59959
rect 29972 59928 30205 59956
rect 29972 59916 29978 59928
rect 30193 59925 30205 59928
rect 30239 59925 30251 59959
rect 30193 59919 30251 59925
rect 35250 59916 35256 59968
rect 35308 59956 35314 59968
rect 35802 59956 35808 59968
rect 35308 59928 35808 59956
rect 35308 59916 35314 59928
rect 35802 59916 35808 59928
rect 35860 59916 35866 59968
rect 1104 59866 38824 59888
rect 1104 59814 4246 59866
rect 4298 59814 4310 59866
rect 4362 59814 4374 59866
rect 4426 59814 4438 59866
rect 4490 59814 34966 59866
rect 35018 59814 35030 59866
rect 35082 59814 35094 59866
rect 35146 59814 35158 59866
rect 35210 59814 38824 59866
rect 1104 59792 38824 59814
rect 17862 59752 17868 59764
rect 17823 59724 17868 59752
rect 17862 59712 17868 59724
rect 17920 59712 17926 59764
rect 19886 59712 19892 59764
rect 19944 59752 19950 59764
rect 22830 59752 22836 59764
rect 19944 59724 22836 59752
rect 19944 59712 19950 59724
rect 22830 59712 22836 59724
rect 22888 59712 22894 59764
rect 25498 59752 25504 59764
rect 25459 59724 25504 59752
rect 25498 59712 25504 59724
rect 25556 59712 25562 59764
rect 18785 59687 18843 59693
rect 18785 59653 18797 59687
rect 18831 59684 18843 59687
rect 19978 59684 19984 59696
rect 18831 59656 19984 59684
rect 18831 59653 18843 59656
rect 18785 59647 18843 59653
rect 19978 59644 19984 59656
rect 20036 59644 20042 59696
rect 22186 59644 22192 59696
rect 22244 59684 22250 59696
rect 22281 59687 22339 59693
rect 22281 59684 22293 59687
rect 22244 59656 22293 59684
rect 22244 59644 22250 59656
rect 22281 59653 22293 59656
rect 22327 59653 22339 59687
rect 27246 59684 27252 59696
rect 27207 59656 27252 59684
rect 22281 59647 22339 59653
rect 27246 59644 27252 59656
rect 27304 59644 27310 59696
rect 19613 59619 19671 59625
rect 19613 59585 19625 59619
rect 19659 59616 19671 59619
rect 20530 59616 20536 59628
rect 19659 59588 20536 59616
rect 19659 59585 19671 59588
rect 19613 59579 19671 59585
rect 20530 59576 20536 59588
rect 20588 59576 20594 59628
rect 20622 59576 20628 59628
rect 20680 59616 20686 59628
rect 21361 59619 21419 59625
rect 20680 59588 20725 59616
rect 20680 59576 20686 59588
rect 21361 59585 21373 59619
rect 21407 59616 21419 59619
rect 21637 59619 21695 59625
rect 21637 59616 21649 59619
rect 21407 59588 21649 59616
rect 21407 59585 21419 59588
rect 21361 59579 21419 59585
rect 21637 59585 21649 59588
rect 21683 59616 21695 59619
rect 22738 59616 22744 59628
rect 21683 59588 22744 59616
rect 21683 59585 21695 59588
rect 21637 59579 21695 59585
rect 22738 59576 22744 59588
rect 22796 59576 22802 59628
rect 23937 59619 23995 59625
rect 23937 59585 23949 59619
rect 23983 59616 23995 59619
rect 24394 59616 24400 59628
rect 23983 59588 24400 59616
rect 23983 59585 23995 59588
rect 23937 59579 23995 59585
rect 24394 59576 24400 59588
rect 24452 59576 24458 59628
rect 25961 59619 26019 59625
rect 25961 59585 25973 59619
rect 26007 59616 26019 59619
rect 26602 59616 26608 59628
rect 26007 59588 26608 59616
rect 26007 59585 26019 59588
rect 25961 59579 26019 59585
rect 26602 59576 26608 59588
rect 26660 59576 26666 59628
rect 30374 59616 30380 59628
rect 30335 59588 30380 59616
rect 30374 59576 30380 59588
rect 30432 59576 30438 59628
rect 32306 59616 32312 59628
rect 31128 59588 32312 59616
rect 18598 59548 18604 59560
rect 18559 59520 18604 59548
rect 18598 59508 18604 59520
rect 18656 59508 18662 59560
rect 20162 59548 20168 59560
rect 20123 59520 20168 59548
rect 20162 59508 20168 59520
rect 20220 59508 20226 59560
rect 20346 59508 20352 59560
rect 20404 59548 20410 59560
rect 20441 59551 20499 59557
rect 20441 59548 20453 59551
rect 20404 59520 20453 59548
rect 20404 59508 20410 59520
rect 20441 59517 20453 59520
rect 20487 59517 20499 59551
rect 21818 59548 21824 59560
rect 21779 59520 21824 59548
rect 20441 59511 20499 59517
rect 21818 59508 21824 59520
rect 21876 59508 21882 59560
rect 22370 59548 22376 59560
rect 22283 59520 22376 59548
rect 22370 59508 22376 59520
rect 22428 59548 22434 59560
rect 24210 59548 24216 59560
rect 22428 59520 23336 59548
rect 24171 59520 24216 59548
rect 22428 59508 22434 59520
rect 19518 59480 19524 59492
rect 18432 59452 19524 59480
rect 18138 59372 18144 59424
rect 18196 59412 18202 59424
rect 18432 59421 18460 59452
rect 19518 59440 19524 59452
rect 19576 59440 19582 59492
rect 19702 59440 19708 59492
rect 19760 59440 19766 59492
rect 18417 59415 18475 59421
rect 18417 59412 18429 59415
rect 18196 59384 18429 59412
rect 18196 59372 18202 59384
rect 18417 59381 18429 59384
rect 18463 59381 18475 59415
rect 18417 59375 18475 59381
rect 19337 59415 19395 59421
rect 19337 59381 19349 59415
rect 19383 59412 19395 59415
rect 19720 59412 19748 59440
rect 23308 59424 23336 59520
rect 24210 59508 24216 59520
rect 24268 59508 24274 59560
rect 26329 59551 26387 59557
rect 26329 59517 26341 59551
rect 26375 59548 26387 59551
rect 26786 59548 26792 59560
rect 26375 59520 26792 59548
rect 26375 59517 26387 59520
rect 26329 59511 26387 59517
rect 26786 59508 26792 59520
rect 26844 59508 26850 59560
rect 27249 59551 27307 59557
rect 27249 59517 27261 59551
rect 27295 59548 27307 59551
rect 27801 59551 27859 59557
rect 27801 59548 27813 59551
rect 27295 59520 27813 59548
rect 27295 59517 27307 59520
rect 27249 59511 27307 59517
rect 27801 59517 27813 59520
rect 27847 59517 27859 59551
rect 27801 59511 27859 59517
rect 26510 59440 26516 59492
rect 26568 59480 26574 59492
rect 27264 59480 27292 59511
rect 28994 59508 29000 59560
rect 29052 59548 29058 59560
rect 31128 59557 31156 59588
rect 32306 59576 32312 59588
rect 32364 59576 32370 59628
rect 30009 59551 30067 59557
rect 30009 59548 30021 59551
rect 29052 59520 30021 59548
rect 29052 59508 29058 59520
rect 30009 59517 30021 59520
rect 30055 59548 30067 59551
rect 30285 59551 30343 59557
rect 30285 59548 30297 59551
rect 30055 59520 30297 59548
rect 30055 59517 30067 59520
rect 30009 59511 30067 59517
rect 30285 59517 30297 59520
rect 30331 59517 30343 59551
rect 30285 59511 30343 59517
rect 31113 59551 31171 59557
rect 31113 59517 31125 59551
rect 31159 59517 31171 59551
rect 31113 59511 31171 59517
rect 31205 59551 31263 59557
rect 31205 59517 31217 59551
rect 31251 59517 31263 59551
rect 31205 59511 31263 59517
rect 26568 59452 27292 59480
rect 29733 59483 29791 59489
rect 26568 59440 26574 59452
rect 29733 59449 29745 59483
rect 29779 59480 29791 59483
rect 31128 59480 31156 59511
rect 29779 59452 31156 59480
rect 29779 59449 29791 59452
rect 29733 59443 29791 59449
rect 20530 59412 20536 59424
rect 19383 59384 20536 59412
rect 19383 59381 19395 59384
rect 19337 59375 19395 59381
rect 20530 59372 20536 59384
rect 20588 59372 20594 59424
rect 20898 59412 20904 59424
rect 20859 59384 20904 59412
rect 20898 59372 20904 59384
rect 20956 59372 20962 59424
rect 23290 59412 23296 59424
rect 23251 59384 23296 59412
rect 23290 59372 23296 59384
rect 23348 59372 23354 59424
rect 28166 59412 28172 59424
rect 28127 59384 28172 59412
rect 28166 59372 28172 59384
rect 28224 59372 28230 59424
rect 29089 59415 29147 59421
rect 29089 59381 29101 59415
rect 29135 59412 29147 59415
rect 29178 59412 29184 59424
rect 29135 59384 29184 59412
rect 29135 59381 29147 59384
rect 29089 59375 29147 59381
rect 29178 59372 29184 59384
rect 29236 59372 29242 59424
rect 29914 59372 29920 59424
rect 29972 59412 29978 59424
rect 31220 59412 31248 59511
rect 29972 59384 31248 59412
rect 29972 59372 29978 59384
rect 1104 59322 38824 59344
rect 1104 59270 19606 59322
rect 19658 59270 19670 59322
rect 19722 59270 19734 59322
rect 19786 59270 19798 59322
rect 19850 59270 38824 59322
rect 1104 59248 38824 59270
rect 1578 59208 1584 59220
rect 1539 59180 1584 59208
rect 1578 59168 1584 59180
rect 1636 59168 1642 59220
rect 21542 59208 21548 59220
rect 21503 59180 21548 59208
rect 21542 59168 21548 59180
rect 21600 59168 21606 59220
rect 22094 59168 22100 59220
rect 22152 59208 22158 59220
rect 22370 59208 22376 59220
rect 22152 59180 22376 59208
rect 22152 59168 22158 59180
rect 22370 59168 22376 59180
rect 22428 59168 22434 59220
rect 19242 59140 19248 59152
rect 19203 59112 19248 59140
rect 19242 59100 19248 59112
rect 19300 59100 19306 59152
rect 19978 59100 19984 59152
rect 20036 59140 20042 59152
rect 20349 59143 20407 59149
rect 20349 59140 20361 59143
rect 20036 59112 20361 59140
rect 20036 59100 20042 59112
rect 20349 59109 20361 59112
rect 20395 59140 20407 59143
rect 21818 59140 21824 59152
rect 20395 59112 21824 59140
rect 20395 59109 20407 59112
rect 20349 59103 20407 59109
rect 21818 59100 21824 59112
rect 21876 59100 21882 59152
rect 24486 59100 24492 59152
rect 24544 59140 24550 59152
rect 26510 59140 26516 59152
rect 24544 59112 25268 59140
rect 26471 59112 26516 59140
rect 24544 59100 24550 59112
rect 16574 59032 16580 59084
rect 16632 59072 16638 59084
rect 16669 59075 16727 59081
rect 16669 59072 16681 59075
rect 16632 59044 16681 59072
rect 16632 59032 16638 59044
rect 16669 59041 16681 59044
rect 16715 59041 16727 59075
rect 16669 59035 16727 59041
rect 17402 59032 17408 59084
rect 17460 59072 17466 59084
rect 17681 59075 17739 59081
rect 17681 59072 17693 59075
rect 17460 59044 17693 59072
rect 17460 59032 17466 59044
rect 17681 59041 17693 59044
rect 17727 59041 17739 59075
rect 20898 59072 20904 59084
rect 20859 59044 20904 59072
rect 17681 59035 17739 59041
rect 20898 59032 20904 59044
rect 20956 59032 20962 59084
rect 23014 59072 23020 59084
rect 22975 59044 23020 59072
rect 23014 59032 23020 59044
rect 23072 59032 23078 59084
rect 23290 59072 23296 59084
rect 23251 59044 23296 59072
rect 23290 59032 23296 59044
rect 23348 59032 23354 59084
rect 23842 59032 23848 59084
rect 23900 59072 23906 59084
rect 24302 59072 24308 59084
rect 23900 59044 24308 59072
rect 23900 59032 23906 59044
rect 24302 59032 24308 59044
rect 24360 59072 24366 59084
rect 25240 59081 25268 59112
rect 26510 59100 26516 59112
rect 26568 59100 26574 59152
rect 26602 59100 26608 59152
rect 26660 59140 26666 59152
rect 29086 59140 29092 59152
rect 26660 59112 27568 59140
rect 29047 59112 29092 59140
rect 26660 59100 26666 59112
rect 24765 59075 24823 59081
rect 24765 59072 24777 59075
rect 24360 59044 24777 59072
rect 24360 59032 24366 59044
rect 24765 59041 24777 59044
rect 24811 59041 24823 59075
rect 24765 59035 24823 59041
rect 25225 59075 25283 59081
rect 25225 59041 25237 59075
rect 25271 59041 25283 59075
rect 25225 59035 25283 59041
rect 27246 59032 27252 59084
rect 27304 59072 27310 59084
rect 27540 59081 27568 59112
rect 29086 59100 29092 59112
rect 29144 59100 29150 59152
rect 27341 59075 27399 59081
rect 27341 59072 27353 59075
rect 27304 59044 27353 59072
rect 27304 59032 27310 59044
rect 27341 59041 27353 59044
rect 27387 59041 27399 59075
rect 27341 59035 27399 59041
rect 27525 59075 27583 59081
rect 27525 59041 27537 59075
rect 27571 59041 27583 59075
rect 29822 59072 29828 59084
rect 29783 59044 29828 59072
rect 27525 59035 27583 59041
rect 29822 59032 29828 59044
rect 29880 59032 29886 59084
rect 35161 59075 35219 59081
rect 35161 59041 35173 59075
rect 35207 59072 35219 59075
rect 35250 59072 35256 59084
rect 35207 59044 35256 59072
rect 35207 59041 35219 59044
rect 35161 59035 35219 59041
rect 35250 59032 35256 59044
rect 35308 59032 35314 59084
rect 35434 59072 35440 59084
rect 35395 59044 35440 59072
rect 35434 59032 35440 59044
rect 35492 59032 35498 59084
rect 17218 58964 17224 59016
rect 17276 59004 17282 59016
rect 17862 59004 17868 59016
rect 17276 58976 17868 59004
rect 17276 58964 17282 58976
rect 17862 58964 17868 58976
rect 17920 59004 17926 59016
rect 18046 59004 18052 59016
rect 17920 58976 18052 59004
rect 17920 58964 17926 58976
rect 18046 58964 18052 58976
rect 18104 58964 18110 59016
rect 18966 58964 18972 59016
rect 19024 59004 19030 59016
rect 19613 59007 19671 59013
rect 19613 59004 19625 59007
rect 19024 58976 19625 59004
rect 19024 58964 19030 58976
rect 19613 58973 19625 58976
rect 19659 58973 19671 59007
rect 19613 58967 19671 58973
rect 20438 58964 20444 59016
rect 20496 59004 20502 59016
rect 20717 59007 20775 59013
rect 20717 59004 20729 59007
rect 20496 58976 20729 59004
rect 20496 58964 20502 58976
rect 20717 58973 20729 58976
rect 20763 59004 20775 59007
rect 21269 59007 21327 59013
rect 21269 59004 21281 59007
rect 20763 58976 21281 59004
rect 20763 58973 20775 58976
rect 20717 58967 20775 58973
rect 21269 58973 21281 58976
rect 21315 58973 21327 59007
rect 21269 58967 21327 58973
rect 22649 59007 22707 59013
rect 22649 58973 22661 59007
rect 22695 59004 22707 59007
rect 22738 59004 22744 59016
rect 22695 58976 22744 59004
rect 22695 58973 22707 58976
rect 22649 58967 22707 58973
rect 22738 58964 22744 58976
rect 22796 58964 22802 59016
rect 24581 59007 24639 59013
rect 24581 58973 24593 59007
rect 24627 59004 24639 59007
rect 25130 59004 25136 59016
rect 24627 58976 25136 59004
rect 24627 58973 24639 58976
rect 24581 58967 24639 58973
rect 25130 58964 25136 58976
rect 25188 58964 25194 59016
rect 27062 59004 27068 59016
rect 27023 58976 27068 59004
rect 27062 58964 27068 58976
rect 27120 58964 27126 59016
rect 28994 59004 29000 59016
rect 28955 58976 29000 59004
rect 28994 58964 29000 58976
rect 29052 58964 29058 59016
rect 29730 58964 29736 59016
rect 29788 59004 29794 59016
rect 29917 59007 29975 59013
rect 29917 59004 29929 59007
rect 29788 58976 29929 59004
rect 29788 58964 29794 58976
rect 29917 58973 29929 58976
rect 29963 58973 29975 59007
rect 29917 58967 29975 58973
rect 19521 58939 19579 58945
rect 19521 58905 19533 58939
rect 19567 58936 19579 58939
rect 19978 58936 19984 58948
rect 19567 58908 19984 58936
rect 19567 58905 19579 58908
rect 19521 58899 19579 58905
rect 19978 58896 19984 58908
rect 20036 58936 20042 58948
rect 21177 58939 21235 58945
rect 21177 58936 21189 58939
rect 20036 58908 21189 58936
rect 20036 58896 20042 58908
rect 21177 58905 21189 58908
rect 21223 58905 21235 58939
rect 23382 58936 23388 58948
rect 23343 58908 23388 58936
rect 21177 58899 21235 58905
rect 23382 58896 23388 58908
rect 23440 58896 23446 58948
rect 25222 58936 25228 58948
rect 25183 58908 25228 58936
rect 25222 58896 25228 58908
rect 25280 58896 25286 58948
rect 26329 58939 26387 58945
rect 26329 58905 26341 58939
rect 26375 58936 26387 58939
rect 27080 58936 27108 58964
rect 26375 58908 27108 58936
rect 26375 58905 26387 58908
rect 26329 58899 26387 58905
rect 16758 58828 16764 58880
rect 16816 58868 16822 58880
rect 16853 58871 16911 58877
rect 16853 58868 16865 58871
rect 16816 58840 16865 58868
rect 16816 58828 16822 58840
rect 16853 58837 16865 58840
rect 16899 58837 16911 58871
rect 16853 58831 16911 58837
rect 17221 58871 17279 58877
rect 17221 58837 17233 58871
rect 17267 58868 17279 58871
rect 17402 58868 17408 58880
rect 17267 58840 17408 58868
rect 17267 58837 17279 58840
rect 17221 58831 17279 58837
rect 17402 58828 17408 58840
rect 17460 58828 17466 58880
rect 17589 58871 17647 58877
rect 17589 58837 17601 58871
rect 17635 58868 17647 58871
rect 17770 58868 17776 58880
rect 17635 58840 17776 58868
rect 17635 58837 17647 58840
rect 17589 58831 17647 58837
rect 17770 58828 17776 58840
rect 17828 58877 17834 58880
rect 17828 58871 17877 58877
rect 17828 58837 17831 58871
rect 17865 58837 17877 58871
rect 17828 58831 17877 58837
rect 17957 58871 18015 58877
rect 17957 58837 17969 58871
rect 18003 58868 18015 58871
rect 18046 58868 18052 58880
rect 18003 58840 18052 58868
rect 18003 58837 18015 58840
rect 17957 58831 18015 58837
rect 17828 58828 17834 58831
rect 18046 58828 18052 58840
rect 18104 58828 18110 58880
rect 18322 58868 18328 58880
rect 18283 58840 18328 58868
rect 18322 58828 18328 58840
rect 18380 58828 18386 58880
rect 18969 58871 19027 58877
rect 18969 58837 18981 58871
rect 19015 58868 19027 58871
rect 19058 58868 19064 58880
rect 19015 58840 19064 58868
rect 19015 58837 19027 58840
rect 18969 58831 19027 58837
rect 19058 58828 19064 58840
rect 19116 58868 19122 58880
rect 19383 58871 19441 58877
rect 19383 58868 19395 58871
rect 19116 58840 19395 58868
rect 19116 58828 19122 58840
rect 19383 58837 19395 58840
rect 19429 58837 19441 58871
rect 19886 58868 19892 58880
rect 19847 58840 19892 58868
rect 19383 58831 19441 58837
rect 19886 58828 19892 58840
rect 19944 58828 19950 58880
rect 20530 58828 20536 58880
rect 20588 58868 20594 58880
rect 21039 58871 21097 58877
rect 21039 58868 21051 58871
rect 20588 58840 21051 58868
rect 20588 58828 20594 58840
rect 21039 58837 21051 58840
rect 21085 58837 21097 58871
rect 21910 58868 21916 58880
rect 21871 58840 21916 58868
rect 21039 58831 21097 58837
rect 21910 58828 21916 58840
rect 21968 58828 21974 58880
rect 24029 58871 24087 58877
rect 24029 58837 24041 58871
rect 24075 58868 24087 58871
rect 24210 58868 24216 58880
rect 24075 58840 24216 58868
rect 24075 58837 24087 58840
rect 24029 58831 24087 58837
rect 24210 58828 24216 58840
rect 24268 58868 24274 58880
rect 24578 58868 24584 58880
rect 24268 58840 24584 58868
rect 24268 58828 24274 58840
rect 24578 58828 24584 58840
rect 24636 58828 24642 58880
rect 35802 58828 35808 58880
rect 35860 58868 35866 58880
rect 36541 58871 36599 58877
rect 36541 58868 36553 58871
rect 35860 58840 36553 58868
rect 35860 58828 35866 58840
rect 36541 58837 36553 58840
rect 36587 58837 36599 58871
rect 36541 58831 36599 58837
rect 1104 58778 38824 58800
rect 1104 58726 4246 58778
rect 4298 58726 4310 58778
rect 4362 58726 4374 58778
rect 4426 58726 4438 58778
rect 4490 58726 34966 58778
rect 35018 58726 35030 58778
rect 35082 58726 35094 58778
rect 35146 58726 35158 58778
rect 35210 58726 38824 58778
rect 1104 58704 38824 58726
rect 16853 58667 16911 58673
rect 16853 58633 16865 58667
rect 16899 58664 16911 58667
rect 17129 58667 17187 58673
rect 17129 58664 17141 58667
rect 16899 58636 17141 58664
rect 16899 58633 16911 58636
rect 16853 58627 16911 58633
rect 17129 58633 17141 58636
rect 17175 58664 17187 58667
rect 17218 58664 17224 58676
rect 17175 58636 17224 58664
rect 17175 58633 17187 58636
rect 17129 58627 17187 58633
rect 17218 58624 17224 58636
rect 17276 58624 17282 58676
rect 19058 58673 19064 58676
rect 19042 58667 19064 58673
rect 19042 58633 19054 58667
rect 19042 58627 19064 58633
rect 19058 58624 19064 58627
rect 19116 58624 19122 58676
rect 19337 58667 19395 58673
rect 19337 58633 19349 58667
rect 19383 58664 19395 58667
rect 19426 58664 19432 58676
rect 19383 58636 19432 58664
rect 19383 58633 19395 58636
rect 19337 58627 19395 58633
rect 19426 58624 19432 58636
rect 19484 58624 19490 58676
rect 22925 58667 22983 58673
rect 22925 58633 22937 58667
rect 22971 58664 22983 58667
rect 23014 58664 23020 58676
rect 22971 58636 23020 58664
rect 22971 58633 22983 58636
rect 22925 58627 22983 58633
rect 23014 58624 23020 58636
rect 23072 58624 23078 58676
rect 25130 58664 25136 58676
rect 25091 58636 25136 58664
rect 25130 58624 25136 58636
rect 25188 58624 25194 58676
rect 35253 58667 35311 58673
rect 35253 58633 35265 58667
rect 35299 58664 35311 58667
rect 35434 58664 35440 58676
rect 35299 58636 35440 58664
rect 35299 58633 35311 58636
rect 35253 58627 35311 58633
rect 35434 58624 35440 58636
rect 35492 58624 35498 58676
rect 18785 58599 18843 58605
rect 18785 58565 18797 58599
rect 18831 58596 18843 58599
rect 19150 58596 19156 58608
rect 18831 58568 19156 58596
rect 18831 58565 18843 58568
rect 18785 58559 18843 58565
rect 19150 58556 19156 58568
rect 19208 58556 19214 58608
rect 24118 58596 24124 58608
rect 23952 58568 24124 58596
rect 1578 58528 1584 58540
rect 1539 58500 1584 58528
rect 1578 58488 1584 58500
rect 1636 58488 1642 58540
rect 1854 58528 1860 58540
rect 1815 58500 1860 58528
rect 1854 58488 1860 58500
rect 1912 58488 1918 58540
rect 19245 58531 19303 58537
rect 19245 58497 19257 58531
rect 19291 58497 19303 58531
rect 21174 58528 21180 58540
rect 21135 58500 21180 58528
rect 19245 58491 19303 58497
rect 16942 58460 16948 58472
rect 16855 58432 16948 58460
rect 16942 58420 16948 58432
rect 17000 58460 17006 58472
rect 17405 58463 17463 58469
rect 17405 58460 17417 58463
rect 17000 58432 17417 58460
rect 17000 58420 17006 58432
rect 17405 58429 17417 58432
rect 17451 58429 17463 58463
rect 17405 58423 17463 58429
rect 18417 58463 18475 58469
rect 18417 58429 18429 58463
rect 18463 58460 18475 58463
rect 18966 58460 18972 58472
rect 18463 58432 18972 58460
rect 18463 58429 18475 58432
rect 18417 58423 18475 58429
rect 18966 58420 18972 58432
rect 19024 58460 19030 58472
rect 19260 58460 19288 58491
rect 21174 58488 21180 58500
rect 21232 58488 21238 58540
rect 21910 58488 21916 58540
rect 21968 58528 21974 58540
rect 23952 58537 23980 58568
rect 24118 58556 24124 58568
rect 24176 58596 24182 58608
rect 25869 58599 25927 58605
rect 25869 58596 25881 58599
rect 24176 58568 25881 58596
rect 24176 58556 24182 58568
rect 25869 58565 25881 58568
rect 25915 58565 25927 58599
rect 25869 58559 25927 58565
rect 26421 58599 26479 58605
rect 26421 58565 26433 58599
rect 26467 58596 26479 58599
rect 27246 58596 27252 58608
rect 26467 58568 27252 58596
rect 26467 58565 26479 58568
rect 26421 58559 26479 58565
rect 27246 58556 27252 58568
rect 27304 58556 27310 58608
rect 27706 58596 27712 58608
rect 27667 58568 27712 58596
rect 27706 58556 27712 58568
rect 27764 58556 27770 58608
rect 23477 58531 23535 58537
rect 21968 58500 22232 58528
rect 21968 58488 21974 58500
rect 19024 58432 19288 58460
rect 19024 58420 19030 58432
rect 21634 58420 21640 58472
rect 21692 58460 21698 58472
rect 21729 58463 21787 58469
rect 21729 58460 21741 58463
rect 21692 58432 21741 58460
rect 21692 58420 21698 58432
rect 21729 58429 21741 58432
rect 21775 58429 21787 58463
rect 21729 58423 21787 58429
rect 21818 58420 21824 58472
rect 21876 58460 21882 58472
rect 22204 58469 22232 58500
rect 23477 58497 23489 58531
rect 23523 58528 23535 58531
rect 23937 58531 23995 58537
rect 23937 58528 23949 58531
rect 23523 58500 23949 58528
rect 23523 58497 23535 58500
rect 23477 58491 23535 58497
rect 23937 58497 23949 58500
rect 23983 58497 23995 58531
rect 24762 58528 24768 58540
rect 24723 58500 24768 58528
rect 23937 58491 23995 58497
rect 24762 58488 24768 58500
rect 24820 58488 24826 58540
rect 22005 58463 22063 58469
rect 22005 58460 22017 58463
rect 21876 58432 22017 58460
rect 21876 58420 21882 58432
rect 22005 58429 22017 58432
rect 22051 58429 22063 58463
rect 22005 58423 22063 58429
rect 22189 58463 22247 58469
rect 22189 58429 22201 58463
rect 22235 58460 22247 58463
rect 22370 58460 22376 58472
rect 22235 58432 22376 58460
rect 22235 58429 22247 58432
rect 22189 58423 22247 58429
rect 22370 58420 22376 58432
rect 22428 58420 22434 58472
rect 24210 58460 24216 58472
rect 24171 58432 24216 58460
rect 24210 58420 24216 58432
rect 24268 58420 24274 58472
rect 24486 58420 24492 58472
rect 24544 58460 24550 58472
rect 24581 58463 24639 58469
rect 24581 58460 24593 58463
rect 24544 58432 24593 58460
rect 24544 58420 24550 58432
rect 24581 58429 24593 58432
rect 24627 58429 24639 58463
rect 25685 58463 25743 58469
rect 25685 58460 25697 58463
rect 24581 58423 24639 58429
rect 25516 58432 25697 58460
rect 18877 58395 18935 58401
rect 18877 58361 18889 58395
rect 18923 58392 18935 58395
rect 19150 58392 19156 58404
rect 18923 58364 19156 58392
rect 18923 58361 18935 58364
rect 18877 58355 18935 58361
rect 19150 58352 19156 58364
rect 19208 58352 19214 58404
rect 20901 58395 20959 58401
rect 20901 58392 20913 58395
rect 19996 58364 20913 58392
rect 19996 58336 20024 58364
rect 20901 58361 20913 58364
rect 20947 58361 20959 58395
rect 20901 58355 20959 58361
rect 23014 58352 23020 58404
rect 23072 58392 23078 58404
rect 25222 58392 25228 58404
rect 23072 58364 25228 58392
rect 23072 58352 23078 58364
rect 25222 58352 25228 58364
rect 25280 58352 25286 58404
rect 2958 58324 2964 58336
rect 2919 58296 2964 58324
rect 2958 58284 2964 58296
rect 3016 58284 3022 58336
rect 16485 58327 16543 58333
rect 16485 58293 16497 58327
rect 16531 58324 16543 58327
rect 16574 58324 16580 58336
rect 16531 58296 16580 58324
rect 16531 58293 16543 58296
rect 16485 58287 16543 58293
rect 16574 58284 16580 58296
rect 16632 58284 16638 58336
rect 17865 58327 17923 58333
rect 17865 58293 17877 58327
rect 17911 58324 17923 58327
rect 18138 58324 18144 58336
rect 17911 58296 18144 58324
rect 17911 58293 17923 58296
rect 17865 58287 17923 58293
rect 18138 58284 18144 58296
rect 18196 58284 18202 58336
rect 19978 58324 19984 58336
rect 19939 58296 19984 58324
rect 19978 58284 19984 58296
rect 20036 58284 20042 58336
rect 20530 58324 20536 58336
rect 20491 58296 20536 58324
rect 20530 58284 20536 58296
rect 20588 58284 20594 58336
rect 22557 58327 22615 58333
rect 22557 58293 22569 58327
rect 22603 58324 22615 58327
rect 22738 58324 22744 58336
rect 22603 58296 22744 58324
rect 22603 58293 22615 58296
rect 22557 58287 22615 58293
rect 22738 58284 22744 58296
rect 22796 58284 22802 58336
rect 25314 58284 25320 58336
rect 25372 58324 25378 58336
rect 25516 58333 25544 58432
rect 25685 58429 25697 58432
rect 25731 58429 25743 58463
rect 26878 58460 26884 58472
rect 26839 58432 26884 58460
rect 25685 58423 25743 58429
rect 26878 58420 26884 58432
rect 26936 58420 26942 58472
rect 27433 58463 27491 58469
rect 27433 58429 27445 58463
rect 27479 58429 27491 58463
rect 27433 58423 27491 58429
rect 25501 58327 25559 58333
rect 25501 58324 25513 58327
rect 25372 58296 25513 58324
rect 25372 58284 25378 58296
rect 25501 58293 25513 58296
rect 25547 58293 25559 58327
rect 26786 58324 26792 58336
rect 26699 58296 26792 58324
rect 25501 58287 25559 58293
rect 26786 58284 26792 58296
rect 26844 58324 26850 58336
rect 27448 58324 27476 58423
rect 27614 58420 27620 58472
rect 27672 58460 27678 58472
rect 27709 58463 27767 58469
rect 27709 58460 27721 58463
rect 27672 58432 27721 58460
rect 27672 58420 27678 58432
rect 27709 58429 27721 58432
rect 27755 58460 27767 58463
rect 28261 58463 28319 58469
rect 28261 58460 28273 58463
rect 27755 58432 28273 58460
rect 27755 58429 27767 58432
rect 27709 58423 27767 58429
rect 28261 58429 28273 58432
rect 28307 58460 28319 58463
rect 28905 58463 28963 58469
rect 28905 58460 28917 58463
rect 28307 58432 28917 58460
rect 28307 58429 28319 58432
rect 28261 58423 28319 58429
rect 28905 58429 28917 58432
rect 28951 58460 28963 58463
rect 28994 58460 29000 58472
rect 28951 58432 29000 58460
rect 28951 58429 28963 58432
rect 28905 58423 28963 58429
rect 28994 58420 29000 58432
rect 29052 58420 29058 58472
rect 27614 58324 27620 58336
rect 26844 58296 27620 58324
rect 26844 58284 26850 58296
rect 27614 58284 27620 58296
rect 27672 58284 27678 58336
rect 29549 58327 29607 58333
rect 29549 58293 29561 58327
rect 29595 58324 29607 58327
rect 29730 58324 29736 58336
rect 29595 58296 29736 58324
rect 29595 58293 29607 58296
rect 29549 58287 29607 58293
rect 29730 58284 29736 58296
rect 29788 58284 29794 58336
rect 35250 58284 35256 58336
rect 35308 58324 35314 58336
rect 35529 58327 35587 58333
rect 35529 58324 35541 58327
rect 35308 58296 35541 58324
rect 35308 58284 35314 58296
rect 35529 58293 35541 58296
rect 35575 58293 35587 58327
rect 35529 58287 35587 58293
rect 1104 58234 38824 58256
rect 1104 58182 19606 58234
rect 19658 58182 19670 58234
rect 19722 58182 19734 58234
rect 19786 58182 19798 58234
rect 19850 58182 38824 58234
rect 1104 58160 38824 58182
rect 1673 58123 1731 58129
rect 1673 58089 1685 58123
rect 1719 58120 1731 58123
rect 1854 58120 1860 58132
rect 1719 58092 1860 58120
rect 1719 58089 1731 58092
rect 1673 58083 1731 58089
rect 1854 58080 1860 58092
rect 1912 58080 1918 58132
rect 15654 58120 15660 58132
rect 15615 58092 15660 58120
rect 15654 58080 15660 58092
rect 15712 58080 15718 58132
rect 19334 58080 19340 58132
rect 19392 58120 19398 58132
rect 19705 58123 19763 58129
rect 19705 58120 19717 58123
rect 19392 58092 19717 58120
rect 19392 58080 19398 58092
rect 19705 58089 19717 58092
rect 19751 58089 19763 58123
rect 19705 58083 19763 58089
rect 24486 58080 24492 58132
rect 24544 58120 24550 58132
rect 25777 58123 25835 58129
rect 25777 58120 25789 58123
rect 24544 58092 25789 58120
rect 24544 58080 24550 58092
rect 25777 58089 25789 58092
rect 25823 58089 25835 58123
rect 25777 58083 25835 58089
rect 26329 58123 26387 58129
rect 26329 58089 26341 58123
rect 26375 58120 26387 58123
rect 26602 58120 26608 58132
rect 26375 58092 26608 58120
rect 26375 58089 26387 58092
rect 26329 58083 26387 58089
rect 26602 58080 26608 58092
rect 26660 58080 26666 58132
rect 28997 58123 29055 58129
rect 28997 58089 29009 58123
rect 29043 58120 29055 58123
rect 29822 58120 29828 58132
rect 29043 58092 29828 58120
rect 29043 58089 29055 58092
rect 28997 58083 29055 58089
rect 29822 58080 29828 58092
rect 29880 58080 29886 58132
rect 17497 58055 17555 58061
rect 17497 58052 17509 58055
rect 15488 58024 17509 58052
rect 15102 57944 15108 57996
rect 15160 57984 15166 57996
rect 15488 57993 15516 58024
rect 17497 58021 17509 58024
rect 17543 58021 17555 58055
rect 17497 58015 17555 58021
rect 20717 58055 20775 58061
rect 20717 58021 20729 58055
rect 20763 58052 20775 58055
rect 20898 58052 20904 58064
rect 20763 58024 20904 58052
rect 20763 58021 20775 58024
rect 20717 58015 20775 58021
rect 20898 58012 20904 58024
rect 20956 58012 20962 58064
rect 23400 58024 23704 58052
rect 15473 57987 15531 57993
rect 15473 57984 15485 57987
rect 15160 57956 15485 57984
rect 15160 57944 15166 57956
rect 15473 57953 15485 57956
rect 15519 57953 15531 57987
rect 16477 57987 16535 57993
rect 16477 57984 16489 57987
rect 15473 57947 15531 57953
rect 16408 57956 16489 57984
rect 9122 57876 9128 57928
rect 9180 57916 9186 57928
rect 9490 57916 9496 57928
rect 9180 57888 9496 57916
rect 9180 57876 9186 57888
rect 9490 57876 9496 57888
rect 9548 57876 9554 57928
rect 13722 57876 13728 57928
rect 13780 57916 13786 57928
rect 13906 57916 13912 57928
rect 13780 57888 13912 57916
rect 13780 57876 13786 57888
rect 13906 57876 13912 57888
rect 13964 57876 13970 57928
rect 16408 57848 16436 57956
rect 16477 57953 16489 57956
rect 16523 57953 16535 57987
rect 16477 57947 16535 57953
rect 17865 57987 17923 57993
rect 17865 57953 17877 57987
rect 17911 57953 17923 57987
rect 17865 57947 17923 57953
rect 19061 57987 19119 57993
rect 19061 57953 19073 57987
rect 19107 57984 19119 57987
rect 19150 57984 19156 57996
rect 19107 57956 19156 57984
rect 19107 57953 19119 57956
rect 19061 57947 19119 57953
rect 17880 57916 17908 57947
rect 19150 57944 19156 57956
rect 19208 57944 19214 57996
rect 18046 57916 18052 57928
rect 17880 57888 18052 57916
rect 18046 57876 18052 57888
rect 18104 57876 18110 57928
rect 18966 57876 18972 57928
rect 19024 57916 19030 57928
rect 19429 57919 19487 57925
rect 19429 57916 19441 57919
rect 19024 57888 19441 57916
rect 19024 57876 19030 57888
rect 19429 57885 19441 57888
rect 19475 57885 19487 57919
rect 20162 57916 20168 57928
rect 20075 57888 20168 57916
rect 19429 57879 19487 57885
rect 20162 57876 20168 57888
rect 20220 57916 20226 57928
rect 20916 57916 20944 58012
rect 23109 57987 23167 57993
rect 23109 57953 23121 57987
rect 23155 57984 23167 57987
rect 23290 57984 23296 57996
rect 23155 57956 23296 57984
rect 23155 57953 23167 57956
rect 23109 57947 23167 57953
rect 23290 57944 23296 57956
rect 23348 57944 23354 57996
rect 20220 57888 20944 57916
rect 21269 57919 21327 57925
rect 20220 57876 20226 57888
rect 21269 57885 21281 57919
rect 21315 57885 21327 57919
rect 22738 57916 22744 57928
rect 22699 57888 22744 57916
rect 21269 57879 21327 57885
rect 18601 57851 18659 57857
rect 16408 57820 17080 57848
rect 16393 57783 16451 57789
rect 16393 57749 16405 57783
rect 16439 57780 16451 57783
rect 16482 57780 16488 57792
rect 16439 57752 16488 57780
rect 16439 57749 16451 57752
rect 16393 57743 16451 57749
rect 16482 57740 16488 57752
rect 16540 57740 16546 57792
rect 16666 57780 16672 57792
rect 16627 57752 16672 57780
rect 16666 57740 16672 57752
rect 16724 57740 16730 57792
rect 17052 57789 17080 57820
rect 18601 57817 18613 57851
rect 18647 57848 18659 57851
rect 19058 57848 19064 57860
rect 18647 57820 19064 57848
rect 18647 57817 18659 57820
rect 18601 57811 18659 57817
rect 19058 57808 19064 57820
rect 19116 57848 19122 57860
rect 19199 57851 19257 57857
rect 19199 57848 19211 57851
rect 19116 57820 19211 57848
rect 19116 57808 19122 57820
rect 19199 57817 19211 57820
rect 19245 57817 19257 57851
rect 19199 57811 19257 57817
rect 20898 57808 20904 57860
rect 20956 57848 20962 57860
rect 21284 57848 21312 57879
rect 22738 57876 22744 57888
rect 22796 57876 22802 57928
rect 22830 57876 22836 57928
rect 22888 57916 22894 57928
rect 23400 57916 23428 58024
rect 23523 57987 23581 57993
rect 23523 57953 23535 57987
rect 23569 57984 23581 57987
rect 23676 57984 23704 58024
rect 28718 58012 28724 58064
rect 28776 58052 28782 58064
rect 28776 58024 28856 58052
rect 28776 58012 28782 58024
rect 28828 57996 28856 58024
rect 23569 57956 23704 57984
rect 23569 57953 23581 57956
rect 23523 57947 23581 57953
rect 24026 57944 24032 57996
rect 24084 57984 24090 57996
rect 24489 57987 24547 57993
rect 24489 57984 24501 57987
rect 24084 57956 24501 57984
rect 24084 57944 24090 57956
rect 24489 57953 24501 57956
rect 24535 57953 24547 57987
rect 24489 57947 24547 57953
rect 25222 57944 25228 57996
rect 25280 57984 25286 57996
rect 25317 57987 25375 57993
rect 25317 57984 25329 57987
rect 25280 57956 25329 57984
rect 25280 57944 25286 57956
rect 25317 57953 25329 57956
rect 25363 57953 25375 57987
rect 28442 57984 28448 57996
rect 28403 57956 28448 57984
rect 25317 57947 25375 57953
rect 28442 57944 28448 57956
rect 28500 57944 28506 57996
rect 28810 57944 28816 57996
rect 28868 57944 28874 57996
rect 22888 57888 23428 57916
rect 25041 57919 25099 57925
rect 22888 57876 22894 57888
rect 25041 57885 25053 57919
rect 25087 57885 25099 57919
rect 25501 57919 25559 57925
rect 25501 57916 25513 57919
rect 25041 57879 25099 57885
rect 25424 57888 25513 57916
rect 20956 57820 21312 57848
rect 20956 57808 20962 57820
rect 22462 57808 22468 57860
rect 22520 57848 22526 57860
rect 23385 57851 23443 57857
rect 23385 57848 23397 57851
rect 22520 57820 23397 57848
rect 22520 57808 22526 57820
rect 23385 57817 23397 57820
rect 23431 57817 23443 57851
rect 24302 57848 24308 57860
rect 24263 57820 24308 57848
rect 23385 57811 23443 57817
rect 24302 57808 24308 57820
rect 24360 57848 24366 57860
rect 25056 57848 25084 57879
rect 24360 57820 25084 57848
rect 24360 57808 24366 57820
rect 17037 57783 17095 57789
rect 17037 57749 17049 57783
rect 17083 57780 17095 57783
rect 17126 57780 17132 57792
rect 17083 57752 17132 57780
rect 17083 57749 17095 57752
rect 17037 57743 17095 57749
rect 17126 57740 17132 57752
rect 17184 57740 17190 57792
rect 17402 57780 17408 57792
rect 17363 57752 17408 57780
rect 17402 57740 17408 57752
rect 17460 57740 17466 57792
rect 18966 57780 18972 57792
rect 18927 57752 18972 57780
rect 18966 57740 18972 57752
rect 19024 57740 19030 57792
rect 19337 57783 19395 57789
rect 19337 57749 19349 57783
rect 19383 57780 19395 57783
rect 19426 57780 19432 57792
rect 19383 57752 19432 57780
rect 19383 57749 19395 57752
rect 19337 57743 19395 57749
rect 19426 57740 19432 57752
rect 19484 57740 19490 57792
rect 20622 57740 20628 57792
rect 20680 57780 20686 57792
rect 21039 57783 21097 57789
rect 21039 57780 21051 57783
rect 20680 57752 21051 57780
rect 20680 57740 20686 57752
rect 21039 57749 21051 57752
rect 21085 57749 21097 57783
rect 21174 57780 21180 57792
rect 21135 57752 21180 57780
rect 21039 57743 21097 57749
rect 21174 57740 21180 57752
rect 21232 57740 21238 57792
rect 21358 57780 21364 57792
rect 21319 57752 21364 57780
rect 21358 57740 21364 57752
rect 21416 57740 21422 57792
rect 22002 57780 22008 57792
rect 21963 57752 22008 57780
rect 22002 57740 22008 57752
rect 22060 57740 22066 57792
rect 22370 57780 22376 57792
rect 22331 57752 22376 57780
rect 22370 57740 22376 57752
rect 22428 57740 22434 57792
rect 23474 57740 23480 57792
rect 23532 57780 23538 57792
rect 23937 57783 23995 57789
rect 23937 57780 23949 57783
rect 23532 57752 23949 57780
rect 23532 57740 23538 57752
rect 23937 57749 23949 57752
rect 23983 57780 23995 57783
rect 24210 57780 24216 57792
rect 23983 57752 24216 57780
rect 23983 57749 23995 57752
rect 23937 57743 23995 57749
rect 24210 57740 24216 57752
rect 24268 57740 24274 57792
rect 24762 57740 24768 57792
rect 24820 57780 24826 57792
rect 25424 57780 25452 57888
rect 25501 57885 25513 57888
rect 25547 57885 25559 57919
rect 25501 57879 25559 57885
rect 27338 57876 27344 57928
rect 27396 57916 27402 57928
rect 27617 57919 27675 57925
rect 27617 57916 27629 57919
rect 27396 57888 27629 57916
rect 27396 57876 27402 57888
rect 27617 57885 27629 57888
rect 27663 57885 27675 57919
rect 27617 57879 27675 57885
rect 28169 57919 28227 57925
rect 28169 57885 28181 57919
rect 28215 57916 28227 57919
rect 28534 57916 28540 57928
rect 28215 57888 28540 57916
rect 28215 57885 28227 57888
rect 28169 57879 28227 57885
rect 28534 57876 28540 57888
rect 28592 57876 28598 57928
rect 28626 57876 28632 57928
rect 28684 57916 28690 57928
rect 28684 57888 28729 57916
rect 28684 57876 28690 57888
rect 30006 57876 30012 57928
rect 30064 57916 30070 57928
rect 30558 57916 30564 57928
rect 30064 57888 30564 57916
rect 30064 57876 30070 57888
rect 30558 57876 30564 57888
rect 30616 57876 30622 57928
rect 24820 57752 25452 57780
rect 24820 57740 24826 57752
rect 26878 57740 26884 57792
rect 26936 57780 26942 57792
rect 26973 57783 27031 57789
rect 26973 57780 26985 57783
rect 26936 57752 26985 57780
rect 26936 57740 26942 57752
rect 26973 57749 26985 57752
rect 27019 57780 27031 57783
rect 27433 57783 27491 57789
rect 27433 57780 27445 57783
rect 27019 57752 27445 57780
rect 27019 57749 27031 57752
rect 26973 57743 27031 57749
rect 27433 57749 27445 57752
rect 27479 57780 27491 57783
rect 28350 57780 28356 57792
rect 27479 57752 28356 57780
rect 27479 57749 27491 57752
rect 27433 57743 27491 57749
rect 28350 57740 28356 57752
rect 28408 57740 28414 57792
rect 1104 57690 38824 57712
rect 1104 57638 4246 57690
rect 4298 57638 4310 57690
rect 4362 57638 4374 57690
rect 4426 57638 4438 57690
rect 4490 57638 34966 57690
rect 35018 57638 35030 57690
rect 35082 57638 35094 57690
rect 35146 57638 35158 57690
rect 35210 57638 38824 57690
rect 1104 57616 38824 57638
rect 14274 57576 14280 57588
rect 14235 57548 14280 57576
rect 14274 57536 14280 57548
rect 14332 57536 14338 57588
rect 14737 57579 14795 57585
rect 14737 57545 14749 57579
rect 14783 57576 14795 57579
rect 15102 57576 15108 57588
rect 14783 57548 15108 57576
rect 14783 57545 14795 57548
rect 14737 57539 14795 57545
rect 15102 57536 15108 57548
rect 15160 57536 15166 57588
rect 17862 57576 17868 57588
rect 17823 57548 17868 57576
rect 17862 57536 17868 57548
rect 17920 57536 17926 57588
rect 19058 57536 19064 57588
rect 19116 57576 19122 57588
rect 19291 57579 19349 57585
rect 19291 57576 19303 57579
rect 19116 57548 19303 57576
rect 19116 57536 19122 57548
rect 19291 57545 19303 57548
rect 19337 57545 19349 57579
rect 19610 57576 19616 57588
rect 19571 57548 19616 57576
rect 19291 57539 19349 57545
rect 19610 57536 19616 57548
rect 19668 57536 19674 57588
rect 20257 57579 20315 57585
rect 20257 57545 20269 57579
rect 20303 57576 20315 57579
rect 21174 57576 21180 57588
rect 20303 57548 21180 57576
rect 20303 57545 20315 57548
rect 20257 57539 20315 57545
rect 14292 57440 14320 57536
rect 18138 57468 18144 57520
rect 18196 57508 18202 57520
rect 18325 57511 18383 57517
rect 18325 57508 18337 57511
rect 18196 57480 18337 57508
rect 18196 57468 18202 57480
rect 18325 57477 18337 57480
rect 18371 57508 18383 57511
rect 18693 57511 18751 57517
rect 18693 57508 18705 57511
rect 18371 57480 18705 57508
rect 18371 57477 18383 57480
rect 18325 57471 18383 57477
rect 18693 57477 18705 57480
rect 18739 57508 18751 57511
rect 19426 57508 19432 57520
rect 18739 57480 19432 57508
rect 18739 57477 18751 57480
rect 18693 57471 18751 57477
rect 19426 57468 19432 57480
rect 19484 57508 19490 57520
rect 20272 57508 20300 57539
rect 21174 57536 21180 57548
rect 21232 57576 21238 57588
rect 21545 57579 21603 57585
rect 21545 57576 21557 57579
rect 21232 57548 21557 57576
rect 21232 57536 21238 57548
rect 21545 57545 21557 57548
rect 21591 57545 21603 57579
rect 24118 57576 24124 57588
rect 24079 57548 24124 57576
rect 21545 57539 21603 57545
rect 24118 57536 24124 57548
rect 24176 57536 24182 57588
rect 25130 57536 25136 57588
rect 25188 57576 25194 57588
rect 25593 57579 25651 57585
rect 25593 57576 25605 57579
rect 25188 57548 25605 57576
rect 25188 57536 25194 57548
rect 25593 57545 25605 57548
rect 25639 57545 25651 57579
rect 28994 57576 29000 57588
rect 28955 57548 29000 57576
rect 25593 57539 25651 57545
rect 19484 57480 20300 57508
rect 20901 57511 20959 57517
rect 19484 57468 19490 57480
rect 20901 57477 20913 57511
rect 20947 57508 20959 57511
rect 22002 57508 22008 57520
rect 20947 57480 22008 57508
rect 20947 57477 20959 57480
rect 20901 57471 20959 57477
rect 22002 57468 22008 57480
rect 22060 57508 22066 57520
rect 25222 57508 25228 57520
rect 22060 57480 22600 57508
rect 25183 57480 25228 57508
rect 22060 57468 22066 57480
rect 15197 57443 15255 57449
rect 15197 57440 15209 57443
rect 14292 57412 15209 57440
rect 15197 57409 15209 57412
rect 15243 57409 15255 57443
rect 15197 57403 15255 57409
rect 19521 57443 19579 57449
rect 19521 57409 19533 57443
rect 19567 57440 19579 57443
rect 20438 57440 20444 57452
rect 19567 57412 20444 57440
rect 19567 57409 19579 57412
rect 19521 57403 19579 57409
rect 15473 57375 15531 57381
rect 15473 57372 15485 57375
rect 15304 57344 15485 57372
rect 15010 57304 15016 57316
rect 14971 57276 15016 57304
rect 15010 57264 15016 57276
rect 15068 57304 15074 57316
rect 15304 57304 15332 57344
rect 15473 57341 15485 57344
rect 15519 57341 15531 57375
rect 15473 57335 15531 57341
rect 16574 57332 16580 57384
rect 16632 57372 16638 57384
rect 16853 57375 16911 57381
rect 16853 57372 16865 57375
rect 16632 57344 16865 57372
rect 16632 57332 16638 57344
rect 16853 57341 16865 57344
rect 16899 57372 16911 57375
rect 18138 57372 18144 57384
rect 16899 57344 18144 57372
rect 16899 57341 16911 57344
rect 16853 57335 16911 57341
rect 18138 57332 18144 57344
rect 18196 57332 18202 57384
rect 19426 57332 19432 57384
rect 19484 57372 19490 57384
rect 19536 57372 19564 57403
rect 20438 57400 20444 57412
rect 20496 57400 20502 57452
rect 21729 57443 21787 57449
rect 21729 57409 21741 57443
rect 21775 57440 21787 57443
rect 21910 57440 21916 57452
rect 21775 57412 21916 57440
rect 21775 57409 21787 57412
rect 21729 57403 21787 57409
rect 21910 57400 21916 57412
rect 21968 57400 21974 57452
rect 20714 57372 20720 57384
rect 19484 57344 19564 57372
rect 20627 57344 20720 57372
rect 19484 57332 19490 57344
rect 20714 57332 20720 57344
rect 20772 57372 20778 57384
rect 21358 57372 21364 57384
rect 20772 57344 21364 57372
rect 20772 57332 20778 57344
rect 21358 57332 21364 57344
rect 21416 57332 21422 57384
rect 22278 57372 22284 57384
rect 22239 57344 22284 57372
rect 22278 57332 22284 57344
rect 22336 57332 22342 57384
rect 22370 57332 22376 57384
rect 22428 57381 22434 57384
rect 22572 57381 22600 57480
rect 25222 57468 25228 57480
rect 25280 57468 25286 57520
rect 22428 57375 22477 57381
rect 22428 57341 22431 57375
rect 22465 57341 22477 57375
rect 22428 57335 22477 57341
rect 22557 57375 22615 57381
rect 22557 57341 22569 57375
rect 22603 57341 22615 57375
rect 22557 57335 22615 57341
rect 22428 57332 22434 57335
rect 15068 57276 15332 57304
rect 15068 57264 15074 57276
rect 17402 57264 17408 57316
rect 17460 57304 17466 57316
rect 17497 57307 17555 57313
rect 17497 57304 17509 57307
rect 17460 57276 17509 57304
rect 17460 57264 17466 57276
rect 17497 57273 17509 57276
rect 17543 57304 17555 57307
rect 17862 57304 17868 57316
rect 17543 57276 17868 57304
rect 17543 57273 17555 57276
rect 17497 57267 17555 57273
rect 17862 57264 17868 57276
rect 17920 57304 17926 57316
rect 19150 57304 19156 57316
rect 17920 57276 19156 57304
rect 17920 57264 17926 57276
rect 19150 57264 19156 57276
rect 19208 57264 19214 57316
rect 22572 57304 22600 57335
rect 22738 57332 22744 57384
rect 22796 57372 22802 57384
rect 23109 57375 23167 57381
rect 23109 57372 23121 57375
rect 22796 57344 23121 57372
rect 22796 57332 22802 57344
rect 23109 57341 23121 57344
rect 23155 57372 23167 57375
rect 23566 57372 23572 57384
rect 23155 57344 23572 57372
rect 23155 57341 23167 57344
rect 23109 57335 23167 57341
rect 23566 57332 23572 57344
rect 23624 57332 23630 57384
rect 24118 57332 24124 57384
rect 24176 57372 24182 57384
rect 24305 57375 24363 57381
rect 24305 57372 24317 57375
rect 24176 57344 24317 57372
rect 24176 57332 24182 57344
rect 24305 57341 24317 57344
rect 24351 57341 24363 57375
rect 25608 57372 25636 57539
rect 28994 57536 29000 57548
rect 29052 57536 29058 57588
rect 27246 57508 27252 57520
rect 27159 57480 27252 57508
rect 27246 57468 27252 57480
rect 27304 57508 27310 57520
rect 27304 57480 28212 57508
rect 27304 57468 27310 57480
rect 27341 57443 27399 57449
rect 27341 57409 27353 57443
rect 27387 57440 27399 57443
rect 27522 57440 27528 57452
rect 27387 57412 27528 57440
rect 27387 57409 27399 57412
rect 27341 57403 27399 57409
rect 27522 57400 27528 57412
rect 27580 57400 27586 57452
rect 28184 57440 28212 57480
rect 28442 57440 28448 57452
rect 28184 57412 28448 57440
rect 25869 57375 25927 57381
rect 25869 57372 25881 57375
rect 25608 57344 25881 57372
rect 24305 57335 24363 57341
rect 25869 57341 25881 57344
rect 25915 57372 25927 57375
rect 26694 57372 26700 57384
rect 25915 57344 26700 57372
rect 25915 57341 25927 57344
rect 25869 57335 25927 57341
rect 26694 57332 26700 57344
rect 26752 57332 26758 57384
rect 28184 57381 28212 57412
rect 28442 57400 28448 57412
rect 28500 57400 28506 57452
rect 28626 57400 28632 57452
rect 28684 57440 28690 57452
rect 29273 57443 29331 57449
rect 29273 57440 29285 57443
rect 28684 57412 29285 57440
rect 28684 57400 28690 57412
rect 29273 57409 29285 57412
rect 29319 57409 29331 57443
rect 29273 57403 29331 57409
rect 35161 57443 35219 57449
rect 35161 57409 35173 57443
rect 35207 57440 35219 57443
rect 35207 57412 35572 57440
rect 35207 57409 35219 57412
rect 35161 57403 35219 57409
rect 27893 57375 27951 57381
rect 27893 57341 27905 57375
rect 27939 57341 27951 57375
rect 27893 57335 27951 57341
rect 28169 57375 28227 57381
rect 28169 57341 28181 57375
rect 28215 57341 28227 57375
rect 28350 57372 28356 57384
rect 28311 57344 28356 57372
rect 28169 57335 28227 57341
rect 22572 57276 23336 57304
rect 23308 57248 23336 57276
rect 25590 57264 25596 57316
rect 25648 57304 25654 57316
rect 25777 57307 25835 57313
rect 25777 57304 25789 57307
rect 25648 57276 25789 57304
rect 25648 57264 25654 57276
rect 25777 57273 25789 57276
rect 25823 57273 25835 57307
rect 25777 57267 25835 57273
rect 26881 57307 26939 57313
rect 26881 57273 26893 57307
rect 26927 57304 26939 57307
rect 27908 57304 27936 57335
rect 28350 57332 28356 57344
rect 28408 57332 28414 57384
rect 28994 57332 29000 57384
rect 29052 57372 29058 57384
rect 29365 57375 29423 57381
rect 29365 57372 29377 57375
rect 29052 57344 29377 57372
rect 29052 57332 29058 57344
rect 29365 57341 29377 57344
rect 29411 57341 29423 57375
rect 35250 57372 35256 57384
rect 35211 57344 35256 57372
rect 29365 57335 29423 57341
rect 35250 57332 35256 57344
rect 35308 57332 35314 57384
rect 35544 57381 35572 57412
rect 35529 57375 35587 57381
rect 35529 57341 35541 57375
rect 35575 57372 35587 57375
rect 35802 57372 35808 57384
rect 35575 57344 35808 57372
rect 35575 57341 35587 57344
rect 35529 57335 35587 57341
rect 35802 57332 35808 57344
rect 35860 57332 35866 57384
rect 28718 57304 28724 57316
rect 26927 57276 28724 57304
rect 26927 57273 26939 57276
rect 26881 57267 26939 57273
rect 28718 57264 28724 57276
rect 28776 57264 28782 57316
rect 18046 57196 18052 57248
rect 18104 57236 18110 57248
rect 18966 57236 18972 57248
rect 18104 57208 18972 57236
rect 18104 57196 18110 57208
rect 18966 57196 18972 57208
rect 19024 57236 19030 57248
rect 19242 57236 19248 57248
rect 19024 57208 19248 57236
rect 19024 57196 19030 57208
rect 19242 57196 19248 57208
rect 19300 57196 19306 57248
rect 20438 57196 20444 57248
rect 20496 57236 20502 57248
rect 20533 57239 20591 57245
rect 20533 57236 20545 57239
rect 20496 57208 20545 57236
rect 20496 57196 20502 57208
rect 20533 57205 20545 57208
rect 20579 57236 20591 57239
rect 20622 57236 20628 57248
rect 20579 57208 20628 57236
rect 20579 57205 20591 57208
rect 20533 57199 20591 57205
rect 20622 57196 20628 57208
rect 20680 57196 20686 57248
rect 20898 57196 20904 57248
rect 20956 57236 20962 57248
rect 21177 57239 21235 57245
rect 21177 57236 21189 57239
rect 20956 57208 21189 57236
rect 20956 57196 20962 57208
rect 21177 57205 21189 57208
rect 21223 57205 21235 57239
rect 21177 57199 21235 57205
rect 23290 57196 23296 57248
rect 23348 57236 23354 57248
rect 23385 57239 23443 57245
rect 23385 57236 23397 57239
rect 23348 57208 23397 57236
rect 23348 57196 23354 57208
rect 23385 57205 23397 57208
rect 23431 57205 23443 57239
rect 23385 57199 23443 57205
rect 24302 57196 24308 57248
rect 24360 57236 24366 57248
rect 24489 57239 24547 57245
rect 24489 57236 24501 57239
rect 24360 57208 24501 57236
rect 24360 57196 24366 57208
rect 24489 57205 24501 57208
rect 24535 57205 24547 57239
rect 24489 57199 24547 57205
rect 28534 57196 28540 57248
rect 28592 57236 28598 57248
rect 28629 57239 28687 57245
rect 28629 57236 28641 57239
rect 28592 57208 28641 57236
rect 28592 57196 28598 57208
rect 28629 57205 28641 57208
rect 28675 57205 28687 57239
rect 28629 57199 28687 57205
rect 35894 57196 35900 57248
rect 35952 57236 35958 57248
rect 36633 57239 36691 57245
rect 36633 57236 36645 57239
rect 35952 57208 36645 57236
rect 35952 57196 35958 57208
rect 36633 57205 36645 57208
rect 36679 57205 36691 57239
rect 36633 57199 36691 57205
rect 1104 57146 38824 57168
rect 1104 57094 19606 57146
rect 19658 57094 19670 57146
rect 19722 57094 19734 57146
rect 19786 57094 19798 57146
rect 19850 57094 38824 57146
rect 1104 57072 38824 57094
rect 18233 57035 18291 57041
rect 18233 57001 18245 57035
rect 18279 57032 18291 57035
rect 18601 57035 18659 57041
rect 18601 57032 18613 57035
rect 18279 57004 18613 57032
rect 18279 57001 18291 57004
rect 18233 56995 18291 57001
rect 18601 57001 18613 57004
rect 18647 57032 18659 57035
rect 18969 57035 19027 57041
rect 18969 57032 18981 57035
rect 18647 57004 18981 57032
rect 18647 57001 18659 57004
rect 18601 56995 18659 57001
rect 18969 57001 18981 57004
rect 19015 57032 19027 57035
rect 19058 57032 19064 57044
rect 19015 57004 19064 57032
rect 19015 57001 19027 57004
rect 18969 56995 19027 57001
rect 19058 56992 19064 57004
rect 19116 56992 19122 57044
rect 20162 57032 20168 57044
rect 20123 57004 20168 57032
rect 20162 56992 20168 57004
rect 20220 56992 20226 57044
rect 20714 57032 20720 57044
rect 20675 57004 20720 57032
rect 20714 56992 20720 57004
rect 20772 56992 20778 57044
rect 22649 57035 22707 57041
rect 22649 57032 22661 57035
rect 22020 57004 22661 57032
rect 19150 56924 19156 56976
rect 19208 56964 19214 56976
rect 19334 56964 19340 56976
rect 19208 56936 19340 56964
rect 19208 56924 19214 56936
rect 19334 56924 19340 56936
rect 19392 56924 19398 56976
rect 20180 56964 20208 56992
rect 21085 56967 21143 56973
rect 21085 56964 21097 56967
rect 20180 56936 21097 56964
rect 21085 56933 21097 56936
rect 21131 56933 21143 56967
rect 21450 56964 21456 56976
rect 21411 56936 21456 56964
rect 21085 56927 21143 56933
rect 21450 56924 21456 56936
rect 21508 56924 21514 56976
rect 14185 56899 14243 56905
rect 14185 56865 14197 56899
rect 14231 56896 14243 56899
rect 14274 56896 14280 56908
rect 14231 56868 14280 56896
rect 14231 56865 14243 56868
rect 14185 56859 14243 56865
rect 14274 56856 14280 56868
rect 14332 56856 14338 56908
rect 15470 56856 15476 56908
rect 15528 56896 15534 56908
rect 15657 56899 15715 56905
rect 15657 56896 15669 56899
rect 15528 56868 15669 56896
rect 15528 56856 15534 56868
rect 15657 56865 15669 56868
rect 15703 56865 15715 56899
rect 15657 56859 15715 56865
rect 16482 56856 16488 56908
rect 16540 56896 16546 56908
rect 17037 56899 17095 56905
rect 17037 56896 17049 56899
rect 16540 56868 17049 56896
rect 16540 56856 16546 56868
rect 17037 56865 17049 56868
rect 17083 56896 17095 56899
rect 18049 56899 18107 56905
rect 18049 56896 18061 56899
rect 17083 56868 18061 56896
rect 17083 56865 17095 56868
rect 17037 56859 17095 56865
rect 18049 56865 18061 56868
rect 18095 56896 18107 56899
rect 18322 56896 18328 56908
rect 18095 56868 18328 56896
rect 18095 56865 18107 56868
rect 18049 56859 18107 56865
rect 18322 56856 18328 56868
rect 18380 56856 18386 56908
rect 19061 56899 19119 56905
rect 19061 56896 19073 56899
rect 18708 56868 19073 56896
rect 18708 56840 18736 56868
rect 19061 56865 19073 56868
rect 19107 56865 19119 56899
rect 20438 56896 20444 56908
rect 19061 56859 19119 56865
rect 19168 56868 20444 56896
rect 15381 56831 15439 56837
rect 15381 56828 15393 56831
rect 14016 56800 15393 56828
rect 14016 56704 14044 56800
rect 15381 56797 15393 56800
rect 15427 56797 15439 56831
rect 17862 56828 17868 56840
rect 17823 56800 17868 56828
rect 15381 56791 15439 56797
rect 17862 56788 17868 56800
rect 17920 56828 17926 56840
rect 18690 56828 18696 56840
rect 17920 56800 18696 56828
rect 17920 56788 17926 56800
rect 18690 56788 18696 56800
rect 18748 56788 18754 56840
rect 18966 56788 18972 56840
rect 19024 56828 19030 56840
rect 19168 56828 19196 56868
rect 20438 56856 20444 56868
rect 20496 56856 20502 56908
rect 21542 56856 21548 56908
rect 21600 56896 21606 56908
rect 22020 56905 22048 57004
rect 22649 57001 22661 57004
rect 22695 57001 22707 57035
rect 22830 57032 22836 57044
rect 22791 57004 22836 57032
rect 22649 56995 22707 57001
rect 22830 56992 22836 57004
rect 22888 56992 22894 57044
rect 26694 57032 26700 57044
rect 26655 57004 26700 57032
rect 26694 56992 26700 57004
rect 26752 56992 26758 57044
rect 27338 56924 27344 56976
rect 27396 56964 27402 56976
rect 28902 56964 28908 56976
rect 27396 56936 28908 56964
rect 27396 56924 27402 56936
rect 22005 56899 22063 56905
rect 22005 56896 22017 56899
rect 21600 56868 22017 56896
rect 21600 56856 21606 56868
rect 22005 56865 22017 56868
rect 22051 56865 22063 56899
rect 22005 56859 22063 56865
rect 22094 56856 22100 56908
rect 22152 56896 22158 56908
rect 22281 56899 22339 56905
rect 22281 56896 22293 56899
rect 22152 56868 22293 56896
rect 22152 56856 22158 56868
rect 22281 56865 22293 56868
rect 22327 56865 22339 56899
rect 22281 56859 22339 56865
rect 22649 56899 22707 56905
rect 22649 56865 22661 56899
rect 22695 56896 22707 56899
rect 22922 56896 22928 56908
rect 22695 56868 22928 56896
rect 22695 56865 22707 56868
rect 22649 56859 22707 56865
rect 22922 56856 22928 56868
rect 22980 56896 22986 56908
rect 23109 56899 23167 56905
rect 23109 56896 23121 56899
rect 22980 56868 23121 56896
rect 22980 56856 22986 56868
rect 23109 56865 23121 56868
rect 23155 56865 23167 56899
rect 23290 56896 23296 56908
rect 23251 56868 23296 56896
rect 23109 56859 23167 56865
rect 23290 56856 23296 56868
rect 23348 56856 23354 56908
rect 23474 56856 23480 56908
rect 23532 56896 23538 56908
rect 23661 56899 23719 56905
rect 23661 56896 23673 56899
rect 23532 56868 23673 56896
rect 23532 56856 23538 56868
rect 23661 56865 23673 56868
rect 23707 56865 23719 56899
rect 23661 56859 23719 56865
rect 24213 56899 24271 56905
rect 24213 56865 24225 56899
rect 24259 56896 24271 56899
rect 24259 56868 24716 56896
rect 24259 56865 24271 56868
rect 24213 56859 24271 56865
rect 24688 56840 24716 56868
rect 24854 56856 24860 56908
rect 24912 56896 24918 56908
rect 25225 56899 25283 56905
rect 25225 56896 25237 56899
rect 24912 56868 25237 56896
rect 24912 56856 24918 56868
rect 25225 56865 25237 56868
rect 25271 56865 25283 56899
rect 26510 56896 26516 56908
rect 26471 56868 26516 56896
rect 25225 56859 25283 56865
rect 26510 56856 26516 56868
rect 26568 56856 26574 56908
rect 27614 56856 27620 56908
rect 27672 56896 27678 56908
rect 28258 56896 28264 56908
rect 27672 56868 28264 56896
rect 27672 56856 27678 56868
rect 28258 56856 28264 56868
rect 28316 56896 28322 56908
rect 28828 56905 28856 56936
rect 28902 56924 28908 56936
rect 28960 56924 28966 56976
rect 28353 56899 28411 56905
rect 28353 56896 28365 56899
rect 28316 56868 28365 56896
rect 28316 56856 28322 56868
rect 28353 56865 28365 56868
rect 28399 56865 28411 56899
rect 28353 56859 28411 56865
rect 28813 56899 28871 56905
rect 28813 56865 28825 56899
rect 28859 56865 28871 56899
rect 28813 56859 28871 56865
rect 19426 56828 19432 56840
rect 19024 56800 19196 56828
rect 19387 56800 19432 56828
rect 19024 56788 19030 56800
rect 19426 56788 19432 56800
rect 19484 56788 19490 56840
rect 22465 56831 22523 56837
rect 22465 56797 22477 56831
rect 22511 56828 22523 56831
rect 22554 56828 22560 56840
rect 22511 56800 22560 56828
rect 22511 56797 22523 56800
rect 22465 56791 22523 56797
rect 22554 56788 22560 56800
rect 22612 56788 22618 56840
rect 24394 56828 24400 56840
rect 24355 56800 24400 56828
rect 24394 56788 24400 56800
rect 24452 56788 24458 56840
rect 24670 56788 24676 56840
rect 24728 56788 24734 56840
rect 27522 56788 27528 56840
rect 27580 56828 27586 56840
rect 27801 56831 27859 56837
rect 27801 56828 27813 56831
rect 27580 56800 27813 56828
rect 27580 56788 27586 56800
rect 27801 56797 27813 56800
rect 27847 56828 27859 56831
rect 28169 56831 28227 56837
rect 28169 56828 28181 56831
rect 27847 56800 28181 56828
rect 27847 56797 27859 56800
rect 27801 56791 27859 56797
rect 28169 56797 28181 56800
rect 28215 56828 28227 56831
rect 28626 56828 28632 56840
rect 28215 56800 28632 56828
rect 28215 56797 28227 56800
rect 28169 56791 28227 56797
rect 28626 56788 28632 56800
rect 28684 56788 28690 56840
rect 17494 56720 17500 56772
rect 17552 56760 17558 56772
rect 17589 56763 17647 56769
rect 17589 56760 17601 56763
rect 17552 56732 17601 56760
rect 17552 56720 17558 56732
rect 17589 56729 17601 56732
rect 17635 56760 17647 56763
rect 18138 56760 18144 56772
rect 17635 56732 18144 56760
rect 17635 56729 17647 56732
rect 17589 56723 17647 56729
rect 18138 56720 18144 56732
rect 18196 56720 18202 56772
rect 19334 56760 19340 56772
rect 19295 56732 19340 56760
rect 19334 56720 19340 56732
rect 19392 56720 19398 56772
rect 21082 56720 21088 56772
rect 21140 56760 21146 56772
rect 22002 56760 22008 56772
rect 21140 56732 22008 56760
rect 21140 56720 21146 56732
rect 22002 56720 22008 56732
rect 22060 56760 22066 56772
rect 25409 56763 25467 56769
rect 25409 56760 25421 56763
rect 22060 56732 25421 56760
rect 22060 56720 22066 56732
rect 25409 56729 25421 56732
rect 25455 56729 25467 56763
rect 25409 56723 25467 56729
rect 27433 56763 27491 56769
rect 27433 56729 27445 56763
rect 27479 56760 27491 56763
rect 28442 56760 28448 56772
rect 27479 56732 28448 56760
rect 27479 56729 27491 56732
rect 27433 56723 27491 56729
rect 28442 56720 28448 56732
rect 28500 56720 28506 56772
rect 28902 56760 28908 56772
rect 28863 56732 28908 56760
rect 28902 56720 28908 56732
rect 28960 56720 28966 56772
rect 13725 56695 13783 56701
rect 13725 56661 13737 56695
rect 13771 56692 13783 56695
rect 13998 56692 14004 56704
rect 13771 56664 14004 56692
rect 13771 56661 13783 56664
rect 13725 56655 13783 56661
rect 13998 56652 14004 56664
rect 14056 56652 14062 56704
rect 14369 56695 14427 56701
rect 14369 56661 14381 56695
rect 14415 56692 14427 56695
rect 14458 56692 14464 56704
rect 14415 56664 14464 56692
rect 14415 56661 14427 56664
rect 14369 56655 14427 56661
rect 14458 56652 14464 56664
rect 14516 56652 14522 56704
rect 14737 56695 14795 56701
rect 14737 56661 14749 56695
rect 14783 56692 14795 56695
rect 15010 56692 15016 56704
rect 14783 56664 15016 56692
rect 14783 56661 14795 56664
rect 14737 56655 14795 56661
rect 15010 56652 15016 56664
rect 15068 56652 15074 56704
rect 15105 56695 15163 56701
rect 15105 56661 15117 56695
rect 15151 56692 15163 56695
rect 16482 56692 16488 56704
rect 15151 56664 16488 56692
rect 15151 56661 15163 56664
rect 15105 56655 15163 56661
rect 16482 56652 16488 56664
rect 16540 56652 16546 56704
rect 19058 56652 19064 56704
rect 19116 56692 19122 56704
rect 19199 56695 19257 56701
rect 19199 56692 19211 56695
rect 19116 56664 19211 56692
rect 19116 56652 19122 56664
rect 19199 56661 19211 56664
rect 19245 56661 19257 56695
rect 19518 56692 19524 56704
rect 19479 56664 19524 56692
rect 19199 56655 19257 56661
rect 19518 56652 19524 56664
rect 19576 56652 19582 56704
rect 22370 56652 22376 56704
rect 22428 56692 22434 56704
rect 24673 56695 24731 56701
rect 24673 56692 24685 56695
rect 22428 56664 24685 56692
rect 22428 56652 22434 56664
rect 24673 56661 24685 56664
rect 24719 56692 24731 56695
rect 24762 56692 24768 56704
rect 24719 56664 24768 56692
rect 24719 56661 24731 56664
rect 24673 56655 24731 56661
rect 24762 56652 24768 56664
rect 24820 56652 24826 56704
rect 25130 56692 25136 56704
rect 25091 56664 25136 56692
rect 25130 56652 25136 56664
rect 25188 56652 25194 56704
rect 25498 56652 25504 56704
rect 25556 56692 25562 56704
rect 25685 56695 25743 56701
rect 25685 56692 25697 56695
rect 25556 56664 25697 56692
rect 25556 56652 25562 56664
rect 25685 56661 25697 56664
rect 25731 56661 25743 56695
rect 25685 56655 25743 56661
rect 25774 56652 25780 56704
rect 25832 56692 25838 56704
rect 26053 56695 26111 56701
rect 26053 56692 26065 56695
rect 25832 56664 26065 56692
rect 25832 56652 25838 56664
rect 26053 56661 26065 56664
rect 26099 56661 26111 56695
rect 26053 56655 26111 56661
rect 34606 56652 34612 56704
rect 34664 56692 34670 56704
rect 35250 56692 35256 56704
rect 34664 56664 35256 56692
rect 34664 56652 34670 56664
rect 35250 56652 35256 56664
rect 35308 56652 35314 56704
rect 1104 56602 38824 56624
rect 1104 56550 4246 56602
rect 4298 56550 4310 56602
rect 4362 56550 4374 56602
rect 4426 56550 4438 56602
rect 4490 56550 34966 56602
rect 35018 56550 35030 56602
rect 35082 56550 35094 56602
rect 35146 56550 35158 56602
rect 35210 56550 38824 56602
rect 1104 56528 38824 56550
rect 13262 56488 13268 56500
rect 13223 56460 13268 56488
rect 13262 56448 13268 56460
rect 13320 56448 13326 56500
rect 15746 56488 15752 56500
rect 15707 56460 15752 56488
rect 15746 56448 15752 56460
rect 15804 56448 15810 56500
rect 16853 56491 16911 56497
rect 16853 56457 16865 56491
rect 16899 56488 16911 56491
rect 17494 56488 17500 56500
rect 16899 56460 17500 56488
rect 16899 56457 16911 56460
rect 16853 56451 16911 56457
rect 17494 56448 17500 56460
rect 17552 56448 17558 56500
rect 17862 56488 17868 56500
rect 17823 56460 17868 56488
rect 17862 56448 17868 56460
rect 17920 56448 17926 56500
rect 18417 56491 18475 56497
rect 18417 56457 18429 56491
rect 18463 56488 18475 56491
rect 19426 56488 19432 56500
rect 18463 56460 19432 56488
rect 18463 56457 18475 56460
rect 18417 56451 18475 56457
rect 19426 56448 19432 56460
rect 19484 56448 19490 56500
rect 19518 56448 19524 56500
rect 19576 56488 19582 56500
rect 19797 56491 19855 56497
rect 19797 56488 19809 56491
rect 19576 56460 19809 56488
rect 19576 56448 19582 56460
rect 19797 56457 19809 56460
rect 19843 56488 19855 56491
rect 19978 56488 19984 56500
rect 19843 56460 19984 56488
rect 19843 56457 19855 56460
rect 19797 56451 19855 56457
rect 19978 56448 19984 56460
rect 20036 56448 20042 56500
rect 21358 56488 21364 56500
rect 21319 56460 21364 56488
rect 21358 56448 21364 56460
rect 21416 56448 21422 56500
rect 21450 56448 21456 56500
rect 21508 56488 21514 56500
rect 21545 56491 21603 56497
rect 21545 56488 21557 56491
rect 21508 56460 21557 56488
rect 21508 56448 21514 56460
rect 21545 56457 21557 56460
rect 21591 56457 21603 56491
rect 23290 56488 23296 56500
rect 23251 56460 23296 56488
rect 21545 56451 21603 56457
rect 23290 56448 23296 56460
rect 23348 56448 23354 56500
rect 27157 56491 27215 56497
rect 27157 56457 27169 56491
rect 27203 56488 27215 56491
rect 27338 56488 27344 56500
rect 27203 56460 27344 56488
rect 27203 56457 27215 56460
rect 27157 56451 27215 56457
rect 27338 56448 27344 56460
rect 27396 56448 27402 56500
rect 27522 56488 27528 56500
rect 27483 56460 27528 56488
rect 27522 56448 27528 56460
rect 27580 56448 27586 56500
rect 17129 56423 17187 56429
rect 17129 56389 17141 56423
rect 17175 56420 17187 56423
rect 18046 56420 18052 56432
rect 17175 56392 18052 56420
rect 17175 56389 17187 56392
rect 17129 56383 17187 56389
rect 18046 56380 18052 56392
rect 18104 56380 18110 56432
rect 18693 56423 18751 56429
rect 18693 56389 18705 56423
rect 18739 56420 18751 56423
rect 18966 56420 18972 56432
rect 18739 56392 18972 56420
rect 18739 56389 18751 56392
rect 18693 56383 18751 56389
rect 18966 56380 18972 56392
rect 19024 56380 19030 56432
rect 19061 56423 19119 56429
rect 19061 56389 19073 56423
rect 19107 56420 19119 56423
rect 19150 56420 19156 56432
rect 19107 56392 19156 56420
rect 19107 56389 19119 56392
rect 19061 56383 19119 56389
rect 19150 56380 19156 56392
rect 19208 56380 19214 56432
rect 19610 56380 19616 56432
rect 19668 56429 19674 56432
rect 19668 56423 19717 56429
rect 19668 56389 19671 56423
rect 19705 56420 19717 56423
rect 20254 56420 20260 56432
rect 19705 56392 20260 56420
rect 19705 56389 19717 56392
rect 19668 56383 19717 56389
rect 19668 56380 19674 56383
rect 20254 56380 20260 56392
rect 20312 56380 20318 56432
rect 20898 56420 20904 56432
rect 20640 56392 20904 56420
rect 14182 56352 14188 56364
rect 14143 56324 14188 56352
rect 14182 56312 14188 56324
rect 14240 56352 14246 56364
rect 14645 56355 14703 56361
rect 14645 56352 14657 56355
rect 14240 56324 14657 56352
rect 14240 56312 14246 56324
rect 14645 56321 14657 56324
rect 14691 56321 14703 56355
rect 14645 56315 14703 56321
rect 19334 56312 19340 56364
rect 19392 56352 19398 56364
rect 19889 56355 19947 56361
rect 19889 56352 19901 56355
rect 19392 56324 19901 56352
rect 19392 56312 19398 56324
rect 19889 56321 19901 56324
rect 19935 56352 19947 56355
rect 20533 56355 20591 56361
rect 20533 56352 20545 56355
rect 19935 56324 20545 56352
rect 19935 56321 19947 56324
rect 19889 56315 19947 56321
rect 20533 56321 20545 56324
rect 20579 56352 20591 56355
rect 20640 56352 20668 56392
rect 20898 56380 20904 56392
rect 20956 56380 20962 56432
rect 21250 56423 21308 56429
rect 21250 56420 21262 56423
rect 21008 56392 21262 56420
rect 21008 56352 21036 56392
rect 21250 56389 21262 56392
rect 21296 56420 21308 56423
rect 21910 56420 21916 56432
rect 21296 56392 21916 56420
rect 21296 56389 21308 56392
rect 21250 56383 21308 56389
rect 21910 56380 21916 56392
rect 21968 56380 21974 56432
rect 24857 56423 24915 56429
rect 24857 56389 24869 56423
rect 24903 56420 24915 56423
rect 24903 56392 26096 56420
rect 24903 56389 24915 56392
rect 24857 56383 24915 56389
rect 26068 56364 26096 56392
rect 21450 56352 21456 56364
rect 20579 56324 20668 56352
rect 20732 56324 21036 56352
rect 21411 56324 21456 56352
rect 20579 56321 20591 56324
rect 20533 56315 20591 56321
rect 13262 56244 13268 56296
rect 13320 56284 13326 56296
rect 13357 56287 13415 56293
rect 13357 56284 13369 56287
rect 13320 56256 13369 56284
rect 13320 56244 13326 56256
rect 13357 56253 13369 56256
rect 13403 56253 13415 56287
rect 13357 56247 13415 56253
rect 13998 56244 14004 56296
rect 14056 56284 14062 56296
rect 14369 56287 14427 56293
rect 14369 56284 14381 56287
rect 14056 56256 14381 56284
rect 14056 56244 14062 56256
rect 14369 56253 14381 56256
rect 14415 56253 14427 56287
rect 16945 56287 17003 56293
rect 16945 56284 16957 56287
rect 14369 56247 14427 56253
rect 14476 56256 16957 56284
rect 13909 56219 13967 56225
rect 13909 56185 13921 56219
rect 13955 56216 13967 56219
rect 14274 56216 14280 56228
rect 13955 56188 14280 56216
rect 13955 56185 13967 56188
rect 13909 56179 13967 56185
rect 14274 56176 14280 56188
rect 14332 56216 14338 56228
rect 14476 56216 14504 56256
rect 16945 56253 16957 56256
rect 16991 56284 17003 56287
rect 18509 56287 18567 56293
rect 16991 56256 17540 56284
rect 16991 56253 17003 56256
rect 16945 56247 17003 56253
rect 14332 56188 14504 56216
rect 14332 56176 14338 56188
rect 13538 56148 13544 56160
rect 13499 56120 13544 56148
rect 13538 56108 13544 56120
rect 13596 56108 13602 56160
rect 16485 56151 16543 56157
rect 16485 56117 16497 56151
rect 16531 56148 16543 56151
rect 17218 56148 17224 56160
rect 16531 56120 17224 56148
rect 16531 56117 16543 56120
rect 16485 56111 16543 56117
rect 17218 56108 17224 56120
rect 17276 56108 17282 56160
rect 17512 56157 17540 56256
rect 18509 56253 18521 56287
rect 18555 56253 18567 56287
rect 18509 56247 18567 56253
rect 19521 56287 19579 56293
rect 19521 56253 19533 56287
rect 19567 56284 19579 56287
rect 20162 56284 20168 56296
rect 19567 56256 20168 56284
rect 19567 56253 19579 56256
rect 19521 56247 19579 56253
rect 18322 56176 18328 56228
rect 18380 56216 18386 56228
rect 18524 56216 18552 56247
rect 20162 56244 20168 56256
rect 20220 56244 20226 56296
rect 20732 56216 20760 56324
rect 21450 56312 21456 56324
rect 21508 56312 21514 56364
rect 24946 56312 24952 56364
rect 25004 56352 25010 56364
rect 25225 56355 25283 56361
rect 25225 56352 25237 56355
rect 25004 56324 25237 56352
rect 25004 56312 25010 56324
rect 25225 56321 25237 56324
rect 25271 56321 25283 56355
rect 26050 56352 26056 56364
rect 26011 56324 26056 56352
rect 25225 56315 25283 56321
rect 26050 56312 26056 56324
rect 26108 56312 26114 56364
rect 28350 56352 28356 56364
rect 28311 56324 28356 56352
rect 28350 56312 28356 56324
rect 28408 56312 28414 56364
rect 21910 56244 21916 56296
rect 21968 56284 21974 56296
rect 22097 56287 22155 56293
rect 22097 56284 22109 56287
rect 21968 56256 22109 56284
rect 21968 56244 21974 56256
rect 22097 56253 22109 56256
rect 22143 56284 22155 56287
rect 22278 56284 22284 56296
rect 22143 56256 22284 56284
rect 22143 56253 22155 56256
rect 22097 56247 22155 56253
rect 22278 56244 22284 56256
rect 22336 56244 22342 56296
rect 23658 56284 23664 56296
rect 23619 56256 23664 56284
rect 23658 56244 23664 56256
rect 23716 56284 23722 56296
rect 24121 56287 24179 56293
rect 24121 56284 24133 56287
rect 23716 56256 24133 56284
rect 23716 56244 23722 56256
rect 24121 56253 24133 56256
rect 24167 56253 24179 56287
rect 25130 56284 25136 56296
rect 25091 56256 25136 56284
rect 24121 56247 24179 56253
rect 25130 56244 25136 56256
rect 25188 56244 25194 56296
rect 25314 56244 25320 56296
rect 25372 56284 25378 56296
rect 25774 56284 25780 56296
rect 25372 56256 25780 56284
rect 25372 56244 25378 56256
rect 25774 56244 25780 56256
rect 25832 56284 25838 56296
rect 25961 56287 26019 56293
rect 25961 56284 25973 56287
rect 25832 56256 25973 56284
rect 25832 56244 25838 56256
rect 25961 56253 25973 56256
rect 26007 56253 26019 56287
rect 27798 56284 27804 56296
rect 27759 56256 27804 56284
rect 25961 56247 26019 56253
rect 27798 56244 27804 56256
rect 27856 56244 27862 56296
rect 20898 56216 20904 56228
rect 18380 56188 20760 56216
rect 20859 56188 20904 56216
rect 18380 56176 18386 56188
rect 20898 56176 20904 56188
rect 20956 56176 20962 56228
rect 21085 56219 21143 56225
rect 21085 56185 21097 56219
rect 21131 56216 21143 56219
rect 21358 56216 21364 56228
rect 21131 56188 21364 56216
rect 21131 56185 21143 56188
rect 21085 56179 21143 56185
rect 21358 56176 21364 56188
rect 21416 56176 21422 56228
rect 25148 56216 25176 56244
rect 26326 56216 26332 56228
rect 25148 56188 26332 56216
rect 26326 56176 26332 56188
rect 26384 56176 26390 56228
rect 17497 56151 17555 56157
rect 17497 56117 17509 56151
rect 17543 56148 17555 56151
rect 17586 56148 17592 56160
rect 17543 56120 17592 56148
rect 17543 56117 17555 56120
rect 17497 56111 17555 56117
rect 17586 56108 17592 56120
rect 17644 56108 17650 56160
rect 19334 56148 19340 56160
rect 19295 56120 19340 56148
rect 19334 56108 19340 56120
rect 19392 56108 19398 56160
rect 19426 56108 19432 56160
rect 19484 56148 19490 56160
rect 20165 56151 20223 56157
rect 20165 56148 20177 56151
rect 19484 56120 20177 56148
rect 19484 56108 19490 56120
rect 20165 56117 20177 56120
rect 20211 56117 20223 56151
rect 20916 56148 20944 56176
rect 22094 56148 22100 56160
rect 20916 56120 22100 56148
rect 20165 56111 20223 56117
rect 22094 56108 22100 56120
rect 22152 56108 22158 56160
rect 22554 56148 22560 56160
rect 22515 56120 22560 56148
rect 22554 56108 22560 56120
rect 22612 56108 22618 56160
rect 23017 56151 23075 56157
rect 23017 56117 23029 56151
rect 23063 56148 23075 56151
rect 23474 56148 23480 56160
rect 23063 56120 23480 56148
rect 23063 56117 23075 56120
rect 23017 56111 23075 56117
rect 23474 56108 23480 56120
rect 23532 56108 23538 56160
rect 23842 56148 23848 56160
rect 23803 56120 23848 56148
rect 23842 56108 23848 56120
rect 23900 56108 23906 56160
rect 24486 56148 24492 56160
rect 24447 56120 24492 56148
rect 24486 56108 24492 56120
rect 24544 56148 24550 56160
rect 24762 56148 24768 56160
rect 24544 56120 24768 56148
rect 24544 56108 24550 56120
rect 24762 56108 24768 56120
rect 24820 56108 24826 56160
rect 26510 56148 26516 56160
rect 26471 56120 26516 56148
rect 26510 56108 26516 56120
rect 26568 56108 26574 56160
rect 28350 56108 28356 56160
rect 28408 56148 28414 56160
rect 28629 56151 28687 56157
rect 28629 56148 28641 56151
rect 28408 56120 28641 56148
rect 28408 56108 28414 56120
rect 28629 56117 28641 56120
rect 28675 56117 28687 56151
rect 28629 56111 28687 56117
rect 1104 56058 38824 56080
rect 1104 56006 19606 56058
rect 19658 56006 19670 56058
rect 19722 56006 19734 56058
rect 19786 56006 19798 56058
rect 19850 56006 38824 56058
rect 1104 55984 38824 56006
rect 14366 55944 14372 55956
rect 14327 55916 14372 55944
rect 14366 55904 14372 55916
rect 14424 55904 14430 55956
rect 17494 55944 17500 55956
rect 17455 55916 17500 55944
rect 17494 55904 17500 55916
rect 17552 55904 17558 55956
rect 18690 55944 18696 55956
rect 18651 55916 18696 55944
rect 18690 55904 18696 55916
rect 18748 55904 18754 55956
rect 19058 55944 19064 55956
rect 19019 55916 19064 55944
rect 19058 55904 19064 55916
rect 19116 55904 19122 55956
rect 20254 55944 20260 55956
rect 20215 55916 20260 55944
rect 20254 55904 20260 55916
rect 20312 55904 20318 55956
rect 22830 55904 22836 55956
rect 22888 55944 22894 55956
rect 24305 55947 24363 55953
rect 24305 55944 24317 55947
rect 22888 55916 24317 55944
rect 22888 55904 22894 55916
rect 24305 55913 24317 55916
rect 24351 55944 24363 55947
rect 24486 55944 24492 55956
rect 24351 55916 24492 55944
rect 24351 55913 24363 55916
rect 24305 55907 24363 55913
rect 24486 55904 24492 55916
rect 24544 55904 24550 55956
rect 26973 55947 27031 55953
rect 26973 55913 26985 55947
rect 27019 55944 27031 55947
rect 27062 55944 27068 55956
rect 27019 55916 27068 55944
rect 27019 55913 27031 55916
rect 26973 55907 27031 55913
rect 27062 55904 27068 55916
rect 27120 55904 27126 55956
rect 28534 55944 28540 55956
rect 28495 55916 28540 55944
rect 28534 55904 28540 55916
rect 28592 55904 28598 55956
rect 12710 55836 12716 55888
rect 12768 55876 12774 55888
rect 13725 55879 13783 55885
rect 13725 55876 13737 55879
rect 12768 55848 13737 55876
rect 12768 55836 12774 55848
rect 13725 55845 13737 55848
rect 13771 55876 13783 55879
rect 15010 55876 15016 55888
rect 13771 55848 15016 55876
rect 13771 55845 13783 55848
rect 13725 55839 13783 55845
rect 15010 55836 15016 55848
rect 15068 55876 15074 55888
rect 16117 55879 16175 55885
rect 16117 55876 16129 55879
rect 15068 55848 16129 55876
rect 15068 55836 15074 55848
rect 16117 55845 16129 55848
rect 16163 55876 16175 55879
rect 19978 55876 19984 55888
rect 16163 55848 19104 55876
rect 19939 55848 19984 55876
rect 16163 55845 16175 55848
rect 16117 55839 16175 55845
rect 19076 55820 19104 55848
rect 19978 55836 19984 55848
rect 20036 55836 20042 55888
rect 12161 55811 12219 55817
rect 12161 55777 12173 55811
rect 12207 55808 12219 55811
rect 12250 55808 12256 55820
rect 12207 55780 12256 55808
rect 12207 55777 12219 55780
rect 12161 55771 12219 55777
rect 12250 55768 12256 55780
rect 12308 55768 12314 55820
rect 13170 55808 13176 55820
rect 13131 55780 13176 55808
rect 13170 55768 13176 55780
rect 13228 55768 13234 55820
rect 14185 55811 14243 55817
rect 14185 55777 14197 55811
rect 14231 55808 14243 55811
rect 14826 55808 14832 55820
rect 14231 55780 14832 55808
rect 14231 55777 14243 55780
rect 14185 55771 14243 55777
rect 14826 55768 14832 55780
rect 14884 55768 14890 55820
rect 16850 55808 16856 55820
rect 16811 55780 16856 55808
rect 16850 55768 16856 55780
rect 16908 55768 16914 55820
rect 18322 55808 18328 55820
rect 18283 55780 18328 55808
rect 18322 55768 18328 55780
rect 18380 55768 18386 55820
rect 19058 55768 19064 55820
rect 19116 55808 19122 55820
rect 19245 55811 19303 55817
rect 19245 55808 19257 55811
rect 19116 55780 19257 55808
rect 19116 55768 19122 55780
rect 19245 55777 19257 55780
rect 19291 55777 19303 55811
rect 19245 55771 19303 55777
rect 20714 55768 20720 55820
rect 20772 55808 20778 55820
rect 20901 55811 20959 55817
rect 20901 55808 20913 55811
rect 20772 55780 20913 55808
rect 20772 55768 20778 55780
rect 20901 55777 20913 55780
rect 20947 55777 20959 55811
rect 21082 55808 21088 55820
rect 21043 55780 21088 55808
rect 20901 55771 20959 55777
rect 21082 55768 21088 55780
rect 21140 55768 21146 55820
rect 22922 55808 22928 55820
rect 22883 55780 22928 55808
rect 22922 55768 22928 55780
rect 22980 55768 22986 55820
rect 23106 55768 23112 55820
rect 23164 55808 23170 55820
rect 23201 55811 23259 55817
rect 23201 55808 23213 55811
rect 23164 55780 23213 55808
rect 23164 55768 23170 55780
rect 23201 55777 23213 55780
rect 23247 55777 23259 55811
rect 23201 55771 23259 55777
rect 23934 55768 23940 55820
rect 23992 55808 23998 55820
rect 24213 55811 24271 55817
rect 24213 55808 24225 55811
rect 23992 55780 24225 55808
rect 23992 55768 23998 55780
rect 24213 55777 24225 55780
rect 24259 55777 24271 55811
rect 24946 55808 24952 55820
rect 24907 55780 24952 55808
rect 24213 55771 24271 55777
rect 24946 55768 24952 55780
rect 25004 55768 25010 55820
rect 25225 55811 25283 55817
rect 25225 55777 25237 55811
rect 25271 55808 25283 55811
rect 25590 55808 25596 55820
rect 25271 55780 25596 55808
rect 25271 55777 25283 55780
rect 25225 55771 25283 55777
rect 13630 55700 13636 55752
rect 13688 55740 13694 55752
rect 15470 55740 15476 55752
rect 13688 55712 14136 55740
rect 15431 55712 15476 55740
rect 13688 55700 13694 55712
rect 14108 55681 14136 55712
rect 15470 55700 15476 55712
rect 15528 55700 15534 55752
rect 16485 55743 16543 55749
rect 16485 55709 16497 55743
rect 16531 55740 16543 55743
rect 16942 55740 16948 55752
rect 16531 55712 16948 55740
rect 16531 55709 16543 55712
rect 16485 55703 16543 55709
rect 16942 55700 16948 55712
rect 17000 55700 17006 55752
rect 17218 55740 17224 55752
rect 17179 55712 17224 55740
rect 17218 55700 17224 55712
rect 17276 55700 17282 55752
rect 18414 55740 18420 55752
rect 18327 55712 18420 55740
rect 18414 55700 18420 55712
rect 18472 55740 18478 55752
rect 18472 55712 19288 55740
rect 18472 55700 18478 55712
rect 14093 55675 14151 55681
rect 14093 55641 14105 55675
rect 14139 55672 14151 55675
rect 14139 55644 15608 55672
rect 14139 55641 14151 55644
rect 14093 55635 14151 55641
rect 12345 55607 12403 55613
rect 12345 55573 12357 55607
rect 12391 55604 12403 55607
rect 12434 55604 12440 55616
rect 12391 55576 12440 55604
rect 12391 55573 12403 55576
rect 12345 55567 12403 55573
rect 12434 55564 12440 55576
rect 12492 55564 12498 55616
rect 13357 55607 13415 55613
rect 13357 55573 13369 55607
rect 13403 55604 13415 55607
rect 13446 55604 13452 55616
rect 13403 55576 13452 55604
rect 13403 55573 13415 55576
rect 13357 55567 13415 55573
rect 13446 55564 13452 55576
rect 13504 55564 13510 55616
rect 13906 55564 13912 55616
rect 13964 55604 13970 55616
rect 14921 55607 14979 55613
rect 14921 55604 14933 55607
rect 13964 55576 14933 55604
rect 13964 55564 13970 55576
rect 14921 55573 14933 55576
rect 14967 55604 14979 55607
rect 15010 55604 15016 55616
rect 14967 55576 15016 55604
rect 14967 55573 14979 55576
rect 14921 55567 14979 55573
rect 15010 55564 15016 55576
rect 15068 55564 15074 55616
rect 15580 55604 15608 55644
rect 15654 55632 15660 55684
rect 15712 55672 15718 55684
rect 16022 55672 16028 55684
rect 15712 55644 16028 55672
rect 15712 55632 15718 55644
rect 16022 55632 16028 55644
rect 16080 55672 16086 55684
rect 16393 55675 16451 55681
rect 16393 55672 16405 55675
rect 16080 55644 16405 55672
rect 16080 55632 16086 55644
rect 16393 55641 16405 55644
rect 16439 55672 16451 55675
rect 19150 55672 19156 55684
rect 16439 55644 19156 55672
rect 16439 55641 16451 55644
rect 16393 55635 16451 55641
rect 19150 55632 19156 55644
rect 19208 55632 19214 55684
rect 19260 55672 19288 55712
rect 19334 55700 19340 55752
rect 19392 55740 19398 55752
rect 19613 55743 19671 55749
rect 19613 55740 19625 55743
rect 19392 55712 19625 55740
rect 19392 55700 19398 55712
rect 19613 55709 19625 55712
rect 19659 55709 19671 55743
rect 19613 55703 19671 55709
rect 21174 55700 21180 55752
rect 21232 55740 21238 55752
rect 21729 55743 21787 55749
rect 21729 55740 21741 55743
rect 21232 55712 21741 55740
rect 21232 55700 21238 55712
rect 21729 55709 21741 55712
rect 21775 55709 21787 55743
rect 21729 55703 21787 55709
rect 22373 55743 22431 55749
rect 22373 55709 22385 55743
rect 22419 55740 22431 55743
rect 22462 55740 22468 55752
rect 22419 55712 22468 55740
rect 22419 55709 22431 55712
rect 22373 55703 22431 55709
rect 22462 55700 22468 55712
rect 22520 55700 22526 55752
rect 23385 55743 23443 55749
rect 23385 55740 23397 55743
rect 23308 55712 23397 55740
rect 20254 55672 20260 55684
rect 19260 55644 20260 55672
rect 16282 55607 16340 55613
rect 16282 55604 16294 55607
rect 15580 55576 16294 55604
rect 16282 55573 16294 55576
rect 16328 55604 16340 55607
rect 16482 55604 16488 55616
rect 16328 55576 16488 55604
rect 16328 55573 16340 55576
rect 16282 55567 16340 55573
rect 16482 55564 16488 55576
rect 16540 55564 16546 55616
rect 19444 55613 19472 55644
rect 20254 55632 20260 55644
rect 20312 55632 20318 55684
rect 23308 55616 23336 55712
rect 23385 55709 23397 55712
rect 23431 55709 23443 55743
rect 23385 55703 23443 55709
rect 24121 55743 24179 55749
rect 24121 55709 24133 55743
rect 24167 55740 24179 55743
rect 25240 55740 25268 55771
rect 25590 55768 25596 55780
rect 25648 55768 25654 55820
rect 26605 55811 26663 55817
rect 26605 55777 26617 55811
rect 26651 55777 26663 55811
rect 28258 55808 28264 55820
rect 28219 55780 28264 55808
rect 26605 55771 26663 55777
rect 24167 55712 25268 55740
rect 24167 55709 24179 55712
rect 24121 55703 24179 55709
rect 26510 55700 26516 55752
rect 26568 55740 26574 55752
rect 26620 55740 26648 55771
rect 28258 55768 28264 55780
rect 28316 55768 28322 55820
rect 33137 55811 33195 55817
rect 33137 55777 33149 55811
rect 33183 55808 33195 55811
rect 33226 55808 33232 55820
rect 33183 55780 33232 55808
rect 33183 55777 33195 55780
rect 33137 55771 33195 55777
rect 33226 55768 33232 55780
rect 33284 55808 33290 55820
rect 34422 55808 34428 55820
rect 33284 55780 34428 55808
rect 33284 55768 33290 55780
rect 34422 55768 34428 55780
rect 34480 55768 34486 55820
rect 26568 55712 26648 55740
rect 32861 55743 32919 55749
rect 26568 55700 26574 55712
rect 32861 55709 32873 55743
rect 32907 55740 32919 55743
rect 33594 55740 33600 55752
rect 32907 55712 33600 55740
rect 32907 55709 32919 55712
rect 32861 55703 32919 55709
rect 33594 55700 33600 55712
rect 33652 55740 33658 55752
rect 34606 55740 34612 55752
rect 33652 55712 34612 55740
rect 33652 55700 33658 55712
rect 34606 55700 34612 55712
rect 34664 55700 34670 55752
rect 19410 55607 19472 55613
rect 19410 55573 19422 55607
rect 19456 55576 19472 55607
rect 19456 55573 19468 55576
rect 19410 55567 19468 55573
rect 19518 55564 19524 55616
rect 19576 55604 19582 55616
rect 20714 55604 20720 55616
rect 19576 55576 19621 55604
rect 20675 55576 20720 55604
rect 19576 55564 19582 55576
rect 20714 55564 20720 55576
rect 20772 55564 20778 55616
rect 20990 55564 20996 55616
rect 21048 55604 21054 55616
rect 21177 55607 21235 55613
rect 21177 55604 21189 55607
rect 21048 55576 21189 55604
rect 21048 55564 21054 55576
rect 21177 55573 21189 55576
rect 21223 55573 21235 55607
rect 21177 55567 21235 55573
rect 22281 55607 22339 55613
rect 22281 55573 22293 55607
rect 22327 55604 22339 55607
rect 22554 55604 22560 55616
rect 22327 55576 22560 55604
rect 22327 55573 22339 55576
rect 22281 55567 22339 55573
rect 22554 55564 22560 55576
rect 22612 55604 22618 55616
rect 23290 55604 23296 55616
rect 22612 55576 23296 55604
rect 22612 55564 22618 55576
rect 23290 55564 23296 55576
rect 23348 55564 23354 55616
rect 23658 55604 23664 55616
rect 23619 55576 23664 55604
rect 23658 55564 23664 55576
rect 23716 55564 23722 55616
rect 24854 55564 24860 55616
rect 24912 55604 24918 55616
rect 25593 55607 25651 55613
rect 25593 55604 25605 55607
rect 24912 55576 25605 55604
rect 24912 55564 24918 55576
rect 25593 55573 25605 55576
rect 25639 55573 25651 55607
rect 25593 55567 25651 55573
rect 25774 55564 25780 55616
rect 25832 55604 25838 55616
rect 25961 55607 26019 55613
rect 25961 55604 25973 55607
rect 25832 55576 25973 55604
rect 25832 55564 25838 55576
rect 25961 55573 25973 55576
rect 26007 55573 26019 55607
rect 25961 55567 26019 55573
rect 27709 55607 27767 55613
rect 27709 55573 27721 55607
rect 27755 55604 27767 55607
rect 27798 55604 27804 55616
rect 27755 55576 27804 55604
rect 27755 55573 27767 55576
rect 27709 55567 27767 55573
rect 27798 55564 27804 55576
rect 27856 55564 27862 55616
rect 31849 55607 31907 55613
rect 31849 55573 31861 55607
rect 31895 55604 31907 55607
rect 32674 55604 32680 55616
rect 31895 55576 32680 55604
rect 31895 55573 31907 55576
rect 31849 55567 31907 55573
rect 32674 55564 32680 55576
rect 32732 55604 32738 55616
rect 34241 55607 34299 55613
rect 34241 55604 34253 55607
rect 32732 55576 34253 55604
rect 32732 55564 32738 55576
rect 34241 55573 34253 55576
rect 34287 55573 34299 55607
rect 34241 55567 34299 55573
rect 1104 55514 38824 55536
rect 1104 55462 4246 55514
rect 4298 55462 4310 55514
rect 4362 55462 4374 55514
rect 4426 55462 4438 55514
rect 4490 55462 34966 55514
rect 35018 55462 35030 55514
rect 35082 55462 35094 55514
rect 35146 55462 35158 55514
rect 35210 55462 38824 55514
rect 1104 55440 38824 55462
rect 12250 55400 12256 55412
rect 12211 55372 12256 55400
rect 12250 55360 12256 55372
rect 12308 55360 12314 55412
rect 12710 55400 12716 55412
rect 12671 55372 12716 55400
rect 12710 55360 12716 55372
rect 12768 55360 12774 55412
rect 13906 55360 13912 55412
rect 13964 55400 13970 55412
rect 14001 55403 14059 55409
rect 14001 55400 14013 55403
rect 13964 55372 14013 55400
rect 13964 55360 13970 55372
rect 14001 55369 14013 55372
rect 14047 55369 14059 55403
rect 14001 55363 14059 55369
rect 14093 55403 14151 55409
rect 14093 55369 14105 55403
rect 14139 55400 14151 55403
rect 14369 55403 14427 55409
rect 14369 55400 14381 55403
rect 14139 55372 14381 55400
rect 14139 55369 14151 55372
rect 14093 55363 14151 55369
rect 14369 55369 14381 55372
rect 14415 55400 14427 55403
rect 14642 55400 14648 55412
rect 14415 55372 14648 55400
rect 14415 55369 14427 55372
rect 14369 55363 14427 55369
rect 14642 55360 14648 55372
rect 14700 55360 14706 55412
rect 15105 55403 15163 55409
rect 15105 55369 15117 55403
rect 15151 55400 15163 55403
rect 15470 55400 15476 55412
rect 15151 55372 15476 55400
rect 15151 55369 15163 55372
rect 15105 55363 15163 55369
rect 15470 55360 15476 55372
rect 15528 55400 15534 55412
rect 16758 55400 16764 55412
rect 15528 55372 16764 55400
rect 15528 55360 15534 55372
rect 16758 55360 16764 55372
rect 16816 55360 16822 55412
rect 16942 55360 16948 55412
rect 17000 55400 17006 55412
rect 17773 55403 17831 55409
rect 17773 55400 17785 55403
rect 17000 55372 17785 55400
rect 17000 55360 17006 55372
rect 17773 55369 17785 55372
rect 17819 55369 17831 55403
rect 17773 55363 17831 55369
rect 19797 55403 19855 55409
rect 19797 55369 19809 55403
rect 19843 55400 19855 55403
rect 20162 55400 20168 55412
rect 19843 55372 20168 55400
rect 19843 55369 19855 55372
rect 19797 55363 19855 55369
rect 20162 55360 20168 55372
rect 20220 55360 20226 55412
rect 22830 55360 22836 55412
rect 22888 55400 22894 55412
rect 23017 55403 23075 55409
rect 23017 55400 23029 55403
rect 22888 55372 23029 55400
rect 22888 55360 22894 55372
rect 23017 55369 23029 55372
rect 23063 55369 23075 55403
rect 23017 55363 23075 55369
rect 24946 55360 24952 55412
rect 25004 55400 25010 55412
rect 25041 55403 25099 55409
rect 25041 55400 25053 55403
rect 25004 55372 25053 55400
rect 25004 55360 25010 55372
rect 25041 55369 25053 55372
rect 25087 55369 25099 55403
rect 33226 55400 33232 55412
rect 33187 55372 33232 55400
rect 25041 55363 25099 55369
rect 33226 55360 33232 55372
rect 33284 55360 33290 55412
rect 15010 55341 15016 55344
rect 13357 55335 13415 55341
rect 13357 55332 13369 55335
rect 12820 55304 13369 55332
rect 12342 55224 12348 55276
rect 12400 55264 12406 55276
rect 12526 55264 12532 55276
rect 12400 55236 12532 55264
rect 12400 55224 12406 55236
rect 12526 55224 12532 55236
rect 12584 55224 12590 55276
rect 12820 55205 12848 55304
rect 13357 55301 13369 55304
rect 13403 55332 13415 55335
rect 14994 55335 15016 55341
rect 13403 55304 14504 55332
rect 13403 55301 13415 55304
rect 13357 55295 13415 55301
rect 14476 55276 14504 55304
rect 14994 55301 15006 55335
rect 14994 55295 15016 55301
rect 15010 55292 15016 55295
rect 15068 55292 15074 55344
rect 15902 55304 16712 55332
rect 13170 55224 13176 55276
rect 13228 55264 13234 55276
rect 13725 55267 13783 55273
rect 13725 55264 13737 55267
rect 13228 55236 13737 55264
rect 13228 55224 13234 55236
rect 13725 55233 13737 55236
rect 13771 55264 13783 55267
rect 13771 55236 13952 55264
rect 13771 55233 13783 55236
rect 13725 55227 13783 55233
rect 12805 55199 12863 55205
rect 12805 55165 12817 55199
rect 12851 55165 12863 55199
rect 12805 55159 12863 55165
rect 13817 55199 13875 55205
rect 13817 55165 13829 55199
rect 13863 55165 13875 55199
rect 13924 55196 13952 55236
rect 14458 55224 14464 55276
rect 14516 55264 14522 55276
rect 14737 55267 14795 55273
rect 14737 55264 14749 55267
rect 14516 55236 14749 55264
rect 14516 55224 14522 55236
rect 14737 55233 14749 55236
rect 14783 55264 14795 55267
rect 15197 55267 15255 55273
rect 15197 55264 15209 55267
rect 14783 55236 15209 55264
rect 14783 55233 14795 55236
rect 14737 55227 14795 55233
rect 15197 55233 15209 55236
rect 15243 55233 15255 55267
rect 15197 55227 15255 55233
rect 14182 55196 14188 55208
rect 13924 55168 14188 55196
rect 13817 55159 13875 55165
rect 13832 55128 13860 55159
rect 14182 55156 14188 55168
rect 14240 55196 14246 55208
rect 15102 55196 15108 55208
rect 14240 55168 15108 55196
rect 14240 55156 14246 55168
rect 15102 55156 15108 55168
rect 15160 55156 15166 55208
rect 15212 55196 15240 55227
rect 15902 55208 15930 55304
rect 15286 55196 15292 55208
rect 15212 55168 15292 55196
rect 15286 55156 15292 55168
rect 15344 55156 15350 55208
rect 15902 55168 15936 55208
rect 15930 55156 15936 55168
rect 15988 55196 15994 55208
rect 16209 55199 16267 55205
rect 16209 55196 16221 55199
rect 15988 55168 16221 55196
rect 15988 55156 15994 55168
rect 16209 55165 16221 55168
rect 16255 55165 16267 55199
rect 16684 55196 16712 55304
rect 24210 55292 24216 55344
rect 24268 55332 24274 55344
rect 24489 55335 24547 55341
rect 24489 55332 24501 55335
rect 24268 55304 24501 55332
rect 24268 55292 24274 55304
rect 24489 55301 24501 55304
rect 24535 55301 24547 55335
rect 24489 55295 24547 55301
rect 26329 55335 26387 55341
rect 26329 55301 26341 55335
rect 26375 55332 26387 55335
rect 26510 55332 26516 55344
rect 26375 55304 26516 55332
rect 26375 55301 26387 55304
rect 26329 55295 26387 55301
rect 26510 55292 26516 55304
rect 26568 55292 26574 55344
rect 17129 55267 17187 55273
rect 17129 55233 17141 55267
rect 17175 55264 17187 55267
rect 17862 55264 17868 55276
rect 17175 55236 17868 55264
rect 17175 55233 17187 55236
rect 17129 55227 17187 55233
rect 17862 55224 17868 55236
rect 17920 55224 17926 55276
rect 20165 55267 20223 55273
rect 20165 55233 20177 55267
rect 20211 55264 20223 55267
rect 20254 55264 20260 55276
rect 20211 55236 20260 55264
rect 20211 55233 20223 55236
rect 20165 55227 20223 55233
rect 20254 55224 20260 55236
rect 20312 55224 20318 55276
rect 20714 55224 20720 55276
rect 20772 55264 20778 55276
rect 21082 55264 21088 55276
rect 20772 55236 21088 55264
rect 20772 55224 20778 55236
rect 21082 55224 21088 55236
rect 21140 55264 21146 55276
rect 21637 55267 21695 55273
rect 21637 55264 21649 55267
rect 21140 55236 21649 55264
rect 21140 55224 21146 55236
rect 21637 55233 21649 55236
rect 21683 55264 21695 55267
rect 22373 55267 22431 55273
rect 22373 55264 22385 55267
rect 21683 55236 22385 55264
rect 21683 55233 21695 55236
rect 21637 55227 21695 55233
rect 22373 55233 22385 55236
rect 22419 55264 22431 55267
rect 22649 55267 22707 55273
rect 22649 55264 22661 55267
rect 22419 55236 22661 55264
rect 22419 55233 22431 55236
rect 22373 55227 22431 55233
rect 22649 55233 22661 55236
rect 22695 55233 22707 55267
rect 22649 55227 22707 55233
rect 25593 55267 25651 55273
rect 25593 55233 25605 55267
rect 25639 55264 25651 55267
rect 26234 55264 26240 55276
rect 25639 55236 26240 55264
rect 25639 55233 25651 55236
rect 25593 55227 25651 55233
rect 26234 55224 26240 55236
rect 26292 55264 26298 55276
rect 28258 55264 28264 55276
rect 26292 55236 26556 55264
rect 26292 55224 26298 55236
rect 16745 55199 16803 55205
rect 16745 55196 16757 55199
rect 16684 55168 16757 55196
rect 16209 55159 16267 55165
rect 16745 55165 16757 55168
rect 16791 55165 16803 55199
rect 16745 55159 16803 55165
rect 18693 55199 18751 55205
rect 18693 55165 18705 55199
rect 18739 55196 18751 55199
rect 19058 55196 19064 55208
rect 18739 55168 19064 55196
rect 18739 55165 18751 55168
rect 18693 55159 18751 55165
rect 19058 55156 19064 55168
rect 19116 55196 19122 55208
rect 19610 55196 19616 55208
rect 19116 55168 19616 55196
rect 19116 55156 19122 55168
rect 19610 55156 19616 55168
rect 19668 55156 19674 55208
rect 21174 55196 21180 55208
rect 21135 55168 21180 55196
rect 21174 55156 21180 55168
rect 21232 55156 21238 55208
rect 21729 55199 21787 55205
rect 21729 55165 21741 55199
rect 21775 55165 21787 55199
rect 23658 55196 23664 55208
rect 23619 55168 23664 55196
rect 21729 55159 21787 55165
rect 14093 55131 14151 55137
rect 14093 55128 14105 55131
rect 13832 55100 14105 55128
rect 14093 55097 14105 55100
rect 14139 55097 14151 55131
rect 14826 55128 14832 55140
rect 14787 55100 14832 55128
rect 14093 55091 14151 55097
rect 14826 55088 14832 55100
rect 14884 55088 14890 55140
rect 15565 55131 15623 55137
rect 15565 55097 15577 55131
rect 15611 55128 15623 55131
rect 16114 55128 16120 55140
rect 15611 55100 16120 55128
rect 15611 55097 15623 55100
rect 15565 55091 15623 55097
rect 16114 55088 16120 55100
rect 16172 55088 16178 55140
rect 16393 55131 16451 55137
rect 16393 55097 16405 55131
rect 16439 55097 16451 55131
rect 18046 55128 18052 55140
rect 18007 55100 18052 55128
rect 16393 55091 16451 55097
rect 12989 55063 13047 55069
rect 12989 55029 13001 55063
rect 13035 55060 13047 55063
rect 15194 55060 15200 55072
rect 13035 55032 15200 55060
rect 13035 55029 13047 55032
rect 12989 55023 13047 55029
rect 15194 55020 15200 55032
rect 15252 55060 15258 55072
rect 15841 55063 15899 55069
rect 15841 55060 15853 55063
rect 15252 55032 15853 55060
rect 15252 55020 15258 55032
rect 15841 55029 15853 55032
rect 15887 55060 15899 55063
rect 16408 55060 16436 55091
rect 18046 55088 18052 55100
rect 18104 55088 18110 55140
rect 21082 55088 21088 55140
rect 21140 55128 21146 55140
rect 21744 55128 21772 55159
rect 23658 55156 23664 55168
rect 23716 55156 23722 55208
rect 23842 55156 23848 55208
rect 23900 55196 23906 55208
rect 24029 55199 24087 55205
rect 24029 55196 24041 55199
rect 23900 55168 24041 55196
rect 23900 55156 23906 55168
rect 24029 55165 24041 55168
rect 24075 55165 24087 55199
rect 24486 55196 24492 55208
rect 24447 55168 24492 55196
rect 24029 55159 24087 55165
rect 24486 55156 24492 55168
rect 24544 55156 24550 55208
rect 26421 55199 26479 55205
rect 26421 55165 26433 55199
rect 26467 55165 26479 55199
rect 26528 55196 26556 55236
rect 27540 55236 28264 55264
rect 26881 55199 26939 55205
rect 26881 55196 26893 55199
rect 26528 55168 26893 55196
rect 26421 55159 26479 55165
rect 26881 55165 26893 55168
rect 26927 55165 26939 55199
rect 27540 55196 27568 55236
rect 28258 55224 28264 55236
rect 28316 55264 28322 55276
rect 28445 55267 28503 55273
rect 28445 55264 28457 55267
rect 28316 55236 28457 55264
rect 28316 55224 28322 55236
rect 28445 55233 28457 55236
rect 28491 55233 28503 55267
rect 31570 55264 31576 55276
rect 31531 55236 31576 55264
rect 28445 55227 28503 55233
rect 31570 55224 31576 55236
rect 31628 55264 31634 55276
rect 31849 55267 31907 55273
rect 31849 55264 31861 55267
rect 31628 55236 31861 55264
rect 31628 55224 31634 55236
rect 31849 55233 31861 55236
rect 31895 55233 31907 55267
rect 32769 55267 32827 55273
rect 32769 55264 32781 55267
rect 31849 55227 31907 55233
rect 31956 55236 32781 55264
rect 27982 55196 27988 55208
rect 26881 55159 26939 55165
rect 27172 55168 27568 55196
rect 27943 55168 27988 55196
rect 21140 55100 21772 55128
rect 25961 55131 26019 55137
rect 21140 55088 21146 55100
rect 25961 55097 25973 55131
rect 26007 55128 26019 55131
rect 26436 55128 26464 55159
rect 26602 55128 26608 55140
rect 26007 55100 26608 55128
rect 26007 55097 26019 55100
rect 25961 55091 26019 55097
rect 26602 55088 26608 55100
rect 26660 55128 26666 55140
rect 27172 55128 27200 55168
rect 27982 55156 27988 55168
rect 28040 55196 28046 55208
rect 28813 55199 28871 55205
rect 28813 55196 28825 55199
rect 28040 55168 28825 55196
rect 28040 55156 28046 55168
rect 28813 55165 28825 55168
rect 28859 55165 28871 55199
rect 28813 55159 28871 55165
rect 31754 55156 31760 55208
rect 31812 55196 31818 55208
rect 31956 55196 31984 55236
rect 32769 55233 32781 55236
rect 32815 55233 32827 55267
rect 33594 55264 33600 55276
rect 33555 55236 33600 55264
rect 32769 55227 32827 55233
rect 33594 55224 33600 55236
rect 33652 55224 33658 55276
rect 32674 55196 32680 55208
rect 31812 55168 31984 55196
rect 32635 55168 32680 55196
rect 31812 55156 31818 55168
rect 32674 55156 32680 55168
rect 32732 55156 32738 55208
rect 31938 55128 31944 55140
rect 26660 55100 27200 55128
rect 31899 55100 31944 55128
rect 26660 55088 26666 55100
rect 31938 55088 31944 55100
rect 31996 55088 32002 55140
rect 16574 55060 16580 55072
rect 15887 55032 16436 55060
rect 16535 55032 16580 55060
rect 15887 55029 15899 55032
rect 15841 55023 15899 55029
rect 16574 55020 16580 55032
rect 16632 55020 16638 55072
rect 16669 55063 16727 55069
rect 16669 55029 16681 55063
rect 16715 55060 16727 55063
rect 17494 55060 17500 55072
rect 16715 55032 17500 55060
rect 16715 55029 16727 55032
rect 16669 55023 16727 55029
rect 17494 55020 17500 55032
rect 17552 55020 17558 55072
rect 19334 55060 19340 55072
rect 19295 55032 19340 55060
rect 19334 55020 19340 55032
rect 19392 55020 19398 55072
rect 19426 55020 19432 55072
rect 19484 55060 19490 55072
rect 20438 55060 20444 55072
rect 19484 55032 20444 55060
rect 19484 55020 19490 55032
rect 20438 55020 20444 55032
rect 20496 55020 20502 55072
rect 21634 55020 21640 55072
rect 21692 55060 21698 55072
rect 21821 55063 21879 55069
rect 21821 55060 21833 55063
rect 21692 55032 21833 55060
rect 21692 55020 21698 55032
rect 21821 55029 21833 55032
rect 21867 55029 21879 55063
rect 21821 55023 21879 55029
rect 23477 55063 23535 55069
rect 23477 55029 23489 55063
rect 23523 55060 23535 55063
rect 23934 55060 23940 55072
rect 23523 55032 23940 55060
rect 23523 55029 23535 55032
rect 23477 55023 23535 55029
rect 23934 55020 23940 55032
rect 23992 55020 23998 55072
rect 26326 55020 26332 55072
rect 26384 55060 26390 55072
rect 26513 55063 26571 55069
rect 26513 55060 26525 55063
rect 26384 55032 26525 55060
rect 26384 55020 26390 55032
rect 26513 55029 26525 55032
rect 26559 55029 26571 55063
rect 26513 55023 26571 55029
rect 26786 55020 26792 55072
rect 26844 55060 26850 55072
rect 28169 55063 28227 55069
rect 28169 55060 28181 55063
rect 26844 55032 28181 55060
rect 26844 55020 26850 55032
rect 28169 55029 28181 55032
rect 28215 55029 28227 55063
rect 28169 55023 28227 55029
rect 1104 54970 38824 54992
rect 1104 54918 19606 54970
rect 19658 54918 19670 54970
rect 19722 54918 19734 54970
rect 19786 54918 19798 54970
rect 19850 54918 38824 54970
rect 1104 54896 38824 54918
rect 13630 54856 13636 54868
rect 13591 54828 13636 54856
rect 13630 54816 13636 54828
rect 13688 54816 13694 54868
rect 14921 54859 14979 54865
rect 14921 54825 14933 54859
rect 14967 54856 14979 54859
rect 15470 54856 15476 54868
rect 14967 54828 15476 54856
rect 14967 54825 14979 54828
rect 14921 54819 14979 54825
rect 15470 54816 15476 54828
rect 15528 54856 15534 54868
rect 15654 54856 15660 54868
rect 15528 54828 15660 54856
rect 15528 54816 15534 54828
rect 15654 54816 15660 54828
rect 15712 54816 15718 54868
rect 16574 54816 16580 54868
rect 16632 54856 16638 54868
rect 16761 54859 16819 54865
rect 16761 54856 16773 54859
rect 16632 54828 16773 54856
rect 16632 54816 16638 54828
rect 16761 54825 16773 54828
rect 16807 54856 16819 54859
rect 17037 54859 17095 54865
rect 17037 54856 17049 54859
rect 16807 54828 17049 54856
rect 16807 54825 16819 54828
rect 16761 54819 16819 54825
rect 17037 54825 17049 54828
rect 17083 54825 17095 54859
rect 17586 54856 17592 54868
rect 17547 54828 17592 54856
rect 17037 54819 17095 54825
rect 17586 54816 17592 54828
rect 17644 54816 17650 54868
rect 19058 54816 19064 54868
rect 19116 54856 19122 54868
rect 19116 54828 19472 54856
rect 19116 54816 19122 54828
rect 19444 54800 19472 54828
rect 21910 54816 21916 54868
rect 21968 54856 21974 54868
rect 22005 54859 22063 54865
rect 22005 54856 22017 54859
rect 21968 54828 22017 54856
rect 21968 54816 21974 54828
rect 22005 54825 22017 54828
rect 22051 54825 22063 54859
rect 22005 54819 22063 54825
rect 23569 54859 23627 54865
rect 23569 54825 23581 54859
rect 23615 54856 23627 54859
rect 23842 54856 23848 54868
rect 23615 54828 23848 54856
rect 23615 54825 23627 54828
rect 23569 54819 23627 54825
rect 23842 54816 23848 54828
rect 23900 54816 23906 54868
rect 23934 54816 23940 54868
rect 23992 54856 23998 54868
rect 27893 54859 27951 54865
rect 23992 54828 24037 54856
rect 23992 54816 23998 54828
rect 27893 54825 27905 54859
rect 27939 54856 27951 54859
rect 28074 54856 28080 54868
rect 27939 54828 28080 54856
rect 27939 54825 27951 54828
rect 27893 54819 27951 54825
rect 14093 54791 14151 54797
rect 14093 54757 14105 54791
rect 14139 54788 14151 54791
rect 14826 54788 14832 54800
rect 14139 54760 14832 54788
rect 14139 54757 14151 54760
rect 14093 54751 14151 54757
rect 14826 54748 14832 54760
rect 14884 54788 14890 54800
rect 15565 54791 15623 54797
rect 15565 54788 15577 54791
rect 14884 54760 15577 54788
rect 14884 54748 14890 54760
rect 15565 54757 15577 54760
rect 15611 54788 15623 54791
rect 15749 54791 15807 54797
rect 15749 54788 15761 54791
rect 15611 54760 15761 54788
rect 15611 54757 15623 54760
rect 15565 54751 15623 54757
rect 15749 54757 15761 54760
rect 15795 54788 15807 54791
rect 18046 54788 18052 54800
rect 15795 54760 18052 54788
rect 15795 54757 15807 54760
rect 15749 54751 15807 54757
rect 18046 54748 18052 54760
rect 18104 54748 18110 54800
rect 19242 54788 19248 54800
rect 18800 54760 19248 54788
rect 13170 54720 13176 54732
rect 13083 54692 13176 54720
rect 13170 54680 13176 54692
rect 13228 54720 13234 54732
rect 13354 54720 13360 54732
rect 13228 54692 13360 54720
rect 13228 54680 13234 54692
rect 13354 54680 13360 54692
rect 13412 54680 13418 54732
rect 14182 54720 14188 54732
rect 14143 54692 14188 54720
rect 14182 54680 14188 54692
rect 14240 54680 14246 54732
rect 17218 54680 17224 54732
rect 17276 54720 17282 54732
rect 17405 54723 17463 54729
rect 17405 54720 17417 54723
rect 17276 54692 17417 54720
rect 17276 54680 17282 54692
rect 17405 54689 17417 54692
rect 17451 54689 17463 54723
rect 17405 54683 17463 54689
rect 18800 54664 18828 54760
rect 19242 54748 19248 54760
rect 19300 54748 19306 54800
rect 19426 54788 19432 54800
rect 19387 54760 19432 54788
rect 19426 54748 19432 54760
rect 19484 54748 19490 54800
rect 19981 54791 20039 54797
rect 19981 54757 19993 54791
rect 20027 54788 20039 54791
rect 20622 54788 20628 54800
rect 20027 54760 20628 54788
rect 20027 54757 20039 54760
rect 19981 54751 20039 54757
rect 20622 54748 20628 54760
rect 20680 54748 20686 54800
rect 22830 54788 22836 54800
rect 22572 54760 22836 54788
rect 19334 54720 19340 54732
rect 19295 54692 19340 54720
rect 19334 54680 19340 54692
rect 19392 54680 19398 54732
rect 19521 54723 19579 54729
rect 19521 54689 19533 54723
rect 19567 54720 19579 54723
rect 19610 54720 19616 54732
rect 19567 54692 19616 54720
rect 19567 54689 19579 54692
rect 19521 54683 19579 54689
rect 19610 54680 19616 54692
rect 19668 54680 19674 54732
rect 20162 54680 20168 54732
rect 20220 54720 20226 54732
rect 21450 54720 21456 54732
rect 20220 54692 21456 54720
rect 20220 54680 20226 54692
rect 21450 54680 21456 54692
rect 21508 54720 21514 54732
rect 21545 54723 21603 54729
rect 21545 54720 21557 54723
rect 21508 54692 21557 54720
rect 21508 54680 21514 54692
rect 21545 54689 21557 54692
rect 21591 54689 21603 54723
rect 21545 54683 21603 54689
rect 21634 54680 21640 54732
rect 21692 54720 21698 54732
rect 22572 54729 22600 54760
rect 22830 54748 22836 54760
rect 22888 54748 22894 54800
rect 24302 54748 24308 54800
rect 24360 54788 24366 54800
rect 25130 54788 25136 54800
rect 24360 54760 25136 54788
rect 24360 54748 24366 54760
rect 25130 54748 25136 54760
rect 25188 54788 25194 54800
rect 25188 54760 25452 54788
rect 25188 54748 25194 54760
rect 21729 54723 21787 54729
rect 21729 54720 21741 54723
rect 21692 54692 21741 54720
rect 21692 54680 21698 54692
rect 21729 54689 21741 54692
rect 21775 54689 21787 54723
rect 21729 54683 21787 54689
rect 22557 54723 22615 54729
rect 22557 54689 22569 54723
rect 22603 54689 22615 54723
rect 22738 54720 22744 54732
rect 22699 54692 22744 54720
rect 22557 54683 22615 54689
rect 22738 54680 22744 54692
rect 22796 54680 22802 54732
rect 23934 54680 23940 54732
rect 23992 54720 23998 54732
rect 25038 54720 25044 54732
rect 23992 54692 25044 54720
rect 23992 54680 23998 54692
rect 25038 54680 25044 54692
rect 25096 54680 25102 54732
rect 25424 54729 25452 54760
rect 26234 54748 26240 54800
rect 26292 54788 26298 54800
rect 26513 54791 26571 54797
rect 26513 54788 26525 54791
rect 26292 54760 26525 54788
rect 26292 54748 26298 54760
rect 26513 54757 26525 54760
rect 26559 54757 26571 54791
rect 26513 54751 26571 54757
rect 25409 54723 25467 54729
rect 25409 54689 25421 54723
rect 25455 54689 25467 54723
rect 25409 54683 25467 54689
rect 25958 54680 25964 54732
rect 26016 54720 26022 54732
rect 26973 54723 27031 54729
rect 26973 54720 26985 54723
rect 26016 54692 26985 54720
rect 26016 54680 26022 54692
rect 26973 54689 26985 54692
rect 27019 54689 27031 54723
rect 26973 54683 27031 54689
rect 27341 54723 27399 54729
rect 27341 54689 27353 54723
rect 27387 54720 27399 54723
rect 27908 54720 27936 54819
rect 28074 54816 28080 54828
rect 28132 54816 28138 54868
rect 27387 54692 27936 54720
rect 28629 54723 28687 54729
rect 27387 54689 27399 54692
rect 27341 54683 27399 54689
rect 28629 54689 28641 54723
rect 28675 54720 28687 54723
rect 28994 54720 29000 54732
rect 28675 54692 29000 54720
rect 28675 54689 28687 54692
rect 28629 54683 28687 54689
rect 28994 54680 29000 54692
rect 29052 54680 29058 54732
rect 15286 54612 15292 54664
rect 15344 54652 15350 54664
rect 16117 54655 16175 54661
rect 16117 54652 16129 54655
rect 15344 54624 16129 54652
rect 15344 54612 15350 54624
rect 16117 54621 16129 54624
rect 16163 54652 16175 54655
rect 16850 54652 16856 54664
rect 16163 54624 16856 54652
rect 16163 54621 16175 54624
rect 16117 54615 16175 54621
rect 16850 54612 16856 54624
rect 16908 54612 16914 54664
rect 17037 54655 17095 54661
rect 17037 54621 17049 54655
rect 17083 54652 17095 54655
rect 18601 54655 18659 54661
rect 18601 54652 18613 54655
rect 17083 54624 18613 54652
rect 17083 54621 17095 54624
rect 17037 54615 17095 54621
rect 18601 54621 18613 54624
rect 18647 54652 18659 54655
rect 18782 54652 18788 54664
rect 18647 54624 18788 54652
rect 18647 54621 18659 54624
rect 18601 54615 18659 54621
rect 18782 54612 18788 54624
rect 18840 54612 18846 54664
rect 19153 54655 19211 54661
rect 19153 54621 19165 54655
rect 19199 54652 19211 54655
rect 22278 54652 22284 54664
rect 19199 54624 22284 54652
rect 19199 54621 19211 54624
rect 19153 54615 19211 54621
rect 22278 54612 22284 54624
rect 22336 54612 22342 54664
rect 22462 54612 22468 54664
rect 22520 54652 22526 54664
rect 23106 54652 23112 54664
rect 22520 54624 23112 54652
rect 22520 54612 22526 54624
rect 23106 54612 23112 54624
rect 23164 54612 23170 54664
rect 25133 54655 25191 54661
rect 25133 54621 25145 54655
rect 25179 54621 25191 54655
rect 25498 54652 25504 54664
rect 25459 54624 25504 54652
rect 25133 54615 25191 54621
rect 14366 54584 14372 54596
rect 14327 54556 14372 54584
rect 14366 54544 14372 54556
rect 14424 54544 14430 54596
rect 16022 54584 16028 54596
rect 15983 54556 16028 54584
rect 16022 54544 16028 54556
rect 16080 54584 16086 54596
rect 16574 54584 16580 54596
rect 16080 54556 16580 54584
rect 16080 54544 16086 54556
rect 16574 54544 16580 54556
rect 16632 54544 16638 54596
rect 17221 54587 17279 54593
rect 17221 54553 17233 54587
rect 17267 54584 17279 54587
rect 17494 54584 17500 54596
rect 17267 54556 17500 54584
rect 17267 54553 17279 54556
rect 17221 54547 17279 54553
rect 17494 54544 17500 54556
rect 17552 54584 17558 54596
rect 18506 54584 18512 54596
rect 17552 54556 18512 54584
rect 17552 54544 17558 54556
rect 18506 54544 18512 54556
rect 18564 54544 18570 54596
rect 20254 54544 20260 54596
rect 20312 54584 20318 54596
rect 20625 54587 20683 54593
rect 20625 54584 20637 54587
rect 20312 54556 20637 54584
rect 20312 54544 20318 54556
rect 20625 54553 20637 54556
rect 20671 54553 20683 54587
rect 20625 54547 20683 54553
rect 24305 54587 24363 54593
rect 24305 54553 24317 54587
rect 24351 54584 24363 54587
rect 25148 54584 25176 54615
rect 25498 54612 25504 54624
rect 25556 54612 25562 54664
rect 27433 54655 27491 54661
rect 27433 54621 27445 54655
rect 27479 54652 27491 54655
rect 27522 54652 27528 54664
rect 27479 54624 27528 54652
rect 27479 54621 27491 54624
rect 27433 54615 27491 54621
rect 27522 54612 27528 54624
rect 27580 54612 27586 54664
rect 28810 54612 28816 54664
rect 28868 54652 28874 54664
rect 28905 54655 28963 54661
rect 28905 54652 28917 54655
rect 28868 54624 28917 54652
rect 28868 54612 28874 54624
rect 28905 54621 28917 54624
rect 28951 54621 28963 54655
rect 28905 54615 28963 54621
rect 25406 54584 25412 54596
rect 24351 54556 25412 54584
rect 24351 54553 24363 54556
rect 24305 54547 24363 54553
rect 25406 54544 25412 54556
rect 25464 54544 25470 54596
rect 13354 54516 13360 54528
rect 13315 54488 13360 54516
rect 13354 54476 13360 54488
rect 13412 54476 13418 54528
rect 15010 54476 15016 54528
rect 15068 54516 15074 54528
rect 15838 54516 15844 54528
rect 15068 54488 15844 54516
rect 15068 54476 15074 54488
rect 15838 54476 15844 54488
rect 15896 54525 15902 54528
rect 15896 54519 15945 54525
rect 15896 54485 15899 54519
rect 15933 54485 15945 54519
rect 15896 54479 15945 54485
rect 16393 54519 16451 54525
rect 16393 54485 16405 54519
rect 16439 54516 16451 54519
rect 16482 54516 16488 54528
rect 16439 54488 16488 54516
rect 16439 54485 16451 54488
rect 16393 54479 16451 54485
rect 15896 54476 15902 54479
rect 16482 54476 16488 54488
rect 16540 54476 16546 54528
rect 20349 54519 20407 54525
rect 20349 54485 20361 54519
rect 20395 54516 20407 54519
rect 20714 54516 20720 54528
rect 20395 54488 20720 54516
rect 20395 54485 20407 54488
rect 20349 54479 20407 54485
rect 20714 54476 20720 54488
rect 20772 54476 20778 54528
rect 21082 54516 21088 54528
rect 21043 54488 21088 54516
rect 21082 54476 21088 54488
rect 21140 54476 21146 54528
rect 24486 54516 24492 54528
rect 24447 54488 24492 54516
rect 24486 54476 24492 54488
rect 24544 54476 24550 54528
rect 25774 54476 25780 54528
rect 25832 54516 25838 54528
rect 25869 54519 25927 54525
rect 25869 54516 25881 54519
rect 25832 54488 25881 54516
rect 25832 54476 25838 54488
rect 25869 54485 25881 54488
rect 25915 54485 25927 54519
rect 25869 54479 25927 54485
rect 26329 54519 26387 54525
rect 26329 54485 26341 54519
rect 26375 54516 26387 54519
rect 26878 54516 26884 54528
rect 26375 54488 26884 54516
rect 26375 54485 26387 54488
rect 26329 54479 26387 54485
rect 26878 54476 26884 54488
rect 26936 54476 26942 54528
rect 29086 54476 29092 54528
rect 29144 54516 29150 54528
rect 30009 54519 30067 54525
rect 30009 54516 30021 54519
rect 29144 54488 30021 54516
rect 29144 54476 29150 54488
rect 30009 54485 30021 54488
rect 30055 54485 30067 54519
rect 30009 54479 30067 54485
rect 31754 54476 31760 54528
rect 31812 54516 31818 54528
rect 31812 54488 31857 54516
rect 31812 54476 31818 54488
rect 1104 54426 38824 54448
rect 1104 54374 4246 54426
rect 4298 54374 4310 54426
rect 4362 54374 4374 54426
rect 4426 54374 4438 54426
rect 4490 54374 34966 54426
rect 35018 54374 35030 54426
rect 35082 54374 35094 54426
rect 35146 54374 35158 54426
rect 35210 54374 38824 54426
rect 1104 54352 38824 54374
rect 13170 54312 13176 54324
rect 13131 54284 13176 54312
rect 13170 54272 13176 54284
rect 13228 54272 13234 54324
rect 14182 54272 14188 54324
rect 14240 54312 14246 54324
rect 14277 54315 14335 54321
rect 14277 54312 14289 54315
rect 14240 54284 14289 54312
rect 14240 54272 14246 54284
rect 14277 54281 14289 54284
rect 14323 54281 14335 54315
rect 16850 54312 16856 54324
rect 16811 54284 16856 54312
rect 14277 54275 14335 54281
rect 16850 54272 16856 54284
rect 16908 54272 16914 54324
rect 17586 54312 17592 54324
rect 17499 54284 17592 54312
rect 17586 54272 17592 54284
rect 17644 54312 17650 54324
rect 18046 54312 18052 54324
rect 17644 54284 18052 54312
rect 17644 54272 17650 54284
rect 18046 54272 18052 54284
rect 18104 54272 18110 54324
rect 19334 54272 19340 54324
rect 19392 54312 19398 54324
rect 19981 54315 20039 54321
rect 19981 54312 19993 54315
rect 19392 54284 19993 54312
rect 19392 54272 19398 54284
rect 19981 54281 19993 54284
rect 20027 54281 20039 54315
rect 19981 54275 20039 54281
rect 22002 54272 22008 54324
rect 22060 54312 22066 54324
rect 22186 54312 22192 54324
rect 22060 54284 22192 54312
rect 22060 54272 22066 54284
rect 22186 54272 22192 54284
rect 22244 54272 22250 54324
rect 23109 54315 23167 54321
rect 23109 54281 23121 54315
rect 23155 54312 23167 54315
rect 23842 54312 23848 54324
rect 23155 54284 23848 54312
rect 23155 54281 23167 54284
rect 23109 54275 23167 54281
rect 15838 54204 15844 54256
rect 15896 54244 15902 54256
rect 17129 54247 17187 54253
rect 17129 54244 17141 54247
rect 15896 54216 17141 54244
rect 15896 54204 15902 54216
rect 17129 54213 17141 54216
rect 17175 54244 17187 54247
rect 17770 54244 17776 54256
rect 17175 54216 17776 54244
rect 17175 54213 17187 54216
rect 17129 54207 17187 54213
rect 17770 54204 17776 54216
rect 17828 54204 17834 54256
rect 19610 54244 19616 54256
rect 19571 54216 19616 54244
rect 19610 54204 19616 54216
rect 19668 54204 19674 54256
rect 13998 54136 14004 54188
rect 14056 54176 14062 54188
rect 14458 54176 14464 54188
rect 14056 54148 14464 54176
rect 14056 54136 14062 54148
rect 14458 54136 14464 54148
rect 14516 54176 14522 54188
rect 14829 54179 14887 54185
rect 14829 54176 14841 54179
rect 14516 54148 14841 54176
rect 14516 54136 14522 54148
rect 14829 54145 14841 54148
rect 14875 54145 14887 54179
rect 14829 54139 14887 54145
rect 16485 54179 16543 54185
rect 16485 54145 16497 54179
rect 16531 54176 16543 54179
rect 17218 54176 17224 54188
rect 16531 54148 17224 54176
rect 16531 54145 16543 54148
rect 16485 54139 16543 54145
rect 17218 54136 17224 54148
rect 17276 54136 17282 54188
rect 19426 54136 19432 54188
rect 19484 54176 19490 54188
rect 20165 54179 20223 54185
rect 20165 54176 20177 54179
rect 19484 54148 20177 54176
rect 19484 54136 19490 54148
rect 20165 54145 20177 54148
rect 20211 54176 20223 54179
rect 20622 54176 20628 54188
rect 20211 54148 20628 54176
rect 20211 54145 20223 54148
rect 20165 54139 20223 54145
rect 20622 54136 20628 54148
rect 20680 54136 20686 54188
rect 20901 54179 20959 54185
rect 20901 54145 20913 54179
rect 20947 54176 20959 54179
rect 21174 54176 21180 54188
rect 20947 54148 21180 54176
rect 20947 54145 20959 54148
rect 20901 54139 20959 54145
rect 21174 54136 21180 54148
rect 21232 54136 21238 54188
rect 21450 54136 21456 54188
rect 21508 54176 21514 54188
rect 22370 54176 22376 54188
rect 21508 54148 22376 54176
rect 21508 54136 21514 54148
rect 22370 54136 22376 54148
rect 22428 54185 22434 54188
rect 22428 54179 22477 54185
rect 22428 54145 22431 54179
rect 22465 54145 22477 54179
rect 22428 54139 22477 54145
rect 22428 54136 22434 54139
rect 12434 54068 12440 54120
rect 12492 54108 12498 54120
rect 13725 54111 13783 54117
rect 13725 54108 13737 54111
rect 12492 54080 13737 54108
rect 12492 54068 12498 54080
rect 13725 54077 13737 54080
rect 13771 54108 13783 54111
rect 13817 54111 13875 54117
rect 13817 54108 13829 54111
rect 13771 54080 13829 54108
rect 13771 54077 13783 54080
rect 13725 54071 13783 54077
rect 13817 54077 13829 54080
rect 13863 54108 13875 54111
rect 14366 54108 14372 54120
rect 13863 54080 14372 54108
rect 13863 54077 13875 54080
rect 13817 54071 13875 54077
rect 14366 54068 14372 54080
rect 14424 54068 14430 54120
rect 15105 54111 15163 54117
rect 15105 54108 15117 54111
rect 14936 54080 15117 54108
rect 14826 54040 14832 54052
rect 14016 54012 14832 54040
rect 14016 53981 14044 54012
rect 14826 54000 14832 54012
rect 14884 54000 14890 54052
rect 14001 53975 14059 53981
rect 14001 53941 14013 53975
rect 14047 53941 14059 53975
rect 14734 53972 14740 53984
rect 14695 53944 14740 53972
rect 14001 53935 14059 53941
rect 14734 53932 14740 53944
rect 14792 53972 14798 53984
rect 14936 53972 14964 54080
rect 15105 54077 15117 54080
rect 15151 54077 15163 54111
rect 18598 54108 18604 54120
rect 18559 54080 18604 54108
rect 15105 54071 15163 54077
rect 18598 54068 18604 54080
rect 18656 54068 18662 54120
rect 18782 54108 18788 54120
rect 18743 54080 18788 54108
rect 18782 54068 18788 54080
rect 18840 54068 18846 54120
rect 18877 54111 18935 54117
rect 18877 54077 18889 54111
rect 18923 54077 18935 54111
rect 18877 54071 18935 54077
rect 19337 54111 19395 54117
rect 19337 54077 19349 54111
rect 19383 54108 19395 54111
rect 21545 54111 21603 54117
rect 21545 54108 21557 54111
rect 19383 54080 21557 54108
rect 19383 54077 19395 54080
rect 19337 54071 19395 54077
rect 21545 54077 21557 54080
rect 21591 54108 21603 54111
rect 21634 54108 21640 54120
rect 21591 54080 21640 54108
rect 21591 54077 21603 54080
rect 21545 54071 21603 54077
rect 18892 54040 18920 54071
rect 21634 54068 21640 54080
rect 21692 54068 21698 54120
rect 22002 54068 22008 54120
rect 22060 54108 22066 54120
rect 22281 54111 22339 54117
rect 22281 54108 22293 54111
rect 22060 54080 22293 54108
rect 22060 54068 22066 54080
rect 22281 54077 22293 54080
rect 22327 54077 22339 54111
rect 22554 54108 22560 54120
rect 22467 54080 22560 54108
rect 22281 54071 22339 54077
rect 19610 54040 19616 54052
rect 18892 54012 19616 54040
rect 14792 53944 14964 53972
rect 18509 53975 18567 53981
rect 14792 53932 14798 53944
rect 18509 53941 18521 53975
rect 18555 53972 18567 53975
rect 18892 53972 18920 54012
rect 19610 54000 19616 54012
rect 19668 54040 19674 54052
rect 20070 54040 20076 54052
rect 19668 54012 20076 54040
rect 19668 54000 19674 54012
rect 20070 54000 20076 54012
rect 20128 54000 20134 54052
rect 20533 54043 20591 54049
rect 20533 54009 20545 54043
rect 20579 54040 20591 54043
rect 20714 54040 20720 54052
rect 20579 54012 20720 54040
rect 20579 54009 20591 54012
rect 20533 54003 20591 54009
rect 20714 54000 20720 54012
rect 20772 54000 20778 54052
rect 21082 54000 21088 54052
rect 21140 54040 21146 54052
rect 21269 54043 21327 54049
rect 21269 54040 21281 54043
rect 21140 54012 21281 54040
rect 21140 54000 21146 54012
rect 21269 54009 21281 54012
rect 21315 54040 21327 54043
rect 21729 54043 21787 54049
rect 21315 54012 21680 54040
rect 21315 54009 21327 54012
rect 21269 54003 21327 54009
rect 18555 53944 18920 53972
rect 18555 53941 18567 53944
rect 18509 53935 18567 53941
rect 19334 53932 19340 53984
rect 19392 53972 19398 53984
rect 20254 53972 20260 53984
rect 19392 53944 20260 53972
rect 19392 53932 19398 53944
rect 20254 53932 20260 53944
rect 20312 53972 20318 53984
rect 20349 53975 20407 53981
rect 20349 53972 20361 53975
rect 20312 53944 20361 53972
rect 20312 53932 20318 53944
rect 20349 53941 20361 53944
rect 20395 53941 20407 53975
rect 20349 53935 20407 53941
rect 20438 53932 20444 53984
rect 20496 53972 20502 53984
rect 21652 53972 21680 54012
rect 21729 54009 21741 54043
rect 21775 54040 21787 54043
rect 21910 54040 21916 54052
rect 21775 54012 21916 54040
rect 21775 54009 21787 54012
rect 21729 54003 21787 54009
rect 21910 54000 21916 54012
rect 21968 54000 21974 54052
rect 22296 54040 22324 54071
rect 22554 54068 22560 54080
rect 22612 54108 22618 54120
rect 23124 54108 23152 54275
rect 23842 54272 23848 54284
rect 23900 54272 23906 54324
rect 24302 54312 24308 54324
rect 24263 54284 24308 54312
rect 24302 54272 24308 54284
rect 24360 54272 24366 54324
rect 27890 54312 27896 54324
rect 27851 54284 27896 54312
rect 27890 54272 27896 54284
rect 27948 54272 27954 54324
rect 28721 54315 28779 54321
rect 28721 54281 28733 54315
rect 28767 54312 28779 54315
rect 28810 54312 28816 54324
rect 28767 54284 28816 54312
rect 28767 54281 28779 54284
rect 28721 54275 28779 54281
rect 28810 54272 28816 54284
rect 28868 54272 28874 54324
rect 28994 54272 29000 54324
rect 29052 54312 29058 54324
rect 29089 54315 29147 54321
rect 29089 54312 29101 54315
rect 29052 54284 29101 54312
rect 29052 54272 29058 54284
rect 29089 54281 29101 54284
rect 29135 54312 29147 54315
rect 29546 54312 29552 54324
rect 29135 54284 29552 54312
rect 29135 54281 29147 54284
rect 29089 54275 29147 54281
rect 29546 54272 29552 54284
rect 29604 54312 29610 54324
rect 30282 54312 30288 54324
rect 29604 54284 30288 54312
rect 29604 54272 29610 54284
rect 30282 54272 30288 54284
rect 30340 54272 30346 54324
rect 23477 54247 23535 54253
rect 23477 54213 23489 54247
rect 23523 54244 23535 54247
rect 23934 54244 23940 54256
rect 23523 54216 23940 54244
rect 23523 54213 23535 54216
rect 23477 54207 23535 54213
rect 23934 54204 23940 54216
rect 23992 54204 23998 54256
rect 24762 54204 24768 54256
rect 24820 54244 24826 54256
rect 24820 54216 25636 54244
rect 24820 54204 24826 54216
rect 25608 54188 25636 54216
rect 25225 54179 25283 54185
rect 25225 54145 25237 54179
rect 25271 54176 25283 54179
rect 25406 54176 25412 54188
rect 25271 54148 25412 54176
rect 25271 54145 25283 54148
rect 25225 54139 25283 54145
rect 25406 54136 25412 54148
rect 25464 54136 25470 54188
rect 25590 54176 25596 54188
rect 25551 54148 25596 54176
rect 25590 54136 25596 54148
rect 25648 54136 25654 54188
rect 26234 54136 26240 54188
rect 26292 54176 26298 54188
rect 27249 54179 27307 54185
rect 27249 54176 27261 54179
rect 26292 54148 27261 54176
rect 26292 54136 26298 54148
rect 27249 54145 27261 54148
rect 27295 54145 27307 54179
rect 27249 54139 27307 54145
rect 22612 54080 23152 54108
rect 24029 54111 24087 54117
rect 22612 54068 22618 54080
rect 24029 54077 24041 54111
rect 24075 54108 24087 54111
rect 24946 54108 24952 54120
rect 24075 54080 24952 54108
rect 24075 54077 24087 54080
rect 24029 54071 24087 54077
rect 24946 54068 24952 54080
rect 25004 54068 25010 54120
rect 25038 54068 25044 54120
rect 25096 54108 25102 54120
rect 25133 54111 25191 54117
rect 25133 54108 25145 54111
rect 25096 54080 25145 54108
rect 25096 54068 25102 54080
rect 25133 54077 25145 54080
rect 25179 54077 25191 54111
rect 25498 54108 25504 54120
rect 25411 54080 25504 54108
rect 25133 54071 25191 54077
rect 25498 54068 25504 54080
rect 25556 54068 25562 54120
rect 26513 54111 26571 54117
rect 26513 54077 26525 54111
rect 26559 54108 26571 54111
rect 26694 54108 26700 54120
rect 26559 54080 26700 54108
rect 26559 54077 26571 54080
rect 26513 54071 26571 54077
rect 26694 54068 26700 54080
rect 26752 54068 26758 54120
rect 26786 54068 26792 54120
rect 26844 54108 26850 54120
rect 27525 54111 27583 54117
rect 27525 54108 27537 54111
rect 26844 54080 27537 54108
rect 26844 54068 26850 54080
rect 27525 54077 27537 54080
rect 27571 54077 27583 54111
rect 27525 54071 27583 54077
rect 27890 54068 27896 54120
rect 27948 54108 27954 54120
rect 28077 54111 28135 54117
rect 28077 54108 28089 54111
rect 27948 54080 28089 54108
rect 27948 54068 27954 54080
rect 28077 54077 28089 54080
rect 28123 54077 28135 54111
rect 28077 54071 28135 54077
rect 22370 54040 22376 54052
rect 22296 54012 22376 54040
rect 22370 54000 22376 54012
rect 22428 54000 22434 54052
rect 24486 54040 24492 54052
rect 24447 54012 24492 54040
rect 24486 54000 24492 54012
rect 24544 54000 24550 54052
rect 24964 54040 24992 54068
rect 25516 54040 25544 54068
rect 24964 54012 25544 54040
rect 26234 54000 26240 54052
rect 26292 54040 26298 54052
rect 26878 54040 26884 54052
rect 26292 54012 26740 54040
rect 26839 54012 26884 54040
rect 26292 54000 26298 54012
rect 22830 53972 22836 53984
rect 20496 53944 20541 53972
rect 21652 53944 22836 53972
rect 20496 53932 20502 53944
rect 22830 53932 22836 53944
rect 22888 53932 22894 53984
rect 25958 53972 25964 53984
rect 25919 53944 25964 53972
rect 25958 53932 25964 53944
rect 26016 53932 26022 53984
rect 26326 53972 26332 53984
rect 26287 53944 26332 53972
rect 26326 53932 26332 53944
rect 26384 53932 26390 53984
rect 26712 53981 26740 54012
rect 26878 54000 26884 54012
rect 26936 54000 26942 54052
rect 26697 53975 26755 53981
rect 26697 53941 26709 53975
rect 26743 53972 26755 53975
rect 28261 53975 28319 53981
rect 28261 53972 28273 53975
rect 26743 53944 28273 53972
rect 26743 53941 26755 53944
rect 26697 53935 26755 53941
rect 28261 53941 28273 53944
rect 28307 53941 28319 53975
rect 28261 53935 28319 53941
rect 1104 53882 38824 53904
rect 1104 53830 19606 53882
rect 19658 53830 19670 53882
rect 19722 53830 19734 53882
rect 19786 53830 19798 53882
rect 19850 53830 38824 53882
rect 1104 53808 38824 53830
rect 14093 53771 14151 53777
rect 14093 53737 14105 53771
rect 14139 53768 14151 53771
rect 14458 53768 14464 53780
rect 14139 53740 14464 53768
rect 14139 53737 14151 53740
rect 14093 53731 14151 53737
rect 14458 53728 14464 53740
rect 14516 53728 14522 53780
rect 14642 53728 14648 53780
rect 14700 53768 14706 53780
rect 15841 53771 15899 53777
rect 15841 53768 15853 53771
rect 14700 53740 15853 53768
rect 14700 53728 14706 53740
rect 15841 53737 15853 53740
rect 15887 53737 15899 53771
rect 15841 53731 15899 53737
rect 16390 53728 16396 53780
rect 16448 53768 16454 53780
rect 17037 53771 17095 53777
rect 17037 53768 17049 53771
rect 16448 53740 17049 53768
rect 16448 53728 16454 53740
rect 17037 53737 17049 53740
rect 17083 53768 17095 53771
rect 17586 53768 17592 53780
rect 17083 53740 17592 53768
rect 17083 53737 17095 53740
rect 17037 53731 17095 53737
rect 17586 53728 17592 53740
rect 17644 53728 17650 53780
rect 19334 53728 19340 53780
rect 19392 53768 19398 53780
rect 19429 53771 19487 53777
rect 19429 53768 19441 53771
rect 19392 53740 19441 53768
rect 19392 53728 19398 53740
rect 19429 53737 19441 53740
rect 19475 53737 19487 53771
rect 19429 53731 19487 53737
rect 19521 53771 19579 53777
rect 19521 53737 19533 53771
rect 19567 53768 19579 53771
rect 19978 53768 19984 53780
rect 19567 53740 19984 53768
rect 19567 53737 19579 53740
rect 19521 53731 19579 53737
rect 19978 53728 19984 53740
rect 20036 53728 20042 53780
rect 20349 53771 20407 53777
rect 20349 53737 20361 53771
rect 20395 53768 20407 53771
rect 20438 53768 20444 53780
rect 20395 53740 20444 53768
rect 20395 53737 20407 53740
rect 20349 53731 20407 53737
rect 20438 53728 20444 53740
rect 20496 53728 20502 53780
rect 20622 53768 20628 53780
rect 20583 53740 20628 53768
rect 20622 53728 20628 53740
rect 20680 53728 20686 53780
rect 21177 53771 21235 53777
rect 21177 53737 21189 53771
rect 21223 53768 21235 53771
rect 22370 53768 22376 53780
rect 21223 53740 22376 53768
rect 21223 53737 21235 53740
rect 21177 53731 21235 53737
rect 22370 53728 22376 53740
rect 22428 53728 22434 53780
rect 22741 53771 22799 53777
rect 22741 53737 22753 53771
rect 22787 53768 22799 53771
rect 22922 53768 22928 53780
rect 22787 53740 22928 53768
rect 22787 53737 22799 53740
rect 22741 53731 22799 53737
rect 22922 53728 22928 53740
rect 22980 53728 22986 53780
rect 15102 53700 15108 53712
rect 15063 53672 15108 53700
rect 15102 53660 15108 53672
rect 15160 53660 15166 53712
rect 15654 53660 15660 53712
rect 15712 53700 15718 53712
rect 15749 53703 15807 53709
rect 15749 53700 15761 53703
rect 15712 53672 15761 53700
rect 15712 53660 15718 53672
rect 15749 53669 15761 53672
rect 15795 53669 15807 53703
rect 15930 53700 15936 53712
rect 15891 53672 15936 53700
rect 15749 53663 15807 53669
rect 15930 53660 15936 53672
rect 15988 53660 15994 53712
rect 16298 53700 16304 53712
rect 16259 53672 16304 53700
rect 16298 53660 16304 53672
rect 16356 53660 16362 53712
rect 16574 53700 16580 53712
rect 16535 53672 16580 53700
rect 16574 53660 16580 53672
rect 16632 53660 16638 53712
rect 16942 53660 16948 53712
rect 17000 53700 17006 53712
rect 17000 53672 18000 53700
rect 17000 53660 17006 53672
rect 14185 53635 14243 53641
rect 14185 53601 14197 53635
rect 14231 53632 14243 53635
rect 14274 53632 14280 53644
rect 14231 53604 14280 53632
rect 14231 53601 14243 53604
rect 14185 53595 14243 53601
rect 14274 53592 14280 53604
rect 14332 53592 14338 53644
rect 14366 53592 14372 53644
rect 14424 53632 14430 53644
rect 15565 53635 15623 53641
rect 15565 53632 15577 53635
rect 14424 53604 15577 53632
rect 14424 53592 14430 53604
rect 15565 53601 15577 53604
rect 15611 53632 15623 53635
rect 16758 53632 16764 53644
rect 15611 53604 16764 53632
rect 15611 53601 15623 53604
rect 15565 53595 15623 53601
rect 16758 53592 16764 53604
rect 16816 53592 16822 53644
rect 16850 53592 16856 53644
rect 16908 53632 16914 53644
rect 17129 53635 17187 53641
rect 17129 53632 17141 53635
rect 16908 53604 17141 53632
rect 16908 53592 16914 53604
rect 17129 53601 17141 53604
rect 17175 53601 17187 53635
rect 17494 53632 17500 53644
rect 17455 53604 17500 53632
rect 17129 53595 17187 53601
rect 17494 53592 17500 53604
rect 17552 53592 17558 53644
rect 17972 53641 18000 53672
rect 18598 53660 18604 53712
rect 18656 53700 18662 53712
rect 19245 53703 19303 53709
rect 19245 53700 19257 53703
rect 18656 53672 19257 53700
rect 18656 53660 18662 53672
rect 19245 53669 19257 53672
rect 19291 53669 19303 53703
rect 19610 53700 19616 53712
rect 19523 53672 19616 53700
rect 19245 53663 19303 53669
rect 19610 53660 19616 53672
rect 19668 53700 19674 53712
rect 20714 53700 20720 53712
rect 19668 53672 20720 53700
rect 19668 53660 19674 53672
rect 20714 53660 20720 53672
rect 20772 53660 20778 53712
rect 21542 53700 21548 53712
rect 21503 53672 21548 53700
rect 21542 53660 21548 53672
rect 21600 53660 21606 53712
rect 23477 53703 23535 53709
rect 23477 53669 23489 53703
rect 23523 53700 23535 53703
rect 23566 53700 23572 53712
rect 23523 53672 23572 53700
rect 23523 53669 23535 53672
rect 23477 53663 23535 53669
rect 23566 53660 23572 53672
rect 23624 53700 23630 53712
rect 23624 53672 24164 53700
rect 23624 53660 23630 53672
rect 24136 53644 24164 53672
rect 17957 53635 18015 53641
rect 17957 53601 17969 53635
rect 18003 53632 18015 53635
rect 18966 53632 18972 53644
rect 18003 53604 18972 53632
rect 18003 53601 18015 53604
rect 17957 53595 18015 53601
rect 18966 53592 18972 53604
rect 19024 53592 19030 53644
rect 19981 53635 20039 53641
rect 19981 53601 19993 53635
rect 20027 53632 20039 53635
rect 21634 53632 21640 53644
rect 20027 53604 21640 53632
rect 20027 53601 20039 53604
rect 19981 53595 20039 53601
rect 21634 53592 21640 53604
rect 21692 53592 21698 53644
rect 22370 53592 22376 53644
rect 22428 53632 22434 53644
rect 22465 53635 22523 53641
rect 22465 53632 22477 53635
rect 22428 53604 22477 53632
rect 22428 53592 22434 53604
rect 22465 53601 22477 53604
rect 22511 53601 22523 53635
rect 22465 53595 22523 53601
rect 23753 53635 23811 53641
rect 23753 53601 23765 53635
rect 23799 53632 23811 53635
rect 23842 53632 23848 53644
rect 23799 53604 23848 53632
rect 23799 53601 23811 53604
rect 23753 53595 23811 53601
rect 23842 53592 23848 53604
rect 23900 53592 23906 53644
rect 24118 53632 24124 53644
rect 24079 53604 24124 53632
rect 24118 53592 24124 53604
rect 24176 53592 24182 53644
rect 24486 53632 24492 53644
rect 24447 53604 24492 53632
rect 24486 53592 24492 53604
rect 24544 53632 24550 53644
rect 24670 53632 24676 53644
rect 24544 53604 24676 53632
rect 24544 53592 24550 53604
rect 24670 53592 24676 53604
rect 24728 53592 24734 53644
rect 27338 53632 27344 53644
rect 27299 53604 27344 53632
rect 27338 53592 27344 53604
rect 27396 53592 27402 53644
rect 27522 53632 27528 53644
rect 27435 53604 27528 53632
rect 27522 53592 27528 53604
rect 27580 53592 27586 53644
rect 27709 53635 27767 53641
rect 27709 53601 27721 53635
rect 27755 53632 27767 53635
rect 28166 53632 28172 53644
rect 27755 53604 28172 53632
rect 27755 53601 27767 53604
rect 27709 53595 27767 53601
rect 28166 53592 28172 53604
rect 28224 53592 28230 53644
rect 19426 53524 19432 53576
rect 19484 53564 19490 53576
rect 20346 53564 20352 53576
rect 19484 53536 20352 53564
rect 19484 53524 19490 53536
rect 20346 53524 20352 53536
rect 20404 53524 20410 53576
rect 21358 53524 21364 53576
rect 21416 53564 21422 53576
rect 22557 53567 22615 53573
rect 22557 53564 22569 53567
rect 21416 53536 22569 53564
rect 21416 53524 21422 53536
rect 22557 53533 22569 53536
rect 22603 53564 22615 53567
rect 22603 53536 23152 53564
rect 22603 53533 22615 53536
rect 22557 53527 22615 53533
rect 14369 53499 14427 53505
rect 14369 53465 14381 53499
rect 14415 53496 14427 53499
rect 14918 53496 14924 53508
rect 14415 53468 14924 53496
rect 14415 53465 14427 53468
rect 14369 53459 14427 53465
rect 14918 53456 14924 53468
rect 14976 53456 14982 53508
rect 17954 53496 17960 53508
rect 17915 53468 17960 53496
rect 17954 53456 17960 53468
rect 18012 53456 18018 53508
rect 19058 53496 19064 53508
rect 18064 53468 19064 53496
rect 14734 53428 14740 53440
rect 14695 53400 14740 53428
rect 14734 53388 14740 53400
rect 14792 53388 14798 53440
rect 15654 53388 15660 53440
rect 15712 53428 15718 53440
rect 18064 53428 18092 53468
rect 19058 53456 19064 53468
rect 19116 53456 19122 53508
rect 18598 53428 18604 53440
rect 15712 53400 18092 53428
rect 18559 53400 18604 53428
rect 15712 53388 15718 53400
rect 18598 53388 18604 53400
rect 18656 53388 18662 53440
rect 23124 53437 23152 53536
rect 23290 53524 23296 53576
rect 23348 53564 23354 53576
rect 23348 53536 23888 53564
rect 23348 53524 23354 53536
rect 23860 53508 23888 53536
rect 26326 53524 26332 53576
rect 26384 53564 26390 53576
rect 27540 53564 27568 53592
rect 26384 53536 27568 53564
rect 26384 53524 26390 53536
rect 23842 53456 23848 53508
rect 23900 53456 23906 53508
rect 24394 53496 24400 53508
rect 24355 53468 24400 53496
rect 24394 53456 24400 53468
rect 24452 53456 24458 53508
rect 25222 53456 25228 53508
rect 25280 53496 25286 53508
rect 25685 53499 25743 53505
rect 25685 53496 25697 53499
rect 25280 53468 25697 53496
rect 25280 53456 25286 53468
rect 25685 53465 25697 53468
rect 25731 53465 25743 53499
rect 27154 53496 27160 53508
rect 27115 53468 27160 53496
rect 25685 53459 25743 53465
rect 27154 53456 27160 53468
rect 27212 53456 27218 53508
rect 23109 53431 23167 53437
rect 23109 53397 23121 53431
rect 23155 53428 23167 53431
rect 23290 53428 23296 53440
rect 23155 53400 23296 53428
rect 23155 53397 23167 53400
rect 23109 53391 23167 53397
rect 23290 53388 23296 53400
rect 23348 53388 23354 53440
rect 24946 53428 24952 53440
rect 24907 53400 24952 53428
rect 24946 53388 24952 53400
rect 25004 53388 25010 53440
rect 25409 53431 25467 53437
rect 25409 53397 25421 53431
rect 25455 53428 25467 53431
rect 25498 53428 25504 53440
rect 25455 53400 25504 53428
rect 25455 53397 25467 53400
rect 25409 53391 25467 53397
rect 25498 53388 25504 53400
rect 25556 53388 25562 53440
rect 26234 53428 26240 53440
rect 26195 53400 26240 53428
rect 26234 53388 26240 53400
rect 26292 53388 26298 53440
rect 26694 53428 26700 53440
rect 26655 53400 26700 53428
rect 26694 53388 26700 53400
rect 26752 53388 26758 53440
rect 1104 53338 38824 53360
rect 1104 53286 4246 53338
rect 4298 53286 4310 53338
rect 4362 53286 4374 53338
rect 4426 53286 4438 53338
rect 4490 53286 34966 53338
rect 35018 53286 35030 53338
rect 35082 53286 35094 53338
rect 35146 53286 35158 53338
rect 35210 53286 38824 53338
rect 1104 53264 38824 53286
rect 13814 53184 13820 53236
rect 13872 53224 13878 53236
rect 15105 53227 15163 53233
rect 15105 53224 15117 53227
rect 13872 53196 15117 53224
rect 13872 53184 13878 53196
rect 15105 53193 15117 53196
rect 15151 53224 15163 53227
rect 15838 53224 15844 53236
rect 15151 53196 15844 53224
rect 15151 53193 15163 53196
rect 15105 53187 15163 53193
rect 15838 53184 15844 53196
rect 15896 53184 15902 53236
rect 16574 53184 16580 53236
rect 16632 53224 16638 53236
rect 16669 53227 16727 53233
rect 16669 53224 16681 53227
rect 16632 53196 16681 53224
rect 16632 53184 16638 53196
rect 16669 53193 16681 53196
rect 16715 53193 16727 53227
rect 16669 53187 16727 53193
rect 16850 53184 16856 53236
rect 16908 53224 16914 53236
rect 17402 53224 17408 53236
rect 16908 53196 17408 53224
rect 16908 53184 16914 53196
rect 17402 53184 17408 53196
rect 17460 53224 17466 53236
rect 17773 53227 17831 53233
rect 17773 53224 17785 53227
rect 17460 53196 17785 53224
rect 17460 53184 17466 53196
rect 17773 53193 17785 53196
rect 17819 53193 17831 53227
rect 17773 53187 17831 53193
rect 18598 53184 18604 53236
rect 18656 53224 18662 53236
rect 19518 53224 19524 53236
rect 18656 53196 19524 53224
rect 18656 53184 18662 53196
rect 19518 53184 19524 53196
rect 19576 53184 19582 53236
rect 22554 53184 22560 53236
rect 22612 53224 22618 53236
rect 22649 53227 22707 53233
rect 22649 53224 22661 53227
rect 22612 53196 22661 53224
rect 22612 53184 22618 53196
rect 22649 53193 22661 53196
rect 22695 53193 22707 53227
rect 23474 53224 23480 53236
rect 23435 53196 23480 53224
rect 22649 53187 22707 53193
rect 23474 53184 23480 53196
rect 23532 53184 23538 53236
rect 24762 53224 24768 53236
rect 24723 53196 24768 53224
rect 24762 53184 24768 53196
rect 24820 53184 24826 53236
rect 29546 53224 29552 53236
rect 29507 53196 29552 53224
rect 29546 53184 29552 53196
rect 29604 53184 29610 53236
rect 14274 53156 14280 53168
rect 14235 53128 14280 53156
rect 14274 53116 14280 53128
rect 14332 53116 14338 53168
rect 14642 53116 14648 53168
rect 14700 53156 14706 53168
rect 14921 53159 14979 53165
rect 14921 53156 14933 53159
rect 14700 53128 14933 53156
rect 14700 53116 14706 53128
rect 14921 53125 14933 53128
rect 14967 53125 14979 53159
rect 14921 53119 14979 53125
rect 18230 53116 18236 53168
rect 18288 53156 18294 53168
rect 18969 53159 19027 53165
rect 18969 53156 18981 53159
rect 18288 53128 18981 53156
rect 18288 53116 18294 53128
rect 18969 53125 18981 53128
rect 19015 53125 19027 53159
rect 19978 53156 19984 53168
rect 19939 53128 19984 53156
rect 18969 53119 19027 53125
rect 19978 53116 19984 53128
rect 20036 53116 20042 53168
rect 20254 53116 20260 53168
rect 20312 53156 20318 53168
rect 20901 53159 20959 53165
rect 20901 53156 20913 53159
rect 20312 53128 20913 53156
rect 20312 53116 20318 53128
rect 20901 53125 20913 53128
rect 20947 53125 20959 53159
rect 20901 53119 20959 53125
rect 21818 53116 21824 53168
rect 21876 53156 21882 53168
rect 22005 53159 22063 53165
rect 22005 53156 22017 53159
rect 21876 53128 22017 53156
rect 21876 53116 21882 53128
rect 22005 53125 22017 53128
rect 22051 53125 22063 53159
rect 22005 53119 22063 53125
rect 14553 53091 14611 53097
rect 14553 53057 14565 53091
rect 14599 53088 14611 53091
rect 15654 53088 15660 53100
rect 14599 53060 15660 53088
rect 14599 53057 14611 53060
rect 14553 53051 14611 53057
rect 15654 53048 15660 53060
rect 15712 53048 15718 53100
rect 16758 53088 16764 53100
rect 16719 53060 16764 53088
rect 16758 53048 16764 53060
rect 16816 53048 16822 53100
rect 17129 53091 17187 53097
rect 17129 53057 17141 53091
rect 17175 53088 17187 53091
rect 20625 53091 20683 53097
rect 17175 53060 20116 53088
rect 17175 53057 17187 53060
rect 17129 53051 17187 53057
rect 13909 53023 13967 53029
rect 13909 52989 13921 53023
rect 13955 53020 13967 53023
rect 15286 53020 15292 53032
rect 13955 52992 15292 53020
rect 13955 52989 13967 52992
rect 13909 52983 13967 52989
rect 15286 52980 15292 52992
rect 15344 52980 15350 53032
rect 15381 53023 15439 53029
rect 15381 52989 15393 53023
rect 15427 53020 15439 53023
rect 15930 53020 15936 53032
rect 15427 52992 15936 53020
rect 15427 52989 15439 52992
rect 15381 52983 15439 52989
rect 15930 52980 15936 52992
rect 15988 52980 15994 53032
rect 16390 53020 16396 53032
rect 16351 52992 16396 53020
rect 16390 52980 16396 52992
rect 16448 52980 16454 53032
rect 16540 53023 16598 53029
rect 16540 52989 16552 53023
rect 16586 53020 16598 53023
rect 17497 53023 17555 53029
rect 17497 53020 17509 53023
rect 16586 52992 17509 53020
rect 16586 52989 16598 52992
rect 16540 52983 16598 52989
rect 17497 52989 17509 52992
rect 17543 53020 17555 53023
rect 17770 53020 17776 53032
rect 17543 52992 17776 53020
rect 17543 52989 17555 52992
rect 17497 52983 17555 52989
rect 17770 52980 17776 52992
rect 17828 52980 17834 53032
rect 18138 53020 18144 53032
rect 18099 52992 18144 53020
rect 18138 52980 18144 52992
rect 18196 52980 18202 53032
rect 18506 53020 18512 53032
rect 18467 52992 18512 53020
rect 18506 52980 18512 52992
rect 18564 52980 18570 53032
rect 18966 53020 18972 53032
rect 18927 52992 18972 53020
rect 18966 52980 18972 52992
rect 19024 52980 19030 53032
rect 20088 53029 20116 53060
rect 20625 53057 20637 53091
rect 20671 53088 20683 53091
rect 20714 53088 20720 53100
rect 20671 53060 20720 53088
rect 20671 53057 20683 53060
rect 20625 53051 20683 53057
rect 20714 53048 20720 53060
rect 20772 53048 20778 53100
rect 23492 53088 23520 53184
rect 23750 53156 23756 53168
rect 23711 53128 23756 53156
rect 23750 53116 23756 53128
rect 23808 53116 23814 53168
rect 23934 53116 23940 53168
rect 23992 53156 23998 53168
rect 23992 53128 24164 53156
rect 23992 53116 23998 53128
rect 24136 53097 24164 53128
rect 24121 53091 24179 53097
rect 23492 53060 23980 53088
rect 20073 53023 20131 53029
rect 20073 52989 20085 53023
rect 20119 53020 20131 53023
rect 20530 53020 20536 53032
rect 20119 52992 20536 53020
rect 20119 52989 20131 52992
rect 20073 52983 20131 52989
rect 20530 52980 20536 52992
rect 20588 52980 20594 53032
rect 21358 53020 21364 53032
rect 21319 52992 21364 53020
rect 21358 52980 21364 52992
rect 21416 52980 21422 53032
rect 22097 53023 22155 53029
rect 22097 52989 22109 53023
rect 22143 52989 22155 53023
rect 22278 53020 22284 53032
rect 22239 52992 22284 53020
rect 22097 52983 22155 52989
rect 15470 52844 15476 52896
rect 15528 52884 15534 52896
rect 15948 52893 15976 52980
rect 22112 52952 22140 52983
rect 22278 52980 22284 52992
rect 22336 52980 22342 53032
rect 23952 53029 23980 53060
rect 24121 53057 24133 53091
rect 24167 53057 24179 53091
rect 24121 53051 24179 53057
rect 25590 53048 25596 53100
rect 25648 53088 25654 53100
rect 25961 53091 26019 53097
rect 25961 53088 25973 53091
rect 25648 53060 25973 53088
rect 25648 53048 25654 53060
rect 25961 53057 25973 53060
rect 26007 53057 26019 53091
rect 25961 53051 26019 53057
rect 23661 53023 23719 53029
rect 23661 53020 23673 53023
rect 23032 52992 23673 53020
rect 22370 52952 22376 52964
rect 22112 52924 22376 52952
rect 22370 52912 22376 52924
rect 22428 52912 22434 52964
rect 15565 52887 15623 52893
rect 15565 52884 15577 52887
rect 15528 52856 15577 52884
rect 15528 52844 15534 52856
rect 15565 52853 15577 52856
rect 15611 52853 15623 52887
rect 15565 52847 15623 52853
rect 15933 52887 15991 52893
rect 15933 52853 15945 52887
rect 15979 52884 15991 52887
rect 16301 52887 16359 52893
rect 16301 52884 16313 52887
rect 15979 52856 16313 52884
rect 15979 52853 15991 52856
rect 15933 52847 15991 52853
rect 16301 52853 16313 52856
rect 16347 52884 16359 52887
rect 17862 52884 17868 52896
rect 16347 52856 17868 52884
rect 16347 52853 16359 52856
rect 16301 52847 16359 52853
rect 17862 52844 17868 52856
rect 17920 52844 17926 52896
rect 18782 52844 18788 52896
rect 18840 52884 18846 52896
rect 20257 52887 20315 52893
rect 20257 52884 20269 52887
rect 18840 52856 20269 52884
rect 18840 52844 18846 52856
rect 20257 52853 20269 52856
rect 20303 52853 20315 52887
rect 20257 52847 20315 52853
rect 22922 52844 22928 52896
rect 22980 52884 22986 52896
rect 23032 52893 23060 52992
rect 23661 52989 23673 52992
rect 23707 52989 23719 53023
rect 23661 52983 23719 52989
rect 23937 53023 23995 53029
rect 23937 52989 23949 53023
rect 23983 52989 23995 53023
rect 25222 53020 25228 53032
rect 23937 52983 23995 52989
rect 24044 52992 25228 53020
rect 24044 52952 24072 52992
rect 25222 52980 25228 52992
rect 25280 52980 25286 53032
rect 26234 53020 26240 53032
rect 25424 52992 26240 53020
rect 23952 52924 24072 52952
rect 23952 52896 23980 52924
rect 23017 52887 23075 52893
rect 23017 52884 23029 52887
rect 22980 52856 23029 52884
rect 22980 52844 22986 52856
rect 23017 52853 23029 52856
rect 23063 52853 23075 52887
rect 23017 52847 23075 52853
rect 23934 52844 23940 52896
rect 23992 52844 23998 52896
rect 24762 52844 24768 52896
rect 24820 52884 24826 52896
rect 25424 52893 25452 52992
rect 26234 52980 26240 52992
rect 26292 52980 26298 53032
rect 26510 52980 26516 53032
rect 26568 53020 26574 53032
rect 26881 53023 26939 53029
rect 26881 53020 26893 53023
rect 26568 52992 26893 53020
rect 26568 52980 26574 52992
rect 26881 52989 26893 52992
rect 26927 53020 26939 53023
rect 27065 53023 27123 53029
rect 27065 53020 27077 53023
rect 26927 52992 27077 53020
rect 26927 52989 26939 52992
rect 26881 52983 26939 52989
rect 27065 52989 27077 52992
rect 27111 52989 27123 53023
rect 27065 52983 27123 52989
rect 27154 52980 27160 53032
rect 27212 53020 27218 53032
rect 27525 53023 27583 53029
rect 27525 53020 27537 53023
rect 27212 52992 27537 53020
rect 27212 52980 27218 52992
rect 27525 52989 27537 52992
rect 27571 53020 27583 53023
rect 28445 53023 28503 53029
rect 28445 53020 28457 53023
rect 27571 52992 28457 53020
rect 27571 52989 27583 52992
rect 27525 52983 27583 52989
rect 28445 52989 28457 52992
rect 28491 52989 28503 53023
rect 28445 52983 28503 52989
rect 25593 52955 25651 52961
rect 25593 52921 25605 52955
rect 25639 52952 25651 52955
rect 25774 52952 25780 52964
rect 25639 52924 25780 52952
rect 25639 52921 25651 52924
rect 25593 52915 25651 52921
rect 25774 52912 25780 52924
rect 25832 52952 25838 52964
rect 26786 52952 26792 52964
rect 25832 52924 26792 52952
rect 25832 52912 25838 52924
rect 26786 52912 26792 52924
rect 26844 52912 26850 52964
rect 25041 52887 25099 52893
rect 25041 52884 25053 52887
rect 24820 52856 25053 52884
rect 24820 52844 24826 52856
rect 25041 52853 25053 52856
rect 25087 52884 25099 52887
rect 25409 52887 25467 52893
rect 25409 52884 25421 52887
rect 25087 52856 25421 52884
rect 25087 52853 25099 52856
rect 25041 52847 25099 52853
rect 25409 52853 25421 52856
rect 25455 52853 25467 52887
rect 25409 52847 25467 52853
rect 25501 52887 25559 52893
rect 25501 52853 25513 52887
rect 25547 52884 25559 52887
rect 26234 52884 26240 52896
rect 25547 52856 26240 52884
rect 25547 52853 25559 52856
rect 25501 52847 25559 52853
rect 26234 52844 26240 52856
rect 26292 52844 26298 52896
rect 26326 52844 26332 52896
rect 26384 52884 26390 52896
rect 26513 52887 26571 52893
rect 26513 52884 26525 52887
rect 26384 52856 26525 52884
rect 26384 52844 26390 52856
rect 26513 52853 26525 52856
rect 26559 52853 26571 52887
rect 27154 52884 27160 52896
rect 27115 52856 27160 52884
rect 26513 52847 26571 52853
rect 27154 52844 27160 52856
rect 27212 52844 27218 52896
rect 27338 52844 27344 52896
rect 27396 52884 27402 52896
rect 28077 52887 28135 52893
rect 28077 52884 28089 52887
rect 27396 52856 28089 52884
rect 27396 52844 27402 52856
rect 28077 52853 28089 52856
rect 28123 52853 28135 52887
rect 28077 52847 28135 52853
rect 1104 52794 38824 52816
rect 1104 52742 19606 52794
rect 19658 52742 19670 52794
rect 19722 52742 19734 52794
rect 19786 52742 19798 52794
rect 19850 52742 38824 52794
rect 1104 52720 38824 52742
rect 14734 52680 14740 52692
rect 14695 52652 14740 52680
rect 14734 52640 14740 52652
rect 14792 52640 14798 52692
rect 16574 52640 16580 52692
rect 16632 52680 16638 52692
rect 16853 52683 16911 52689
rect 16853 52680 16865 52683
rect 16632 52652 16865 52680
rect 16632 52640 16638 52652
rect 16853 52649 16865 52652
rect 16899 52649 16911 52683
rect 18322 52680 18328 52692
rect 18283 52652 18328 52680
rect 16853 52643 16911 52649
rect 18322 52640 18328 52652
rect 18380 52640 18386 52692
rect 20622 52640 20628 52692
rect 20680 52680 20686 52692
rect 21085 52683 21143 52689
rect 21085 52680 21097 52683
rect 20680 52652 21097 52680
rect 20680 52640 20686 52652
rect 21085 52649 21097 52652
rect 21131 52649 21143 52683
rect 21634 52680 21640 52692
rect 21595 52652 21640 52680
rect 21085 52643 21143 52649
rect 21634 52640 21640 52652
rect 21692 52640 21698 52692
rect 23106 52640 23112 52692
rect 23164 52680 23170 52692
rect 23750 52680 23756 52692
rect 23164 52652 23244 52680
rect 23711 52652 23756 52680
rect 23164 52640 23170 52652
rect 15470 52572 15476 52624
rect 15528 52612 15534 52624
rect 15841 52615 15899 52621
rect 15841 52612 15853 52615
rect 15528 52584 15853 52612
rect 15528 52572 15534 52584
rect 15841 52581 15853 52584
rect 15887 52581 15899 52615
rect 16206 52612 16212 52624
rect 16167 52584 16212 52612
rect 15841 52575 15899 52581
rect 16206 52572 16212 52584
rect 16264 52572 16270 52624
rect 16942 52572 16948 52624
rect 17000 52612 17006 52624
rect 17037 52615 17095 52621
rect 17037 52612 17049 52615
rect 17000 52584 17049 52612
rect 17000 52572 17006 52584
rect 17037 52581 17049 52584
rect 17083 52581 17095 52615
rect 17037 52575 17095 52581
rect 20349 52615 20407 52621
rect 20349 52581 20361 52615
rect 20395 52612 20407 52615
rect 20438 52612 20444 52624
rect 20395 52584 20444 52612
rect 20395 52581 20407 52584
rect 20349 52575 20407 52581
rect 20438 52572 20444 52584
rect 20496 52612 20502 52624
rect 20990 52612 20996 52624
rect 20496 52584 20996 52612
rect 20496 52572 20502 52584
rect 20990 52572 20996 52584
rect 21048 52572 21054 52624
rect 22094 52572 22100 52624
rect 22152 52612 22158 52624
rect 22152 52584 23152 52612
rect 22152 52572 22158 52584
rect 9950 52504 9956 52556
rect 10008 52544 10014 52556
rect 10505 52547 10563 52553
rect 10505 52544 10517 52547
rect 10008 52516 10517 52544
rect 10008 52504 10014 52516
rect 10505 52513 10517 52516
rect 10551 52513 10563 52547
rect 10505 52507 10563 52513
rect 10778 52504 10784 52556
rect 10836 52504 10842 52556
rect 15654 52544 15660 52556
rect 15615 52516 15660 52544
rect 15654 52504 15660 52516
rect 15712 52504 15718 52556
rect 15746 52504 15752 52556
rect 15804 52544 15810 52556
rect 16577 52547 16635 52553
rect 15804 52516 15849 52544
rect 15804 52504 15810 52516
rect 16577 52513 16589 52547
rect 16623 52544 16635 52547
rect 16758 52544 16764 52556
rect 16623 52516 16764 52544
rect 16623 52513 16635 52516
rect 16577 52507 16635 52513
rect 10229 52479 10287 52485
rect 10229 52445 10241 52479
rect 10275 52476 10287 52479
rect 10796 52476 10824 52504
rect 11882 52476 11888 52488
rect 10275 52448 10824 52476
rect 11843 52448 11888 52476
rect 10275 52445 10287 52448
rect 10229 52439 10287 52445
rect 11882 52436 11888 52448
rect 11940 52436 11946 52488
rect 15194 52436 15200 52488
rect 15252 52476 15258 52488
rect 15473 52479 15531 52485
rect 15473 52476 15485 52479
rect 15252 52448 15485 52476
rect 15252 52436 15258 52448
rect 15473 52445 15485 52448
rect 15519 52445 15531 52479
rect 15473 52439 15531 52445
rect 15105 52411 15163 52417
rect 15105 52377 15117 52411
rect 15151 52408 15163 52411
rect 16592 52408 16620 52507
rect 16758 52504 16764 52516
rect 16816 52504 16822 52556
rect 17954 52553 17960 52556
rect 17911 52547 17960 52553
rect 17911 52513 17923 52547
rect 17957 52513 17960 52547
rect 17911 52507 17960 52513
rect 17954 52504 17960 52507
rect 18012 52504 18018 52556
rect 18690 52504 18696 52556
rect 18748 52544 18754 52556
rect 18877 52547 18935 52553
rect 18877 52544 18889 52547
rect 18748 52516 18889 52544
rect 18748 52504 18754 52516
rect 18877 52513 18889 52516
rect 18923 52513 18935 52547
rect 19426 52544 19432 52556
rect 19387 52516 19432 52544
rect 18877 52507 18935 52513
rect 19426 52504 19432 52516
rect 19484 52504 19490 52556
rect 19797 52547 19855 52553
rect 19797 52513 19809 52547
rect 19843 52544 19855 52547
rect 19886 52544 19892 52556
rect 19843 52516 19892 52544
rect 19843 52513 19855 52516
rect 19797 52507 19855 52513
rect 19886 52504 19892 52516
rect 19944 52504 19950 52556
rect 20530 52504 20536 52556
rect 20588 52544 20594 52556
rect 20625 52547 20683 52553
rect 20625 52544 20637 52547
rect 20588 52516 20637 52544
rect 20588 52504 20594 52516
rect 20625 52513 20637 52516
rect 20671 52513 20683 52547
rect 20898 52544 20904 52556
rect 20859 52516 20904 52544
rect 20625 52507 20683 52513
rect 20898 52504 20904 52516
rect 20956 52504 20962 52556
rect 22186 52504 22192 52556
rect 22244 52544 22250 52556
rect 23124 52553 23152 52584
rect 22649 52547 22707 52553
rect 22649 52544 22661 52547
rect 22244 52516 22661 52544
rect 22244 52504 22250 52516
rect 22649 52513 22661 52516
rect 22695 52513 22707 52547
rect 22649 52507 22707 52513
rect 23109 52547 23167 52553
rect 23109 52513 23121 52547
rect 23155 52513 23167 52547
rect 23109 52507 23167 52513
rect 17586 52476 17592 52488
rect 17547 52448 17592 52476
rect 17586 52436 17592 52448
rect 17644 52436 17650 52488
rect 17770 52485 17776 52488
rect 17727 52479 17776 52485
rect 17727 52445 17739 52479
rect 17773 52445 17776 52479
rect 17727 52439 17776 52445
rect 17770 52436 17776 52439
rect 17828 52436 17834 52488
rect 19978 52476 19984 52488
rect 19260 52448 19984 52476
rect 15151 52380 16620 52408
rect 15151 52377 15163 52380
rect 15105 52371 15163 52377
rect 18966 52368 18972 52420
rect 19024 52408 19030 52420
rect 19260 52408 19288 52448
rect 19978 52436 19984 52448
rect 20036 52436 20042 52488
rect 20254 52436 20260 52488
rect 20312 52476 20318 52488
rect 20714 52476 20720 52488
rect 20312 52448 20720 52476
rect 20312 52436 20318 52448
rect 20714 52436 20720 52448
rect 20772 52436 20778 52488
rect 22465 52479 22523 52485
rect 22465 52445 22477 52479
rect 22511 52476 22523 52479
rect 23216 52476 23244 52652
rect 23750 52640 23756 52652
rect 23808 52640 23814 52692
rect 23934 52640 23940 52692
rect 23992 52680 23998 52692
rect 24029 52683 24087 52689
rect 24029 52680 24041 52683
rect 23992 52652 24041 52680
rect 23992 52640 23998 52652
rect 24029 52649 24041 52652
rect 24075 52649 24087 52683
rect 24029 52643 24087 52649
rect 25685 52683 25743 52689
rect 25685 52649 25697 52683
rect 25731 52680 25743 52683
rect 25774 52680 25780 52692
rect 25731 52652 25780 52680
rect 25731 52649 25743 52652
rect 25685 52643 25743 52649
rect 25774 52640 25780 52652
rect 25832 52640 25838 52692
rect 28721 52683 28779 52689
rect 28721 52649 28733 52683
rect 28767 52680 28779 52683
rect 29086 52680 29092 52692
rect 28767 52652 29092 52680
rect 28767 52649 28779 52652
rect 28721 52643 28779 52649
rect 24946 52612 24952 52624
rect 24907 52584 24952 52612
rect 24946 52572 24952 52584
rect 25004 52572 25010 52624
rect 27430 52612 27436 52624
rect 27391 52584 27436 52612
rect 27430 52572 27436 52584
rect 27488 52572 27494 52624
rect 24670 52544 24676 52556
rect 24631 52516 24676 52544
rect 24670 52504 24676 52516
rect 24728 52504 24734 52556
rect 25774 52504 25780 52556
rect 25832 52544 25838 52556
rect 25961 52547 26019 52553
rect 25961 52544 25973 52547
rect 25832 52516 25973 52544
rect 25832 52504 25838 52516
rect 25961 52513 25973 52516
rect 26007 52513 26019 52547
rect 25961 52507 26019 52513
rect 27522 52504 27528 52556
rect 27580 52544 27586 52556
rect 28169 52547 28227 52553
rect 28169 52544 28181 52547
rect 27580 52516 28181 52544
rect 27580 52504 27586 52516
rect 28169 52513 28181 52516
rect 28215 52544 28227 52547
rect 28736 52544 28764 52643
rect 29086 52640 29092 52652
rect 29144 52640 29150 52692
rect 29454 52544 29460 52556
rect 28215 52516 28764 52544
rect 29415 52516 29460 52544
rect 28215 52513 28227 52516
rect 28169 52507 28227 52513
rect 29454 52504 29460 52516
rect 29512 52504 29518 52556
rect 29546 52504 29552 52556
rect 29604 52504 29610 52556
rect 22511 52448 23244 52476
rect 22511 52445 22523 52448
rect 22465 52439 22523 52445
rect 24486 52436 24492 52488
rect 24544 52476 24550 52488
rect 24544 52448 24900 52476
rect 24544 52436 24550 52448
rect 19024 52380 19288 52408
rect 19024 52368 19030 52380
rect 19334 52368 19340 52420
rect 19392 52408 19398 52420
rect 19705 52411 19763 52417
rect 19705 52408 19717 52411
rect 19392 52380 19717 52408
rect 19392 52368 19398 52380
rect 19705 52377 19717 52380
rect 19751 52377 19763 52411
rect 19996 52408 20024 52436
rect 19996 52380 22324 52408
rect 19705 52371 19763 52377
rect 16942 52300 16948 52352
rect 17000 52340 17006 52352
rect 18138 52340 18144 52352
rect 17000 52312 18144 52340
rect 17000 52300 17006 52312
rect 18138 52300 18144 52312
rect 18196 52340 18202 52352
rect 18693 52343 18751 52349
rect 18693 52340 18705 52343
rect 18196 52312 18705 52340
rect 18196 52300 18202 52312
rect 18693 52309 18705 52312
rect 18739 52340 18751 52343
rect 18782 52340 18788 52352
rect 18739 52312 18788 52340
rect 18739 52309 18751 52312
rect 18693 52303 18751 52309
rect 18782 52300 18788 52312
rect 18840 52300 18846 52352
rect 22094 52300 22100 52352
rect 22152 52340 22158 52352
rect 22296 52340 22324 52380
rect 22830 52368 22836 52420
rect 22888 52408 22894 52420
rect 23109 52411 23167 52417
rect 23109 52408 23121 52411
rect 22888 52380 23121 52408
rect 22888 52368 22894 52380
rect 23109 52377 23121 52380
rect 23155 52377 23167 52411
rect 24872 52408 24900 52448
rect 27154 52436 27160 52488
rect 27212 52476 27218 52488
rect 27341 52479 27399 52485
rect 27341 52476 27353 52479
rect 27212 52448 27353 52476
rect 27212 52436 27218 52448
rect 27341 52445 27353 52448
rect 27387 52476 27399 52479
rect 28258 52476 28264 52488
rect 27387 52448 27660 52476
rect 28219 52448 28264 52476
rect 27387 52445 27399 52448
rect 27341 52439 27399 52445
rect 24946 52408 24952 52420
rect 24872 52380 24952 52408
rect 23109 52371 23167 52377
rect 24946 52368 24952 52380
rect 25004 52368 25010 52420
rect 27632 52408 27660 52448
rect 28258 52436 28264 52448
rect 28316 52436 28322 52488
rect 29181 52479 29239 52485
rect 29181 52445 29193 52479
rect 29227 52476 29239 52479
rect 29564 52476 29592 52504
rect 30282 52476 30288 52488
rect 29227 52448 30288 52476
rect 29227 52445 29239 52448
rect 29181 52439 29239 52445
rect 30282 52436 30288 52448
rect 30340 52436 30346 52488
rect 30742 52476 30748 52488
rect 30703 52448 30748 52476
rect 30742 52436 30748 52448
rect 30800 52436 30806 52488
rect 34698 52436 34704 52488
rect 34756 52476 34762 52488
rect 35802 52476 35808 52488
rect 34756 52448 35808 52476
rect 34756 52436 34762 52448
rect 35802 52436 35808 52448
rect 35860 52436 35866 52488
rect 28350 52408 28356 52420
rect 27632 52380 28356 52408
rect 28350 52368 28356 52380
rect 28408 52368 28414 52420
rect 25225 52343 25283 52349
rect 25225 52340 25237 52343
rect 22152 52312 22197 52340
rect 22296 52312 25237 52340
rect 22152 52300 22158 52312
rect 25225 52309 25237 52312
rect 25271 52340 25283 52343
rect 26234 52340 26240 52352
rect 25271 52312 26240 52340
rect 25271 52309 25283 52312
rect 25225 52303 25283 52309
rect 26234 52300 26240 52312
rect 26292 52300 26298 52352
rect 26786 52340 26792 52352
rect 26747 52312 26792 52340
rect 26786 52300 26792 52312
rect 26844 52300 26850 52352
rect 26878 52300 26884 52352
rect 26936 52340 26942 52352
rect 27065 52343 27123 52349
rect 27065 52340 27077 52343
rect 26936 52312 27077 52340
rect 26936 52300 26942 52312
rect 27065 52309 27077 52312
rect 27111 52309 27123 52343
rect 27065 52303 27123 52309
rect 1104 52250 38824 52272
rect 1104 52198 4246 52250
rect 4298 52198 4310 52250
rect 4362 52198 4374 52250
rect 4426 52198 4438 52250
rect 4490 52198 34966 52250
rect 35018 52198 35030 52250
rect 35082 52198 35094 52250
rect 35146 52198 35158 52250
rect 35210 52198 38824 52250
rect 1104 52176 38824 52198
rect 9950 52096 9956 52148
rect 10008 52136 10014 52148
rect 10229 52139 10287 52145
rect 10229 52136 10241 52139
rect 10008 52108 10241 52136
rect 10008 52096 10014 52108
rect 10229 52105 10241 52108
rect 10275 52105 10287 52139
rect 10229 52099 10287 52105
rect 10689 52139 10747 52145
rect 10689 52105 10701 52139
rect 10735 52136 10747 52139
rect 10778 52136 10784 52148
rect 10735 52108 10784 52136
rect 10735 52105 10747 52108
rect 10689 52099 10747 52105
rect 10778 52096 10784 52108
rect 10836 52096 10842 52148
rect 15194 52096 15200 52148
rect 15252 52136 15258 52148
rect 15473 52139 15531 52145
rect 15473 52136 15485 52139
rect 15252 52108 15485 52136
rect 15252 52096 15258 52108
rect 15473 52105 15485 52108
rect 15519 52105 15531 52139
rect 15473 52099 15531 52105
rect 15654 52096 15660 52148
rect 15712 52136 15718 52148
rect 15841 52139 15899 52145
rect 15841 52136 15853 52139
rect 15712 52108 15853 52136
rect 15712 52096 15718 52108
rect 15841 52105 15853 52108
rect 15887 52105 15899 52139
rect 15841 52099 15899 52105
rect 18690 52096 18696 52148
rect 18748 52136 18754 52148
rect 19058 52136 19064 52148
rect 18748 52108 19064 52136
rect 18748 52096 18754 52108
rect 19058 52096 19064 52108
rect 19116 52096 19122 52148
rect 20898 52096 20904 52148
rect 20956 52136 20962 52148
rect 20993 52139 21051 52145
rect 20993 52136 21005 52139
rect 20956 52108 21005 52136
rect 20956 52096 20962 52108
rect 20993 52105 21005 52108
rect 21039 52105 21051 52139
rect 20993 52099 21051 52105
rect 23017 52139 23075 52145
rect 23017 52105 23029 52139
rect 23063 52136 23075 52139
rect 23106 52136 23112 52148
rect 23063 52108 23112 52136
rect 23063 52105 23075 52108
rect 23017 52099 23075 52105
rect 23106 52096 23112 52108
rect 23164 52096 23170 52148
rect 23290 52096 23296 52148
rect 23348 52136 23354 52148
rect 24121 52139 24179 52145
rect 24121 52136 24133 52139
rect 23348 52108 24133 52136
rect 23348 52096 23354 52108
rect 24121 52105 24133 52108
rect 24167 52105 24179 52139
rect 25130 52136 25136 52148
rect 25091 52108 25136 52136
rect 24121 52099 24179 52105
rect 25130 52096 25136 52108
rect 25188 52096 25194 52148
rect 25498 52136 25504 52148
rect 25459 52108 25504 52136
rect 25498 52096 25504 52108
rect 25556 52096 25562 52148
rect 27706 52136 27712 52148
rect 27619 52108 27712 52136
rect 27706 52096 27712 52108
rect 27764 52136 27770 52148
rect 28258 52136 28264 52148
rect 27764 52108 28264 52136
rect 27764 52096 27770 52108
rect 28258 52096 28264 52108
rect 28316 52096 28322 52148
rect 29454 52096 29460 52148
rect 29512 52136 29518 52148
rect 29733 52139 29791 52145
rect 29733 52136 29745 52139
rect 29512 52108 29745 52136
rect 29512 52096 29518 52108
rect 29733 52105 29745 52108
rect 29779 52105 29791 52139
rect 29733 52099 29791 52105
rect 14461 52071 14519 52077
rect 14461 52037 14473 52071
rect 14507 52068 14519 52071
rect 17954 52068 17960 52080
rect 14507 52040 17960 52068
rect 14507 52037 14519 52040
rect 14461 52031 14519 52037
rect 17954 52028 17960 52040
rect 18012 52028 18018 52080
rect 22278 52068 22284 52080
rect 22239 52040 22284 52068
rect 22278 52028 22284 52040
rect 22336 52028 22342 52080
rect 23661 52071 23719 52077
rect 23661 52037 23673 52071
rect 23707 52068 23719 52071
rect 23934 52068 23940 52080
rect 23707 52040 23940 52068
rect 23707 52037 23719 52040
rect 23661 52031 23719 52037
rect 23934 52028 23940 52040
rect 23992 52028 23998 52080
rect 16114 52000 16120 52012
rect 16075 51972 16120 52000
rect 16114 51960 16120 51972
rect 16172 51960 16178 52012
rect 16666 52000 16672 52012
rect 16627 51972 16672 52000
rect 16666 51960 16672 51972
rect 16724 51960 16730 52012
rect 18049 52003 18107 52009
rect 18049 51969 18061 52003
rect 18095 52000 18107 52003
rect 18322 52000 18328 52012
rect 18095 51972 18328 52000
rect 18095 51969 18107 51972
rect 18049 51963 18107 51969
rect 18322 51960 18328 51972
rect 18380 51960 18386 52012
rect 18785 52003 18843 52009
rect 18785 51969 18797 52003
rect 18831 52000 18843 52003
rect 22296 52000 22324 52028
rect 24118 52000 24124 52012
rect 18831 51972 21588 52000
rect 22296 51972 24124 52000
rect 18831 51969 18843 51972
rect 18785 51963 18843 51969
rect 21560 51944 21588 51972
rect 24118 51960 24124 51972
rect 24176 51960 24182 52012
rect 24854 51960 24860 52012
rect 24912 51960 24918 52012
rect 25148 52000 25176 52096
rect 27614 52028 27620 52080
rect 27672 52068 27678 52080
rect 28353 52071 28411 52077
rect 28353 52068 28365 52071
rect 27672 52040 28365 52068
rect 27672 52028 27678 52040
rect 28353 52037 28365 52040
rect 28399 52037 28411 52071
rect 28353 52031 28411 52037
rect 27338 52000 27344 52012
rect 25148 51972 25360 52000
rect 27299 51972 27344 52000
rect 14829 51935 14887 51941
rect 14829 51901 14841 51935
rect 14875 51932 14887 51935
rect 16942 51932 16948 51944
rect 14875 51904 16948 51932
rect 14875 51901 14887 51904
rect 14829 51895 14887 51901
rect 16942 51892 16948 51904
rect 17000 51892 17006 51944
rect 17129 51935 17187 51941
rect 17129 51901 17141 51935
rect 17175 51932 17187 51935
rect 17770 51932 17776 51944
rect 17175 51904 17776 51932
rect 17175 51901 17187 51904
rect 17129 51895 17187 51901
rect 17770 51892 17776 51904
rect 17828 51892 17834 51944
rect 18233 51935 18291 51941
rect 18233 51901 18245 51935
rect 18279 51932 18291 51935
rect 18598 51932 18604 51944
rect 18279 51904 18604 51932
rect 18279 51901 18291 51904
rect 18233 51895 18291 51901
rect 18598 51892 18604 51904
rect 18656 51932 18662 51944
rect 19150 51932 19156 51944
rect 18656 51904 19156 51932
rect 18656 51892 18662 51904
rect 19150 51892 19156 51904
rect 19208 51892 19214 51944
rect 19521 51935 19579 51941
rect 19521 51901 19533 51935
rect 19567 51932 19579 51935
rect 19889 51935 19947 51941
rect 19889 51932 19901 51935
rect 19567 51904 19901 51932
rect 19567 51901 19579 51904
rect 19521 51895 19579 51901
rect 19889 51901 19901 51904
rect 19935 51932 19947 51935
rect 19978 51932 19984 51944
rect 19935 51904 19984 51932
rect 19935 51901 19947 51904
rect 19889 51895 19947 51901
rect 19978 51892 19984 51904
rect 20036 51892 20042 51944
rect 20254 51932 20260 51944
rect 20215 51904 20260 51932
rect 20254 51892 20260 51904
rect 20312 51892 20318 51944
rect 20438 51932 20444 51944
rect 20399 51904 20444 51932
rect 20438 51892 20444 51904
rect 20496 51892 20502 51944
rect 21542 51932 21548 51944
rect 21455 51904 21548 51932
rect 21542 51892 21548 51904
rect 21600 51892 21606 51944
rect 22370 51932 22376 51944
rect 22331 51904 22376 51932
rect 22370 51892 22376 51904
rect 22428 51892 22434 51944
rect 22554 51932 22560 51944
rect 22515 51904 22560 51932
rect 22554 51892 22560 51904
rect 22612 51892 22618 51944
rect 23474 51932 23480 51944
rect 23387 51904 23480 51932
rect 23474 51892 23480 51904
rect 23532 51932 23538 51944
rect 23937 51935 23995 51941
rect 23937 51932 23949 51935
rect 23532 51904 23949 51932
rect 23532 51892 23538 51904
rect 23937 51901 23949 51904
rect 23983 51901 23995 51935
rect 24872 51932 24900 51960
rect 25332 51941 25360 51972
rect 27338 51960 27344 51972
rect 27396 51960 27402 52012
rect 30193 52003 30251 52009
rect 30193 51969 30205 52003
rect 30239 52000 30251 52003
rect 30558 52000 30564 52012
rect 30239 51972 30564 52000
rect 30239 51969 30251 51972
rect 30193 51963 30251 51969
rect 30558 51960 30564 51972
rect 30616 51960 30622 52012
rect 25225 51935 25283 51941
rect 25225 51932 25237 51935
rect 24872 51904 25237 51932
rect 23937 51895 23995 51901
rect 25225 51901 25237 51904
rect 25271 51901 25283 51935
rect 25225 51895 25283 51901
rect 25317 51935 25375 51941
rect 25317 51901 25329 51935
rect 25363 51901 25375 51935
rect 26786 51932 26792 51944
rect 26747 51904 26792 51932
rect 25317 51895 25375 51901
rect 17862 51864 17868 51876
rect 17775 51836 17868 51864
rect 17862 51824 17868 51836
rect 17920 51864 17926 51876
rect 18414 51864 18420 51876
rect 17920 51836 18420 51864
rect 17920 51824 17926 51836
rect 18414 51824 18420 51836
rect 18472 51824 18478 51876
rect 19242 51824 19248 51876
rect 19300 51864 19306 51876
rect 19300 51836 19748 51864
rect 19300 51824 19306 51836
rect 15197 51799 15255 51805
rect 15197 51765 15209 51799
rect 15243 51796 15255 51799
rect 15746 51796 15752 51808
rect 15243 51768 15752 51796
rect 15243 51765 15255 51768
rect 15197 51759 15255 51765
rect 15746 51756 15752 51768
rect 15804 51796 15810 51808
rect 17497 51799 17555 51805
rect 17497 51796 17509 51799
rect 15804 51768 17509 51796
rect 15804 51756 15810 51768
rect 17497 51765 17509 51768
rect 17543 51796 17555 51799
rect 18325 51799 18383 51805
rect 18325 51796 18337 51799
rect 17543 51768 18337 51796
rect 17543 51765 17555 51768
rect 17497 51759 17555 51765
rect 18325 51765 18337 51768
rect 18371 51796 18383 51799
rect 18966 51796 18972 51808
rect 18371 51768 18972 51796
rect 18371 51765 18383 51768
rect 18325 51759 18383 51765
rect 18966 51756 18972 51768
rect 19024 51756 19030 51808
rect 19720 51805 19748 51836
rect 21634 51824 21640 51876
rect 21692 51864 21698 51876
rect 22572 51864 22600 51892
rect 21692 51836 22600 51864
rect 21692 51824 21698 51836
rect 23290 51824 23296 51876
rect 23348 51864 23354 51876
rect 23845 51867 23903 51873
rect 23845 51864 23857 51867
rect 23348 51836 23857 51864
rect 23348 51824 23354 51836
rect 23845 51833 23857 51836
rect 23891 51833 23903 51867
rect 23952 51864 23980 51895
rect 25240 51864 25268 51895
rect 26786 51892 26792 51904
rect 26844 51892 26850 51944
rect 26878 51892 26884 51944
rect 26936 51932 26942 51944
rect 26936 51904 26981 51932
rect 26936 51892 26942 51904
rect 28074 51892 28080 51944
rect 28132 51932 28138 51944
rect 28169 51935 28227 51941
rect 28169 51932 28181 51935
rect 28132 51904 28181 51932
rect 28132 51892 28138 51904
rect 28169 51901 28181 51904
rect 28215 51932 28227 51935
rect 28629 51935 28687 51941
rect 28629 51932 28641 51935
rect 28215 51904 28641 51932
rect 28215 51901 28227 51904
rect 28169 51895 28227 51901
rect 28629 51901 28641 51904
rect 28675 51901 28687 51935
rect 29086 51932 29092 51944
rect 28999 51904 29092 51932
rect 28629 51895 28687 51901
rect 29086 51892 29092 51904
rect 29144 51932 29150 51944
rect 29273 51935 29331 51941
rect 29273 51932 29285 51935
rect 29144 51904 29285 51932
rect 29144 51892 29150 51904
rect 29273 51901 29285 51904
rect 29319 51901 29331 51935
rect 30282 51932 30288 51944
rect 30243 51904 30288 51932
rect 29273 51895 29331 51901
rect 30282 51892 30288 51904
rect 30340 51892 30346 51944
rect 25774 51864 25780 51876
rect 23952 51836 25176 51864
rect 25240 51836 25780 51864
rect 23845 51827 23903 51833
rect 19705 51799 19763 51805
rect 19705 51765 19717 51799
rect 19751 51765 19763 51799
rect 21450 51796 21456 51808
rect 21363 51768 21456 51796
rect 19705 51759 19763 51765
rect 21450 51756 21456 51768
rect 21508 51796 21514 51808
rect 22186 51796 22192 51808
rect 21508 51768 22192 51796
rect 21508 51756 21514 51768
rect 22186 51756 22192 51768
rect 22244 51756 22250 51808
rect 24670 51796 24676 51808
rect 24631 51768 24676 51796
rect 24670 51756 24676 51768
rect 24728 51756 24734 51808
rect 25148 51796 25176 51836
rect 25774 51824 25780 51836
rect 25832 51864 25838 51876
rect 26053 51867 26111 51873
rect 26053 51864 26065 51867
rect 25832 51836 26065 51864
rect 25832 51824 25838 51836
rect 26053 51833 26065 51836
rect 26099 51833 26111 51867
rect 26053 51827 26111 51833
rect 26605 51867 26663 51873
rect 26605 51833 26617 51867
rect 26651 51833 26663 51867
rect 26605 51827 26663 51833
rect 26973 51867 27031 51873
rect 26973 51833 26985 51867
rect 27019 51864 27031 51867
rect 27522 51864 27528 51876
rect 27019 51836 27528 51864
rect 27019 51833 27031 51836
rect 26973 51827 27031 51833
rect 25314 51796 25320 51808
rect 25148 51768 25320 51796
rect 25314 51756 25320 51768
rect 25372 51756 25378 51808
rect 26234 51756 26240 51808
rect 26292 51796 26298 51808
rect 26421 51799 26479 51805
rect 26421 51796 26433 51799
rect 26292 51768 26433 51796
rect 26292 51756 26298 51768
rect 26421 51765 26433 51768
rect 26467 51796 26479 51799
rect 26620 51796 26648 51827
rect 27522 51824 27528 51836
rect 27580 51824 27586 51876
rect 26467 51768 26648 51796
rect 28077 51799 28135 51805
rect 26467 51765 26479 51768
rect 26421 51759 26479 51765
rect 28077 51765 28089 51799
rect 28123 51796 28135 51799
rect 28258 51796 28264 51808
rect 28123 51768 28264 51796
rect 28123 51765 28135 51768
rect 28077 51759 28135 51765
rect 28258 51756 28264 51768
rect 28316 51756 28322 51808
rect 28994 51756 29000 51808
rect 29052 51796 29058 51808
rect 29457 51799 29515 51805
rect 29457 51796 29469 51799
rect 29052 51768 29469 51796
rect 29052 51756 29058 51768
rect 29457 51765 29469 51768
rect 29503 51765 29515 51799
rect 29457 51759 29515 51765
rect 31754 51756 31760 51808
rect 31812 51796 31818 51808
rect 31849 51799 31907 51805
rect 31849 51796 31861 51799
rect 31812 51768 31861 51796
rect 31812 51756 31818 51768
rect 31849 51765 31861 51768
rect 31895 51765 31907 51799
rect 31849 51759 31907 51765
rect 1104 51706 38824 51728
rect 1104 51654 19606 51706
rect 19658 51654 19670 51706
rect 19722 51654 19734 51706
rect 19786 51654 19798 51706
rect 19850 51654 38824 51706
rect 1104 51632 38824 51654
rect 15102 51592 15108 51604
rect 15063 51564 15108 51592
rect 15102 51552 15108 51564
rect 15160 51552 15166 51604
rect 15470 51592 15476 51604
rect 15431 51564 15476 51592
rect 15470 51552 15476 51564
rect 15528 51552 15534 51604
rect 18509 51595 18567 51601
rect 18509 51561 18521 51595
rect 18555 51592 18567 51595
rect 18598 51592 18604 51604
rect 18555 51564 18604 51592
rect 18555 51561 18567 51564
rect 18509 51555 18567 51561
rect 18598 51552 18604 51564
rect 18656 51552 18662 51604
rect 18782 51592 18788 51604
rect 18743 51564 18788 51592
rect 18782 51552 18788 51564
rect 18840 51552 18846 51604
rect 20254 51592 20260 51604
rect 20215 51564 20260 51592
rect 20254 51552 20260 51564
rect 20312 51592 20318 51604
rect 20530 51592 20536 51604
rect 20312 51564 20536 51592
rect 20312 51552 20318 51564
rect 20530 51552 20536 51564
rect 20588 51552 20594 51604
rect 21358 51592 21364 51604
rect 21319 51564 21364 51592
rect 21358 51552 21364 51564
rect 21416 51552 21422 51604
rect 21818 51592 21824 51604
rect 21779 51564 21824 51592
rect 21818 51552 21824 51564
rect 21876 51592 21882 51604
rect 22002 51592 22008 51604
rect 21876 51564 22008 51592
rect 21876 51552 21882 51564
rect 22002 51552 22008 51564
rect 22060 51552 22066 51604
rect 23290 51592 23296 51604
rect 23251 51564 23296 51592
rect 23290 51552 23296 51564
rect 23348 51552 23354 51604
rect 24854 51552 24860 51604
rect 24912 51592 24918 51604
rect 25869 51595 25927 51601
rect 25869 51592 25881 51595
rect 24912 51564 25881 51592
rect 24912 51552 24918 51564
rect 25869 51561 25881 51564
rect 25915 51561 25927 51595
rect 25869 51555 25927 51561
rect 26878 51552 26884 51604
rect 26936 51592 26942 51604
rect 27893 51595 27951 51601
rect 27893 51592 27905 51595
rect 26936 51564 27905 51592
rect 26936 51552 26942 51564
rect 27893 51561 27905 51564
rect 27939 51592 27951 51595
rect 27982 51592 27988 51604
rect 27939 51564 27988 51592
rect 27939 51561 27951 51564
rect 27893 51555 27951 51561
rect 27982 51552 27988 51564
rect 28040 51552 28046 51604
rect 30282 51552 30288 51604
rect 30340 51592 30346 51604
rect 30650 51592 30656 51604
rect 30340 51564 30656 51592
rect 30340 51552 30346 51564
rect 30650 51552 30656 51564
rect 30708 51552 30714 51604
rect 14918 51484 14924 51536
rect 14976 51524 14982 51536
rect 15841 51527 15899 51533
rect 15841 51524 15853 51527
rect 14976 51496 15853 51524
rect 14976 51484 14982 51496
rect 15841 51493 15853 51496
rect 15887 51493 15899 51527
rect 16577 51527 16635 51533
rect 16577 51524 16589 51527
rect 15841 51487 15899 51493
rect 16040 51496 16589 51524
rect 15856 51388 15884 51487
rect 16040 51468 16068 51496
rect 16577 51493 16589 51496
rect 16623 51524 16635 51527
rect 16945 51527 17003 51533
rect 16945 51524 16957 51527
rect 16623 51496 16957 51524
rect 16623 51493 16635 51496
rect 16577 51487 16635 51493
rect 16945 51493 16957 51496
rect 16991 51524 17003 51527
rect 17770 51524 17776 51536
rect 16991 51496 17776 51524
rect 16991 51493 17003 51496
rect 16945 51487 17003 51493
rect 17770 51484 17776 51496
rect 17828 51484 17834 51536
rect 20070 51484 20076 51536
rect 20128 51524 20134 51536
rect 21174 51524 21180 51536
rect 20128 51496 21180 51524
rect 20128 51484 20134 51496
rect 21174 51484 21180 51496
rect 21232 51484 21238 51536
rect 22370 51524 22376 51536
rect 21376 51496 22376 51524
rect 16022 51456 16028 51468
rect 15935 51428 16028 51456
rect 16022 51416 16028 51428
rect 16080 51416 16086 51468
rect 17402 51456 17408 51468
rect 17363 51428 17408 51456
rect 17402 51416 17408 51428
rect 17460 51416 17466 51468
rect 17862 51456 17868 51468
rect 17823 51428 17868 51456
rect 17862 51416 17868 51428
rect 17920 51416 17926 51468
rect 19797 51459 19855 51465
rect 19797 51425 19809 51459
rect 19843 51456 19855 51459
rect 20898 51456 20904 51468
rect 19843 51428 19932 51456
rect 20859 51428 20904 51456
rect 19843 51425 19855 51428
rect 19797 51419 19855 51425
rect 16574 51388 16580 51400
rect 15856 51360 16580 51388
rect 16574 51348 16580 51360
rect 16632 51348 16638 51400
rect 17221 51391 17279 51397
rect 17221 51357 17233 51391
rect 17267 51388 17279 51391
rect 17494 51388 17500 51400
rect 17267 51360 17500 51388
rect 17267 51357 17279 51360
rect 17221 51351 17279 51357
rect 17494 51348 17500 51360
rect 17552 51348 17558 51400
rect 18966 51388 18972 51400
rect 18927 51360 18972 51388
rect 18966 51348 18972 51360
rect 19024 51348 19030 51400
rect 19518 51388 19524 51400
rect 19479 51360 19524 51388
rect 19518 51348 19524 51360
rect 19576 51348 19582 51400
rect 17954 51320 17960 51332
rect 17915 51292 17960 51320
rect 17954 51280 17960 51292
rect 18012 51280 18018 51332
rect 19794 51280 19800 51332
rect 19852 51320 19858 51332
rect 19904 51320 19932 51428
rect 20898 51416 20904 51428
rect 20956 51416 20962 51468
rect 21376 51400 21404 51496
rect 22370 51484 22376 51496
rect 22428 51484 22434 51536
rect 22554 51484 22560 51536
rect 22612 51524 22618 51536
rect 24581 51527 24639 51533
rect 24581 51524 24593 51527
rect 22612 51496 24593 51524
rect 22612 51484 22618 51496
rect 24581 51493 24593 51496
rect 24627 51524 24639 51527
rect 26237 51527 26295 51533
rect 26237 51524 26249 51527
rect 24627 51496 26249 51524
rect 24627 51493 24639 51496
rect 24581 51487 24639 51493
rect 26237 51493 26249 51496
rect 26283 51493 26295 51527
rect 27246 51524 27252 51536
rect 27207 51496 27252 51524
rect 26237 51487 26295 51493
rect 27246 51484 27252 51496
rect 27304 51484 27310 51536
rect 29086 51484 29092 51536
rect 29144 51524 29150 51536
rect 29144 51496 30236 51524
rect 29144 51484 29150 51496
rect 30208 51468 30236 51496
rect 21726 51416 21732 51468
rect 21784 51456 21790 51468
rect 21913 51459 21971 51465
rect 21913 51456 21925 51459
rect 21784 51428 21925 51456
rect 21784 51416 21790 51428
rect 21913 51425 21925 51428
rect 21959 51425 21971 51459
rect 21913 51419 21971 51425
rect 19978 51348 19984 51400
rect 20036 51388 20042 51400
rect 20717 51391 20775 51397
rect 20036 51360 20081 51388
rect 20036 51348 20042 51360
rect 20717 51357 20729 51391
rect 20763 51388 20775 51391
rect 21358 51388 21364 51400
rect 20763 51360 21364 51388
rect 20763 51357 20775 51360
rect 20717 51351 20775 51357
rect 21358 51348 21364 51360
rect 21416 51348 21422 51400
rect 21085 51323 21143 51329
rect 21085 51320 21097 51323
rect 19852 51292 21097 51320
rect 19852 51280 19858 51292
rect 21085 51289 21097 51292
rect 21131 51289 21143 51323
rect 21928 51320 21956 51419
rect 22002 51416 22008 51468
rect 22060 51456 22066 51468
rect 22281 51459 22339 51465
rect 22281 51456 22293 51459
rect 22060 51428 22293 51456
rect 22060 51416 22066 51428
rect 22281 51425 22293 51428
rect 22327 51425 22339 51459
rect 22281 51419 22339 51425
rect 22741 51459 22799 51465
rect 22741 51425 22753 51459
rect 22787 51425 22799 51459
rect 23934 51456 23940 51468
rect 23895 51428 23940 51456
rect 22741 51419 22799 51425
rect 22094 51348 22100 51400
rect 22152 51388 22158 51400
rect 22756 51388 22784 51419
rect 23934 51416 23940 51428
rect 23992 51416 23998 51468
rect 24029 51459 24087 51465
rect 24029 51425 24041 51459
rect 24075 51425 24087 51459
rect 24029 51419 24087 51425
rect 24121 51459 24179 51465
rect 24121 51425 24133 51459
rect 24167 51456 24179 51459
rect 24302 51456 24308 51468
rect 24167 51428 24308 51456
rect 24167 51425 24179 51428
rect 24121 51419 24179 51425
rect 22152 51360 22784 51388
rect 23017 51391 23075 51397
rect 22152 51348 22158 51360
rect 23017 51357 23029 51391
rect 23063 51388 23075 51391
rect 23106 51388 23112 51400
rect 23063 51360 23112 51388
rect 23063 51357 23075 51360
rect 23017 51351 23075 51357
rect 23106 51348 23112 51360
rect 23164 51348 23170 51400
rect 24044 51388 24072 51419
rect 24302 51416 24308 51428
rect 24360 51416 24366 51468
rect 24946 51456 24952 51468
rect 24907 51428 24952 51456
rect 24946 51416 24952 51428
rect 25004 51416 25010 51468
rect 25038 51416 25044 51468
rect 25096 51456 25102 51468
rect 25225 51459 25283 51465
rect 25225 51456 25237 51459
rect 25096 51428 25237 51456
rect 25096 51416 25102 51428
rect 25225 51425 25237 51428
rect 25271 51425 25283 51459
rect 25225 51419 25283 51425
rect 25314 51416 25320 51468
rect 25372 51456 25378 51468
rect 25409 51459 25467 51465
rect 25409 51456 25421 51459
rect 25372 51428 25421 51456
rect 25372 51416 25378 51428
rect 25409 51425 25421 51428
rect 25455 51425 25467 51459
rect 25409 51419 25467 51425
rect 26789 51459 26847 51465
rect 26789 51425 26801 51459
rect 26835 51425 26847 51459
rect 26970 51456 26976 51468
rect 26931 51428 26976 51456
rect 26789 51419 26847 51425
rect 24762 51388 24768 51400
rect 23676 51360 24768 51388
rect 22278 51320 22284 51332
rect 21928 51292 22284 51320
rect 21085 51283 21143 51289
rect 22278 51280 22284 51292
rect 22336 51280 22342 51332
rect 14734 51252 14740 51264
rect 14695 51224 14740 51252
rect 14734 51212 14740 51224
rect 14792 51212 14798 51264
rect 16206 51252 16212 51264
rect 16167 51224 16212 51252
rect 16206 51212 16212 51224
rect 16264 51212 16270 51264
rect 21726 51212 21732 51264
rect 21784 51252 21790 51264
rect 23676 51261 23704 51360
rect 24762 51348 24768 51360
rect 24820 51348 24826 51400
rect 26804 51388 26832 51419
rect 26970 51416 26976 51428
rect 27028 51416 27034 51468
rect 29181 51459 29239 51465
rect 29181 51425 29193 51459
rect 29227 51425 29239 51459
rect 29181 51419 29239 51425
rect 29273 51459 29331 51465
rect 29273 51425 29285 51459
rect 29319 51456 29331 51459
rect 29546 51456 29552 51468
rect 29319 51428 29552 51456
rect 29319 51425 29331 51428
rect 29273 51419 29331 51425
rect 26878 51388 26884 51400
rect 26804 51360 26884 51388
rect 26878 51348 26884 51360
rect 26936 51348 26942 51400
rect 28350 51388 28356 51400
rect 28311 51360 28356 51388
rect 28350 51348 28356 51360
rect 28408 51348 28414 51400
rect 28442 51348 28448 51400
rect 28500 51388 28506 51400
rect 28500 51360 28545 51388
rect 28500 51348 28506 51360
rect 29196 51320 29224 51419
rect 29546 51416 29552 51428
rect 29604 51416 29610 51468
rect 30190 51456 30196 51468
rect 30103 51428 30196 51456
rect 30190 51416 30196 51428
rect 30248 51416 30254 51468
rect 31386 51456 31392 51468
rect 31347 51428 31392 51456
rect 31386 51416 31392 51428
rect 31444 51416 31450 51468
rect 33686 51416 33692 51468
rect 33744 51456 33750 51468
rect 33873 51459 33931 51465
rect 33873 51456 33885 51459
rect 33744 51428 33885 51456
rect 33744 51416 33750 51428
rect 33873 51425 33885 51428
rect 33919 51425 33931 51459
rect 33873 51419 33931 51425
rect 29733 51323 29791 51329
rect 29733 51320 29745 51323
rect 29196 51292 29745 51320
rect 29733 51289 29745 51292
rect 29779 51320 29791 51323
rect 30282 51320 30288 51332
rect 29779 51292 30288 51320
rect 29779 51289 29791 51292
rect 29733 51283 29791 51289
rect 30282 51280 30288 51292
rect 30340 51280 30346 51332
rect 23661 51255 23719 51261
rect 23661 51252 23673 51255
rect 21784 51224 23673 51252
rect 21784 51212 21790 51224
rect 23661 51221 23673 51224
rect 23707 51221 23719 51255
rect 23661 51215 23719 51221
rect 25593 51255 25651 51261
rect 25593 51221 25605 51255
rect 25639 51252 25651 51255
rect 26326 51252 26332 51264
rect 25639 51224 26332 51252
rect 25639 51221 25651 51224
rect 25593 51215 25651 51221
rect 26326 51212 26332 51224
rect 26384 51212 26390 51264
rect 27522 51252 27528 51264
rect 27483 51224 27528 51252
rect 27522 51212 27528 51224
rect 27580 51212 27586 51264
rect 28902 51212 28908 51264
rect 28960 51252 28966 51264
rect 29546 51252 29552 51264
rect 28960 51224 29552 51252
rect 28960 51212 28966 51224
rect 29546 51212 29552 51224
rect 29604 51212 29610 51264
rect 30098 51252 30104 51264
rect 30059 51224 30104 51252
rect 30098 51212 30104 51224
rect 30156 51212 30162 51264
rect 30374 51252 30380 51264
rect 30335 51224 30380 51252
rect 30374 51212 30380 51224
rect 30432 51212 30438 51264
rect 31205 51255 31263 51261
rect 31205 51221 31217 51255
rect 31251 51252 31263 51255
rect 31478 51252 31484 51264
rect 31251 51224 31484 51252
rect 31251 51221 31263 51224
rect 31205 51215 31263 51221
rect 31478 51212 31484 51224
rect 31536 51212 31542 51264
rect 33594 51212 33600 51264
rect 33652 51252 33658 51264
rect 33689 51255 33747 51261
rect 33689 51252 33701 51255
rect 33652 51224 33701 51252
rect 33652 51212 33658 51224
rect 33689 51221 33701 51224
rect 33735 51252 33747 51255
rect 34146 51252 34152 51264
rect 33735 51224 34152 51252
rect 33735 51221 33747 51224
rect 33689 51215 33747 51221
rect 34146 51212 34152 51224
rect 34204 51212 34210 51264
rect 1104 51162 38824 51184
rect 1104 51110 4246 51162
rect 4298 51110 4310 51162
rect 4362 51110 4374 51162
rect 4426 51110 4438 51162
rect 4490 51110 34966 51162
rect 35018 51110 35030 51162
rect 35082 51110 35094 51162
rect 35146 51110 35158 51162
rect 35210 51110 38824 51162
rect 1104 51088 38824 51110
rect 15010 51008 15016 51060
rect 15068 51048 15074 51060
rect 15289 51051 15347 51057
rect 15289 51048 15301 51051
rect 15068 51020 15301 51048
rect 15068 51008 15074 51020
rect 15289 51017 15301 51020
rect 15335 51017 15347 51051
rect 16022 51048 16028 51060
rect 15983 51020 16028 51048
rect 15289 51011 15347 51017
rect 16022 51008 16028 51020
rect 16080 51008 16086 51060
rect 18598 51008 18604 51060
rect 18656 51048 18662 51060
rect 19794 51048 19800 51060
rect 18656 51020 19800 51048
rect 18656 51008 18662 51020
rect 19794 51008 19800 51020
rect 19852 51008 19858 51060
rect 20346 51048 20352 51060
rect 20307 51020 20352 51048
rect 20346 51008 20352 51020
rect 20404 51008 20410 51060
rect 22002 51048 22008 51060
rect 21963 51020 22008 51048
rect 22002 51008 22008 51020
rect 22060 51008 22066 51060
rect 22278 51048 22284 51060
rect 22239 51020 22284 51048
rect 22278 51008 22284 51020
rect 22336 51008 22342 51060
rect 22649 51051 22707 51057
rect 22649 51017 22661 51051
rect 22695 51048 22707 51051
rect 23382 51048 23388 51060
rect 22695 51020 23388 51048
rect 22695 51017 22707 51020
rect 22649 51011 22707 51017
rect 23382 51008 23388 51020
rect 23440 51008 23446 51060
rect 24302 51048 24308 51060
rect 24044 51020 24308 51048
rect 15657 50983 15715 50989
rect 15657 50949 15669 50983
rect 15703 50980 15715 50983
rect 16206 50980 16212 50992
rect 15703 50952 16212 50980
rect 15703 50949 15715 50952
rect 15657 50943 15715 50949
rect 16206 50940 16212 50952
rect 16264 50980 16270 50992
rect 18874 50980 18880 50992
rect 16264 50952 17172 50980
rect 18835 50952 18880 50980
rect 16264 50940 16270 50952
rect 16574 50872 16580 50924
rect 16632 50912 16638 50924
rect 17144 50921 17172 50952
rect 18874 50940 18880 50952
rect 18932 50940 18938 50992
rect 24044 50980 24072 51020
rect 24302 51008 24308 51020
rect 24360 51008 24366 51060
rect 24854 51048 24860 51060
rect 24815 51020 24860 51048
rect 24854 51008 24860 51020
rect 24912 51008 24918 51060
rect 28074 51008 28080 51060
rect 28132 51008 28138 51060
rect 28350 51008 28356 51060
rect 28408 51048 28414 51060
rect 28445 51051 28503 51057
rect 28445 51048 28457 51051
rect 28408 51020 28457 51048
rect 28408 51008 28414 51020
rect 28445 51017 28457 51020
rect 28491 51017 28503 51051
rect 28445 51011 28503 51017
rect 30190 51008 30196 51060
rect 30248 51048 30254 51060
rect 30377 51051 30435 51057
rect 30377 51048 30389 51051
rect 30248 51020 30389 51048
rect 30248 51008 30254 51020
rect 30377 51017 30389 51020
rect 30423 51017 30435 51051
rect 30377 51011 30435 51017
rect 31386 51008 31392 51060
rect 31444 51048 31450 51060
rect 31757 51051 31815 51057
rect 31757 51048 31769 51051
rect 31444 51020 31769 51048
rect 31444 51008 31450 51020
rect 31757 51017 31769 51020
rect 31803 51017 31815 51051
rect 31757 51011 31815 51017
rect 23400 50952 24072 50980
rect 24121 50983 24179 50989
rect 17129 50915 17187 50921
rect 16632 50884 16988 50912
rect 16632 50872 16638 50884
rect 14645 50847 14703 50853
rect 14645 50813 14657 50847
rect 14691 50844 14703 50847
rect 15102 50844 15108 50856
rect 14691 50816 15108 50844
rect 14691 50813 14703 50816
rect 14645 50807 14703 50813
rect 15102 50804 15108 50816
rect 15160 50804 15166 50856
rect 16666 50844 16672 50856
rect 15488 50816 16672 50844
rect 15013 50779 15071 50785
rect 15013 50745 15025 50779
rect 15059 50776 15071 50779
rect 15488 50776 15516 50816
rect 16666 50804 16672 50816
rect 16724 50804 16730 50856
rect 16960 50853 16988 50884
rect 17129 50881 17141 50915
rect 17175 50912 17187 50915
rect 17218 50912 17224 50924
rect 17175 50884 17224 50912
rect 17175 50881 17187 50884
rect 17129 50875 17187 50881
rect 17218 50872 17224 50884
rect 17276 50872 17282 50924
rect 17862 50872 17868 50924
rect 17920 50912 17926 50924
rect 21634 50912 21640 50924
rect 17920 50884 19012 50912
rect 17920 50872 17926 50884
rect 16945 50847 17003 50853
rect 16945 50813 16957 50847
rect 16991 50813 17003 50847
rect 16945 50807 17003 50813
rect 18049 50847 18107 50853
rect 18049 50813 18061 50847
rect 18095 50844 18107 50847
rect 18601 50847 18659 50853
rect 18095 50816 18129 50844
rect 18095 50813 18107 50816
rect 18049 50807 18107 50813
rect 18601 50813 18613 50847
rect 18647 50844 18659 50847
rect 18782 50844 18788 50856
rect 18647 50816 18788 50844
rect 18647 50813 18659 50816
rect 18601 50807 18659 50813
rect 15059 50748 15516 50776
rect 16117 50779 16175 50785
rect 15059 50745 15071 50748
rect 15013 50739 15071 50745
rect 16117 50745 16129 50779
rect 16163 50776 16175 50779
rect 17310 50776 17316 50788
rect 16163 50748 17316 50776
rect 16163 50745 16175 50748
rect 16117 50739 16175 50745
rect 17310 50736 17316 50748
rect 17368 50736 17374 50788
rect 17494 50776 17500 50788
rect 17407 50748 17500 50776
rect 17494 50736 17500 50748
rect 17552 50776 17558 50788
rect 17865 50779 17923 50785
rect 17865 50776 17877 50779
rect 17552 50748 17877 50776
rect 17552 50736 17558 50748
rect 17865 50745 17877 50748
rect 17911 50776 17923 50779
rect 18064 50776 18092 50807
rect 18782 50804 18788 50816
rect 18840 50804 18846 50856
rect 18984 50853 19012 50884
rect 20824 50884 21640 50912
rect 18969 50847 19027 50853
rect 18969 50813 18981 50847
rect 19015 50844 19027 50847
rect 19242 50844 19248 50856
rect 19015 50816 19248 50844
rect 19015 50813 19027 50816
rect 18969 50807 19027 50813
rect 19242 50804 19248 50816
rect 19300 50804 19306 50856
rect 20714 50804 20720 50856
rect 20772 50844 20778 50856
rect 20824 50853 20852 50884
rect 21634 50872 21640 50884
rect 21692 50872 21698 50924
rect 22002 50872 22008 50924
rect 22060 50872 22066 50924
rect 20809 50847 20867 50853
rect 20809 50844 20821 50847
rect 20772 50816 20821 50844
rect 20772 50804 20778 50816
rect 20809 50813 20821 50816
rect 20855 50813 20867 50847
rect 20809 50807 20867 50813
rect 20993 50847 21051 50853
rect 20993 50813 21005 50847
rect 21039 50813 21051 50847
rect 21358 50844 21364 50856
rect 21319 50816 21364 50844
rect 20993 50807 21051 50813
rect 18230 50776 18236 50788
rect 17911 50748 18236 50776
rect 17911 50745 17923 50748
rect 17865 50739 17923 50745
rect 18230 50736 18236 50748
rect 18288 50736 18294 50788
rect 20438 50736 20444 50788
rect 20496 50776 20502 50788
rect 21008 50776 21036 50807
rect 21358 50804 21364 50816
rect 21416 50804 21422 50856
rect 22020 50776 22048 50872
rect 23400 50853 23428 50952
rect 24121 50949 24133 50983
rect 24167 50980 24179 50983
rect 24762 50980 24768 50992
rect 24167 50952 24768 50980
rect 24167 50949 24179 50952
rect 24121 50943 24179 50949
rect 24762 50940 24768 50952
rect 24820 50940 24826 50992
rect 24872 50912 24900 51008
rect 27614 50940 27620 50992
rect 27672 50980 27678 50992
rect 28092 50980 28120 51008
rect 27672 50952 28120 50980
rect 27672 50940 27678 50952
rect 25225 50915 25283 50921
rect 25225 50912 25237 50915
rect 24872 50884 25237 50912
rect 25225 50881 25237 50884
rect 25271 50881 25283 50915
rect 25225 50875 25283 50881
rect 26605 50915 26663 50921
rect 26605 50881 26617 50915
rect 26651 50912 26663 50915
rect 27338 50912 27344 50924
rect 26651 50884 27344 50912
rect 26651 50881 26663 50884
rect 26605 50875 26663 50881
rect 27338 50872 27344 50884
rect 27396 50872 27402 50924
rect 28718 50872 28724 50924
rect 28776 50912 28782 50924
rect 29273 50915 29331 50921
rect 29273 50912 29285 50915
rect 28776 50884 29285 50912
rect 28776 50872 28782 50884
rect 29273 50881 29285 50884
rect 29319 50881 29331 50915
rect 29273 50875 29331 50881
rect 30006 50872 30012 50924
rect 30064 50912 30070 50924
rect 30558 50912 30564 50924
rect 30064 50884 30564 50912
rect 30064 50872 30070 50884
rect 30558 50872 30564 50884
rect 30616 50872 30622 50924
rect 22465 50847 22523 50853
rect 22465 50813 22477 50847
rect 22511 50844 22523 50847
rect 22925 50847 22983 50853
rect 22925 50844 22937 50847
rect 22511 50816 22937 50844
rect 22511 50813 22523 50816
rect 22465 50807 22523 50813
rect 22925 50813 22937 50816
rect 22971 50844 22983 50847
rect 23385 50847 23443 50853
rect 23385 50844 23397 50847
rect 22971 50816 23397 50844
rect 22971 50813 22983 50816
rect 22925 50807 22983 50813
rect 23385 50813 23397 50816
rect 23431 50813 23443 50847
rect 23385 50807 23443 50813
rect 23937 50847 23995 50853
rect 23937 50813 23949 50847
rect 23983 50844 23995 50847
rect 23983 50816 24348 50844
rect 23983 50813 23995 50816
rect 23937 50807 23995 50813
rect 20496 50748 22048 50776
rect 20496 50736 20502 50748
rect 17954 50668 17960 50720
rect 18012 50708 18018 50720
rect 18138 50708 18144 50720
rect 18012 50680 18144 50708
rect 18012 50668 18018 50680
rect 18138 50668 18144 50680
rect 18196 50668 18202 50720
rect 19521 50711 19579 50717
rect 19521 50677 19533 50711
rect 19567 50708 19579 50711
rect 19978 50708 19984 50720
rect 19567 50680 19984 50708
rect 19567 50677 19579 50680
rect 19521 50671 19579 50677
rect 19978 50668 19984 50680
rect 20036 50708 20042 50720
rect 20346 50708 20352 50720
rect 20036 50680 20352 50708
rect 20036 50668 20042 50680
rect 20346 50668 20352 50680
rect 20404 50668 20410 50720
rect 20809 50711 20867 50717
rect 20809 50677 20821 50711
rect 20855 50708 20867 50711
rect 20898 50708 20904 50720
rect 20855 50680 20904 50708
rect 20855 50677 20867 50680
rect 20809 50671 20867 50677
rect 20898 50668 20904 50680
rect 20956 50668 20962 50720
rect 21174 50668 21180 50720
rect 21232 50708 21238 50720
rect 22002 50708 22008 50720
rect 21232 50680 22008 50708
rect 21232 50668 21238 50680
rect 22002 50668 22008 50680
rect 22060 50708 22066 50720
rect 22480 50708 22508 50807
rect 24320 50720 24348 50816
rect 24854 50804 24860 50856
rect 24912 50844 24918 50856
rect 24949 50847 25007 50853
rect 24949 50844 24961 50847
rect 24912 50816 24961 50844
rect 24912 50804 24918 50816
rect 24949 50813 24961 50816
rect 24995 50844 25007 50847
rect 25498 50844 25504 50856
rect 24995 50816 25504 50844
rect 24995 50813 25007 50816
rect 24949 50807 25007 50813
rect 25498 50804 25504 50816
rect 25556 50804 25562 50856
rect 27062 50804 27068 50856
rect 27120 50844 27126 50856
rect 27785 50847 27843 50853
rect 27785 50844 27797 50847
rect 27120 50816 27797 50844
rect 27120 50804 27126 50816
rect 27785 50813 27797 50816
rect 27831 50844 27843 50847
rect 29365 50847 29423 50853
rect 29365 50844 29377 50847
rect 27831 50816 28396 50844
rect 27831 50813 27843 50816
rect 27785 50807 27843 50813
rect 26418 50736 26424 50788
rect 26476 50776 26482 50788
rect 27249 50779 27307 50785
rect 27249 50776 27261 50779
rect 26476 50748 27261 50776
rect 26476 50736 26482 50748
rect 27249 50745 27261 50748
rect 27295 50776 27307 50779
rect 27433 50779 27491 50785
rect 27433 50776 27445 50779
rect 27295 50748 27445 50776
rect 27295 50745 27307 50748
rect 27249 50739 27307 50745
rect 27433 50745 27445 50748
rect 27479 50745 27491 50779
rect 27433 50739 27491 50745
rect 27709 50779 27767 50785
rect 27709 50745 27721 50779
rect 27755 50776 27767 50779
rect 27982 50776 27988 50788
rect 27755 50748 27988 50776
rect 27755 50745 27767 50748
rect 27709 50739 27767 50745
rect 27982 50736 27988 50748
rect 28040 50736 28046 50788
rect 28166 50776 28172 50788
rect 28127 50748 28172 50776
rect 28166 50736 28172 50748
rect 28224 50736 28230 50788
rect 28368 50720 28396 50816
rect 29012 50816 29377 50844
rect 29012 50720 29040 50816
rect 29365 50813 29377 50816
rect 29411 50813 29423 50847
rect 30834 50844 30840 50856
rect 30795 50816 30840 50844
rect 29365 50807 29423 50813
rect 30834 50804 30840 50816
rect 30892 50844 30898 50856
rect 31297 50847 31355 50853
rect 31297 50844 31309 50847
rect 30892 50816 31309 50844
rect 30892 50804 30898 50816
rect 31297 50813 31309 50816
rect 31343 50813 31355 50847
rect 33686 50844 33692 50856
rect 33647 50816 33692 50844
rect 31297 50807 31355 50813
rect 33686 50804 33692 50816
rect 33744 50804 33750 50856
rect 22060 50680 22508 50708
rect 22060 50668 22066 50680
rect 24302 50668 24308 50720
rect 24360 50708 24366 50720
rect 24397 50711 24455 50717
rect 24397 50708 24409 50711
rect 24360 50680 24409 50708
rect 24360 50668 24366 50680
rect 24397 50677 24409 50680
rect 24443 50677 24455 50711
rect 26878 50708 26884 50720
rect 26839 50680 26884 50708
rect 24397 50671 24455 50677
rect 26878 50668 26884 50680
rect 26936 50668 26942 50720
rect 27522 50668 27528 50720
rect 27580 50708 27586 50720
rect 27617 50711 27675 50717
rect 27617 50708 27629 50711
rect 27580 50680 27629 50708
rect 27580 50668 27586 50680
rect 27617 50677 27629 50680
rect 27663 50708 27675 50711
rect 27798 50708 27804 50720
rect 27663 50680 27804 50708
rect 27663 50677 27675 50680
rect 27617 50671 27675 50677
rect 27798 50668 27804 50680
rect 27856 50668 27862 50720
rect 28350 50668 28356 50720
rect 28408 50668 28414 50720
rect 28994 50708 29000 50720
rect 28955 50680 29000 50708
rect 28994 50668 29000 50680
rect 29052 50668 29058 50720
rect 29454 50668 29460 50720
rect 29512 50708 29518 50720
rect 29730 50708 29736 50720
rect 29512 50680 29736 50708
rect 29512 50668 29518 50680
rect 29730 50668 29736 50680
rect 29788 50668 29794 50720
rect 30745 50711 30803 50717
rect 30745 50677 30757 50711
rect 30791 50708 30803 50711
rect 30926 50708 30932 50720
rect 30791 50680 30932 50708
rect 30791 50677 30803 50680
rect 30745 50671 30803 50677
rect 30926 50668 30932 50680
rect 30984 50668 30990 50720
rect 31018 50668 31024 50720
rect 31076 50708 31082 50720
rect 31076 50680 31121 50708
rect 31076 50668 31082 50680
rect 34790 50668 34796 50720
rect 34848 50708 34854 50720
rect 35434 50708 35440 50720
rect 34848 50680 35440 50708
rect 34848 50668 34854 50680
rect 35434 50668 35440 50680
rect 35492 50668 35498 50720
rect 1104 50618 38824 50640
rect 1104 50566 19606 50618
rect 19658 50566 19670 50618
rect 19722 50566 19734 50618
rect 19786 50566 19798 50618
rect 19850 50566 38824 50618
rect 1104 50544 38824 50566
rect 17681 50507 17739 50513
rect 17681 50473 17693 50507
rect 17727 50504 17739 50507
rect 17862 50504 17868 50516
rect 17727 50476 17868 50504
rect 17727 50473 17739 50476
rect 17681 50467 17739 50473
rect 17862 50464 17868 50476
rect 17920 50504 17926 50516
rect 18049 50507 18107 50513
rect 18049 50504 18061 50507
rect 17920 50476 18061 50504
rect 17920 50464 17926 50476
rect 18049 50473 18061 50476
rect 18095 50473 18107 50507
rect 18049 50467 18107 50473
rect 20625 50507 20683 50513
rect 20625 50473 20637 50507
rect 20671 50504 20683 50507
rect 21358 50504 21364 50516
rect 20671 50476 21364 50504
rect 20671 50473 20683 50476
rect 20625 50467 20683 50473
rect 21358 50464 21364 50476
rect 21416 50464 21422 50516
rect 23569 50507 23627 50513
rect 23569 50473 23581 50507
rect 23615 50504 23627 50507
rect 23934 50504 23940 50516
rect 23615 50476 23940 50504
rect 23615 50473 23627 50476
rect 23569 50467 23627 50473
rect 23934 50464 23940 50476
rect 23992 50464 23998 50516
rect 26789 50507 26847 50513
rect 26789 50473 26801 50507
rect 26835 50504 26847 50507
rect 26970 50504 26976 50516
rect 26835 50476 26976 50504
rect 26835 50473 26847 50476
rect 26789 50467 26847 50473
rect 26970 50464 26976 50476
rect 27028 50464 27034 50516
rect 27157 50507 27215 50513
rect 27157 50473 27169 50507
rect 27203 50504 27215 50507
rect 27522 50504 27528 50516
rect 27203 50476 27528 50504
rect 27203 50473 27215 50476
rect 27157 50467 27215 50473
rect 27522 50464 27528 50476
rect 27580 50504 27586 50516
rect 28166 50504 28172 50516
rect 27580 50476 28172 50504
rect 27580 50464 27586 50476
rect 28166 50464 28172 50476
rect 28224 50464 28230 50516
rect 30466 50464 30472 50516
rect 30524 50504 30530 50516
rect 30929 50507 30987 50513
rect 30929 50504 30941 50507
rect 30524 50476 30941 50504
rect 30524 50464 30530 50476
rect 30929 50473 30941 50476
rect 30975 50473 30987 50507
rect 30929 50467 30987 50473
rect 18506 50396 18512 50448
rect 18564 50396 18570 50448
rect 21082 50396 21088 50448
rect 21140 50436 21146 50448
rect 21177 50439 21235 50445
rect 21177 50436 21189 50439
rect 21140 50408 21189 50436
rect 21140 50396 21146 50408
rect 21177 50405 21189 50408
rect 21223 50405 21235 50439
rect 21177 50399 21235 50405
rect 22833 50439 22891 50445
rect 22833 50405 22845 50439
rect 22879 50436 22891 50439
rect 22922 50436 22928 50448
rect 22879 50408 22928 50436
rect 22879 50405 22891 50408
rect 22833 50399 22891 50405
rect 15565 50371 15623 50377
rect 15565 50368 15577 50371
rect 15028 50340 15577 50368
rect 14826 50124 14832 50176
rect 14884 50164 14890 50176
rect 15028 50173 15056 50340
rect 15565 50337 15577 50340
rect 15611 50368 15623 50371
rect 15654 50368 15660 50380
rect 15611 50340 15660 50368
rect 15611 50337 15623 50340
rect 15565 50331 15623 50337
rect 15654 50328 15660 50340
rect 15712 50328 15718 50380
rect 17954 50328 17960 50380
rect 18012 50368 18018 50380
rect 18524 50368 18552 50396
rect 18785 50371 18843 50377
rect 18785 50368 18797 50371
rect 18012 50340 18797 50368
rect 18012 50328 18018 50340
rect 18785 50337 18797 50340
rect 18831 50337 18843 50371
rect 18785 50331 18843 50337
rect 18966 50328 18972 50380
rect 19024 50368 19030 50380
rect 19245 50371 19303 50377
rect 19245 50368 19257 50371
rect 19024 50340 19257 50368
rect 19024 50328 19030 50340
rect 19245 50337 19257 50340
rect 19291 50337 19303 50371
rect 19981 50371 20039 50377
rect 19981 50368 19993 50371
rect 19245 50331 19303 50337
rect 19352 50340 19993 50368
rect 19352 50312 19380 50340
rect 19981 50337 19993 50340
rect 20027 50368 20039 50371
rect 20622 50368 20628 50380
rect 20027 50340 20628 50368
rect 20027 50337 20039 50340
rect 19981 50331 20039 50337
rect 20622 50328 20628 50340
rect 20680 50328 20686 50380
rect 21726 50368 21732 50380
rect 21687 50340 21732 50368
rect 21726 50328 21732 50340
rect 21784 50328 21790 50380
rect 22278 50368 22284 50380
rect 22239 50340 22284 50368
rect 22278 50328 22284 50340
rect 22336 50328 22342 50380
rect 22646 50368 22652 50380
rect 22607 50340 22652 50368
rect 22646 50328 22652 50340
rect 22704 50328 22710 50380
rect 15286 50300 15292 50312
rect 15247 50272 15292 50300
rect 15286 50260 15292 50272
rect 15344 50260 15350 50312
rect 17313 50303 17371 50309
rect 17313 50269 17325 50303
rect 17359 50300 17371 50303
rect 17402 50300 17408 50312
rect 17359 50272 17408 50300
rect 17359 50269 17371 50272
rect 17313 50263 17371 50269
rect 17402 50260 17408 50272
rect 17460 50260 17466 50312
rect 18046 50260 18052 50312
rect 18104 50300 18110 50312
rect 18509 50303 18567 50309
rect 18509 50300 18521 50303
rect 18104 50272 18521 50300
rect 18104 50260 18110 50272
rect 18509 50269 18521 50272
rect 18555 50300 18567 50303
rect 19334 50300 19340 50312
rect 18555 50272 19340 50300
rect 18555 50269 18567 50272
rect 18509 50263 18567 50269
rect 19334 50260 19340 50272
rect 19392 50260 19398 50312
rect 19521 50303 19579 50309
rect 19521 50269 19533 50303
rect 19567 50300 19579 50303
rect 20162 50300 20168 50312
rect 19567 50272 20168 50300
rect 19567 50269 19579 50272
rect 19521 50263 19579 50269
rect 20162 50260 20168 50272
rect 20220 50260 20226 50312
rect 21637 50235 21695 50241
rect 21637 50201 21649 50235
rect 21683 50232 21695 50235
rect 22186 50232 22192 50244
rect 21683 50204 22192 50232
rect 21683 50201 21695 50204
rect 21637 50195 21695 50201
rect 22186 50192 22192 50204
rect 22244 50232 22250 50244
rect 22848 50232 22876 50399
rect 22922 50396 22928 50408
rect 22980 50396 22986 50448
rect 26329 50439 26387 50445
rect 26329 50405 26341 50439
rect 26375 50436 26387 50439
rect 27062 50436 27068 50448
rect 26375 50408 27068 50436
rect 26375 50405 26387 50408
rect 26329 50399 26387 50405
rect 27062 50396 27068 50408
rect 27120 50396 27126 50448
rect 27706 50396 27712 50448
rect 27764 50436 27770 50448
rect 27764 50408 28488 50436
rect 27764 50396 27770 50408
rect 24118 50328 24124 50380
rect 24176 50368 24182 50380
rect 24213 50371 24271 50377
rect 24213 50368 24225 50371
rect 24176 50340 24225 50368
rect 24176 50328 24182 50340
rect 24213 50337 24225 50340
rect 24259 50337 24271 50371
rect 24486 50368 24492 50380
rect 24447 50340 24492 50368
rect 24213 50331 24271 50337
rect 24486 50328 24492 50340
rect 24544 50368 24550 50380
rect 24949 50371 25007 50377
rect 24949 50368 24961 50371
rect 24544 50340 24961 50368
rect 24544 50328 24550 50340
rect 24949 50337 24961 50340
rect 24995 50337 25007 50371
rect 24949 50331 25007 50337
rect 27246 50328 27252 50380
rect 27304 50368 27310 50380
rect 27525 50371 27583 50377
rect 27525 50368 27537 50371
rect 27304 50340 27537 50368
rect 27304 50328 27310 50340
rect 27525 50337 27537 50340
rect 27571 50337 27583 50371
rect 28350 50368 28356 50380
rect 28311 50340 28356 50368
rect 27525 50331 27583 50337
rect 28350 50328 28356 50340
rect 28408 50328 28414 50380
rect 28460 50377 28488 50408
rect 28445 50371 28503 50377
rect 28445 50337 28457 50371
rect 28491 50337 28503 50371
rect 28445 50331 28503 50337
rect 29086 50328 29092 50380
rect 29144 50368 29150 50380
rect 31478 50368 31484 50380
rect 29144 50340 31484 50368
rect 29144 50328 29150 50340
rect 31478 50328 31484 50340
rect 31536 50328 31542 50380
rect 23658 50300 23664 50312
rect 23619 50272 23664 50300
rect 23658 50260 23664 50272
rect 23716 50260 23722 50312
rect 23842 50260 23848 50312
rect 23900 50300 23906 50312
rect 24673 50303 24731 50309
rect 24673 50300 24685 50303
rect 23900 50272 24685 50300
rect 23900 50260 23906 50272
rect 24673 50269 24685 50272
rect 24719 50300 24731 50303
rect 25777 50303 25835 50309
rect 25777 50300 25789 50303
rect 24719 50272 25789 50300
rect 24719 50269 24731 50272
rect 24673 50263 24731 50269
rect 25777 50269 25789 50272
rect 25823 50269 25835 50303
rect 25777 50263 25835 50269
rect 27617 50303 27675 50309
rect 27617 50269 27629 50303
rect 27663 50300 27675 50303
rect 28258 50300 28264 50312
rect 27663 50272 28264 50300
rect 27663 50269 27675 50272
rect 27617 50263 27675 50269
rect 28258 50260 28264 50272
rect 28316 50260 28322 50312
rect 29546 50300 29552 50312
rect 29507 50272 29552 50300
rect 29546 50260 29552 50272
rect 29604 50260 29610 50312
rect 29730 50260 29736 50312
rect 29788 50300 29794 50312
rect 29825 50303 29883 50309
rect 29825 50300 29837 50303
rect 29788 50272 29837 50300
rect 29788 50260 29794 50272
rect 29825 50269 29837 50272
rect 29871 50269 29883 50303
rect 29825 50263 29883 50269
rect 22244 50204 22876 50232
rect 22244 50192 22250 50204
rect 27798 50192 27804 50244
rect 27856 50232 27862 50244
rect 28534 50232 28540 50244
rect 27856 50204 28540 50232
rect 27856 50192 27862 50204
rect 28534 50192 28540 50204
rect 28592 50192 28598 50244
rect 15013 50167 15071 50173
rect 15013 50164 15025 50167
rect 14884 50136 15025 50164
rect 14884 50124 14890 50136
rect 15013 50133 15025 50136
rect 15059 50133 15071 50167
rect 15013 50127 15071 50133
rect 15194 50124 15200 50176
rect 15252 50164 15258 50176
rect 16298 50164 16304 50176
rect 15252 50136 16304 50164
rect 15252 50124 15258 50136
rect 16298 50124 16304 50136
rect 16356 50164 16362 50176
rect 16669 50167 16727 50173
rect 16669 50164 16681 50167
rect 16356 50136 16681 50164
rect 16356 50124 16362 50136
rect 16669 50133 16681 50136
rect 16715 50133 16727 50167
rect 16669 50127 16727 50133
rect 22462 50124 22468 50176
rect 22520 50164 22526 50176
rect 23109 50167 23167 50173
rect 23109 50164 23121 50167
rect 22520 50136 23121 50164
rect 22520 50124 22526 50136
rect 23109 50133 23121 50136
rect 23155 50133 23167 50167
rect 23109 50127 23167 50133
rect 25314 50124 25320 50176
rect 25372 50164 25378 50176
rect 25501 50167 25559 50173
rect 25501 50164 25513 50167
rect 25372 50136 25513 50164
rect 25372 50124 25378 50136
rect 25501 50133 25513 50136
rect 25547 50164 25559 50167
rect 25590 50164 25596 50176
rect 25547 50136 25596 50164
rect 25547 50133 25559 50136
rect 25501 50127 25559 50133
rect 25590 50124 25596 50136
rect 25648 50124 25654 50176
rect 28902 50164 28908 50176
rect 28863 50136 28908 50164
rect 28902 50124 28908 50136
rect 28960 50124 28966 50176
rect 29270 50164 29276 50176
rect 29231 50136 29276 50164
rect 29270 50124 29276 50136
rect 29328 50124 29334 50176
rect 1104 50074 38824 50096
rect 1104 50022 4246 50074
rect 4298 50022 4310 50074
rect 4362 50022 4374 50074
rect 4426 50022 4438 50074
rect 4490 50022 34966 50074
rect 35018 50022 35030 50074
rect 35082 50022 35094 50074
rect 35146 50022 35158 50074
rect 35210 50022 38824 50074
rect 1104 50000 38824 50022
rect 17129 49963 17187 49969
rect 17129 49929 17141 49963
rect 17175 49960 17187 49963
rect 17218 49960 17224 49972
rect 17175 49932 17224 49960
rect 17175 49929 17187 49932
rect 17129 49923 17187 49929
rect 17218 49920 17224 49932
rect 17276 49920 17282 49972
rect 17310 49920 17316 49972
rect 17368 49960 17374 49972
rect 17405 49963 17463 49969
rect 17405 49960 17417 49963
rect 17368 49932 17417 49960
rect 17368 49920 17374 49932
rect 17405 49929 17417 49932
rect 17451 49929 17463 49963
rect 17405 49923 17463 49929
rect 17865 49963 17923 49969
rect 17865 49929 17877 49963
rect 17911 49960 17923 49963
rect 18230 49960 18236 49972
rect 17911 49932 18236 49960
rect 17911 49929 17923 49932
rect 17865 49923 17923 49929
rect 14461 49895 14519 49901
rect 14461 49861 14473 49895
rect 14507 49892 14519 49895
rect 15194 49892 15200 49904
rect 14507 49864 15200 49892
rect 14507 49861 14519 49864
rect 14461 49855 14519 49861
rect 15194 49852 15200 49864
rect 15252 49852 15258 49904
rect 15654 49852 15660 49904
rect 15712 49852 15718 49904
rect 15378 49824 15384 49836
rect 15339 49796 15384 49824
rect 15378 49784 15384 49796
rect 15436 49784 15442 49836
rect 15672 49824 15700 49852
rect 15749 49827 15807 49833
rect 15749 49824 15761 49827
rect 15672 49796 15761 49824
rect 15749 49793 15761 49796
rect 15795 49793 15807 49827
rect 16209 49827 16267 49833
rect 16209 49824 16221 49827
rect 15749 49787 15807 49793
rect 15856 49796 16221 49824
rect 13814 49716 13820 49768
rect 13872 49756 13878 49768
rect 14737 49759 14795 49765
rect 14737 49756 14749 49759
rect 13872 49728 14749 49756
rect 13872 49716 13878 49728
rect 14737 49725 14749 49728
rect 14783 49756 14795 49759
rect 15197 49759 15255 49765
rect 14783 49728 15148 49756
rect 14783 49725 14795 49728
rect 14737 49719 14795 49725
rect 15120 49688 15148 49728
rect 15197 49725 15209 49759
rect 15243 49756 15255 49759
rect 15654 49756 15660 49768
rect 15243 49728 15660 49756
rect 15243 49725 15255 49728
rect 15197 49719 15255 49725
rect 15654 49716 15660 49728
rect 15712 49756 15718 49768
rect 15856 49756 15884 49796
rect 16209 49793 16221 49796
rect 16255 49793 16267 49827
rect 17420 49824 17448 49923
rect 18230 49920 18236 49932
rect 18288 49960 18294 49972
rect 18288 49932 19012 49960
rect 18288 49920 18294 49932
rect 18138 49852 18144 49904
rect 18196 49892 18202 49904
rect 18877 49895 18935 49901
rect 18877 49892 18889 49895
rect 18196 49864 18889 49892
rect 18196 49852 18202 49864
rect 18877 49861 18889 49864
rect 18923 49861 18935 49895
rect 18984 49892 19012 49932
rect 19334 49920 19340 49972
rect 19392 49960 19398 49972
rect 19429 49963 19487 49969
rect 19429 49960 19441 49963
rect 19392 49932 19441 49960
rect 19392 49920 19398 49932
rect 19429 49929 19441 49932
rect 19475 49929 19487 49963
rect 19429 49923 19487 49929
rect 21453 49963 21511 49969
rect 21453 49929 21465 49963
rect 21499 49960 21511 49963
rect 21726 49960 21732 49972
rect 21499 49932 21732 49960
rect 21499 49929 21511 49932
rect 21453 49923 21511 49929
rect 18984 49864 19380 49892
rect 18877 49855 18935 49861
rect 17420 49796 18920 49824
rect 16209 49787 16267 49793
rect 15712 49728 15884 49756
rect 15933 49759 15991 49765
rect 15712 49716 15718 49728
rect 15933 49725 15945 49759
rect 15979 49725 15991 49759
rect 16298 49756 16304 49768
rect 16259 49728 16304 49756
rect 15933 49719 15991 49725
rect 15948 49688 15976 49719
rect 16298 49716 16304 49728
rect 16356 49716 16362 49768
rect 18230 49756 18236 49768
rect 18191 49728 18236 49756
rect 18230 49716 18236 49728
rect 18288 49716 18294 49768
rect 18598 49756 18604 49768
rect 18559 49728 18604 49756
rect 18598 49716 18604 49728
rect 18656 49716 18662 49768
rect 18892 49765 18920 49796
rect 18877 49759 18935 49765
rect 18877 49725 18889 49759
rect 18923 49756 18935 49759
rect 19352 49756 19380 49864
rect 19444 49824 19472 49923
rect 21726 49920 21732 49932
rect 21784 49920 21790 49972
rect 22554 49920 22560 49972
rect 22612 49960 22618 49972
rect 22922 49960 22928 49972
rect 22612 49932 22928 49960
rect 22612 49920 22618 49932
rect 22922 49920 22928 49932
rect 22980 49920 22986 49972
rect 24118 49920 24124 49972
rect 24176 49960 24182 49972
rect 26421 49963 26479 49969
rect 26421 49960 26433 49963
rect 24176 49932 26433 49960
rect 24176 49920 24182 49932
rect 26421 49929 26433 49932
rect 26467 49929 26479 49963
rect 28350 49960 28356 49972
rect 28311 49932 28356 49960
rect 26421 49923 26479 49929
rect 28350 49920 28356 49932
rect 28408 49920 28414 49972
rect 28905 49963 28963 49969
rect 28905 49929 28917 49963
rect 28951 49960 28963 49963
rect 29546 49960 29552 49972
rect 28951 49932 29552 49960
rect 28951 49929 28963 49932
rect 28905 49923 28963 49929
rect 29546 49920 29552 49932
rect 29604 49960 29610 49972
rect 30650 49960 30656 49972
rect 29604 49932 30656 49960
rect 29604 49920 29610 49932
rect 30650 49920 30656 49932
rect 30708 49920 30714 49972
rect 31938 49920 31944 49972
rect 31996 49960 32002 49972
rect 32214 49960 32220 49972
rect 31996 49932 32220 49960
rect 31996 49920 32002 49932
rect 32214 49920 32220 49932
rect 32272 49920 32278 49972
rect 21082 49852 21088 49904
rect 21140 49892 21146 49904
rect 21140 49864 22416 49892
rect 21140 49852 21146 49864
rect 19444 49796 20392 49824
rect 19889 49759 19947 49765
rect 19889 49756 19901 49759
rect 18923 49728 19288 49756
rect 19352 49728 19901 49756
rect 18923 49725 18935 49728
rect 18877 49719 18935 49725
rect 15120 49660 15976 49688
rect 19260 49688 19288 49728
rect 19889 49725 19901 49728
rect 19935 49756 19947 49759
rect 20070 49756 20076 49768
rect 19935 49728 20076 49756
rect 19935 49725 19947 49728
rect 19889 49719 19947 49725
rect 20070 49716 20076 49728
rect 20128 49716 20134 49768
rect 20364 49765 20392 49796
rect 20349 49759 20407 49765
rect 20349 49725 20361 49759
rect 20395 49725 20407 49759
rect 20809 49759 20867 49765
rect 20809 49756 20821 49759
rect 20349 49719 20407 49725
rect 20640 49728 20821 49756
rect 20254 49688 20260 49700
rect 19260 49660 20260 49688
rect 20254 49648 20260 49660
rect 20312 49688 20318 49700
rect 20640 49688 20668 49728
rect 20809 49725 20821 49728
rect 20855 49725 20867 49759
rect 21082 49756 21088 49768
rect 21043 49728 21088 49756
rect 20809 49719 20867 49725
rect 21082 49716 21088 49728
rect 21140 49716 21146 49768
rect 22186 49756 22192 49768
rect 22147 49728 22192 49756
rect 22186 49716 22192 49728
rect 22244 49716 22250 49768
rect 22388 49765 22416 49864
rect 23934 49852 23940 49904
rect 23992 49892 23998 49904
rect 24302 49892 24308 49904
rect 23992 49864 24308 49892
rect 23992 49852 23998 49864
rect 24302 49852 24308 49864
rect 24360 49892 24366 49904
rect 24857 49895 24915 49901
rect 24857 49892 24869 49895
rect 24360 49864 24869 49892
rect 24360 49852 24366 49864
rect 24857 49861 24869 49864
rect 24903 49861 24915 49895
rect 26234 49892 26240 49904
rect 24857 49855 24915 49861
rect 25424 49864 26240 49892
rect 23474 49824 23480 49836
rect 23387 49796 23480 49824
rect 23474 49784 23480 49796
rect 23532 49824 23538 49836
rect 23532 49796 24164 49824
rect 23532 49784 23538 49796
rect 22373 49759 22431 49765
rect 22373 49725 22385 49759
rect 22419 49725 22431 49759
rect 22373 49719 22431 49725
rect 23109 49759 23167 49765
rect 23109 49725 23121 49759
rect 23155 49756 23167 49759
rect 23382 49756 23388 49768
rect 23155 49728 23388 49756
rect 23155 49725 23167 49728
rect 23109 49719 23167 49725
rect 23382 49716 23388 49728
rect 23440 49756 23446 49768
rect 23845 49759 23903 49765
rect 23845 49756 23857 49759
rect 23440 49728 23857 49756
rect 23440 49716 23446 49728
rect 23845 49725 23857 49728
rect 23891 49725 23903 49759
rect 23845 49719 23903 49725
rect 23934 49716 23940 49768
rect 23992 49756 23998 49768
rect 24136 49765 24164 49796
rect 25130 49784 25136 49836
rect 25188 49824 25194 49836
rect 25424 49833 25452 49864
rect 26234 49852 26240 49864
rect 26292 49852 26298 49904
rect 26326 49852 26332 49904
rect 26384 49892 26390 49904
rect 26881 49895 26939 49901
rect 26881 49892 26893 49895
rect 26384 49864 26893 49892
rect 26384 49852 26390 49864
rect 26881 49861 26893 49864
rect 26927 49892 26939 49895
rect 29822 49892 29828 49904
rect 26927 49864 27568 49892
rect 26927 49861 26939 49864
rect 26881 49855 26939 49861
rect 25225 49827 25283 49833
rect 25225 49824 25237 49827
rect 25188 49796 25237 49824
rect 25188 49784 25194 49796
rect 25225 49793 25237 49796
rect 25271 49824 25283 49827
rect 25409 49827 25467 49833
rect 25409 49824 25421 49827
rect 25271 49796 25421 49824
rect 25271 49793 25283 49796
rect 25225 49787 25283 49793
rect 25409 49793 25421 49796
rect 25455 49793 25467 49827
rect 25409 49787 25467 49793
rect 25958 49784 25964 49836
rect 26016 49824 26022 49836
rect 26145 49827 26203 49833
rect 26145 49824 26157 49827
rect 26016 49796 26157 49824
rect 26016 49784 26022 49796
rect 26145 49793 26157 49796
rect 26191 49793 26203 49827
rect 26145 49787 26203 49793
rect 26970 49784 26976 49836
rect 27028 49824 27034 49836
rect 27065 49827 27123 49833
rect 27065 49824 27077 49827
rect 27028 49796 27077 49824
rect 27028 49784 27034 49796
rect 27065 49793 27077 49796
rect 27111 49793 27123 49827
rect 27540 49824 27568 49864
rect 28736 49864 29828 49892
rect 27540 49796 27752 49824
rect 27065 49787 27123 49793
rect 24121 49759 24179 49765
rect 23992 49728 24037 49756
rect 23992 49716 23998 49728
rect 24121 49725 24133 49759
rect 24167 49725 24179 49759
rect 24121 49719 24179 49725
rect 25590 49716 25596 49768
rect 25648 49756 25654 49768
rect 27522 49756 27528 49768
rect 25648 49728 26188 49756
rect 27483 49728 27528 49756
rect 25648 49716 25654 49728
rect 20312 49660 20668 49688
rect 21821 49691 21879 49697
rect 20312 49648 20318 49660
rect 21821 49657 21833 49691
rect 21867 49688 21879 49691
rect 22278 49688 22284 49700
rect 21867 49660 22284 49688
rect 21867 49657 21879 49660
rect 21821 49651 21879 49657
rect 22278 49648 22284 49660
rect 22336 49648 22342 49700
rect 25222 49648 25228 49700
rect 25280 49688 25286 49700
rect 25498 49688 25504 49700
rect 25280 49660 25504 49688
rect 25280 49648 25286 49660
rect 25498 49648 25504 49660
rect 25556 49688 25562 49700
rect 25777 49691 25835 49697
rect 25777 49688 25789 49691
rect 25556 49660 25789 49688
rect 25556 49648 25562 49660
rect 25777 49657 25789 49660
rect 25823 49657 25835 49691
rect 26160 49688 26188 49728
rect 27522 49716 27528 49728
rect 27580 49716 27586 49768
rect 27724 49765 27752 49796
rect 27709 49759 27767 49765
rect 27709 49725 27721 49759
rect 27755 49756 27767 49759
rect 27798 49756 27804 49768
rect 27755 49728 27804 49756
rect 27755 49725 27767 49728
rect 27709 49719 27767 49725
rect 27798 49716 27804 49728
rect 27856 49716 27862 49768
rect 27890 49716 27896 49768
rect 27948 49756 27954 49768
rect 27948 49728 27993 49756
rect 27948 49716 27954 49728
rect 28626 49716 28632 49768
rect 28684 49756 28690 49768
rect 28736 49765 28764 49864
rect 29822 49852 29828 49864
rect 29880 49892 29886 49904
rect 29880 49864 30328 49892
rect 29880 49852 29886 49864
rect 29457 49827 29515 49833
rect 29457 49793 29469 49827
rect 29503 49824 29515 49827
rect 30098 49824 30104 49836
rect 29503 49796 30104 49824
rect 29503 49793 29515 49796
rect 29457 49787 29515 49793
rect 30098 49784 30104 49796
rect 30156 49784 30162 49836
rect 30300 49833 30328 49864
rect 30285 49827 30343 49833
rect 30285 49793 30297 49827
rect 30331 49793 30343 49827
rect 30285 49787 30343 49793
rect 30558 49784 30564 49836
rect 30616 49824 30622 49836
rect 30653 49827 30711 49833
rect 30653 49824 30665 49827
rect 30616 49796 30665 49824
rect 30616 49784 30622 49796
rect 30653 49793 30665 49796
rect 30699 49793 30711 49827
rect 31202 49824 31208 49836
rect 31163 49796 31208 49824
rect 30653 49787 30711 49793
rect 31202 49784 31208 49796
rect 31260 49784 31266 49836
rect 28721 49759 28779 49765
rect 28721 49756 28733 49759
rect 28684 49728 28733 49756
rect 28684 49716 28690 49728
rect 28721 49725 28733 49728
rect 28767 49725 28779 49759
rect 29086 49756 29092 49768
rect 29047 49728 29092 49756
rect 28721 49719 28779 49725
rect 29086 49716 29092 49728
rect 29144 49716 29150 49768
rect 29270 49716 29276 49768
rect 29328 49756 29334 49768
rect 29365 49759 29423 49765
rect 29365 49756 29377 49759
rect 29328 49728 29377 49756
rect 29328 49716 29334 49728
rect 29365 49725 29377 49728
rect 29411 49756 29423 49759
rect 29822 49756 29828 49768
rect 29411 49728 29828 49756
rect 29411 49725 29423 49728
rect 29365 49719 29423 49725
rect 29822 49716 29828 49728
rect 29880 49716 29886 49768
rect 30193 49759 30251 49765
rect 30193 49725 30205 49759
rect 30239 49725 30251 49759
rect 31018 49756 31024 49768
rect 30979 49728 31024 49756
rect 30193 49719 30251 49725
rect 26326 49688 26332 49700
rect 26160 49660 26332 49688
rect 25777 49651 25835 49657
rect 26326 49648 26332 49660
rect 26384 49648 26390 49700
rect 30208 49688 30236 49719
rect 31018 49716 31024 49728
rect 31076 49756 31082 49768
rect 31297 49759 31355 49765
rect 31297 49756 31309 49759
rect 31076 49728 31309 49756
rect 31076 49716 31082 49728
rect 31297 49725 31309 49728
rect 31343 49725 31355 49759
rect 31297 49719 31355 49725
rect 30374 49688 30380 49700
rect 30208 49660 30380 49688
rect 30374 49648 30380 49660
rect 30432 49648 30438 49700
rect 22186 49620 22192 49632
rect 22147 49592 22192 49620
rect 22186 49580 22192 49592
rect 22244 49580 22250 49632
rect 23750 49580 23756 49632
rect 23808 49620 23814 49632
rect 24305 49623 24363 49629
rect 24305 49620 24317 49623
rect 23808 49592 24317 49620
rect 23808 49580 23814 49592
rect 24305 49589 24317 49592
rect 24351 49589 24363 49623
rect 25590 49620 25596 49632
rect 25551 49592 25596 49620
rect 24305 49583 24363 49589
rect 25590 49580 25596 49592
rect 25648 49580 25654 49632
rect 25685 49623 25743 49629
rect 25685 49589 25697 49623
rect 25731 49620 25743 49623
rect 25958 49620 25964 49632
rect 25731 49592 25964 49620
rect 25731 49589 25743 49592
rect 25685 49583 25743 49589
rect 25958 49580 25964 49592
rect 26016 49580 26022 49632
rect 1104 49530 38824 49552
rect 1104 49478 19606 49530
rect 19658 49478 19670 49530
rect 19722 49478 19734 49530
rect 19786 49478 19798 49530
rect 19850 49478 38824 49530
rect 1104 49456 38824 49478
rect 17405 49419 17463 49425
rect 17405 49385 17417 49419
rect 17451 49416 17463 49419
rect 17862 49416 17868 49428
rect 17451 49388 17868 49416
rect 17451 49385 17463 49388
rect 17405 49379 17463 49385
rect 17862 49376 17868 49388
rect 17920 49376 17926 49428
rect 19337 49419 19395 49425
rect 19337 49385 19349 49419
rect 19383 49416 19395 49419
rect 19426 49416 19432 49428
rect 19383 49388 19432 49416
rect 19383 49385 19395 49388
rect 19337 49379 19395 49385
rect 19426 49376 19432 49388
rect 19484 49416 19490 49428
rect 19613 49419 19671 49425
rect 19613 49416 19625 49419
rect 19484 49388 19625 49416
rect 19484 49376 19490 49388
rect 19613 49385 19625 49388
rect 19659 49385 19671 49419
rect 20254 49416 20260 49428
rect 20215 49388 20260 49416
rect 19613 49379 19671 49385
rect 20254 49376 20260 49388
rect 20312 49376 20318 49428
rect 20714 49416 20720 49428
rect 20675 49388 20720 49416
rect 20714 49376 20720 49388
rect 20772 49376 20778 49428
rect 21269 49419 21327 49425
rect 21269 49385 21281 49419
rect 21315 49416 21327 49419
rect 21542 49416 21548 49428
rect 21315 49388 21548 49416
rect 21315 49385 21327 49388
rect 21269 49379 21327 49385
rect 21542 49376 21548 49388
rect 21600 49376 21606 49428
rect 22554 49376 22560 49428
rect 22612 49416 22618 49428
rect 23201 49419 23259 49425
rect 23201 49416 23213 49419
rect 22612 49388 23213 49416
rect 22612 49376 22618 49388
rect 23201 49385 23213 49388
rect 23247 49416 23259 49419
rect 23569 49419 23627 49425
rect 23569 49416 23581 49419
rect 23247 49388 23581 49416
rect 23247 49385 23259 49388
rect 23201 49379 23259 49385
rect 23569 49385 23581 49388
rect 23615 49416 23627 49419
rect 24026 49416 24032 49428
rect 23615 49388 24032 49416
rect 23615 49385 23627 49388
rect 23569 49379 23627 49385
rect 24026 49376 24032 49388
rect 24084 49376 24090 49428
rect 24762 49376 24768 49428
rect 24820 49416 24826 49428
rect 25038 49416 25044 49428
rect 24820 49388 25044 49416
rect 24820 49376 24826 49388
rect 25038 49376 25044 49388
rect 25096 49416 25102 49428
rect 25133 49419 25191 49425
rect 25133 49416 25145 49419
rect 25096 49388 25145 49416
rect 25096 49376 25102 49388
rect 25133 49385 25145 49388
rect 25179 49416 25191 49419
rect 25501 49419 25559 49425
rect 25501 49416 25513 49419
rect 25179 49388 25513 49416
rect 25179 49385 25191 49388
rect 25133 49379 25191 49385
rect 25501 49385 25513 49388
rect 25547 49416 25559 49419
rect 25590 49416 25596 49428
rect 25547 49388 25596 49416
rect 25547 49385 25559 49388
rect 25501 49379 25559 49385
rect 25590 49376 25596 49388
rect 25648 49416 25654 49428
rect 26694 49416 26700 49428
rect 25648 49388 26700 49416
rect 25648 49376 25654 49388
rect 26694 49376 26700 49388
rect 26752 49376 26758 49428
rect 27246 49376 27252 49428
rect 27304 49416 27310 49428
rect 27801 49419 27859 49425
rect 27801 49416 27813 49419
rect 27304 49388 27813 49416
rect 27304 49376 27310 49388
rect 27801 49385 27813 49388
rect 27847 49385 27859 49419
rect 27801 49379 27859 49385
rect 29641 49419 29699 49425
rect 29641 49385 29653 49419
rect 29687 49416 29699 49419
rect 29730 49416 29736 49428
rect 29687 49388 29736 49416
rect 29687 49385 29699 49388
rect 29641 49379 29699 49385
rect 29730 49376 29736 49388
rect 29788 49376 29794 49428
rect 30374 49376 30380 49428
rect 30432 49416 30438 49428
rect 30929 49419 30987 49425
rect 30929 49416 30941 49419
rect 30432 49388 30941 49416
rect 30432 49376 30438 49388
rect 30929 49385 30941 49388
rect 30975 49416 30987 49419
rect 31662 49416 31668 49428
rect 30975 49388 31668 49416
rect 30975 49385 30987 49388
rect 30929 49379 30987 49385
rect 31662 49376 31668 49388
rect 31720 49376 31726 49428
rect 13262 49348 13268 49360
rect 13223 49320 13268 49348
rect 13262 49308 13268 49320
rect 13320 49308 13326 49360
rect 15010 49348 15016 49360
rect 14108 49320 15016 49348
rect 13722 49280 13728 49292
rect 13683 49252 13728 49280
rect 13722 49240 13728 49252
rect 13780 49240 13786 49292
rect 13909 49283 13967 49289
rect 13909 49249 13921 49283
rect 13955 49249 13967 49283
rect 13909 49243 13967 49249
rect 13538 49172 13544 49224
rect 13596 49212 13602 49224
rect 13924 49212 13952 49243
rect 13998 49240 14004 49292
rect 14056 49280 14062 49292
rect 14108 49289 14136 49320
rect 15010 49308 15016 49320
rect 15068 49308 15074 49360
rect 14093 49283 14151 49289
rect 14093 49280 14105 49283
rect 14056 49252 14105 49280
rect 14056 49240 14062 49252
rect 14093 49249 14105 49252
rect 14139 49249 14151 49283
rect 14093 49243 14151 49249
rect 14737 49283 14795 49289
rect 14737 49249 14749 49283
rect 14783 49280 14795 49283
rect 15286 49280 15292 49292
rect 14783 49252 15292 49280
rect 14783 49249 14795 49252
rect 14737 49243 14795 49249
rect 13596 49184 13952 49212
rect 13596 49172 13602 49184
rect 13173 49147 13231 49153
rect 13173 49113 13185 49147
rect 13219 49144 13231 49147
rect 13262 49144 13268 49156
rect 13219 49116 13268 49144
rect 13219 49113 13231 49116
rect 13173 49107 13231 49113
rect 13262 49104 13268 49116
rect 13320 49144 13326 49156
rect 14752 49144 14780 49243
rect 15286 49240 15292 49252
rect 15344 49280 15350 49292
rect 15381 49283 15439 49289
rect 15381 49280 15393 49283
rect 15344 49252 15393 49280
rect 15344 49240 15350 49252
rect 15381 49249 15393 49252
rect 15427 49249 15439 49283
rect 15381 49243 15439 49249
rect 15470 49240 15476 49292
rect 15528 49280 15534 49292
rect 15657 49283 15715 49289
rect 15657 49280 15669 49283
rect 15528 49252 15669 49280
rect 15528 49240 15534 49252
rect 15657 49249 15669 49252
rect 15703 49249 15715 49283
rect 15657 49243 15715 49249
rect 17402 49240 17408 49292
rect 17460 49280 17466 49292
rect 18233 49283 18291 49289
rect 18233 49280 18245 49283
rect 17460 49252 18245 49280
rect 17460 49240 17466 49252
rect 18233 49249 18245 49252
rect 18279 49280 18291 49283
rect 18785 49283 18843 49289
rect 18279 49252 18736 49280
rect 18279 49249 18291 49252
rect 18233 49243 18291 49249
rect 17773 49215 17831 49221
rect 17773 49181 17785 49215
rect 17819 49212 17831 49215
rect 17862 49212 17868 49224
rect 17819 49184 17868 49212
rect 17819 49181 17831 49184
rect 17773 49175 17831 49181
rect 17862 49172 17868 49184
rect 17920 49212 17926 49224
rect 18049 49215 18107 49221
rect 18049 49212 18061 49215
rect 17920 49184 18061 49212
rect 17920 49172 17926 49184
rect 18049 49181 18061 49184
rect 18095 49212 18107 49215
rect 18598 49212 18604 49224
rect 18095 49184 18604 49212
rect 18095 49181 18107 49184
rect 18049 49175 18107 49181
rect 18598 49172 18604 49184
rect 18656 49172 18662 49224
rect 18708 49212 18736 49252
rect 18785 49249 18797 49283
rect 18831 49280 18843 49283
rect 18966 49280 18972 49292
rect 18831 49252 18972 49280
rect 18831 49249 18843 49252
rect 18785 49243 18843 49249
rect 18966 49240 18972 49252
rect 19024 49240 19030 49292
rect 19797 49283 19855 49289
rect 19797 49249 19809 49283
rect 19843 49280 19855 49283
rect 20622 49280 20628 49292
rect 19843 49252 20628 49280
rect 19843 49249 19855 49252
rect 19797 49243 19855 49249
rect 20622 49240 20628 49252
rect 20680 49240 20686 49292
rect 21560 49280 21588 49376
rect 21637 49351 21695 49357
rect 21637 49317 21649 49351
rect 21683 49348 21695 49351
rect 24044 49348 24072 49376
rect 26513 49351 26571 49357
rect 21683 49320 22692 49348
rect 24044 49320 24532 49348
rect 21683 49317 21695 49320
rect 21637 49311 21695 49317
rect 22664 49292 22692 49320
rect 21729 49283 21787 49289
rect 21729 49280 21741 49283
rect 21560 49252 21741 49280
rect 21729 49249 21741 49252
rect 21775 49249 21787 49283
rect 22278 49280 22284 49292
rect 22239 49252 22284 49280
rect 21729 49243 21787 49249
rect 22278 49240 22284 49252
rect 22336 49240 22342 49292
rect 22646 49280 22652 49292
rect 22607 49252 22652 49280
rect 22646 49240 22652 49252
rect 22704 49240 22710 49292
rect 23566 49240 23572 49292
rect 23624 49280 23630 49292
rect 23661 49283 23719 49289
rect 23661 49280 23673 49283
rect 23624 49252 23673 49280
rect 23624 49240 23630 49252
rect 23661 49249 23673 49252
rect 23707 49249 23719 49283
rect 24026 49280 24032 49292
rect 23987 49252 24032 49280
rect 23661 49243 23719 49249
rect 24026 49240 24032 49252
rect 24084 49240 24090 49292
rect 24504 49289 24532 49320
rect 26513 49317 26525 49351
rect 26559 49348 26571 49351
rect 26786 49348 26792 49360
rect 26559 49320 26792 49348
rect 26559 49317 26571 49320
rect 26513 49311 26571 49317
rect 26786 49308 26792 49320
rect 26844 49308 26850 49360
rect 27522 49348 27528 49360
rect 27483 49320 27528 49348
rect 27522 49308 27528 49320
rect 27580 49308 27586 49360
rect 27985 49351 28043 49357
rect 27985 49317 27997 49351
rect 28031 49348 28043 49351
rect 29270 49348 29276 49360
rect 28031 49320 29276 49348
rect 28031 49317 28043 49320
rect 27985 49311 28043 49317
rect 29270 49308 29276 49320
rect 29328 49308 29334 49360
rect 24489 49283 24547 49289
rect 24489 49249 24501 49283
rect 24535 49249 24547 49283
rect 26694 49280 26700 49292
rect 26655 49252 26700 49280
rect 24489 49243 24547 49249
rect 26694 49240 26700 49252
rect 26752 49240 26758 49292
rect 28537 49283 28595 49289
rect 28537 49249 28549 49283
rect 28583 49280 28595 49283
rect 28718 49280 28724 49292
rect 28583 49252 28724 49280
rect 28583 49249 28595 49252
rect 28537 49243 28595 49249
rect 28718 49240 28724 49252
rect 28776 49240 28782 49292
rect 28810 49240 28816 49292
rect 28868 49280 28874 49292
rect 29914 49280 29920 49292
rect 28868 49252 28961 49280
rect 29875 49252 29920 49280
rect 28868 49240 28874 49252
rect 29914 49240 29920 49252
rect 29972 49240 29978 49292
rect 19702 49212 19708 49224
rect 18708 49184 19708 49212
rect 19702 49172 19708 49184
rect 19760 49172 19766 49224
rect 24762 49212 24768 49224
rect 24723 49184 24768 49212
rect 24762 49172 24768 49184
rect 24820 49172 24826 49224
rect 27062 49212 27068 49224
rect 27023 49184 27068 49212
rect 27062 49172 27068 49184
rect 27120 49172 27126 49224
rect 27982 49172 27988 49224
rect 28040 49212 28046 49224
rect 28828 49212 28856 49240
rect 28040 49184 28856 49212
rect 28997 49215 29055 49221
rect 28040 49172 28046 49184
rect 28997 49181 29009 49215
rect 29043 49212 29055 49215
rect 29454 49212 29460 49224
rect 29043 49184 29460 49212
rect 29043 49181 29055 49184
rect 28997 49175 29055 49181
rect 29454 49172 29460 49184
rect 29512 49212 29518 49224
rect 29825 49215 29883 49221
rect 29825 49212 29837 49215
rect 29512 49184 29837 49212
rect 29512 49172 29518 49184
rect 29825 49181 29837 49184
rect 29871 49181 29883 49215
rect 29825 49175 29883 49181
rect 18690 49144 18696 49156
rect 13320 49116 14780 49144
rect 18651 49116 18696 49144
rect 13320 49104 13326 49116
rect 18690 49104 18696 49116
rect 18748 49104 18754 49156
rect 22370 49104 22376 49156
rect 22428 49144 22434 49156
rect 22557 49147 22615 49153
rect 22557 49144 22569 49147
rect 22428 49116 22569 49144
rect 22428 49104 22434 49116
rect 22557 49113 22569 49116
rect 22603 49113 22615 49147
rect 22557 49107 22615 49113
rect 14826 49036 14832 49088
rect 14884 49076 14890 49088
rect 15013 49079 15071 49085
rect 15013 49076 15025 49079
rect 14884 49048 15025 49076
rect 14884 49036 14890 49048
rect 15013 49045 15025 49048
rect 15059 49045 15071 49079
rect 15013 49039 15071 49045
rect 16945 49079 17003 49085
rect 16945 49045 16957 49079
rect 16991 49076 17003 49079
rect 17770 49076 17776 49088
rect 16991 49048 17776 49076
rect 16991 49045 17003 49048
rect 16945 49039 17003 49045
rect 17770 49036 17776 49048
rect 17828 49036 17834 49088
rect 19981 49079 20039 49085
rect 19981 49045 19993 49079
rect 20027 49076 20039 49079
rect 23842 49076 23848 49088
rect 20027 49048 23848 49076
rect 20027 49045 20039 49048
rect 19981 49039 20039 49045
rect 23842 49036 23848 49048
rect 23900 49036 23906 49088
rect 25869 49079 25927 49085
rect 25869 49045 25881 49079
rect 25915 49076 25927 49079
rect 25958 49076 25964 49088
rect 25915 49048 25964 49076
rect 25915 49045 25927 49048
rect 25869 49039 25927 49045
rect 25958 49036 25964 49048
rect 26016 49036 26022 49088
rect 26234 49076 26240 49088
rect 26195 49048 26240 49076
rect 26234 49036 26240 49048
rect 26292 49036 26298 49088
rect 31202 49076 31208 49088
rect 31163 49048 31208 49076
rect 31202 49036 31208 49048
rect 31260 49036 31266 49088
rect 1104 48986 38824 49008
rect 1104 48934 4246 48986
rect 4298 48934 4310 48986
rect 4362 48934 4374 48986
rect 4426 48934 4438 48986
rect 4490 48934 34966 48986
rect 35018 48934 35030 48986
rect 35082 48934 35094 48986
rect 35146 48934 35158 48986
rect 35210 48934 38824 48986
rect 1104 48912 38824 48934
rect 13173 48875 13231 48881
rect 13173 48841 13185 48875
rect 13219 48872 13231 48875
rect 13998 48872 14004 48884
rect 13219 48844 14004 48872
rect 13219 48841 13231 48844
rect 13173 48835 13231 48841
rect 13998 48832 14004 48844
rect 14056 48832 14062 48884
rect 15286 48832 15292 48884
rect 15344 48872 15350 48884
rect 15749 48875 15807 48881
rect 15749 48872 15761 48875
rect 15344 48844 15761 48872
rect 15344 48832 15350 48844
rect 15749 48841 15761 48844
rect 15795 48841 15807 48875
rect 17402 48872 17408 48884
rect 17363 48844 17408 48872
rect 15749 48835 15807 48841
rect 17402 48832 17408 48844
rect 17460 48832 17466 48884
rect 17862 48872 17868 48884
rect 17823 48844 17868 48872
rect 17862 48832 17868 48844
rect 17920 48832 17926 48884
rect 18230 48872 18236 48884
rect 18191 48844 18236 48872
rect 18230 48832 18236 48844
rect 18288 48832 18294 48884
rect 18601 48875 18659 48881
rect 18601 48841 18613 48875
rect 18647 48872 18659 48875
rect 20070 48872 20076 48884
rect 18647 48844 20076 48872
rect 18647 48841 18659 48844
rect 18601 48835 18659 48841
rect 15378 48804 15384 48816
rect 15339 48776 15384 48804
rect 15378 48764 15384 48776
rect 15436 48764 15442 48816
rect 12805 48739 12863 48745
rect 12805 48705 12817 48739
rect 12851 48736 12863 48739
rect 12851 48708 13584 48736
rect 12851 48705 12863 48708
rect 12805 48699 12863 48705
rect 13556 48680 13584 48708
rect 13262 48668 13268 48680
rect 13223 48640 13268 48668
rect 13262 48628 13268 48640
rect 13320 48628 13326 48680
rect 13538 48668 13544 48680
rect 13499 48640 13544 48668
rect 13538 48628 13544 48640
rect 13596 48628 13602 48680
rect 18049 48671 18107 48677
rect 18049 48637 18061 48671
rect 18095 48668 18107 48671
rect 18616 48668 18644 48835
rect 20070 48832 20076 48844
rect 20128 48872 20134 48884
rect 20533 48875 20591 48881
rect 20533 48872 20545 48875
rect 20128 48844 20545 48872
rect 20128 48832 20134 48844
rect 20533 48841 20545 48844
rect 20579 48872 20591 48875
rect 20622 48872 20628 48884
rect 20579 48844 20628 48872
rect 20579 48841 20591 48844
rect 20533 48835 20591 48841
rect 20622 48832 20628 48844
rect 20680 48832 20686 48884
rect 20990 48872 20996 48884
rect 20951 48844 20996 48872
rect 20990 48832 20996 48844
rect 21048 48832 21054 48884
rect 24946 48832 24952 48884
rect 25004 48872 25010 48884
rect 25406 48872 25412 48884
rect 25004 48844 25412 48872
rect 25004 48832 25010 48844
rect 25406 48832 25412 48844
rect 25464 48872 25470 48884
rect 25777 48875 25835 48881
rect 25777 48872 25789 48875
rect 25464 48844 25789 48872
rect 25464 48832 25470 48844
rect 25777 48841 25789 48844
rect 25823 48872 25835 48875
rect 26694 48872 26700 48884
rect 25823 48844 26700 48872
rect 25823 48841 25835 48844
rect 25777 48835 25835 48841
rect 26694 48832 26700 48844
rect 26752 48832 26758 48884
rect 28718 48872 28724 48884
rect 28679 48844 28724 48872
rect 28718 48832 28724 48844
rect 28776 48832 28782 48884
rect 29914 48832 29920 48884
rect 29972 48872 29978 48884
rect 30742 48872 30748 48884
rect 29972 48844 30748 48872
rect 29972 48832 29978 48844
rect 30742 48832 30748 48844
rect 30800 48872 30806 48884
rect 31021 48875 31079 48881
rect 31021 48872 31033 48875
rect 30800 48844 31033 48872
rect 30800 48832 30806 48844
rect 31021 48841 31033 48844
rect 31067 48872 31079 48875
rect 31202 48872 31208 48884
rect 31067 48844 31208 48872
rect 31067 48841 31079 48844
rect 31021 48835 31079 48841
rect 31202 48832 31208 48844
rect 31260 48832 31266 48884
rect 31386 48872 31392 48884
rect 31347 48844 31392 48872
rect 31386 48832 31392 48844
rect 31444 48832 31450 48884
rect 23109 48807 23167 48813
rect 23109 48804 23121 48807
rect 22112 48776 23121 48804
rect 22112 48748 22140 48776
rect 23109 48773 23121 48776
rect 23155 48804 23167 48807
rect 23566 48804 23572 48816
rect 23155 48776 23572 48804
rect 23155 48773 23167 48776
rect 23109 48767 23167 48773
rect 23566 48764 23572 48776
rect 23624 48764 23630 48816
rect 26605 48807 26663 48813
rect 26605 48773 26617 48807
rect 26651 48804 26663 48807
rect 27614 48804 27620 48816
rect 26651 48776 27620 48804
rect 26651 48773 26663 48776
rect 26605 48767 26663 48773
rect 27614 48764 27620 48776
rect 27672 48764 27678 48816
rect 18969 48739 19027 48745
rect 18969 48705 18981 48739
rect 19015 48736 19027 48739
rect 19242 48736 19248 48748
rect 19015 48708 19248 48736
rect 19015 48705 19027 48708
rect 18969 48699 19027 48705
rect 19242 48696 19248 48708
rect 19300 48696 19306 48748
rect 19518 48696 19524 48748
rect 19576 48736 19582 48748
rect 19889 48739 19947 48745
rect 19889 48736 19901 48739
rect 19576 48708 19901 48736
rect 19576 48696 19582 48708
rect 19889 48705 19901 48708
rect 19935 48705 19947 48739
rect 22094 48736 22100 48748
rect 19889 48699 19947 48705
rect 21652 48708 22100 48736
rect 19426 48668 19432 48680
rect 18095 48640 18644 48668
rect 19387 48640 19432 48668
rect 18095 48637 18107 48640
rect 18049 48631 18107 48637
rect 19426 48628 19432 48640
rect 19484 48628 19490 48680
rect 19978 48668 19984 48680
rect 19939 48640 19984 48668
rect 19978 48628 19984 48640
rect 20036 48628 20042 48680
rect 20346 48628 20352 48680
rect 20404 48668 20410 48680
rect 21652 48677 21680 48708
rect 22094 48696 22100 48708
rect 22152 48696 22158 48748
rect 22370 48736 22376 48748
rect 22204 48708 22376 48736
rect 22204 48677 22232 48708
rect 22370 48696 22376 48708
rect 22428 48736 22434 48748
rect 23014 48736 23020 48748
rect 22428 48708 23020 48736
rect 22428 48696 22434 48708
rect 23014 48696 23020 48708
rect 23072 48696 23078 48748
rect 23477 48739 23535 48745
rect 23477 48705 23489 48739
rect 23523 48736 23535 48739
rect 25501 48739 25559 48745
rect 23523 48708 24900 48736
rect 23523 48705 23535 48708
rect 23477 48699 23535 48705
rect 21177 48671 21235 48677
rect 21177 48668 21189 48671
rect 20404 48640 21189 48668
rect 20404 48628 20410 48640
rect 21177 48637 21189 48640
rect 21223 48637 21235 48671
rect 21177 48631 21235 48637
rect 21637 48671 21695 48677
rect 21637 48637 21649 48671
rect 21683 48637 21695 48671
rect 21637 48631 21695 48637
rect 22189 48671 22247 48677
rect 22189 48637 22201 48671
rect 22235 48637 22247 48671
rect 22554 48668 22560 48680
rect 22515 48640 22560 48668
rect 22189 48631 22247 48637
rect 21652 48600 21680 48631
rect 22554 48628 22560 48640
rect 22612 48628 22618 48680
rect 22738 48668 22744 48680
rect 22699 48640 22744 48668
rect 22738 48628 22744 48640
rect 22796 48628 22802 48680
rect 23753 48671 23811 48677
rect 23753 48637 23765 48671
rect 23799 48668 23811 48671
rect 23799 48640 24348 48668
rect 23799 48637 23811 48640
rect 23753 48631 23811 48637
rect 20916 48572 21680 48600
rect 20916 48544 20944 48572
rect 14642 48532 14648 48544
rect 14603 48504 14648 48532
rect 14642 48492 14648 48504
rect 14700 48492 14706 48544
rect 17129 48535 17187 48541
rect 17129 48501 17141 48535
rect 17175 48532 17187 48535
rect 17218 48532 17224 48544
rect 17175 48504 17224 48532
rect 17175 48501 17187 48504
rect 17129 48495 17187 48501
rect 17218 48492 17224 48504
rect 17276 48492 17282 48544
rect 20898 48532 20904 48544
rect 20859 48504 20904 48532
rect 20898 48492 20904 48504
rect 20956 48492 20962 48544
rect 21545 48535 21603 48541
rect 21545 48501 21557 48535
rect 21591 48532 21603 48535
rect 22278 48532 22284 48544
rect 21591 48504 22284 48532
rect 21591 48501 21603 48504
rect 21545 48495 21603 48501
rect 22278 48492 22284 48504
rect 22336 48532 22342 48544
rect 22554 48532 22560 48544
rect 22336 48504 22560 48532
rect 22336 48492 22342 48504
rect 22554 48492 22560 48504
rect 22612 48492 22618 48544
rect 23937 48535 23995 48541
rect 23937 48501 23949 48535
rect 23983 48532 23995 48535
rect 24118 48532 24124 48544
rect 23983 48504 24124 48532
rect 23983 48501 23995 48504
rect 23937 48495 23995 48501
rect 24118 48492 24124 48504
rect 24176 48492 24182 48544
rect 24320 48541 24348 48640
rect 24765 48603 24823 48609
rect 24765 48569 24777 48603
rect 24811 48569 24823 48603
rect 24872 48600 24900 48708
rect 25501 48705 25513 48739
rect 25547 48736 25559 48739
rect 26234 48736 26240 48748
rect 25547 48708 26240 48736
rect 25547 48705 25559 48708
rect 25501 48699 25559 48705
rect 26234 48696 26240 48708
rect 26292 48736 26298 48748
rect 27709 48739 27767 48745
rect 26292 48708 26832 48736
rect 26292 48696 26298 48708
rect 24949 48671 25007 48677
rect 24949 48637 24961 48671
rect 24995 48668 25007 48671
rect 25038 48668 25044 48680
rect 24995 48640 25044 48668
rect 24995 48637 25007 48640
rect 24949 48631 25007 48637
rect 25038 48628 25044 48640
rect 25096 48628 25102 48680
rect 26804 48677 26832 48708
rect 27709 48705 27721 48739
rect 27755 48736 27767 48739
rect 29454 48736 29460 48748
rect 27755 48708 29460 48736
rect 27755 48705 27767 48708
rect 27709 48699 27767 48705
rect 29454 48696 29460 48708
rect 29512 48696 29518 48748
rect 30282 48736 30288 48748
rect 30243 48708 30288 48736
rect 30282 48696 30288 48708
rect 30340 48696 30346 48748
rect 26789 48671 26847 48677
rect 26789 48637 26801 48671
rect 26835 48637 26847 48671
rect 26789 48631 26847 48637
rect 26973 48671 27031 48677
rect 26973 48637 26985 48671
rect 27019 48637 27031 48671
rect 27154 48668 27160 48680
rect 27115 48640 27160 48668
rect 26973 48631 27031 48637
rect 25133 48603 25191 48609
rect 24872 48572 25084 48600
rect 24765 48563 24823 48569
rect 24305 48535 24363 48541
rect 24305 48501 24317 48535
rect 24351 48532 24363 48535
rect 24673 48535 24731 48541
rect 24673 48532 24685 48535
rect 24351 48504 24685 48532
rect 24351 48501 24363 48504
rect 24305 48495 24363 48501
rect 24673 48501 24685 48504
rect 24719 48532 24731 48535
rect 24780 48532 24808 48563
rect 24946 48532 24952 48544
rect 24719 48504 24952 48532
rect 24719 48501 24731 48504
rect 24673 48495 24731 48501
rect 24946 48492 24952 48504
rect 25004 48492 25010 48544
rect 25056 48541 25084 48572
rect 25133 48569 25145 48603
rect 25179 48600 25191 48603
rect 25222 48600 25228 48612
rect 25179 48572 25228 48600
rect 25179 48569 25191 48572
rect 25133 48563 25191 48569
rect 25222 48560 25228 48572
rect 25280 48560 25286 48612
rect 26326 48560 26332 48612
rect 26384 48600 26390 48612
rect 26988 48600 27016 48631
rect 27154 48628 27160 48640
rect 27212 48628 27218 48680
rect 28166 48668 28172 48680
rect 28127 48640 28172 48668
rect 28166 48628 28172 48640
rect 28224 48628 28230 48680
rect 29641 48671 29699 48677
rect 29641 48668 29653 48671
rect 29288 48640 29653 48668
rect 26384 48572 27016 48600
rect 26384 48560 26390 48572
rect 29288 48544 29316 48640
rect 29641 48637 29653 48640
rect 29687 48637 29699 48671
rect 29641 48631 29699 48637
rect 29822 48628 29828 48680
rect 29880 48668 29886 48680
rect 30101 48671 30159 48677
rect 30101 48668 30113 48671
rect 29880 48640 30113 48668
rect 29880 48628 29886 48640
rect 30101 48637 30113 48640
rect 30147 48637 30159 48671
rect 31202 48668 31208 48680
rect 31115 48640 31208 48668
rect 30101 48631 30159 48637
rect 31202 48628 31208 48640
rect 31260 48668 31266 48680
rect 31665 48671 31723 48677
rect 31665 48668 31677 48671
rect 31260 48640 31677 48668
rect 31260 48628 31266 48640
rect 31665 48637 31677 48640
rect 31711 48637 31723 48671
rect 31665 48631 31723 48637
rect 25041 48535 25099 48541
rect 25041 48501 25053 48535
rect 25087 48532 25099 48535
rect 25774 48532 25780 48544
rect 25087 48504 25780 48532
rect 25087 48501 25099 48504
rect 25041 48495 25099 48501
rect 25774 48492 25780 48504
rect 25832 48532 25838 48544
rect 25958 48532 25964 48544
rect 25832 48504 25964 48532
rect 25832 48492 25838 48504
rect 25958 48492 25964 48504
rect 26016 48492 26022 48544
rect 26237 48535 26295 48541
rect 26237 48501 26249 48535
rect 26283 48532 26295 48535
rect 26786 48532 26792 48544
rect 26283 48504 26792 48532
rect 26283 48501 26295 48504
rect 26237 48495 26295 48501
rect 26786 48492 26792 48504
rect 26844 48532 26850 48544
rect 27430 48532 27436 48544
rect 26844 48504 27436 48532
rect 26844 48492 26850 48504
rect 27430 48492 27436 48504
rect 27488 48492 27494 48544
rect 27982 48532 27988 48544
rect 27943 48504 27988 48532
rect 27982 48492 27988 48504
rect 28040 48492 28046 48544
rect 28353 48535 28411 48541
rect 28353 48501 28365 48535
rect 28399 48532 28411 48535
rect 28534 48532 28540 48544
rect 28399 48504 28540 48532
rect 28399 48501 28411 48504
rect 28353 48495 28411 48501
rect 28534 48492 28540 48504
rect 28592 48532 28598 48544
rect 28810 48532 28816 48544
rect 28592 48504 28816 48532
rect 28592 48492 28598 48504
rect 28810 48492 28816 48504
rect 28868 48492 28874 48544
rect 29089 48535 29147 48541
rect 29089 48501 29101 48535
rect 29135 48532 29147 48535
rect 29270 48532 29276 48544
rect 29135 48504 29276 48532
rect 29135 48501 29147 48504
rect 29089 48495 29147 48501
rect 29270 48492 29276 48504
rect 29328 48492 29334 48544
rect 30650 48532 30656 48544
rect 30611 48504 30656 48532
rect 30650 48492 30656 48504
rect 30708 48492 30714 48544
rect 1104 48442 38824 48464
rect 1104 48390 19606 48442
rect 19658 48390 19670 48442
rect 19722 48390 19734 48442
rect 19786 48390 19798 48442
rect 19850 48390 38824 48442
rect 1104 48368 38824 48390
rect 9122 48288 9128 48340
rect 9180 48328 9186 48340
rect 9398 48328 9404 48340
rect 9180 48300 9404 48328
rect 9180 48288 9186 48300
rect 9398 48288 9404 48300
rect 9456 48288 9462 48340
rect 13538 48288 13544 48340
rect 13596 48328 13602 48340
rect 13725 48331 13783 48337
rect 13725 48328 13737 48331
rect 13596 48300 13737 48328
rect 13596 48288 13602 48300
rect 13725 48297 13737 48300
rect 13771 48328 13783 48331
rect 15470 48328 15476 48340
rect 13771 48300 15476 48328
rect 13771 48297 13783 48300
rect 13725 48291 13783 48297
rect 15470 48288 15476 48300
rect 15528 48288 15534 48340
rect 17218 48288 17224 48340
rect 17276 48328 17282 48340
rect 17957 48331 18015 48337
rect 17957 48328 17969 48331
rect 17276 48300 17969 48328
rect 17276 48288 17282 48300
rect 17957 48297 17969 48300
rect 18003 48328 18015 48331
rect 18966 48328 18972 48340
rect 18003 48300 18972 48328
rect 18003 48297 18015 48300
rect 17957 48291 18015 48297
rect 18966 48288 18972 48300
rect 19024 48288 19030 48340
rect 22005 48331 22063 48337
rect 22005 48297 22017 48331
rect 22051 48328 22063 48331
rect 22646 48328 22652 48340
rect 22051 48300 22652 48328
rect 22051 48297 22063 48300
rect 22005 48291 22063 48297
rect 22646 48288 22652 48300
rect 22704 48328 22710 48340
rect 22704 48300 23428 48328
rect 22704 48288 22710 48300
rect 11606 48260 11612 48272
rect 11567 48232 11612 48260
rect 11606 48220 11612 48232
rect 11664 48220 11670 48272
rect 15102 48260 15108 48272
rect 15063 48232 15108 48260
rect 15102 48220 15108 48232
rect 15160 48220 15166 48272
rect 18414 48260 18420 48272
rect 18375 48232 18420 48260
rect 18414 48220 18420 48232
rect 18472 48220 18478 48272
rect 18598 48220 18604 48272
rect 18656 48260 18662 48272
rect 18785 48263 18843 48269
rect 18785 48260 18797 48263
rect 18656 48232 18797 48260
rect 18656 48220 18662 48232
rect 18785 48229 18797 48232
rect 18831 48260 18843 48263
rect 19978 48260 19984 48272
rect 18831 48232 19984 48260
rect 18831 48229 18843 48232
rect 18785 48223 18843 48229
rect 19978 48220 19984 48232
rect 20036 48220 20042 48272
rect 20438 48220 20444 48272
rect 20496 48260 20502 48272
rect 20533 48263 20591 48269
rect 20533 48260 20545 48263
rect 20496 48232 20545 48260
rect 20496 48220 20502 48232
rect 20533 48229 20545 48232
rect 20579 48229 20591 48263
rect 22370 48260 22376 48272
rect 22331 48232 22376 48260
rect 20533 48223 20591 48229
rect 22370 48220 22376 48232
rect 22428 48220 22434 48272
rect 23014 48260 23020 48272
rect 22975 48232 23020 48260
rect 23014 48220 23020 48232
rect 23072 48220 23078 48272
rect 23400 48260 23428 48300
rect 25038 48288 25044 48340
rect 25096 48328 25102 48340
rect 25590 48328 25596 48340
rect 25096 48300 25596 48328
rect 25096 48288 25102 48300
rect 25590 48288 25596 48300
rect 25648 48328 25654 48340
rect 28166 48328 28172 48340
rect 25648 48300 28172 48328
rect 25648 48288 25654 48300
rect 28166 48288 28172 48300
rect 28224 48288 28230 48340
rect 28629 48331 28687 48337
rect 28629 48297 28641 48331
rect 28675 48328 28687 48331
rect 28718 48328 28724 48340
rect 28675 48300 28724 48328
rect 28675 48297 28687 48300
rect 28629 48291 28687 48297
rect 28718 48288 28724 48300
rect 28776 48288 28782 48340
rect 29454 48328 29460 48340
rect 29415 48300 29460 48328
rect 29454 48288 29460 48300
rect 29512 48288 29518 48340
rect 29822 48328 29828 48340
rect 29783 48300 29828 48328
rect 29822 48288 29828 48300
rect 29880 48288 29886 48340
rect 23566 48260 23572 48272
rect 23400 48232 23572 48260
rect 23566 48220 23572 48232
rect 23624 48220 23630 48272
rect 24118 48220 24124 48272
rect 24176 48260 24182 48272
rect 26418 48260 26424 48272
rect 24176 48232 26424 48260
rect 24176 48220 24182 48232
rect 10962 48152 10968 48204
rect 11020 48192 11026 48204
rect 12250 48192 12256 48204
rect 11020 48164 12256 48192
rect 11020 48152 11026 48164
rect 12250 48152 12256 48164
rect 12308 48152 12314 48204
rect 12621 48195 12679 48201
rect 12621 48161 12633 48195
rect 12667 48161 12679 48195
rect 12802 48192 12808 48204
rect 12763 48164 12808 48192
rect 12621 48155 12679 48161
rect 12158 48124 12164 48136
rect 12119 48096 12164 48124
rect 12158 48084 12164 48096
rect 12216 48084 12222 48136
rect 11422 47988 11428 48000
rect 11383 47960 11428 47988
rect 11422 47948 11428 47960
rect 11480 47988 11486 48000
rect 12636 47988 12664 48155
rect 12802 48152 12808 48164
rect 12860 48152 12866 48204
rect 13909 48195 13967 48201
rect 13909 48161 13921 48195
rect 13955 48192 13967 48195
rect 14274 48192 14280 48204
rect 13955 48164 14280 48192
rect 13955 48161 13967 48164
rect 13909 48155 13967 48161
rect 14274 48152 14280 48164
rect 14332 48192 14338 48204
rect 14642 48192 14648 48204
rect 14332 48164 14648 48192
rect 14332 48152 14338 48164
rect 14642 48152 14648 48164
rect 14700 48152 14706 48204
rect 15749 48195 15807 48201
rect 15749 48161 15761 48195
rect 15795 48192 15807 48195
rect 15838 48192 15844 48204
rect 15795 48164 15844 48192
rect 15795 48161 15807 48164
rect 15749 48155 15807 48161
rect 15838 48152 15844 48164
rect 15896 48152 15902 48204
rect 15933 48195 15991 48201
rect 15933 48161 15945 48195
rect 15979 48161 15991 48195
rect 16114 48192 16120 48204
rect 16075 48164 16120 48192
rect 15933 48155 15991 48161
rect 13817 48127 13875 48133
rect 13817 48093 13829 48127
rect 13863 48124 13875 48127
rect 13998 48124 14004 48136
rect 13863 48096 14004 48124
rect 13863 48093 13875 48096
rect 13817 48087 13875 48093
rect 13998 48084 14004 48096
rect 14056 48084 14062 48136
rect 15948 48124 15976 48155
rect 16114 48152 16120 48164
rect 16172 48152 16178 48204
rect 19058 48192 19064 48204
rect 19019 48164 19064 48192
rect 19058 48152 19064 48164
rect 19116 48152 19122 48204
rect 19426 48192 19432 48204
rect 19387 48164 19432 48192
rect 19426 48152 19432 48164
rect 19484 48152 19490 48204
rect 19797 48195 19855 48201
rect 19797 48161 19809 48195
rect 19843 48192 19855 48195
rect 19996 48192 20024 48220
rect 21174 48192 21180 48204
rect 19843 48164 20024 48192
rect 21135 48164 21180 48192
rect 19843 48161 19855 48164
rect 19797 48155 19855 48161
rect 21174 48152 21180 48164
rect 21232 48152 21238 48204
rect 21450 48192 21456 48204
rect 21411 48164 21456 48192
rect 21450 48152 21456 48164
rect 21508 48152 21514 48204
rect 22554 48192 22560 48204
rect 22515 48164 22560 48192
rect 22554 48152 22560 48164
rect 22612 48192 22618 48204
rect 23293 48195 23351 48201
rect 23293 48192 23305 48195
rect 22612 48164 23305 48192
rect 22612 48152 22618 48164
rect 23293 48161 23305 48164
rect 23339 48161 23351 48195
rect 23842 48192 23848 48204
rect 23803 48164 23848 48192
rect 23293 48155 23351 48161
rect 23842 48152 23848 48164
rect 23900 48152 23906 48204
rect 24213 48195 24271 48201
rect 24213 48161 24225 48195
rect 24259 48161 24271 48195
rect 24486 48192 24492 48204
rect 24213 48155 24271 48161
rect 24320 48164 24492 48192
rect 16666 48124 16672 48136
rect 14660 48096 16672 48124
rect 13357 48059 13415 48065
rect 13357 48025 13369 48059
rect 13403 48056 13415 48059
rect 13722 48056 13728 48068
rect 13403 48028 13728 48056
rect 13403 48025 13415 48028
rect 13357 48019 13415 48025
rect 13722 48016 13728 48028
rect 13780 48056 13786 48068
rect 13780 48028 14136 48056
rect 13780 48016 13786 48028
rect 14108 47997 14136 48028
rect 14660 48000 14688 48096
rect 16666 48084 16672 48096
rect 16724 48084 16730 48136
rect 19978 48124 19984 48136
rect 19939 48096 19984 48124
rect 19978 48084 19984 48096
rect 20036 48084 20042 48136
rect 20714 48084 20720 48136
rect 20772 48124 20778 48136
rect 21361 48127 21419 48133
rect 21361 48124 21373 48127
rect 20772 48096 21373 48124
rect 20772 48084 20778 48096
rect 21361 48093 21373 48096
rect 21407 48093 21419 48127
rect 21361 48087 21419 48093
rect 22465 48127 22523 48133
rect 22465 48093 22477 48127
rect 22511 48093 22523 48127
rect 22465 48087 22523 48093
rect 15562 48056 15568 48068
rect 15523 48028 15568 48056
rect 15562 48016 15568 48028
rect 15620 48016 15626 48068
rect 19886 48016 19892 48068
rect 19944 48056 19950 48068
rect 20254 48056 20260 48068
rect 19944 48028 20260 48056
rect 19944 48016 19950 48028
rect 20254 48016 20260 48028
rect 20312 48016 20318 48068
rect 21082 48016 21088 48068
rect 21140 48056 21146 48068
rect 22480 48056 22508 48087
rect 23382 48084 23388 48136
rect 23440 48124 23446 48136
rect 24228 48124 24256 48155
rect 24320 48136 24348 48164
rect 24486 48152 24492 48164
rect 24544 48192 24550 48204
rect 25148 48201 25176 48232
rect 26418 48220 26424 48232
rect 26476 48220 26482 48272
rect 26513 48263 26571 48269
rect 26513 48229 26525 48263
rect 26559 48260 26571 48263
rect 26602 48260 26608 48272
rect 26559 48232 26608 48260
rect 26559 48229 26571 48232
rect 26513 48223 26571 48229
rect 26602 48220 26608 48232
rect 26660 48220 26666 48272
rect 27614 48220 27620 48272
rect 27672 48260 27678 48272
rect 28442 48260 28448 48272
rect 27672 48232 28448 48260
rect 27672 48220 27678 48232
rect 28442 48220 28448 48232
rect 28500 48260 28506 48272
rect 30745 48263 30803 48269
rect 30745 48260 30757 48263
rect 28500 48232 28856 48260
rect 28500 48220 28506 48232
rect 24581 48195 24639 48201
rect 24581 48192 24593 48195
rect 24544 48164 24593 48192
rect 24544 48152 24550 48164
rect 24581 48161 24593 48164
rect 24627 48161 24639 48195
rect 24581 48155 24639 48161
rect 25133 48195 25191 48201
rect 25133 48161 25145 48195
rect 25179 48161 25191 48195
rect 25133 48155 25191 48161
rect 26786 48152 26792 48204
rect 26844 48192 26850 48204
rect 26973 48195 27031 48201
rect 26973 48192 26985 48195
rect 26844 48164 26985 48192
rect 26844 48152 26850 48164
rect 26973 48161 26985 48164
rect 27019 48161 27031 48195
rect 26973 48155 27031 48161
rect 27062 48152 27068 48204
rect 27120 48192 27126 48204
rect 27157 48195 27215 48201
rect 27157 48192 27169 48195
rect 27120 48164 27169 48192
rect 27120 48152 27126 48164
rect 27157 48161 27169 48164
rect 27203 48161 27215 48195
rect 27157 48155 27215 48161
rect 27341 48195 27399 48201
rect 27341 48161 27353 48195
rect 27387 48192 27399 48195
rect 27522 48192 27528 48204
rect 27387 48164 27528 48192
rect 27387 48161 27399 48164
rect 27341 48155 27399 48161
rect 27522 48152 27528 48164
rect 27580 48152 27586 48204
rect 27798 48192 27804 48204
rect 27759 48164 27804 48192
rect 27798 48152 27804 48164
rect 27856 48152 27862 48204
rect 28534 48192 28540 48204
rect 28495 48164 28540 48192
rect 28534 48152 28540 48164
rect 28592 48152 28598 48204
rect 28828 48201 28856 48232
rect 29932 48232 30757 48260
rect 29932 48204 29960 48232
rect 30745 48229 30757 48232
rect 30791 48229 30803 48263
rect 30745 48223 30803 48229
rect 28813 48195 28871 48201
rect 28813 48161 28825 48195
rect 28859 48161 28871 48195
rect 29546 48192 29552 48204
rect 29507 48164 29552 48192
rect 28813 48155 28871 48161
rect 29546 48152 29552 48164
rect 29604 48152 29610 48204
rect 29914 48192 29920 48204
rect 29875 48164 29920 48192
rect 29914 48152 29920 48164
rect 29972 48152 29978 48204
rect 30009 48195 30067 48201
rect 30009 48161 30021 48195
rect 30055 48192 30067 48195
rect 30374 48192 30380 48204
rect 30055 48164 30380 48192
rect 30055 48161 30067 48164
rect 30009 48155 30067 48161
rect 30374 48152 30380 48164
rect 30432 48152 30438 48204
rect 23440 48096 24256 48124
rect 23440 48084 23446 48096
rect 24302 48084 24308 48136
rect 24360 48084 24366 48136
rect 24670 48124 24676 48136
rect 24631 48096 24676 48124
rect 24670 48084 24676 48096
rect 24728 48084 24734 48136
rect 27540 48124 27568 48152
rect 31113 48127 31171 48133
rect 31113 48124 31125 48127
rect 27540 48096 31125 48124
rect 31113 48093 31125 48096
rect 31159 48124 31171 48127
rect 31386 48124 31392 48136
rect 31159 48096 31392 48124
rect 31159 48093 31171 48096
rect 31113 48087 31171 48093
rect 31386 48084 31392 48096
rect 31444 48084 31450 48136
rect 23658 48056 23664 48068
rect 21140 48028 23664 48056
rect 21140 48016 21146 48028
rect 23658 48016 23664 48028
rect 23716 48016 23722 48068
rect 28074 48016 28080 48068
rect 28132 48056 28138 48068
rect 28902 48056 28908 48068
rect 28132 48028 28908 48056
rect 28132 48016 28138 48028
rect 28902 48016 28908 48028
rect 28960 48016 28966 48068
rect 29086 48016 29092 48068
rect 29144 48056 29150 48068
rect 29454 48056 29460 48068
rect 29144 48028 29460 48056
rect 29144 48016 29150 48028
rect 29454 48016 29460 48028
rect 29512 48016 29518 48068
rect 29549 48059 29607 48065
rect 29549 48025 29561 48059
rect 29595 48056 29607 48059
rect 29638 48056 29644 48068
rect 29595 48028 29644 48056
rect 29595 48025 29607 48028
rect 29549 48019 29607 48025
rect 29638 48016 29644 48028
rect 29696 48016 29702 48068
rect 11480 47960 12664 47988
rect 14093 47991 14151 47997
rect 11480 47948 11486 47960
rect 14093 47957 14105 47991
rect 14139 47957 14151 47991
rect 14642 47988 14648 48000
rect 14603 47960 14648 47988
rect 14093 47951 14151 47957
rect 14642 47948 14648 47960
rect 14700 47948 14706 48000
rect 23753 47991 23811 47997
rect 23753 47957 23765 47991
rect 23799 47988 23811 47991
rect 24026 47988 24032 48000
rect 23799 47960 24032 47988
rect 23799 47957 23811 47960
rect 23753 47951 23811 47957
rect 24026 47948 24032 47960
rect 24084 47948 24090 48000
rect 26234 47988 26240 48000
rect 26195 47960 26240 47988
rect 26234 47948 26240 47960
rect 26292 47948 26298 48000
rect 28994 47948 29000 48000
rect 29052 47988 29058 48000
rect 30193 47991 30251 47997
rect 30193 47988 30205 47991
rect 29052 47960 30205 47988
rect 29052 47948 29058 47960
rect 30193 47957 30205 47960
rect 30239 47957 30251 47991
rect 30193 47951 30251 47957
rect 30834 47948 30840 48000
rect 30892 47988 30898 48000
rect 31481 47991 31539 47997
rect 31481 47988 31493 47991
rect 30892 47960 31493 47988
rect 30892 47948 30898 47960
rect 31481 47957 31493 47960
rect 31527 47957 31539 47991
rect 31481 47951 31539 47957
rect 1104 47898 38824 47920
rect 1104 47846 4246 47898
rect 4298 47846 4310 47898
rect 4362 47846 4374 47898
rect 4426 47846 4438 47898
rect 4490 47846 34966 47898
rect 35018 47846 35030 47898
rect 35082 47846 35094 47898
rect 35146 47846 35158 47898
rect 35210 47846 38824 47898
rect 1104 47824 38824 47846
rect 10962 47784 10968 47796
rect 10923 47756 10968 47784
rect 10962 47744 10968 47756
rect 11020 47744 11026 47796
rect 11333 47787 11391 47793
rect 11333 47753 11345 47787
rect 11379 47784 11391 47787
rect 12802 47784 12808 47796
rect 11379 47756 12808 47784
rect 11379 47753 11391 47756
rect 11333 47747 11391 47753
rect 12802 47744 12808 47756
rect 12860 47784 12866 47796
rect 13170 47784 13176 47796
rect 12860 47756 13176 47784
rect 12860 47744 12866 47756
rect 13170 47744 13176 47756
rect 13228 47784 13234 47796
rect 13814 47784 13820 47796
rect 13228 47756 13820 47784
rect 13228 47744 13234 47756
rect 13814 47744 13820 47756
rect 13872 47744 13878 47796
rect 14274 47784 14280 47796
rect 14235 47756 14280 47784
rect 14274 47744 14280 47756
rect 14332 47744 14338 47796
rect 16666 47784 16672 47796
rect 16627 47756 16672 47784
rect 16666 47744 16672 47756
rect 16724 47744 16730 47796
rect 18598 47784 18604 47796
rect 18559 47756 18604 47784
rect 18598 47744 18604 47756
rect 18656 47744 18662 47796
rect 18969 47787 19027 47793
rect 18969 47753 18981 47787
rect 19015 47784 19027 47787
rect 19058 47784 19064 47796
rect 19015 47756 19064 47784
rect 19015 47753 19027 47756
rect 18969 47747 19027 47753
rect 19058 47744 19064 47756
rect 19116 47744 19122 47796
rect 19337 47787 19395 47793
rect 19337 47753 19349 47787
rect 19383 47784 19395 47787
rect 19426 47784 19432 47796
rect 19383 47756 19432 47784
rect 19383 47753 19395 47756
rect 19337 47747 19395 47753
rect 19426 47744 19432 47756
rect 19484 47744 19490 47796
rect 19613 47787 19671 47793
rect 19613 47753 19625 47787
rect 19659 47784 19671 47787
rect 20070 47784 20076 47796
rect 19659 47756 20076 47784
rect 19659 47753 19671 47756
rect 19613 47747 19671 47753
rect 20070 47744 20076 47756
rect 20128 47744 20134 47796
rect 21174 47744 21180 47796
rect 21232 47784 21238 47796
rect 21453 47787 21511 47793
rect 21453 47784 21465 47787
rect 21232 47756 21465 47784
rect 21232 47744 21238 47756
rect 21453 47753 21465 47756
rect 21499 47753 21511 47787
rect 21453 47747 21511 47753
rect 22738 47744 22744 47796
rect 22796 47784 22802 47796
rect 23382 47784 23388 47796
rect 22796 47756 23388 47784
rect 22796 47744 22802 47756
rect 23382 47744 23388 47756
rect 23440 47784 23446 47796
rect 23477 47787 23535 47793
rect 23477 47784 23489 47787
rect 23440 47756 23489 47784
rect 23440 47744 23446 47756
rect 23477 47753 23489 47756
rect 23523 47753 23535 47787
rect 23477 47747 23535 47753
rect 26973 47787 27031 47793
rect 26973 47753 26985 47787
rect 27019 47784 27031 47787
rect 27062 47784 27068 47796
rect 27019 47756 27068 47784
rect 27019 47753 27031 47756
rect 26973 47747 27031 47753
rect 27062 47744 27068 47756
rect 27120 47744 27126 47796
rect 29086 47784 29092 47796
rect 29047 47756 29092 47784
rect 29086 47744 29092 47756
rect 29144 47744 29150 47796
rect 31110 47784 31116 47796
rect 31071 47756 31116 47784
rect 31110 47744 31116 47756
rect 31168 47744 31174 47796
rect 11701 47719 11759 47725
rect 11701 47685 11713 47719
rect 11747 47716 11759 47719
rect 12158 47716 12164 47728
rect 11747 47688 12164 47716
rect 11747 47685 11759 47688
rect 11701 47679 11759 47685
rect 12158 47676 12164 47688
rect 12216 47716 12222 47728
rect 23109 47719 23167 47725
rect 12216 47688 13308 47716
rect 12216 47676 12222 47688
rect 12529 47651 12587 47657
rect 12529 47617 12541 47651
rect 12575 47648 12587 47651
rect 12618 47648 12624 47660
rect 12575 47620 12624 47648
rect 12575 47617 12587 47620
rect 12529 47611 12587 47617
rect 12618 47608 12624 47620
rect 12676 47608 12682 47660
rect 13280 47592 13308 47688
rect 23109 47685 23121 47719
rect 23155 47716 23167 47719
rect 23934 47716 23940 47728
rect 23155 47688 23940 47716
rect 23155 47685 23167 47688
rect 23109 47679 23167 47685
rect 23934 47676 23940 47688
rect 23992 47716 23998 47728
rect 27525 47719 27583 47725
rect 23992 47688 24716 47716
rect 23992 47676 23998 47688
rect 14369 47651 14427 47657
rect 14369 47617 14381 47651
rect 14415 47648 14427 47651
rect 15102 47648 15108 47660
rect 14415 47620 15108 47648
rect 14415 47617 14427 47620
rect 14369 47611 14427 47617
rect 15102 47608 15108 47620
rect 15160 47608 15166 47660
rect 21177 47651 21235 47657
rect 21177 47617 21189 47651
rect 21223 47648 21235 47651
rect 22002 47648 22008 47660
rect 21223 47620 22008 47648
rect 21223 47617 21235 47620
rect 21177 47611 21235 47617
rect 22002 47608 22008 47620
rect 22060 47608 22066 47660
rect 22741 47651 22799 47657
rect 22741 47617 22753 47651
rect 22787 47648 22799 47651
rect 23658 47648 23664 47660
rect 22787 47620 23664 47648
rect 22787 47617 22799 47620
rect 22741 47611 22799 47617
rect 23658 47608 23664 47620
rect 23716 47608 23722 47660
rect 24688 47592 24716 47688
rect 27525 47685 27537 47719
rect 27571 47685 27583 47719
rect 27525 47679 27583 47685
rect 24946 47608 24952 47660
rect 25004 47648 25010 47660
rect 25409 47651 25467 47657
rect 25409 47648 25421 47651
rect 25004 47620 25421 47648
rect 25004 47608 25010 47620
rect 25409 47617 25421 47620
rect 25455 47648 25467 47651
rect 25501 47651 25559 47657
rect 25501 47648 25513 47651
rect 25455 47620 25513 47648
rect 25455 47617 25467 47620
rect 25409 47611 25467 47617
rect 25501 47617 25513 47620
rect 25547 47648 25559 47651
rect 26326 47648 26332 47660
rect 25547 47620 26332 47648
rect 25547 47617 25559 47620
rect 25501 47611 25559 47617
rect 26326 47608 26332 47620
rect 26384 47608 26390 47660
rect 27540 47648 27568 47679
rect 29270 47676 29276 47728
rect 29328 47716 29334 47728
rect 32398 47716 32404 47728
rect 29328 47688 29960 47716
rect 32359 47688 32404 47716
rect 29328 47676 29334 47688
rect 29932 47660 29960 47688
rect 32398 47676 32404 47688
rect 32456 47676 32462 47728
rect 27540 47620 29776 47648
rect 12986 47580 12992 47592
rect 12947 47552 12992 47580
rect 12986 47540 12992 47552
rect 13044 47540 13050 47592
rect 13262 47540 13268 47592
rect 13320 47580 13326 47592
rect 13357 47583 13415 47589
rect 13357 47580 13369 47583
rect 13320 47552 13369 47580
rect 13320 47540 13326 47552
rect 13357 47549 13369 47552
rect 13403 47549 13415 47583
rect 13357 47543 13415 47549
rect 13446 47540 13452 47592
rect 13504 47580 13510 47592
rect 14642 47580 14648 47592
rect 13504 47552 13549 47580
rect 14603 47552 14648 47580
rect 13504 47540 13510 47552
rect 14642 47540 14648 47552
rect 14700 47540 14706 47592
rect 15286 47540 15292 47592
rect 15344 47580 15350 47592
rect 16114 47580 16120 47592
rect 15344 47552 16120 47580
rect 15344 47540 15350 47552
rect 16114 47540 16120 47552
rect 16172 47580 16178 47592
rect 16301 47583 16359 47589
rect 16301 47580 16313 47583
rect 16172 47552 16313 47580
rect 16172 47540 16178 47552
rect 16301 47549 16313 47552
rect 16347 47549 16359 47583
rect 16850 47580 16856 47592
rect 16811 47552 16856 47580
rect 16301 47543 16359 47549
rect 13909 47447 13967 47453
rect 13909 47413 13921 47447
rect 13955 47444 13967 47447
rect 13998 47444 14004 47456
rect 13955 47416 14004 47444
rect 13955 47413 13967 47416
rect 13909 47407 13967 47413
rect 13998 47404 14004 47416
rect 14056 47404 14062 47456
rect 15746 47444 15752 47456
rect 15707 47416 15752 47444
rect 15746 47404 15752 47416
rect 15804 47404 15810 47456
rect 16316 47444 16344 47543
rect 16850 47540 16856 47552
rect 16908 47580 16914 47592
rect 17313 47583 17371 47589
rect 17313 47580 17325 47583
rect 16908 47552 17325 47580
rect 16908 47540 16914 47552
rect 17313 47549 17325 47552
rect 17359 47549 17371 47583
rect 17313 47543 17371 47549
rect 19429 47583 19487 47589
rect 19429 47549 19441 47583
rect 19475 47580 19487 47583
rect 20349 47583 20407 47589
rect 19475 47552 20024 47580
rect 19475 47549 19487 47552
rect 19429 47543 19487 47549
rect 19996 47453 20024 47552
rect 20349 47549 20361 47583
rect 20395 47580 20407 47583
rect 21082 47580 21088 47592
rect 20395 47552 21088 47580
rect 20395 47549 20407 47552
rect 20349 47543 20407 47549
rect 21082 47540 21088 47552
rect 21140 47540 21146 47592
rect 21634 47540 21640 47592
rect 21692 47580 21698 47592
rect 21913 47583 21971 47589
rect 21913 47580 21925 47583
rect 21692 47552 21925 47580
rect 21692 47540 21698 47552
rect 21913 47549 21925 47552
rect 21959 47580 21971 47583
rect 22649 47583 22707 47589
rect 22649 47580 22661 47583
rect 21959 47552 22661 47580
rect 21959 47549 21971 47552
rect 21913 47543 21971 47549
rect 22649 47549 22661 47552
rect 22695 47580 22707 47583
rect 23382 47580 23388 47592
rect 22695 47552 23388 47580
rect 22695 47549 22707 47552
rect 22649 47543 22707 47549
rect 23382 47540 23388 47552
rect 23440 47540 23446 47592
rect 24026 47540 24032 47592
rect 24084 47580 24090 47592
rect 24213 47583 24271 47589
rect 24213 47580 24225 47583
rect 24084 47552 24225 47580
rect 24084 47540 24090 47552
rect 24213 47549 24225 47552
rect 24259 47549 24271 47583
rect 24486 47580 24492 47592
rect 24447 47552 24492 47580
rect 24213 47543 24271 47549
rect 24486 47540 24492 47552
rect 24544 47540 24550 47592
rect 24670 47580 24676 47592
rect 24631 47552 24676 47580
rect 24670 47540 24676 47552
rect 24728 47540 24734 47592
rect 25590 47540 25596 47592
rect 25648 47580 25654 47592
rect 25685 47583 25743 47589
rect 25685 47580 25697 47583
rect 25648 47552 25697 47580
rect 25648 47540 25654 47552
rect 25685 47549 25697 47552
rect 25731 47549 25743 47583
rect 27706 47580 27712 47592
rect 27667 47552 27712 47580
rect 25685 47543 25743 47549
rect 27706 47540 27712 47552
rect 27764 47540 27770 47592
rect 27798 47540 27804 47592
rect 27856 47580 27862 47592
rect 27893 47583 27951 47589
rect 27893 47580 27905 47583
rect 27856 47552 27905 47580
rect 27856 47540 27862 47552
rect 27893 47549 27905 47552
rect 27939 47580 27951 47583
rect 27982 47580 27988 47592
rect 27939 47552 27988 47580
rect 27939 47549 27951 47552
rect 27893 47543 27951 47549
rect 27982 47540 27988 47552
rect 28040 47540 28046 47592
rect 28077 47583 28135 47589
rect 28077 47549 28089 47583
rect 28123 47549 28135 47583
rect 28077 47543 28135 47549
rect 23566 47472 23572 47524
rect 23624 47512 23630 47524
rect 23661 47515 23719 47521
rect 23661 47512 23673 47515
rect 23624 47484 23673 47512
rect 23624 47472 23630 47484
rect 23661 47481 23673 47484
rect 23707 47481 23719 47515
rect 24504 47512 24532 47540
rect 24949 47515 25007 47521
rect 24949 47512 24961 47515
rect 24504 47484 24961 47512
rect 23661 47475 23719 47481
rect 24949 47481 24961 47484
rect 24995 47481 25007 47515
rect 24949 47475 25007 47481
rect 25314 47472 25320 47524
rect 25372 47512 25378 47524
rect 25869 47515 25927 47521
rect 25869 47512 25881 47515
rect 25372 47484 25881 47512
rect 25372 47472 25378 47484
rect 25869 47481 25881 47484
rect 25915 47481 25927 47515
rect 25869 47475 25927 47481
rect 25958 47472 25964 47524
rect 26016 47512 26022 47524
rect 26237 47515 26295 47521
rect 26237 47512 26249 47515
rect 26016 47484 26249 47512
rect 26016 47472 26022 47484
rect 26237 47481 26249 47484
rect 26283 47481 26295 47515
rect 26237 47475 26295 47481
rect 27522 47472 27528 47524
rect 27580 47512 27586 47524
rect 28092 47512 28120 47543
rect 29086 47540 29092 47592
rect 29144 47580 29150 47592
rect 29748 47589 29776 47620
rect 29914 47608 29920 47660
rect 29972 47648 29978 47660
rect 29972 47620 32260 47648
rect 29972 47608 29978 47620
rect 29273 47583 29331 47589
rect 29273 47580 29285 47583
rect 29144 47552 29285 47580
rect 29144 47540 29150 47552
rect 29273 47549 29285 47552
rect 29319 47549 29331 47583
rect 29273 47543 29331 47549
rect 29733 47583 29791 47589
rect 29733 47549 29745 47583
rect 29779 47580 29791 47583
rect 29822 47580 29828 47592
rect 29779 47552 29828 47580
rect 29779 47549 29791 47552
rect 29733 47543 29791 47549
rect 29822 47540 29828 47552
rect 29880 47540 29886 47592
rect 30834 47580 30840 47592
rect 30795 47552 30840 47580
rect 30834 47540 30840 47552
rect 30892 47540 30898 47592
rect 30926 47540 30932 47592
rect 30984 47580 30990 47592
rect 32232 47589 32260 47620
rect 31665 47583 31723 47589
rect 31665 47580 31677 47583
rect 30984 47552 31677 47580
rect 30984 47540 30990 47552
rect 31665 47549 31677 47552
rect 31711 47549 31723 47583
rect 31665 47543 31723 47549
rect 32217 47583 32275 47589
rect 32217 47549 32229 47583
rect 32263 47580 32275 47583
rect 32677 47583 32735 47589
rect 32677 47580 32689 47583
rect 32263 47552 32689 47580
rect 32263 47549 32275 47552
rect 32217 47543 32275 47549
rect 32677 47549 32689 47552
rect 32723 47549 32735 47583
rect 32677 47543 32735 47549
rect 30374 47512 30380 47524
rect 27580 47484 28120 47512
rect 30287 47484 30380 47512
rect 27580 47472 27586 47484
rect 30374 47472 30380 47484
rect 30432 47512 30438 47524
rect 31018 47512 31024 47524
rect 30432 47484 31024 47512
rect 30432 47472 30438 47484
rect 31018 47472 31024 47484
rect 31076 47472 31082 47524
rect 17037 47447 17095 47453
rect 17037 47444 17049 47447
rect 16316 47416 17049 47444
rect 17037 47413 17049 47416
rect 17083 47413 17095 47447
rect 17037 47407 17095 47413
rect 19981 47447 20039 47453
rect 19981 47413 19993 47447
rect 20027 47444 20039 47447
rect 20070 47444 20076 47456
rect 20027 47416 20076 47444
rect 20027 47413 20039 47416
rect 19981 47407 20039 47413
rect 20070 47404 20076 47416
rect 20128 47404 20134 47456
rect 25590 47404 25596 47456
rect 25648 47444 25654 47456
rect 25777 47447 25835 47453
rect 25777 47444 25789 47447
rect 25648 47416 25789 47444
rect 25648 47404 25654 47416
rect 25777 47413 25789 47416
rect 25823 47413 25835 47447
rect 25777 47407 25835 47413
rect 26605 47447 26663 47453
rect 26605 47413 26617 47447
rect 26651 47444 26663 47447
rect 26786 47444 26792 47456
rect 26651 47416 26792 47444
rect 26651 47413 26663 47416
rect 26605 47407 26663 47413
rect 26786 47404 26792 47416
rect 26844 47404 26850 47456
rect 28534 47444 28540 47456
rect 28495 47416 28540 47444
rect 28534 47404 28540 47416
rect 28592 47404 28598 47456
rect 29362 47444 29368 47456
rect 29323 47416 29368 47444
rect 29362 47404 29368 47416
rect 29420 47404 29426 47456
rect 30650 47444 30656 47456
rect 30611 47416 30656 47444
rect 30650 47404 30656 47416
rect 30708 47404 30714 47456
rect 1104 47354 38824 47376
rect 1104 47302 19606 47354
rect 19658 47302 19670 47354
rect 19722 47302 19734 47354
rect 19786 47302 19798 47354
rect 19850 47302 38824 47354
rect 1104 47280 38824 47302
rect 12250 47200 12256 47252
rect 12308 47240 12314 47252
rect 12713 47243 12771 47249
rect 12713 47240 12725 47243
rect 12308 47212 12725 47240
rect 12308 47200 12314 47212
rect 12713 47209 12725 47212
rect 12759 47209 12771 47243
rect 12713 47203 12771 47209
rect 13446 47200 13452 47252
rect 13504 47240 13510 47252
rect 13633 47243 13691 47249
rect 13633 47240 13645 47243
rect 13504 47212 13645 47240
rect 13504 47200 13510 47212
rect 13633 47209 13645 47212
rect 13679 47209 13691 47243
rect 13633 47203 13691 47209
rect 19426 47200 19432 47252
rect 19484 47240 19490 47252
rect 19981 47243 20039 47249
rect 19981 47240 19993 47243
rect 19484 47212 19993 47240
rect 19484 47200 19490 47212
rect 19981 47209 19993 47212
rect 20027 47209 20039 47243
rect 21174 47240 21180 47252
rect 21135 47212 21180 47240
rect 19981 47203 20039 47209
rect 21174 47200 21180 47212
rect 21232 47200 21238 47252
rect 21450 47240 21456 47252
rect 21411 47212 21456 47240
rect 21450 47200 21456 47212
rect 21508 47200 21514 47252
rect 22465 47243 22523 47249
rect 22465 47209 22477 47243
rect 22511 47240 22523 47243
rect 22554 47240 22560 47252
rect 22511 47212 22560 47240
rect 22511 47209 22523 47212
rect 22465 47203 22523 47209
rect 22554 47200 22560 47212
rect 22612 47200 22618 47252
rect 23109 47243 23167 47249
rect 23109 47209 23121 47243
rect 23155 47240 23167 47243
rect 23750 47240 23756 47252
rect 23155 47212 23756 47240
rect 23155 47209 23167 47212
rect 23109 47203 23167 47209
rect 23750 47200 23756 47212
rect 23808 47200 23814 47252
rect 24118 47200 24124 47252
rect 24176 47240 24182 47252
rect 24581 47243 24639 47249
rect 24581 47240 24593 47243
rect 24176 47212 24593 47240
rect 24176 47200 24182 47212
rect 24581 47209 24593 47212
rect 24627 47209 24639 47243
rect 25406 47240 25412 47252
rect 25367 47212 25412 47240
rect 24581 47203 24639 47209
rect 25406 47200 25412 47212
rect 25464 47200 25470 47252
rect 25774 47240 25780 47252
rect 25735 47212 25780 47240
rect 25774 47200 25780 47212
rect 25832 47200 25838 47252
rect 26237 47243 26295 47249
rect 26237 47209 26249 47243
rect 26283 47240 26295 47243
rect 27062 47240 27068 47252
rect 26283 47212 27068 47240
rect 26283 47209 26295 47212
rect 26237 47203 26295 47209
rect 27062 47200 27068 47212
rect 27120 47200 27126 47252
rect 28442 47240 28448 47252
rect 28403 47212 28448 47240
rect 28442 47200 28448 47212
rect 28500 47200 28506 47252
rect 29822 47240 29828 47252
rect 29783 47212 29828 47240
rect 29822 47200 29828 47212
rect 29880 47200 29886 47252
rect 30190 47240 30196 47252
rect 30151 47212 30196 47240
rect 30190 47200 30196 47212
rect 30248 47240 30254 47252
rect 30653 47243 30711 47249
rect 30653 47240 30665 47243
rect 30248 47212 30665 47240
rect 30248 47200 30254 47212
rect 30653 47209 30665 47212
rect 30699 47209 30711 47243
rect 31386 47240 31392 47252
rect 31347 47212 31392 47240
rect 30653 47203 30711 47209
rect 31386 47200 31392 47212
rect 31444 47240 31450 47252
rect 31757 47243 31815 47249
rect 31757 47240 31769 47243
rect 31444 47212 31769 47240
rect 31444 47200 31450 47212
rect 31757 47209 31769 47212
rect 31803 47209 31815 47243
rect 31757 47203 31815 47209
rect 12986 47132 12992 47184
rect 13044 47172 13050 47184
rect 13357 47175 13415 47181
rect 13357 47172 13369 47175
rect 13044 47144 13369 47172
rect 13044 47132 13050 47144
rect 13357 47141 13369 47144
rect 13403 47172 13415 47175
rect 14369 47175 14427 47181
rect 14369 47172 14381 47175
rect 13403 47144 14381 47172
rect 13403 47141 13415 47144
rect 13357 47135 13415 47141
rect 14369 47141 14381 47144
rect 14415 47141 14427 47175
rect 15838 47172 15844 47184
rect 15799 47144 15844 47172
rect 14369 47135 14427 47141
rect 15838 47132 15844 47144
rect 15896 47172 15902 47184
rect 16117 47175 16175 47181
rect 16117 47172 16129 47175
rect 15896 47144 16129 47172
rect 15896 47132 15902 47144
rect 16117 47141 16129 47144
rect 16163 47141 16175 47175
rect 23014 47172 23020 47184
rect 16117 47135 16175 47141
rect 20732 47144 23020 47172
rect 11422 47064 11428 47116
rect 11480 47104 11486 47116
rect 11609 47107 11667 47113
rect 11609 47104 11621 47107
rect 11480 47076 11621 47104
rect 11480 47064 11486 47076
rect 11609 47073 11621 47076
rect 11655 47073 11667 47107
rect 13906 47104 13912 47116
rect 13867 47076 13912 47104
rect 11609 47067 11667 47073
rect 13906 47064 13912 47076
rect 13964 47064 13970 47116
rect 15381 47107 15439 47113
rect 15381 47073 15393 47107
rect 15427 47104 15439 47107
rect 15746 47104 15752 47116
rect 15427 47076 15752 47104
rect 15427 47073 15439 47076
rect 15381 47067 15439 47073
rect 15746 47064 15752 47076
rect 15804 47064 15810 47116
rect 16669 47107 16727 47113
rect 16669 47073 16681 47107
rect 16715 47104 16727 47107
rect 17310 47104 17316 47116
rect 16715 47076 17316 47104
rect 16715 47073 16727 47076
rect 16669 47067 16727 47073
rect 17310 47064 17316 47076
rect 17368 47064 17374 47116
rect 19797 47107 19855 47113
rect 19797 47073 19809 47107
rect 19843 47104 19855 47107
rect 19886 47104 19892 47116
rect 19843 47076 19892 47104
rect 19843 47073 19855 47076
rect 19797 47067 19855 47073
rect 19886 47064 19892 47076
rect 19944 47064 19950 47116
rect 11333 47039 11391 47045
rect 11333 47005 11345 47039
rect 11379 47036 11391 47039
rect 11698 47036 11704 47048
rect 11379 47008 11704 47036
rect 11379 47005 11391 47008
rect 11333 46999 11391 47005
rect 11698 46996 11704 47008
rect 11756 46996 11762 47048
rect 13817 47039 13875 47045
rect 13817 47005 13829 47039
rect 13863 47036 13875 47039
rect 13998 47036 14004 47048
rect 13863 47008 14004 47036
rect 13863 47005 13875 47008
rect 13817 46999 13875 47005
rect 13998 46996 14004 47008
rect 14056 47036 14062 47048
rect 15289 47039 15347 47045
rect 15289 47036 15301 47039
rect 14056 47008 15301 47036
rect 14056 46996 14062 47008
rect 15289 47005 15301 47008
rect 15335 47005 15347 47039
rect 16942 47036 16948 47048
rect 16903 47008 16948 47036
rect 15289 46999 15347 47005
rect 16942 46996 16948 47008
rect 17000 46996 17006 47048
rect 20732 47045 20760 47144
rect 23014 47132 23020 47144
rect 23072 47172 23078 47184
rect 23569 47175 23627 47181
rect 23569 47172 23581 47175
rect 23072 47144 23581 47172
rect 23072 47132 23078 47144
rect 23569 47141 23581 47144
rect 23615 47172 23627 47175
rect 23842 47172 23848 47184
rect 23615 47144 23848 47172
rect 23615 47141 23627 47144
rect 23569 47135 23627 47141
rect 23842 47132 23848 47144
rect 23900 47132 23906 47184
rect 24210 47132 24216 47184
rect 24268 47172 24274 47184
rect 24305 47175 24363 47181
rect 24305 47172 24317 47175
rect 24268 47144 24317 47172
rect 24268 47132 24274 47144
rect 24305 47141 24317 47144
rect 24351 47141 24363 47175
rect 24305 47135 24363 47141
rect 25041 47175 25099 47181
rect 25041 47141 25053 47175
rect 25087 47172 25099 47175
rect 25590 47172 25596 47184
rect 25087 47144 25596 47172
rect 25087 47141 25099 47144
rect 25041 47135 25099 47141
rect 20993 47107 21051 47113
rect 20993 47073 21005 47107
rect 21039 47104 21051 47107
rect 22005 47107 22063 47113
rect 21039 47076 21956 47104
rect 21039 47073 21051 47076
rect 20993 47067 21051 47073
rect 18325 47039 18383 47045
rect 18325 47005 18337 47039
rect 18371 47036 18383 47039
rect 20717 47039 20775 47045
rect 20717 47036 20729 47039
rect 18371 47008 20729 47036
rect 18371 47005 18383 47008
rect 18325 46999 18383 47005
rect 20717 47005 20729 47008
rect 20763 47005 20775 47039
rect 20717 46999 20775 47005
rect 21928 46980 21956 47076
rect 22005 47073 22017 47107
rect 22051 47073 22063 47107
rect 22005 47067 22063 47073
rect 20346 46968 20352 46980
rect 20307 46940 20352 46968
rect 20346 46928 20352 46940
rect 20404 46928 20410 46980
rect 21910 46968 21916 46980
rect 21871 46940 21916 46968
rect 21910 46928 21916 46940
rect 21968 46928 21974 46980
rect 1394 46860 1400 46912
rect 1452 46900 1458 46912
rect 1581 46903 1639 46909
rect 1581 46900 1593 46903
rect 1452 46872 1593 46900
rect 1452 46860 1458 46872
rect 1581 46869 1593 46872
rect 1627 46869 1639 46903
rect 14918 46900 14924 46912
rect 14879 46872 14924 46900
rect 1581 46863 1639 46869
rect 14918 46860 14924 46872
rect 14976 46860 14982 46912
rect 22020 46900 22048 47067
rect 22094 47064 22100 47116
rect 22152 47104 22158 47116
rect 22281 47107 22339 47113
rect 22281 47104 22293 47107
rect 22152 47076 22293 47104
rect 22152 47064 22158 47076
rect 22281 47073 22293 47076
rect 22327 47104 22339 47107
rect 23477 47107 23535 47113
rect 22327 47076 22876 47104
rect 22327 47073 22339 47076
rect 22281 47067 22339 47073
rect 22848 47036 22876 47076
rect 23477 47073 23489 47107
rect 23523 47104 23535 47107
rect 23523 47076 24348 47104
rect 23523 47073 23535 47076
rect 23477 47067 23535 47073
rect 24320 47048 24348 47076
rect 23658 47036 23664 47048
rect 22848 47008 23664 47036
rect 23658 46996 23664 47008
rect 23716 47036 23722 47048
rect 23937 47039 23995 47045
rect 23937 47036 23949 47039
rect 23716 47008 23949 47036
rect 23716 46996 23722 47008
rect 23937 47005 23949 47008
rect 23983 47005 23995 47039
rect 23937 46999 23995 47005
rect 24302 46996 24308 47048
rect 24360 46996 24366 47048
rect 22097 46971 22155 46977
rect 22097 46937 22109 46971
rect 22143 46968 22155 46971
rect 22186 46968 22192 46980
rect 22143 46940 22192 46968
rect 22143 46937 22155 46940
rect 22097 46931 22155 46937
rect 22186 46928 22192 46940
rect 22244 46928 22250 46980
rect 23566 46928 23572 46980
rect 23624 46968 23630 46980
rect 25056 46968 25084 47135
rect 25590 47132 25596 47144
rect 25648 47172 25654 47184
rect 25792 47172 25820 47200
rect 25648 47144 25820 47172
rect 26513 47175 26571 47181
rect 25648 47132 25654 47144
rect 26513 47141 26525 47175
rect 26559 47172 26571 47175
rect 26878 47172 26884 47184
rect 26559 47144 26884 47172
rect 26559 47141 26571 47144
rect 26513 47135 26571 47141
rect 26878 47132 26884 47144
rect 26936 47172 26942 47184
rect 28534 47172 28540 47184
rect 26936 47144 28540 47172
rect 26936 47132 26942 47144
rect 28534 47132 28540 47144
rect 28592 47132 28598 47184
rect 30742 47172 30748 47184
rect 30703 47144 30748 47172
rect 30742 47132 30748 47144
rect 30800 47172 30806 47184
rect 31846 47172 31852 47184
rect 30800 47144 31852 47172
rect 30800 47132 30806 47144
rect 31846 47132 31852 47144
rect 31904 47132 31910 47184
rect 25222 47104 25228 47116
rect 25183 47076 25228 47104
rect 25222 47064 25228 47076
rect 25280 47064 25286 47116
rect 27154 47104 27160 47116
rect 27115 47076 27160 47104
rect 27154 47064 27160 47076
rect 27212 47064 27218 47116
rect 27522 47104 27528 47116
rect 27483 47076 27528 47104
rect 27522 47064 27528 47076
rect 27580 47064 27586 47116
rect 28994 47104 29000 47116
rect 28955 47076 29000 47104
rect 28994 47064 29000 47076
rect 29052 47064 29058 47116
rect 29270 47064 29276 47116
rect 29328 47104 29334 47116
rect 29365 47107 29423 47113
rect 29365 47104 29377 47107
rect 29328 47076 29377 47104
rect 29328 47064 29334 47076
rect 29365 47073 29377 47076
rect 29411 47073 29423 47107
rect 29365 47067 29423 47073
rect 29457 47107 29515 47113
rect 29457 47073 29469 47107
rect 29503 47104 29515 47107
rect 29914 47104 29920 47116
rect 29503 47076 29920 47104
rect 29503 47073 29515 47076
rect 29457 47067 29515 47073
rect 26878 46996 26884 47048
rect 26936 47036 26942 47048
rect 27065 47039 27123 47045
rect 27065 47036 27077 47039
rect 26936 47008 27077 47036
rect 26936 46996 26942 47008
rect 27065 47005 27077 47008
rect 27111 47005 27123 47039
rect 27065 46999 27123 47005
rect 27430 46996 27436 47048
rect 27488 47036 27494 47048
rect 27617 47039 27675 47045
rect 27617 47036 27629 47039
rect 27488 47008 27629 47036
rect 27488 46996 27494 47008
rect 27617 47005 27629 47008
rect 27663 47005 27675 47039
rect 27617 46999 27675 47005
rect 27706 46996 27712 47048
rect 27764 47036 27770 47048
rect 28077 47039 28135 47045
rect 28077 47036 28089 47039
rect 27764 47008 28089 47036
rect 27764 46996 27770 47008
rect 28077 47005 28089 47008
rect 28123 47036 28135 47039
rect 28902 47036 28908 47048
rect 28123 47008 28908 47036
rect 28123 47005 28135 47008
rect 28077 46999 28135 47005
rect 28902 46996 28908 47008
rect 28960 46996 28966 47048
rect 29086 46996 29092 47048
rect 29144 47036 29150 47048
rect 29472 47036 29500 47067
rect 29914 47064 29920 47076
rect 29972 47064 29978 47116
rect 30558 47104 30564 47116
rect 30519 47076 30564 47104
rect 30558 47064 30564 47076
rect 30616 47064 30622 47116
rect 31018 47064 31024 47116
rect 31076 47104 31082 47116
rect 32122 47104 32128 47116
rect 31076 47076 32128 47104
rect 31076 47064 31082 47076
rect 32122 47064 32128 47076
rect 32180 47064 32186 47116
rect 30374 47036 30380 47048
rect 29144 47008 29500 47036
rect 30335 47008 30380 47036
rect 29144 46996 29150 47008
rect 30374 46996 30380 47008
rect 30432 46996 30438 47048
rect 31110 47036 31116 47048
rect 31071 47008 31116 47036
rect 31110 46996 31116 47008
rect 31168 46996 31174 47048
rect 28810 46968 28816 46980
rect 23624 46940 25084 46968
rect 28771 46940 28816 46968
rect 23624 46928 23630 46940
rect 22278 46900 22284 46912
rect 22020 46872 22284 46900
rect 22278 46860 22284 46872
rect 22336 46900 22342 46912
rect 22738 46900 22744 46912
rect 22336 46872 22744 46900
rect 22336 46860 22342 46872
rect 22738 46860 22744 46872
rect 22796 46860 22802 46912
rect 23676 46900 23704 46940
rect 28810 46928 28816 46940
rect 28868 46928 28874 46980
rect 23734 46903 23792 46909
rect 23734 46900 23746 46903
rect 23676 46872 23746 46900
rect 23734 46869 23746 46872
rect 23780 46869 23792 46903
rect 23734 46863 23792 46869
rect 23845 46903 23903 46909
rect 23845 46869 23857 46903
rect 23891 46900 23903 46903
rect 24026 46900 24032 46912
rect 23891 46872 24032 46900
rect 23891 46869 23903 46872
rect 23845 46863 23903 46869
rect 24026 46860 24032 46872
rect 24084 46860 24090 46912
rect 29638 46860 29644 46912
rect 29696 46900 29702 46912
rect 32309 46903 32367 46909
rect 32309 46900 32321 46903
rect 29696 46872 32321 46900
rect 29696 46860 29702 46872
rect 32309 46869 32321 46872
rect 32355 46869 32367 46903
rect 32309 46863 32367 46869
rect 1104 46810 38824 46832
rect 1104 46758 4246 46810
rect 4298 46758 4310 46810
rect 4362 46758 4374 46810
rect 4426 46758 4438 46810
rect 4490 46758 34966 46810
rect 35018 46758 35030 46810
rect 35082 46758 35094 46810
rect 35146 46758 35158 46810
rect 35210 46758 38824 46810
rect 1104 46736 38824 46758
rect 11698 46696 11704 46708
rect 11659 46668 11704 46696
rect 11698 46656 11704 46668
rect 11756 46656 11762 46708
rect 13817 46699 13875 46705
rect 13817 46665 13829 46699
rect 13863 46696 13875 46699
rect 13906 46696 13912 46708
rect 13863 46668 13912 46696
rect 13863 46665 13875 46668
rect 13817 46659 13875 46665
rect 13906 46656 13912 46668
rect 13964 46656 13970 46708
rect 19886 46696 19892 46708
rect 19847 46668 19892 46696
rect 19886 46656 19892 46668
rect 19944 46656 19950 46708
rect 20898 46656 20904 46708
rect 20956 46696 20962 46708
rect 21177 46699 21235 46705
rect 21177 46696 21189 46699
rect 20956 46668 21189 46696
rect 20956 46656 20962 46668
rect 21177 46665 21189 46668
rect 21223 46665 21235 46699
rect 21177 46659 21235 46665
rect 21545 46699 21603 46705
rect 21545 46665 21557 46699
rect 21591 46696 21603 46699
rect 22002 46696 22008 46708
rect 21591 46668 22008 46696
rect 21591 46665 21603 46668
rect 21545 46659 21603 46665
rect 22002 46656 22008 46668
rect 22060 46656 22066 46708
rect 25222 46696 25228 46708
rect 25183 46668 25228 46696
rect 25222 46656 25228 46668
rect 25280 46656 25286 46708
rect 27154 46656 27160 46708
rect 27212 46696 27218 46708
rect 27433 46699 27491 46705
rect 27433 46696 27445 46699
rect 27212 46668 27445 46696
rect 27212 46656 27218 46668
rect 27433 46665 27445 46668
rect 27479 46665 27491 46699
rect 29086 46696 29092 46708
rect 29047 46668 29092 46696
rect 27433 46659 27491 46665
rect 29086 46656 29092 46668
rect 29144 46656 29150 46708
rect 29546 46656 29552 46708
rect 29604 46696 29610 46708
rect 29641 46699 29699 46705
rect 29641 46696 29653 46699
rect 29604 46668 29653 46696
rect 29604 46656 29610 46668
rect 29641 46665 29653 46668
rect 29687 46665 29699 46699
rect 32122 46696 32128 46708
rect 32083 46668 32128 46696
rect 29641 46659 29699 46665
rect 21913 46631 21971 46637
rect 21913 46597 21925 46631
rect 21959 46628 21971 46631
rect 22186 46628 22192 46640
rect 21959 46600 22192 46628
rect 21959 46597 21971 46600
rect 21913 46591 21971 46597
rect 22186 46588 22192 46600
rect 22244 46628 22250 46640
rect 22244 46600 22600 46628
rect 22244 46588 22250 46600
rect 1670 46560 1676 46572
rect 1631 46532 1676 46560
rect 1670 46520 1676 46532
rect 1728 46520 1734 46572
rect 12710 46560 12716 46572
rect 12623 46532 12716 46560
rect 12710 46520 12716 46532
rect 12768 46560 12774 46572
rect 13446 46560 13452 46572
rect 12768 46532 13452 46560
rect 12768 46520 12774 46532
rect 13446 46520 13452 46532
rect 13504 46520 13510 46572
rect 14550 46520 14556 46572
rect 14608 46560 14614 46572
rect 14921 46563 14979 46569
rect 14921 46560 14933 46563
rect 14608 46532 14933 46560
rect 14608 46520 14614 46532
rect 14921 46529 14933 46532
rect 14967 46529 14979 46563
rect 14921 46523 14979 46529
rect 20901 46563 20959 46569
rect 20901 46529 20913 46563
rect 20947 46560 20959 46563
rect 22462 46560 22468 46572
rect 20947 46532 21956 46560
rect 22423 46532 22468 46560
rect 20947 46529 20959 46532
rect 20901 46523 20959 46529
rect 21928 46504 21956 46532
rect 22462 46520 22468 46532
rect 22520 46520 22526 46572
rect 22572 46560 22600 46600
rect 28166 46588 28172 46640
rect 28224 46628 28230 46640
rect 28626 46628 28632 46640
rect 28224 46600 28632 46628
rect 28224 46588 28230 46600
rect 28626 46588 28632 46600
rect 28684 46588 28690 46640
rect 24670 46560 24676 46572
rect 22572 46532 23152 46560
rect 24631 46532 24676 46560
rect 1394 46492 1400 46504
rect 1355 46464 1400 46492
rect 1394 46452 1400 46464
rect 1452 46452 1458 46504
rect 11698 46452 11704 46504
rect 11756 46492 11762 46504
rect 12434 46492 12440 46504
rect 11756 46464 12440 46492
rect 11756 46452 11762 46464
rect 12434 46452 12440 46464
rect 12492 46492 12498 46504
rect 12492 46464 12537 46492
rect 12492 46452 12498 46464
rect 15010 46452 15016 46504
rect 15068 46492 15074 46504
rect 15381 46495 15439 46501
rect 15381 46492 15393 46495
rect 15068 46464 15393 46492
rect 15068 46452 15074 46464
rect 15381 46461 15393 46464
rect 15427 46461 15439 46495
rect 15562 46492 15568 46504
rect 15523 46464 15568 46492
rect 15381 46455 15439 46461
rect 15562 46452 15568 46464
rect 15620 46452 15626 46504
rect 15654 46452 15660 46504
rect 15712 46492 15718 46504
rect 15749 46495 15807 46501
rect 15749 46492 15761 46495
rect 15712 46464 15761 46492
rect 15712 46452 15718 46464
rect 15749 46461 15761 46464
rect 15795 46461 15807 46495
rect 15749 46455 15807 46461
rect 20533 46495 20591 46501
rect 20533 46461 20545 46495
rect 20579 46492 20591 46495
rect 20990 46492 20996 46504
rect 20579 46464 20996 46492
rect 20579 46461 20591 46464
rect 20533 46455 20591 46461
rect 20990 46452 20996 46464
rect 21048 46452 21054 46504
rect 21910 46452 21916 46504
rect 21968 46492 21974 46504
rect 22005 46495 22063 46501
rect 22005 46492 22017 46495
rect 21968 46464 22017 46492
rect 21968 46452 21974 46464
rect 22005 46461 22017 46464
rect 22051 46461 22063 46495
rect 22005 46455 22063 46461
rect 22094 46452 22100 46504
rect 22152 46492 22158 46504
rect 22281 46495 22339 46501
rect 22152 46464 22197 46492
rect 22152 46452 22158 46464
rect 22281 46461 22293 46495
rect 22327 46492 22339 46495
rect 22922 46492 22928 46504
rect 22327 46464 22928 46492
rect 22327 46461 22339 46464
rect 22281 46455 22339 46461
rect 22922 46452 22928 46464
rect 22980 46452 22986 46504
rect 23124 46501 23152 46532
rect 24670 46520 24676 46532
rect 24728 46520 24734 46572
rect 26145 46563 26203 46569
rect 26145 46529 26157 46563
rect 26191 46560 26203 46563
rect 26510 46560 26516 46572
rect 26191 46532 26516 46560
rect 26191 46529 26203 46532
rect 26145 46523 26203 46529
rect 26510 46520 26516 46532
rect 26568 46520 26574 46572
rect 26697 46563 26755 46569
rect 26697 46529 26709 46563
rect 26743 46560 26755 46563
rect 29656 46560 29684 46659
rect 32122 46656 32128 46668
rect 32180 46656 32186 46708
rect 31846 46588 31852 46640
rect 31904 46628 31910 46640
rect 32493 46631 32551 46637
rect 32493 46628 32505 46631
rect 31904 46600 32505 46628
rect 31904 46588 31910 46600
rect 32493 46597 32505 46600
rect 32539 46597 32551 46631
rect 32493 46591 32551 46597
rect 30101 46563 30159 46569
rect 30101 46560 30113 46563
rect 26743 46532 28764 46560
rect 29656 46532 30113 46560
rect 26743 46529 26755 46532
rect 26697 46523 26755 46529
rect 23109 46495 23167 46501
rect 23109 46461 23121 46495
rect 23155 46492 23167 46495
rect 23477 46495 23535 46501
rect 23477 46492 23489 46495
rect 23155 46464 23489 46492
rect 23155 46461 23167 46464
rect 23109 46455 23167 46461
rect 23477 46461 23489 46464
rect 23523 46492 23535 46495
rect 24026 46492 24032 46504
rect 23523 46464 24032 46492
rect 23523 46461 23535 46464
rect 23477 46455 23535 46461
rect 24026 46452 24032 46464
rect 24084 46492 24090 46504
rect 24581 46495 24639 46501
rect 24581 46492 24593 46495
rect 24084 46464 24593 46492
rect 24084 46452 24090 46464
rect 24581 46461 24593 46464
rect 24627 46492 24639 46495
rect 24854 46492 24860 46504
rect 24627 46464 24860 46492
rect 24627 46461 24639 46464
rect 24581 46455 24639 46461
rect 24854 46452 24860 46464
rect 24912 46452 24918 46504
rect 26053 46495 26111 46501
rect 26053 46461 26065 46495
rect 26099 46492 26111 46495
rect 26602 46492 26608 46504
rect 26099 46464 26608 46492
rect 26099 46461 26111 46464
rect 26053 46455 26111 46461
rect 26602 46452 26608 46464
rect 26660 46492 26666 46504
rect 26712 46492 26740 46523
rect 26660 46464 26740 46492
rect 26973 46495 27031 46501
rect 26660 46452 26666 46464
rect 26973 46461 26985 46495
rect 27019 46492 27031 46495
rect 27062 46492 27068 46504
rect 27019 46464 27068 46492
rect 27019 46461 27031 46464
rect 26973 46455 27031 46461
rect 27062 46452 27068 46464
rect 27120 46452 27126 46504
rect 27157 46495 27215 46501
rect 27157 46461 27169 46495
rect 27203 46461 27215 46495
rect 27157 46455 27215 46461
rect 28077 46495 28135 46501
rect 28077 46461 28089 46495
rect 28123 46492 28135 46495
rect 28166 46492 28172 46504
rect 28123 46464 28172 46492
rect 28123 46461 28135 46464
rect 28077 46455 28135 46461
rect 3050 46424 3056 46436
rect 3011 46396 3056 46424
rect 3050 46384 3056 46396
rect 3108 46384 3114 46436
rect 15580 46424 15608 46452
rect 16209 46427 16267 46433
rect 16209 46424 16221 46427
rect 15580 46396 16221 46424
rect 16209 46393 16221 46396
rect 16255 46393 16267 46427
rect 16209 46387 16267 46393
rect 16761 46427 16819 46433
rect 16761 46393 16773 46427
rect 16807 46424 16819 46427
rect 16942 46424 16948 46436
rect 16807 46396 16948 46424
rect 16807 46393 16819 46396
rect 16761 46387 16819 46393
rect 16942 46384 16948 46396
rect 17000 46424 17006 46436
rect 17494 46424 17500 46436
rect 17000 46396 17500 46424
rect 17000 46384 17006 46396
rect 17494 46384 17500 46396
rect 17552 46384 17558 46436
rect 26418 46384 26424 46436
rect 26476 46424 26482 46436
rect 27172 46424 27200 46455
rect 28166 46452 28172 46464
rect 28224 46452 28230 46504
rect 26476 46396 27200 46424
rect 26476 46384 26482 46396
rect 11422 46356 11428 46368
rect 11383 46328 11428 46356
rect 11422 46316 11428 46328
rect 11480 46316 11486 46368
rect 12253 46359 12311 46365
rect 12253 46325 12265 46359
rect 12299 46356 12311 46359
rect 12342 46356 12348 46368
rect 12299 46328 12348 46356
rect 12299 46325 12311 46328
rect 12253 46319 12311 46325
rect 12342 46316 12348 46328
rect 12400 46356 12406 46368
rect 12710 46356 12716 46368
rect 12400 46328 12716 46356
rect 12400 46316 12406 46328
rect 12710 46316 12716 46328
rect 12768 46316 12774 46368
rect 13998 46316 14004 46368
rect 14056 46356 14062 46368
rect 14369 46359 14427 46365
rect 14369 46356 14381 46359
rect 14056 46328 14381 46356
rect 14056 46316 14062 46328
rect 14369 46325 14381 46328
rect 14415 46356 14427 46359
rect 14737 46359 14795 46365
rect 14737 46356 14749 46359
rect 14415 46328 14749 46356
rect 14415 46325 14427 46328
rect 14369 46319 14427 46325
rect 14737 46325 14749 46328
rect 14783 46325 14795 46359
rect 14737 46319 14795 46325
rect 17129 46359 17187 46365
rect 17129 46325 17141 46359
rect 17175 46356 17187 46359
rect 17310 46356 17316 46368
rect 17175 46328 17316 46356
rect 17175 46325 17187 46328
rect 17129 46319 17187 46325
rect 17310 46316 17316 46328
rect 17368 46316 17374 46368
rect 25685 46359 25743 46365
rect 25685 46325 25697 46359
rect 25731 46356 25743 46359
rect 25774 46356 25780 46368
rect 25731 46328 25780 46356
rect 25731 46325 25743 46328
rect 25685 46319 25743 46325
rect 25774 46316 25780 46328
rect 25832 46316 25838 46368
rect 27798 46316 27804 46368
rect 27856 46356 27862 46368
rect 28074 46356 28080 46368
rect 27856 46328 28080 46356
rect 27856 46316 27862 46328
rect 28074 46316 28080 46328
rect 28132 46356 28138 46368
rect 28736 46365 28764 46532
rect 30101 46529 30113 46532
rect 30147 46529 30159 46563
rect 30101 46523 30159 46529
rect 31938 46520 31944 46572
rect 31996 46560 32002 46572
rect 32861 46563 32919 46569
rect 32861 46560 32873 46563
rect 31996 46532 32873 46560
rect 31996 46520 32002 46532
rect 32861 46529 32873 46532
rect 32907 46529 32919 46563
rect 32861 46523 32919 46529
rect 29546 46452 29552 46504
rect 29604 46492 29610 46504
rect 29825 46495 29883 46501
rect 29825 46492 29837 46495
rect 29604 46464 29837 46492
rect 29604 46452 29610 46464
rect 29825 46461 29837 46464
rect 29871 46492 29883 46495
rect 31956 46492 31984 46520
rect 29871 46464 31984 46492
rect 29871 46461 29883 46464
rect 29825 46455 29883 46461
rect 28353 46359 28411 46365
rect 28353 46356 28365 46359
rect 28132 46328 28365 46356
rect 28132 46316 28138 46328
rect 28353 46325 28365 46328
rect 28399 46325 28411 46359
rect 28353 46319 28411 46325
rect 28721 46359 28779 46365
rect 28721 46325 28733 46359
rect 28767 46356 28779 46359
rect 28902 46356 28908 46368
rect 28767 46328 28908 46356
rect 28767 46325 28779 46328
rect 28721 46319 28779 46325
rect 28902 46316 28908 46328
rect 28960 46316 28966 46368
rect 31202 46356 31208 46368
rect 31163 46328 31208 46356
rect 31202 46316 31208 46328
rect 31260 46316 31266 46368
rect 31754 46316 31760 46368
rect 31812 46356 31818 46368
rect 31812 46328 31857 46356
rect 31812 46316 31818 46328
rect 1104 46266 38824 46288
rect 1104 46214 19606 46266
rect 19658 46214 19670 46266
rect 19722 46214 19734 46266
rect 19786 46214 19798 46266
rect 19850 46214 38824 46266
rect 1104 46192 38824 46214
rect 1670 46152 1676 46164
rect 1631 46124 1676 46152
rect 1670 46112 1676 46124
rect 1728 46112 1734 46164
rect 8846 46152 8852 46164
rect 8807 46124 8852 46152
rect 8846 46112 8852 46124
rect 8904 46152 8910 46164
rect 9674 46152 9680 46164
rect 8904 46124 9680 46152
rect 8904 46112 8910 46124
rect 9674 46112 9680 46124
rect 9732 46112 9738 46164
rect 12434 46112 12440 46164
rect 12492 46152 12498 46164
rect 12529 46155 12587 46161
rect 12529 46152 12541 46155
rect 12492 46124 12541 46152
rect 12492 46112 12498 46124
rect 12529 46121 12541 46124
rect 12575 46152 12587 46155
rect 13354 46152 13360 46164
rect 12575 46124 13360 46152
rect 12575 46121 12587 46124
rect 12529 46115 12587 46121
rect 13354 46112 13360 46124
rect 13412 46112 13418 46164
rect 13725 46155 13783 46161
rect 13725 46121 13737 46155
rect 13771 46152 13783 46155
rect 13906 46152 13912 46164
rect 13771 46124 13912 46152
rect 13771 46121 13783 46124
rect 13725 46115 13783 46121
rect 13906 46112 13912 46124
rect 13964 46112 13970 46164
rect 15565 46155 15623 46161
rect 15565 46121 15577 46155
rect 15611 46152 15623 46155
rect 15746 46152 15752 46164
rect 15611 46124 15752 46152
rect 15611 46121 15623 46124
rect 15565 46115 15623 46121
rect 15746 46112 15752 46124
rect 15804 46112 15810 46164
rect 21361 46155 21419 46161
rect 21361 46121 21373 46155
rect 21407 46152 21419 46155
rect 22094 46152 22100 46164
rect 21407 46124 22100 46152
rect 21407 46121 21419 46124
rect 21361 46115 21419 46121
rect 22094 46112 22100 46124
rect 22152 46152 22158 46164
rect 22370 46152 22376 46164
rect 22152 46124 22376 46152
rect 22152 46112 22158 46124
rect 22370 46112 22376 46124
rect 22428 46112 22434 46164
rect 23658 46152 23664 46164
rect 23619 46124 23664 46152
rect 23658 46112 23664 46124
rect 23716 46112 23722 46164
rect 25777 46155 25835 46161
rect 25777 46121 25789 46155
rect 25823 46152 25835 46155
rect 25958 46152 25964 46164
rect 25823 46124 25964 46152
rect 25823 46121 25835 46124
rect 25777 46115 25835 46121
rect 25958 46112 25964 46124
rect 26016 46112 26022 46164
rect 27157 46155 27215 46161
rect 27157 46121 27169 46155
rect 27203 46152 27215 46155
rect 27246 46152 27252 46164
rect 27203 46124 27252 46152
rect 27203 46121 27215 46124
rect 27157 46115 27215 46121
rect 27246 46112 27252 46124
rect 27304 46112 27310 46164
rect 27430 46112 27436 46164
rect 27488 46112 27494 46164
rect 28353 46155 28411 46161
rect 28353 46121 28365 46155
rect 28399 46152 28411 46155
rect 28626 46152 28632 46164
rect 28399 46124 28488 46152
rect 28587 46124 28632 46152
rect 28399 46121 28411 46124
rect 28353 46115 28411 46121
rect 14369 46087 14427 46093
rect 14369 46053 14381 46087
rect 14415 46084 14427 46087
rect 14918 46084 14924 46096
rect 14415 46056 14924 46084
rect 14415 46053 14427 46056
rect 14369 46047 14427 46053
rect 14918 46044 14924 46056
rect 14976 46044 14982 46096
rect 22922 46084 22928 46096
rect 22756 46056 22928 46084
rect 22756 46028 22784 46056
rect 22922 46044 22928 46056
rect 22980 46044 22986 46096
rect 26789 46087 26847 46093
rect 26789 46053 26801 46087
rect 26835 46084 26847 46087
rect 27448 46084 27476 46112
rect 26835 46056 27476 46084
rect 28460 46084 28488 46124
rect 28626 46112 28632 46124
rect 28684 46112 28690 46164
rect 29089 46155 29147 46161
rect 29089 46121 29101 46155
rect 29135 46152 29147 46155
rect 29270 46152 29276 46164
rect 29135 46124 29276 46152
rect 29135 46121 29147 46124
rect 29089 46115 29147 46121
rect 29270 46112 29276 46124
rect 29328 46152 29334 46164
rect 29454 46152 29460 46164
rect 29328 46124 29460 46152
rect 29328 46112 29334 46124
rect 29454 46112 29460 46124
rect 29512 46152 29518 46164
rect 30374 46152 30380 46164
rect 29512 46124 30380 46152
rect 29512 46112 29518 46124
rect 30374 46112 30380 46124
rect 30432 46112 30438 46164
rect 30558 46112 30564 46164
rect 30616 46152 30622 46164
rect 30926 46152 30932 46164
rect 30616 46124 30932 46152
rect 30616 46112 30622 46124
rect 30926 46112 30932 46124
rect 30984 46152 30990 46164
rect 31205 46155 31263 46161
rect 31205 46152 31217 46155
rect 30984 46124 31217 46152
rect 30984 46112 30990 46124
rect 31205 46121 31217 46124
rect 31251 46152 31263 46155
rect 31754 46152 31760 46164
rect 31251 46124 31760 46152
rect 31251 46121 31263 46124
rect 31205 46115 31263 46121
rect 31754 46112 31760 46124
rect 31812 46112 31818 46164
rect 28534 46084 28540 46096
rect 28460 46056 28540 46084
rect 26835 46053 26847 46056
rect 26789 46047 26847 46053
rect 28534 46044 28540 46056
rect 28592 46044 28598 46096
rect 28644 46084 28672 46112
rect 29178 46084 29184 46096
rect 28644 46056 29184 46084
rect 29178 46044 29184 46056
rect 29236 46044 29242 46096
rect 12802 46016 12808 46028
rect 12763 45988 12808 46016
rect 12802 45976 12808 45988
rect 12860 45976 12866 46028
rect 13909 46019 13967 46025
rect 13909 45985 13921 46019
rect 13955 46016 13967 46019
rect 14734 46016 14740 46028
rect 13955 45988 14740 46016
rect 13955 45985 13967 45988
rect 13909 45979 13967 45985
rect 14734 45976 14740 45988
rect 14792 45976 14798 46028
rect 21174 45976 21180 46028
rect 21232 46016 21238 46028
rect 21453 46019 21511 46025
rect 21453 46016 21465 46019
rect 21232 45988 21465 46016
rect 21232 45976 21238 45988
rect 21453 45985 21465 45988
rect 21499 45985 21511 46019
rect 21453 45979 21511 45985
rect 22097 46019 22155 46025
rect 22097 45985 22109 46019
rect 22143 46016 22155 46019
rect 22278 46016 22284 46028
rect 22143 45988 22284 46016
rect 22143 45985 22155 45988
rect 22097 45979 22155 45985
rect 22278 45976 22284 45988
rect 22336 46016 22342 46028
rect 22465 46019 22523 46025
rect 22465 46016 22477 46019
rect 22336 45988 22477 46016
rect 22336 45976 22342 45988
rect 22465 45985 22477 45988
rect 22511 45985 22523 46019
rect 22738 46016 22744 46028
rect 22651 45988 22744 46016
rect 22465 45979 22523 45985
rect 13817 45951 13875 45957
rect 13817 45917 13829 45951
rect 13863 45948 13875 45951
rect 13998 45948 14004 45960
rect 13863 45920 14004 45948
rect 13863 45917 13875 45920
rect 13817 45911 13875 45917
rect 13998 45908 14004 45920
rect 14056 45908 14062 45960
rect 22480 45948 22508 45979
rect 22738 45976 22744 45988
rect 22796 45976 22802 46028
rect 24854 46016 24860 46028
rect 24815 45988 24860 46016
rect 24854 45976 24860 45988
rect 24912 45976 24918 46028
rect 27522 46016 27528 46028
rect 27483 45988 27528 46016
rect 27522 45976 27528 45988
rect 27580 45976 27586 46028
rect 27614 45976 27620 46028
rect 27672 46016 27678 46028
rect 28077 46019 28135 46025
rect 28077 46016 28089 46019
rect 27672 45988 28089 46016
rect 27672 45976 27678 45988
rect 28077 45985 28089 45988
rect 28123 45985 28135 46019
rect 28077 45979 28135 45985
rect 28261 46019 28319 46025
rect 28261 45985 28273 46019
rect 28307 46016 28319 46019
rect 28350 46016 28356 46028
rect 28307 45988 28356 46016
rect 28307 45985 28319 45988
rect 28261 45979 28319 45985
rect 28350 45976 28356 45988
rect 28408 45976 28414 46028
rect 29086 45976 29092 46028
rect 29144 46016 29150 46028
rect 29273 46019 29331 46025
rect 29273 46016 29285 46019
rect 29144 45988 29285 46016
rect 29144 45976 29150 45988
rect 29273 45985 29285 45988
rect 29319 45985 29331 46019
rect 29273 45979 29331 45985
rect 29917 46019 29975 46025
rect 29917 45985 29929 46019
rect 29963 46016 29975 46019
rect 30745 46019 30803 46025
rect 30745 46016 30757 46019
rect 29963 45988 30757 46016
rect 29963 45985 29975 45988
rect 29917 45979 29975 45985
rect 30745 45985 30757 45988
rect 30791 46016 30803 46019
rect 31018 46016 31024 46028
rect 30791 45988 31024 46016
rect 30791 45985 30803 45988
rect 30745 45979 30803 45985
rect 31018 45976 31024 45988
rect 31076 45976 31082 46028
rect 32122 46016 32128 46028
rect 32083 45988 32128 46016
rect 32122 45976 32128 45988
rect 32180 45976 32186 46028
rect 32214 45976 32220 46028
rect 32272 46016 32278 46028
rect 32272 45988 32317 46016
rect 32272 45976 32278 45988
rect 22922 45948 22928 45960
rect 22480 45920 22784 45948
rect 22883 45920 22928 45948
rect 21634 45880 21640 45892
rect 21595 45852 21640 45880
rect 21634 45840 21640 45852
rect 21692 45880 21698 45892
rect 21692 45852 22324 45880
rect 21692 45840 21698 45852
rect 12989 45815 13047 45821
rect 12989 45781 13001 45815
rect 13035 45812 13047 45815
rect 13262 45812 13268 45824
rect 13035 45784 13268 45812
rect 13035 45781 13047 45784
rect 12989 45775 13047 45781
rect 13262 45772 13268 45784
rect 13320 45812 13326 45824
rect 14921 45815 14979 45821
rect 14921 45812 14933 45815
rect 13320 45784 14933 45812
rect 13320 45772 13326 45784
rect 14921 45781 14933 45784
rect 14967 45812 14979 45815
rect 15654 45812 15660 45824
rect 14967 45784 15660 45812
rect 14967 45781 14979 45784
rect 14921 45775 14979 45781
rect 15654 45772 15660 45784
rect 15712 45772 15718 45824
rect 22296 45812 22324 45852
rect 22370 45840 22376 45892
rect 22428 45880 22434 45892
rect 22557 45883 22615 45889
rect 22557 45880 22569 45883
rect 22428 45852 22569 45880
rect 22428 45840 22434 45852
rect 22557 45849 22569 45852
rect 22603 45849 22615 45883
rect 22756 45880 22784 45920
rect 22922 45908 22928 45920
rect 22980 45908 22986 45960
rect 24026 45948 24032 45960
rect 23987 45920 24032 45948
rect 24026 45908 24032 45920
rect 24084 45908 24090 45960
rect 24581 45951 24639 45957
rect 24581 45917 24593 45951
rect 24627 45917 24639 45951
rect 24581 45911 24639 45917
rect 23382 45880 23388 45892
rect 22756 45852 23388 45880
rect 22557 45843 22615 45849
rect 23382 45840 23388 45852
rect 23440 45880 23446 45892
rect 24302 45880 24308 45892
rect 23440 45852 24308 45880
rect 23440 45840 23446 45852
rect 24302 45840 24308 45852
rect 24360 45880 24366 45892
rect 24596 45880 24624 45911
rect 24670 45908 24676 45960
rect 24728 45948 24734 45960
rect 25041 45951 25099 45957
rect 25041 45948 25053 45951
rect 24728 45920 25053 45948
rect 24728 45908 24734 45920
rect 25041 45917 25053 45920
rect 25087 45917 25099 45951
rect 25041 45911 25099 45917
rect 24360 45852 24624 45880
rect 24360 45840 24366 45852
rect 23474 45812 23480 45824
rect 22296 45784 23480 45812
rect 23474 45772 23480 45784
rect 23532 45772 23538 45824
rect 25406 45812 25412 45824
rect 25367 45784 25412 45812
rect 25406 45772 25412 45784
rect 25464 45772 25470 45824
rect 26237 45815 26295 45821
rect 26237 45781 26249 45815
rect 26283 45812 26295 45815
rect 26418 45812 26424 45824
rect 26283 45784 26424 45812
rect 26283 45781 26295 45784
rect 26237 45775 26295 45781
rect 26418 45772 26424 45784
rect 26476 45772 26482 45824
rect 30466 45772 30472 45824
rect 30524 45812 30530 45824
rect 30929 45815 30987 45821
rect 30929 45812 30941 45815
rect 30524 45784 30941 45812
rect 30524 45772 30530 45784
rect 30929 45781 30941 45784
rect 30975 45781 30987 45815
rect 30929 45775 30987 45781
rect 31386 45772 31392 45824
rect 31444 45812 31450 45824
rect 31573 45815 31631 45821
rect 31573 45812 31585 45815
rect 31444 45784 31585 45812
rect 31444 45772 31450 45784
rect 31573 45781 31585 45784
rect 31619 45781 31631 45815
rect 32398 45812 32404 45824
rect 32359 45784 32404 45812
rect 31573 45775 31631 45781
rect 32398 45772 32404 45784
rect 32456 45772 32462 45824
rect 1104 45722 38824 45744
rect 1104 45670 4246 45722
rect 4298 45670 4310 45722
rect 4362 45670 4374 45722
rect 4426 45670 4438 45722
rect 4490 45670 34966 45722
rect 35018 45670 35030 45722
rect 35082 45670 35094 45722
rect 35146 45670 35158 45722
rect 35210 45670 38824 45722
rect 1104 45648 38824 45670
rect 14734 45608 14740 45620
rect 14695 45580 14740 45608
rect 14734 45568 14740 45580
rect 14792 45568 14798 45620
rect 22465 45611 22523 45617
rect 22465 45577 22477 45611
rect 22511 45608 22523 45611
rect 22922 45608 22928 45620
rect 22511 45580 22928 45608
rect 22511 45577 22523 45580
rect 22465 45571 22523 45577
rect 8754 45500 8760 45552
rect 8812 45540 8818 45552
rect 8812 45512 9904 45540
rect 8812 45500 8818 45512
rect 9876 45484 9904 45512
rect 9858 45472 9864 45484
rect 9771 45444 9864 45472
rect 9858 45432 9864 45444
rect 9916 45432 9922 45484
rect 13354 45472 13360 45484
rect 13315 45444 13360 45472
rect 13354 45432 13360 45444
rect 13412 45432 13418 45484
rect 8757 45407 8815 45413
rect 8757 45373 8769 45407
rect 8803 45404 8815 45407
rect 8941 45407 8999 45413
rect 8941 45404 8953 45407
rect 8803 45376 8953 45404
rect 8803 45373 8815 45376
rect 8757 45367 8815 45373
rect 8941 45373 8953 45376
rect 8987 45404 8999 45407
rect 9122 45404 9128 45416
rect 8987 45376 9128 45404
rect 8987 45373 8999 45376
rect 8941 45367 8999 45373
rect 9122 45364 9128 45376
rect 9180 45364 9186 45416
rect 9674 45364 9680 45416
rect 9732 45404 9738 45416
rect 9769 45407 9827 45413
rect 9769 45404 9781 45407
rect 9732 45376 9781 45404
rect 9732 45364 9738 45376
rect 9769 45373 9781 45376
rect 9815 45373 9827 45407
rect 9769 45367 9827 45373
rect 13446 45364 13452 45416
rect 13504 45404 13510 45416
rect 22572 45413 22600 45580
rect 22922 45568 22928 45580
rect 22980 45568 22986 45620
rect 23109 45611 23167 45617
rect 23109 45577 23121 45611
rect 23155 45608 23167 45611
rect 23382 45608 23388 45620
rect 23155 45580 23388 45608
rect 23155 45577 23167 45580
rect 23109 45571 23167 45577
rect 23382 45568 23388 45580
rect 23440 45568 23446 45620
rect 25958 45608 25964 45620
rect 24780 45580 25964 45608
rect 22741 45543 22799 45549
rect 22741 45509 22753 45543
rect 22787 45509 22799 45543
rect 22741 45503 22799 45509
rect 22756 45472 22784 45503
rect 23474 45500 23480 45552
rect 23532 45540 23538 45552
rect 24029 45543 24087 45549
rect 24029 45540 24041 45543
rect 23532 45512 24041 45540
rect 23532 45500 23538 45512
rect 24029 45509 24041 45512
rect 24075 45540 24087 45543
rect 24670 45540 24676 45552
rect 24075 45512 24676 45540
rect 24075 45509 24087 45512
rect 24029 45503 24087 45509
rect 24670 45500 24676 45512
rect 24728 45500 24734 45552
rect 23934 45472 23940 45484
rect 22756 45444 23940 45472
rect 23934 45432 23940 45444
rect 23992 45432 23998 45484
rect 24780 45413 24808 45580
rect 25958 45568 25964 45580
rect 26016 45568 26022 45620
rect 26510 45568 26516 45620
rect 26568 45608 26574 45620
rect 27614 45608 27620 45620
rect 26568 45580 27620 45608
rect 26568 45568 26574 45580
rect 27614 45568 27620 45580
rect 27672 45568 27678 45620
rect 28166 45568 28172 45620
rect 28224 45608 28230 45620
rect 28721 45611 28779 45617
rect 28721 45608 28733 45611
rect 28224 45580 28733 45608
rect 28224 45568 28230 45580
rect 28721 45577 28733 45580
rect 28767 45608 28779 45611
rect 30745 45611 30803 45617
rect 30745 45608 30757 45611
rect 28767 45580 30757 45608
rect 28767 45577 28779 45580
rect 28721 45571 28779 45577
rect 30745 45577 30757 45580
rect 30791 45608 30803 45611
rect 31018 45608 31024 45620
rect 30791 45580 31024 45608
rect 30791 45577 30803 45580
rect 30745 45571 30803 45577
rect 31018 45568 31024 45580
rect 31076 45568 31082 45620
rect 32122 45608 32128 45620
rect 32083 45580 32128 45608
rect 32122 45568 32128 45580
rect 32180 45568 32186 45620
rect 32214 45568 32220 45620
rect 32272 45608 32278 45620
rect 32493 45611 32551 45617
rect 32493 45608 32505 45611
rect 32272 45580 32505 45608
rect 32272 45568 32278 45580
rect 32493 45577 32505 45580
rect 32539 45577 32551 45611
rect 32493 45571 32551 45577
rect 28074 45540 28080 45552
rect 28035 45512 28080 45540
rect 28074 45500 28080 45512
rect 28132 45500 28138 45552
rect 29086 45540 29092 45552
rect 29047 45512 29092 45540
rect 29086 45500 29092 45512
rect 29144 45500 29150 45552
rect 29454 45500 29460 45552
rect 29512 45540 29518 45552
rect 29730 45540 29736 45552
rect 29512 45512 29736 45540
rect 29512 45500 29518 45512
rect 29730 45500 29736 45512
rect 29788 45500 29794 45552
rect 25225 45475 25283 45481
rect 25225 45441 25237 45475
rect 25271 45472 25283 45475
rect 25406 45472 25412 45484
rect 25271 45444 25412 45472
rect 25271 45441 25283 45444
rect 25225 45435 25283 45441
rect 25406 45432 25412 45444
rect 25464 45432 25470 45484
rect 26053 45475 26111 45481
rect 26053 45441 26065 45475
rect 26099 45472 26111 45475
rect 26602 45472 26608 45484
rect 26099 45444 26608 45472
rect 26099 45441 26111 45444
rect 26053 45435 26111 45441
rect 26602 45432 26608 45444
rect 26660 45472 26666 45484
rect 26660 45444 27200 45472
rect 26660 45432 26666 45444
rect 13633 45407 13691 45413
rect 13633 45404 13645 45407
rect 13504 45376 13645 45404
rect 13504 45364 13510 45376
rect 13633 45373 13645 45376
rect 13679 45373 13691 45407
rect 13633 45367 13691 45373
rect 22557 45407 22615 45413
rect 22557 45373 22569 45407
rect 22603 45373 22615 45407
rect 22557 45367 22615 45373
rect 24765 45407 24823 45413
rect 24765 45373 24777 45407
rect 24811 45373 24823 45407
rect 24765 45367 24823 45373
rect 25038 45364 25044 45416
rect 25096 45404 25102 45416
rect 25133 45407 25191 45413
rect 25133 45404 25145 45407
rect 25096 45376 25145 45404
rect 25096 45364 25102 45376
rect 25133 45373 25145 45376
rect 25179 45373 25191 45407
rect 25133 45367 25191 45373
rect 26145 45407 26203 45413
rect 26145 45373 26157 45407
rect 26191 45404 26203 45407
rect 26510 45404 26516 45416
rect 26191 45376 26516 45404
rect 26191 45373 26203 45376
rect 26145 45367 26203 45373
rect 26510 45364 26516 45376
rect 26568 45364 26574 45416
rect 26786 45404 26792 45416
rect 26747 45376 26792 45404
rect 26786 45364 26792 45376
rect 26844 45364 26850 45416
rect 26878 45364 26884 45416
rect 26936 45404 26942 45416
rect 27172 45413 27200 45444
rect 27982 45432 27988 45484
rect 28040 45432 28046 45484
rect 28994 45432 29000 45484
rect 29052 45472 29058 45484
rect 30009 45475 30067 45481
rect 30009 45472 30021 45475
rect 29052 45444 30021 45472
rect 29052 45432 29058 45444
rect 30009 45441 30021 45444
rect 30055 45441 30067 45475
rect 30009 45435 30067 45441
rect 27157 45407 27215 45413
rect 26936 45376 26981 45404
rect 26936 45364 26942 45376
rect 27157 45373 27169 45407
rect 27203 45373 27215 45407
rect 27338 45404 27344 45416
rect 27299 45376 27344 45404
rect 27157 45367 27215 45373
rect 27338 45364 27344 45376
rect 27396 45364 27402 45416
rect 8570 45296 8576 45348
rect 8628 45336 8634 45348
rect 9033 45339 9091 45345
rect 9033 45336 9045 45339
rect 8628 45308 9045 45336
rect 8628 45296 8634 45308
rect 9033 45305 9045 45308
rect 9079 45305 9091 45339
rect 9033 45299 9091 45305
rect 22462 45296 22468 45348
rect 22520 45336 22526 45348
rect 22520 45308 23520 45336
rect 22520 45296 22526 45308
rect 12802 45268 12808 45280
rect 12763 45240 12808 45268
rect 12802 45228 12808 45240
rect 12860 45228 12866 45280
rect 13265 45271 13323 45277
rect 13265 45237 13277 45271
rect 13311 45268 13323 45271
rect 13998 45268 14004 45280
rect 13311 45240 14004 45268
rect 13311 45237 13323 45240
rect 13265 45231 13323 45237
rect 13998 45228 14004 45240
rect 14056 45228 14062 45280
rect 21174 45228 21180 45280
rect 21232 45268 21238 45280
rect 21453 45271 21511 45277
rect 21453 45268 21465 45271
rect 21232 45240 21465 45268
rect 21232 45228 21238 45240
rect 21453 45237 21465 45240
rect 21499 45268 21511 45271
rect 22005 45271 22063 45277
rect 22005 45268 22017 45271
rect 21499 45240 22017 45268
rect 21499 45237 21511 45240
rect 21453 45231 21511 45237
rect 22005 45237 22017 45240
rect 22051 45268 22063 45271
rect 22738 45268 22744 45280
rect 22051 45240 22744 45268
rect 22051 45237 22063 45240
rect 22005 45231 22063 45237
rect 22738 45228 22744 45240
rect 22796 45228 22802 45280
rect 23492 45277 23520 45308
rect 24118 45296 24124 45348
rect 24176 45336 24182 45348
rect 24305 45339 24363 45345
rect 24305 45336 24317 45339
rect 24176 45308 24317 45336
rect 24176 45296 24182 45308
rect 24305 45305 24317 45308
rect 24351 45305 24363 45339
rect 24305 45299 24363 45305
rect 25685 45339 25743 45345
rect 25685 45305 25697 45339
rect 25731 45336 25743 45339
rect 27356 45336 27384 45364
rect 25731 45308 27384 45336
rect 25731 45305 25743 45308
rect 25685 45299 25743 45305
rect 28000 45280 28028 45432
rect 28166 45404 28172 45416
rect 28127 45376 28172 45404
rect 28166 45364 28172 45376
rect 28224 45364 28230 45416
rect 28902 45364 28908 45416
rect 28960 45404 28966 45416
rect 29549 45407 29607 45413
rect 29549 45404 29561 45407
rect 28960 45376 29561 45404
rect 28960 45364 28966 45376
rect 29549 45373 29561 45376
rect 29595 45404 29607 45407
rect 30190 45404 30196 45416
rect 29595 45376 30196 45404
rect 29595 45373 29607 45376
rect 29549 45367 29607 45373
rect 30190 45364 30196 45376
rect 30248 45404 30254 45416
rect 31113 45407 31171 45413
rect 31113 45404 31125 45407
rect 30248 45376 31125 45404
rect 30248 45364 30254 45376
rect 31113 45373 31125 45376
rect 31159 45404 31171 45407
rect 31478 45404 31484 45416
rect 31159 45376 31484 45404
rect 31159 45373 31171 45376
rect 31113 45367 31171 45373
rect 31478 45364 31484 45376
rect 31536 45364 31542 45416
rect 29270 45336 29276 45348
rect 29231 45308 29276 45336
rect 29270 45296 29276 45308
rect 29328 45336 29334 45348
rect 29641 45339 29699 45345
rect 29328 45308 29592 45336
rect 29328 45296 29334 45308
rect 23477 45271 23535 45277
rect 23477 45237 23489 45271
rect 23523 45268 23535 45271
rect 24854 45268 24860 45280
rect 23523 45240 24860 45268
rect 23523 45237 23535 45240
rect 23477 45231 23535 45237
rect 24854 45228 24860 45240
rect 24912 45228 24918 45280
rect 27982 45228 27988 45280
rect 28040 45228 28046 45280
rect 28353 45271 28411 45277
rect 28353 45237 28365 45271
rect 28399 45268 28411 45271
rect 28442 45268 28448 45280
rect 28399 45240 28448 45268
rect 28399 45237 28411 45240
rect 28353 45231 28411 45237
rect 28442 45228 28448 45240
rect 28500 45228 28506 45280
rect 29178 45228 29184 45280
rect 29236 45268 29242 45280
rect 29457 45271 29515 45277
rect 29457 45268 29469 45271
rect 29236 45240 29469 45268
rect 29236 45228 29242 45240
rect 29457 45237 29469 45240
rect 29503 45237 29515 45271
rect 29564 45268 29592 45308
rect 29641 45305 29653 45339
rect 29687 45336 29699 45339
rect 29730 45336 29736 45348
rect 29687 45308 29736 45336
rect 29687 45305 29699 45308
rect 29641 45299 29699 45305
rect 29730 45296 29736 45308
rect 29788 45296 29794 45348
rect 30837 45339 30895 45345
rect 30837 45305 30849 45339
rect 30883 45305 30895 45339
rect 30837 45299 30895 45305
rect 30285 45271 30343 45277
rect 30285 45268 30297 45271
rect 29564 45240 30297 45268
rect 29457 45231 29515 45237
rect 30285 45237 30297 45240
rect 30331 45268 30343 45271
rect 30852 45268 30880 45299
rect 30926 45296 30932 45348
rect 30984 45336 30990 45348
rect 31021 45339 31079 45345
rect 31021 45336 31033 45339
rect 30984 45308 31033 45336
rect 30984 45296 30990 45308
rect 31021 45305 31033 45308
rect 31067 45305 31079 45339
rect 31021 45299 31079 45305
rect 31205 45339 31263 45345
rect 31205 45305 31217 45339
rect 31251 45336 31263 45339
rect 31386 45336 31392 45348
rect 31251 45308 31392 45336
rect 31251 45305 31263 45308
rect 31205 45299 31263 45305
rect 31386 45296 31392 45308
rect 31444 45296 31450 45348
rect 31570 45336 31576 45348
rect 31531 45308 31576 45336
rect 31570 45296 31576 45308
rect 31628 45296 31634 45348
rect 30331 45240 30880 45268
rect 30331 45237 30343 45240
rect 30285 45231 30343 45237
rect 1104 45178 38824 45200
rect 1104 45126 19606 45178
rect 19658 45126 19670 45178
rect 19722 45126 19734 45178
rect 19786 45126 19798 45178
rect 19850 45126 38824 45178
rect 1104 45104 38824 45126
rect 8754 45024 8760 45076
rect 8812 45064 8818 45076
rect 8849 45067 8907 45073
rect 8849 45064 8861 45067
rect 8812 45036 8861 45064
rect 8812 45024 8818 45036
rect 8849 45033 8861 45036
rect 8895 45033 8907 45067
rect 8849 45027 8907 45033
rect 13354 45024 13360 45076
rect 13412 45064 13418 45076
rect 13541 45067 13599 45073
rect 13541 45064 13553 45067
rect 13412 45036 13553 45064
rect 13412 45024 13418 45036
rect 13541 45033 13553 45036
rect 13587 45033 13599 45067
rect 13541 45027 13599 45033
rect 14369 45067 14427 45073
rect 14369 45033 14381 45067
rect 14415 45064 14427 45067
rect 14734 45064 14740 45076
rect 14415 45036 14740 45064
rect 14415 45033 14427 45036
rect 14369 45027 14427 45033
rect 14734 45024 14740 45036
rect 14792 45024 14798 45076
rect 22462 45064 22468 45076
rect 22423 45036 22468 45064
rect 22462 45024 22468 45036
rect 22520 45024 22526 45076
rect 22738 45024 22744 45076
rect 22796 45064 22802 45076
rect 22796 45036 22841 45064
rect 22796 45024 22802 45036
rect 23014 45024 23020 45076
rect 23072 45064 23078 45076
rect 23109 45067 23167 45073
rect 23109 45064 23121 45067
rect 23072 45036 23121 45064
rect 23072 45024 23078 45036
rect 23109 45033 23121 45036
rect 23155 45033 23167 45067
rect 23750 45064 23756 45076
rect 23711 45036 23756 45064
rect 23109 45027 23167 45033
rect 23750 45024 23756 45036
rect 23808 45064 23814 45076
rect 24673 45067 24731 45073
rect 24673 45064 24685 45067
rect 23808 45036 24685 45064
rect 23808 45024 23814 45036
rect 24673 45033 24685 45036
rect 24719 45064 24731 45067
rect 24719 45036 25176 45064
rect 24719 45033 24731 45036
rect 24673 45027 24731 45033
rect 24302 44996 24308 45008
rect 24263 44968 24308 44996
rect 24302 44956 24308 44968
rect 24360 44956 24366 45008
rect 1762 44928 1768 44940
rect 1723 44900 1768 44928
rect 1762 44888 1768 44900
rect 1820 44888 1826 44940
rect 13722 44928 13728 44940
rect 13683 44900 13728 44928
rect 13722 44888 13728 44900
rect 13780 44888 13786 44940
rect 13817 44931 13875 44937
rect 13817 44897 13829 44931
rect 13863 44928 13875 44931
rect 14090 44928 14096 44940
rect 13863 44900 14096 44928
rect 13863 44897 13875 44900
rect 13817 44891 13875 44897
rect 14090 44888 14096 44900
rect 14148 44888 14154 44940
rect 22281 44931 22339 44937
rect 22281 44897 22293 44931
rect 22327 44897 22339 44931
rect 23842 44928 23848 44940
rect 23803 44900 23848 44928
rect 22281 44891 22339 44897
rect 1394 44820 1400 44872
rect 1452 44860 1458 44872
rect 1489 44863 1547 44869
rect 1489 44860 1501 44863
rect 1452 44832 1501 44860
rect 1452 44820 1458 44832
rect 1489 44829 1501 44832
rect 1535 44860 1547 44863
rect 1946 44860 1952 44872
rect 1535 44832 1952 44860
rect 1535 44829 1547 44832
rect 1489 44823 1547 44829
rect 1946 44820 1952 44832
rect 2004 44820 2010 44872
rect 12529 44795 12587 44801
rect 12529 44761 12541 44795
rect 12575 44792 12587 44795
rect 13078 44792 13084 44804
rect 12575 44764 13084 44792
rect 12575 44761 12587 44764
rect 12529 44755 12587 44761
rect 13078 44752 13084 44764
rect 13136 44752 13142 44804
rect 13446 44792 13452 44804
rect 13359 44764 13452 44792
rect 13446 44752 13452 44764
rect 13504 44792 13510 44804
rect 14458 44792 14464 44804
rect 13504 44764 14464 44792
rect 13504 44752 13510 44764
rect 14458 44752 14464 44764
rect 14516 44752 14522 44804
rect 3050 44724 3056 44736
rect 3011 44696 3056 44724
rect 3050 44684 3056 44696
rect 3108 44684 3114 44736
rect 12894 44724 12900 44736
rect 12855 44696 12900 44724
rect 12894 44684 12900 44696
rect 12952 44684 12958 44736
rect 13998 44724 14004 44736
rect 13911 44696 14004 44724
rect 13998 44684 14004 44696
rect 14056 44724 14062 44736
rect 15102 44724 15108 44736
rect 14056 44696 15108 44724
rect 14056 44684 14062 44696
rect 15102 44684 15108 44696
rect 15160 44684 15166 44736
rect 22189 44727 22247 44733
rect 22189 44693 22201 44727
rect 22235 44724 22247 44727
rect 22296 44724 22324 44891
rect 23842 44888 23848 44900
rect 23900 44888 23906 44940
rect 24670 44888 24676 44940
rect 24728 44928 24734 44940
rect 24857 44931 24915 44937
rect 24857 44928 24869 44931
rect 24728 44900 24869 44928
rect 24728 44888 24734 44900
rect 24857 44897 24869 44900
rect 24903 44897 24915 44931
rect 24857 44891 24915 44897
rect 24872 44860 24900 44891
rect 24946 44888 24952 44940
rect 25004 44928 25010 44940
rect 25148 44937 25176 45036
rect 26326 45024 26332 45076
rect 26384 45064 26390 45076
rect 26697 45067 26755 45073
rect 26697 45064 26709 45067
rect 26384 45036 26709 45064
rect 26384 45024 26390 45036
rect 26697 45033 26709 45036
rect 26743 45033 26755 45067
rect 27430 45064 27436 45076
rect 27391 45036 27436 45064
rect 26697 45027 26755 45033
rect 27430 45024 27436 45036
rect 27488 45024 27494 45076
rect 28350 45024 28356 45076
rect 28408 45064 28414 45076
rect 28534 45064 28540 45076
rect 28408 45036 28540 45064
rect 28408 45024 28414 45036
rect 28534 45024 28540 45036
rect 28592 45024 28598 45076
rect 29365 45067 29423 45073
rect 29365 45033 29377 45067
rect 29411 45064 29423 45067
rect 29914 45064 29920 45076
rect 29411 45036 29920 45064
rect 29411 45033 29423 45036
rect 29365 45027 29423 45033
rect 25041 44931 25099 44937
rect 25041 44928 25053 44931
rect 25004 44900 25053 44928
rect 25004 44888 25010 44900
rect 25041 44897 25053 44900
rect 25087 44897 25099 44931
rect 25041 44891 25099 44897
rect 25133 44931 25191 44937
rect 25133 44897 25145 44931
rect 25179 44897 25191 44931
rect 25133 44891 25191 44897
rect 26513 44931 26571 44937
rect 26513 44897 26525 44931
rect 26559 44897 26571 44931
rect 26513 44891 26571 44897
rect 26528 44860 26556 44891
rect 27614 44888 27620 44940
rect 27672 44928 27678 44940
rect 28169 44931 28227 44937
rect 28169 44928 28181 44931
rect 27672 44900 28181 44928
rect 27672 44888 27678 44900
rect 28169 44897 28181 44900
rect 28215 44897 28227 44931
rect 28534 44928 28540 44940
rect 28495 44900 28540 44928
rect 28169 44891 28227 44897
rect 28534 44888 28540 44900
rect 28592 44888 28598 44940
rect 28721 44931 28779 44937
rect 28721 44897 28733 44931
rect 28767 44928 28779 44931
rect 29380 44928 29408 45027
rect 29914 45024 29920 45036
rect 29972 45064 29978 45076
rect 30466 45064 30472 45076
rect 29972 45036 30472 45064
rect 29972 45024 29978 45036
rect 30466 45024 30472 45036
rect 30524 45024 30530 45076
rect 30834 45024 30840 45076
rect 30892 45064 30898 45076
rect 30929 45067 30987 45073
rect 30929 45064 30941 45067
rect 30892 45036 30941 45064
rect 30892 45024 30898 45036
rect 30929 45033 30941 45036
rect 30975 45033 30987 45067
rect 31478 45064 31484 45076
rect 31439 45036 31484 45064
rect 30929 45027 30987 45033
rect 31478 45024 31484 45036
rect 31536 45024 31542 45076
rect 29546 44928 29552 44940
rect 28767 44900 29408 44928
rect 29507 44900 29552 44928
rect 28767 44897 28779 44900
rect 28721 44891 28779 44897
rect 29546 44888 29552 44900
rect 29604 44888 29610 44940
rect 26694 44860 26700 44872
rect 24872 44832 26700 44860
rect 26694 44820 26700 44832
rect 26752 44820 26758 44872
rect 28261 44863 28319 44869
rect 28261 44829 28273 44863
rect 28307 44860 28319 44863
rect 28626 44860 28632 44872
rect 28307 44832 28632 44860
rect 28307 44829 28319 44832
rect 28261 44823 28319 44829
rect 28626 44820 28632 44832
rect 28684 44820 28690 44872
rect 29822 44860 29828 44872
rect 29783 44832 29828 44860
rect 29822 44820 29828 44832
rect 29880 44820 29886 44872
rect 26329 44795 26387 44801
rect 26329 44761 26341 44795
rect 26375 44792 26387 44795
rect 26878 44792 26884 44804
rect 26375 44764 26884 44792
rect 26375 44761 26387 44764
rect 26329 44755 26387 44761
rect 26878 44752 26884 44764
rect 26936 44752 26942 44804
rect 27706 44752 27712 44804
rect 27764 44792 27770 44804
rect 28074 44792 28080 44804
rect 27764 44764 28080 44792
rect 27764 44752 27770 44764
rect 28074 44752 28080 44764
rect 28132 44752 28138 44804
rect 22370 44724 22376 44736
rect 22235 44696 22376 44724
rect 22235 44693 22247 44696
rect 22189 44687 22247 44693
rect 22370 44684 22376 44696
rect 22428 44684 22434 44736
rect 25222 44684 25228 44736
rect 25280 44724 25286 44736
rect 25317 44727 25375 44733
rect 25317 44724 25329 44727
rect 25280 44696 25329 44724
rect 25280 44684 25286 44696
rect 25317 44693 25329 44696
rect 25363 44724 25375 44727
rect 25774 44724 25780 44736
rect 25363 44696 25780 44724
rect 25363 44693 25375 44696
rect 25317 44687 25375 44693
rect 25774 44684 25780 44696
rect 25832 44684 25838 44736
rect 25958 44724 25964 44736
rect 25919 44696 25964 44724
rect 25958 44684 25964 44696
rect 26016 44684 26022 44736
rect 26786 44684 26792 44736
rect 26844 44724 26850 44736
rect 27065 44727 27123 44733
rect 27065 44724 27077 44727
rect 26844 44696 27077 44724
rect 26844 44684 26850 44696
rect 27065 44693 27077 44696
rect 27111 44724 27123 44727
rect 27246 44724 27252 44736
rect 27111 44696 27252 44724
rect 27111 44693 27123 44696
rect 27065 44687 27123 44693
rect 27246 44684 27252 44696
rect 27304 44684 27310 44736
rect 27617 44727 27675 44733
rect 27617 44693 27629 44727
rect 27663 44724 27675 44727
rect 27798 44724 27804 44736
rect 27663 44696 27804 44724
rect 27663 44693 27675 44696
rect 27617 44687 27675 44693
rect 27798 44684 27804 44696
rect 27856 44684 27862 44736
rect 31846 44724 31852 44736
rect 31807 44696 31852 44724
rect 31846 44684 31852 44696
rect 31904 44684 31910 44736
rect 1104 44634 38824 44656
rect 1104 44582 4246 44634
rect 4298 44582 4310 44634
rect 4362 44582 4374 44634
rect 4426 44582 4438 44634
rect 4490 44582 34966 44634
rect 35018 44582 35030 44634
rect 35082 44582 35094 44634
rect 35146 44582 35158 44634
rect 35210 44582 38824 44634
rect 1104 44560 38824 44582
rect 1673 44523 1731 44529
rect 1673 44489 1685 44523
rect 1719 44520 1731 44523
rect 1762 44520 1768 44532
rect 1719 44492 1768 44520
rect 1719 44489 1731 44492
rect 1673 44483 1731 44489
rect 1762 44480 1768 44492
rect 1820 44480 1826 44532
rect 8110 44520 8116 44532
rect 8071 44492 8116 44520
rect 8110 44480 8116 44492
rect 8168 44480 8174 44532
rect 13722 44480 13728 44532
rect 13780 44520 13786 44532
rect 14277 44523 14335 44529
rect 14277 44520 14289 44523
rect 13780 44492 14289 44520
rect 13780 44480 13786 44492
rect 14277 44489 14289 44492
rect 14323 44520 14335 44523
rect 15473 44523 15531 44529
rect 15473 44520 15485 44523
rect 14323 44492 15485 44520
rect 14323 44489 14335 44492
rect 14277 44483 14335 44489
rect 15473 44489 15485 44492
rect 15519 44489 15531 44523
rect 15930 44520 15936 44532
rect 15891 44492 15936 44520
rect 15473 44483 15531 44489
rect 8128 44384 8156 44480
rect 13814 44412 13820 44464
rect 13872 44452 13878 44464
rect 14001 44455 14059 44461
rect 14001 44452 14013 44455
rect 13872 44424 14013 44452
rect 13872 44412 13878 44424
rect 14001 44421 14013 44424
rect 14047 44452 14059 44455
rect 14090 44452 14096 44464
rect 14047 44424 14096 44452
rect 14047 44421 14059 44424
rect 14001 44415 14059 44421
rect 14090 44412 14096 44424
rect 14148 44412 14154 44464
rect 15488 44452 15516 44483
rect 15930 44480 15936 44492
rect 15988 44480 15994 44532
rect 24670 44480 24676 44532
rect 24728 44520 24734 44532
rect 24857 44523 24915 44529
rect 24857 44520 24869 44523
rect 24728 44492 24869 44520
rect 24728 44480 24734 44492
rect 24857 44489 24869 44492
rect 24903 44489 24915 44523
rect 24857 44483 24915 44489
rect 26694 44480 26700 44532
rect 26752 44520 26758 44532
rect 26789 44523 26847 44529
rect 26789 44520 26801 44523
rect 26752 44492 26801 44520
rect 26752 44480 26758 44492
rect 26789 44489 26801 44492
rect 26835 44489 26847 44523
rect 26789 44483 26847 44489
rect 26878 44480 26884 44532
rect 26936 44520 26942 44532
rect 27249 44523 27307 44529
rect 27249 44520 27261 44523
rect 26936 44492 27261 44520
rect 26936 44480 26942 44492
rect 27249 44489 27261 44492
rect 27295 44520 27307 44523
rect 28626 44520 28632 44532
rect 27295 44492 28632 44520
rect 27295 44489 27307 44492
rect 27249 44483 27307 44489
rect 28626 44480 28632 44492
rect 28684 44480 28690 44532
rect 28721 44523 28779 44529
rect 28721 44489 28733 44523
rect 28767 44520 28779 44523
rect 28902 44520 28908 44532
rect 28767 44492 28908 44520
rect 28767 44489 28779 44492
rect 28721 44483 28779 44489
rect 28902 44480 28908 44492
rect 28960 44480 28966 44532
rect 31110 44520 31116 44532
rect 31071 44492 31116 44520
rect 31110 44480 31116 44492
rect 31168 44480 31174 44532
rect 37642 44520 37648 44532
rect 37603 44492 37648 44520
rect 37642 44480 37648 44492
rect 37700 44480 37706 44532
rect 16574 44452 16580 44464
rect 15488 44424 16580 44452
rect 16574 44412 16580 44424
rect 16632 44412 16638 44464
rect 25317 44455 25375 44461
rect 25317 44421 25329 44455
rect 25363 44452 25375 44455
rect 27890 44452 27896 44464
rect 25363 44424 26372 44452
rect 25363 44421 25375 44424
rect 25317 44415 25375 44421
rect 8573 44387 8631 44393
rect 8573 44384 8585 44387
rect 8128 44356 8585 44384
rect 8573 44353 8585 44356
rect 8619 44353 8631 44387
rect 12526 44384 12532 44396
rect 12487 44356 12532 44384
rect 8573 44347 8631 44353
rect 12526 44344 12532 44356
rect 12584 44344 12590 44396
rect 12894 44384 12900 44396
rect 12855 44356 12900 44384
rect 12894 44344 12900 44356
rect 12952 44344 12958 44396
rect 24581 44387 24639 44393
rect 24581 44353 24593 44387
rect 24627 44384 24639 44387
rect 25501 44387 25559 44393
rect 25501 44384 25513 44387
rect 24627 44356 25513 44384
rect 24627 44353 24639 44356
rect 24581 44347 24639 44353
rect 25501 44353 25513 44356
rect 25547 44384 25559 44387
rect 25958 44384 25964 44396
rect 25547 44356 25964 44384
rect 25547 44353 25559 44356
rect 25501 44347 25559 44353
rect 25958 44344 25964 44356
rect 26016 44344 26022 44396
rect 26344 44384 26372 44424
rect 27632 44424 27896 44452
rect 26602 44384 26608 44396
rect 26344 44356 26608 44384
rect 2038 44316 2044 44328
rect 1999 44288 2044 44316
rect 2038 44276 2044 44288
rect 2096 44276 2102 44328
rect 8294 44316 8300 44328
rect 8255 44288 8300 44316
rect 8294 44276 8300 44288
rect 8352 44276 8358 44328
rect 12250 44276 12256 44328
rect 12308 44316 12314 44328
rect 12912 44316 12940 44344
rect 13078 44316 13084 44328
rect 12308 44288 12940 44316
rect 13039 44288 13084 44316
rect 12308 44276 12314 44288
rect 13078 44276 13084 44288
rect 13136 44276 13142 44328
rect 13449 44319 13507 44325
rect 13449 44285 13461 44319
rect 13495 44285 13507 44319
rect 13449 44279 13507 44285
rect 13541 44319 13599 44325
rect 13541 44285 13553 44319
rect 13587 44285 13599 44319
rect 13541 44279 13599 44285
rect 15657 44319 15715 44325
rect 15657 44285 15669 44319
rect 15703 44316 15715 44319
rect 15930 44316 15936 44328
rect 15703 44288 15936 44316
rect 15703 44285 15715 44288
rect 15657 44279 15715 44285
rect 9953 44251 10011 44257
rect 9953 44217 9965 44251
rect 9999 44248 10011 44251
rect 10962 44248 10968 44260
rect 9999 44220 10968 44248
rect 9999 44217 10011 44220
rect 9953 44211 10011 44217
rect 10962 44208 10968 44220
rect 11020 44208 11026 44260
rect 11885 44251 11943 44257
rect 11885 44217 11897 44251
rect 11931 44248 11943 44251
rect 12526 44248 12532 44260
rect 11931 44220 12532 44248
rect 11931 44217 11943 44220
rect 11885 44211 11943 44217
rect 12526 44208 12532 44220
rect 12584 44248 12590 44260
rect 13464 44248 13492 44279
rect 12584 44220 13492 44248
rect 12584 44208 12590 44220
rect 11790 44140 11796 44192
rect 11848 44180 11854 44192
rect 12161 44183 12219 44189
rect 12161 44180 12173 44183
rect 11848 44152 12173 44180
rect 11848 44140 11854 44152
rect 12161 44149 12173 44152
rect 12207 44180 12219 44183
rect 12802 44180 12808 44192
rect 12207 44152 12808 44180
rect 12207 44149 12219 44152
rect 12161 44143 12219 44149
rect 12802 44140 12808 44152
rect 12860 44180 12866 44192
rect 13556 44180 13584 44279
rect 15930 44276 15936 44288
rect 15988 44276 15994 44328
rect 23385 44319 23443 44325
rect 23385 44285 23397 44319
rect 23431 44316 23443 44319
rect 23842 44316 23848 44328
rect 23431 44288 23848 44316
rect 23431 44285 23443 44288
rect 23385 44279 23443 44285
rect 23842 44276 23848 44288
rect 23900 44276 23906 44328
rect 23937 44319 23995 44325
rect 23937 44285 23949 44319
rect 23983 44316 23995 44319
rect 24026 44316 24032 44328
rect 23983 44288 24032 44316
rect 23983 44285 23995 44288
rect 23937 44279 23995 44285
rect 24026 44276 24032 44288
rect 24084 44276 24090 44328
rect 24210 44316 24216 44328
rect 24171 44288 24216 44316
rect 24210 44276 24216 44288
rect 24268 44276 24274 44328
rect 25593 44319 25651 44325
rect 25593 44285 25605 44319
rect 25639 44316 25651 44319
rect 26142 44316 26148 44328
rect 25639 44288 26148 44316
rect 25639 44285 25651 44288
rect 25593 44279 25651 44285
rect 26142 44276 26148 44288
rect 26200 44276 26206 44328
rect 26344 44325 26372 44356
rect 26602 44344 26608 44356
rect 26660 44384 26666 44396
rect 27522 44384 27528 44396
rect 26660 44356 27528 44384
rect 26660 44344 26666 44356
rect 27522 44344 27528 44356
rect 27580 44344 27586 44396
rect 26329 44319 26387 44325
rect 26329 44285 26341 44319
rect 26375 44285 26387 44319
rect 26329 44279 26387 44285
rect 26418 44276 26424 44328
rect 26476 44316 26482 44328
rect 27632 44316 27660 44424
rect 27890 44412 27896 44424
rect 27948 44412 27954 44464
rect 27982 44412 27988 44464
rect 28040 44452 28046 44464
rect 28040 44424 28304 44452
rect 28040 44412 28046 44424
rect 27706 44344 27712 44396
rect 27764 44384 27770 44396
rect 28276 44393 28304 44424
rect 28261 44387 28319 44393
rect 27764 44356 28212 44384
rect 27764 44344 27770 44356
rect 28184 44325 28212 44356
rect 28261 44353 28273 44387
rect 28307 44353 28319 44387
rect 30834 44384 30840 44396
rect 30747 44356 30840 44384
rect 28261 44347 28319 44353
rect 30834 44344 30840 44356
rect 30892 44384 30898 44396
rect 31665 44387 31723 44393
rect 31665 44384 31677 44387
rect 30892 44356 31677 44384
rect 30892 44344 30898 44356
rect 31665 44353 31677 44356
rect 31711 44353 31723 44387
rect 31665 44347 31723 44353
rect 35989 44387 36047 44393
rect 35989 44353 36001 44387
rect 36035 44384 36047 44387
rect 36035 44356 36400 44384
rect 36035 44353 36047 44356
rect 35989 44347 36047 44353
rect 36372 44328 36400 44356
rect 27801 44319 27859 44325
rect 27801 44316 27813 44319
rect 26476 44288 26521 44316
rect 27632 44288 27813 44316
rect 26476 44276 26482 44288
rect 27801 44285 27813 44288
rect 27847 44285 27859 44319
rect 27801 44279 27859 44285
rect 28169 44319 28227 44325
rect 28169 44285 28181 44319
rect 28215 44316 28227 44319
rect 28902 44316 28908 44328
rect 28215 44288 28908 44316
rect 28215 44285 28227 44288
rect 28169 44279 28227 44285
rect 28902 44276 28908 44288
rect 28960 44276 28966 44328
rect 29086 44316 29092 44328
rect 28999 44288 29092 44316
rect 29086 44276 29092 44288
rect 29144 44316 29150 44328
rect 29273 44319 29331 44325
rect 29273 44316 29285 44319
rect 29144 44288 29285 44316
rect 29144 44276 29150 44288
rect 29273 44285 29285 44288
rect 29319 44285 29331 44319
rect 29273 44279 29331 44285
rect 29733 44319 29791 44325
rect 29733 44285 29745 44319
rect 29779 44316 29791 44319
rect 29914 44316 29920 44328
rect 29779 44288 29920 44316
rect 29779 44285 29791 44288
rect 29733 44279 29791 44285
rect 29914 44276 29920 44288
rect 29972 44276 29978 44328
rect 30742 44316 30748 44328
rect 30655 44288 30748 44316
rect 30742 44276 30748 44288
rect 30800 44316 30806 44328
rect 30929 44319 30987 44325
rect 30929 44316 30941 44319
rect 30800 44288 30941 44316
rect 30800 44276 30806 44288
rect 30929 44285 30941 44288
rect 30975 44285 30987 44319
rect 30929 44279 30987 44285
rect 34146 44276 34152 44328
rect 34204 44316 34210 44328
rect 36078 44316 36084 44328
rect 34204 44288 36084 44316
rect 34204 44276 34210 44288
rect 36078 44276 36084 44288
rect 36136 44276 36142 44328
rect 36354 44316 36360 44328
rect 36315 44288 36360 44316
rect 36354 44276 36360 44288
rect 36412 44276 36418 44328
rect 24946 44208 24952 44260
rect 25004 44248 25010 44260
rect 25498 44248 25504 44260
rect 25004 44220 25504 44248
rect 25004 44208 25010 44220
rect 25498 44208 25504 44220
rect 25556 44208 25562 44260
rect 27338 44248 27344 44260
rect 27299 44220 27344 44248
rect 27338 44208 27344 44220
rect 27396 44208 27402 44260
rect 27614 44208 27620 44260
rect 27672 44248 27678 44260
rect 27672 44220 29408 44248
rect 27672 44208 27678 44220
rect 22370 44180 22376 44192
rect 12860 44152 13584 44180
rect 22331 44152 22376 44180
rect 12860 44140 12866 44152
rect 22370 44140 22376 44152
rect 22428 44140 22434 44192
rect 29380 44189 29408 44220
rect 29822 44208 29828 44260
rect 29880 44248 29886 44260
rect 30377 44251 30435 44257
rect 30377 44248 30389 44251
rect 29880 44220 30389 44248
rect 29880 44208 29886 44220
rect 30377 44217 30389 44220
rect 30423 44248 30435 44251
rect 31110 44248 31116 44260
rect 30423 44220 31116 44248
rect 30423 44217 30435 44220
rect 30377 44211 30435 44217
rect 31110 44208 31116 44220
rect 31168 44208 31174 44260
rect 29365 44183 29423 44189
rect 29365 44149 29377 44183
rect 29411 44149 29423 44183
rect 29365 44143 29423 44149
rect 1104 44090 38824 44112
rect 1104 44038 19606 44090
rect 19658 44038 19670 44090
rect 19722 44038 19734 44090
rect 19786 44038 19798 44090
rect 19850 44038 38824 44090
rect 1104 44016 38824 44038
rect 8294 43976 8300 43988
rect 8255 43948 8300 43976
rect 8294 43936 8300 43948
rect 8352 43936 8358 43988
rect 12526 43976 12532 43988
rect 12487 43948 12532 43976
rect 12526 43936 12532 43948
rect 12584 43936 12590 43988
rect 13173 43979 13231 43985
rect 13173 43945 13185 43979
rect 13219 43976 13231 43979
rect 13354 43976 13360 43988
rect 13219 43948 13360 43976
rect 13219 43945 13231 43948
rect 13173 43939 13231 43945
rect 8312 43840 8340 43936
rect 10965 43843 11023 43849
rect 10965 43840 10977 43843
rect 8312 43812 10977 43840
rect 10965 43809 10977 43812
rect 11011 43840 11023 43843
rect 11330 43840 11336 43852
rect 11011 43812 11336 43840
rect 11011 43809 11023 43812
rect 10965 43803 11023 43809
rect 11330 43800 11336 43812
rect 11388 43840 11394 43852
rect 13078 43840 13084 43852
rect 11388 43812 13084 43840
rect 11388 43800 11394 43812
rect 13078 43800 13084 43812
rect 13136 43840 13142 43852
rect 13188 43840 13216 43939
rect 13354 43936 13360 43948
rect 13412 43936 13418 43988
rect 17310 43936 17316 43988
rect 17368 43976 17374 43988
rect 17773 43979 17831 43985
rect 17773 43976 17785 43979
rect 17368 43948 17785 43976
rect 17368 43936 17374 43948
rect 17773 43945 17785 43948
rect 17819 43976 17831 43979
rect 23845 43979 23903 43985
rect 17819 43948 20852 43976
rect 17819 43945 17831 43948
rect 17773 43939 17831 43945
rect 15378 43840 15384 43852
rect 13136 43812 13216 43840
rect 15339 43812 15384 43840
rect 13136 43800 13142 43812
rect 15378 43800 15384 43812
rect 15436 43800 15442 43852
rect 16574 43800 16580 43852
rect 16632 43840 16638 43852
rect 17770 43840 17776 43852
rect 16632 43812 17776 43840
rect 16632 43800 16638 43812
rect 17770 43800 17776 43812
rect 17828 43840 17834 43852
rect 17957 43843 18015 43849
rect 17957 43840 17969 43843
rect 17828 43812 17969 43840
rect 17828 43800 17834 43812
rect 17957 43809 17969 43812
rect 18003 43809 18015 43843
rect 20824 43840 20852 43948
rect 23845 43945 23857 43979
rect 23891 43976 23903 43979
rect 24302 43976 24308 43988
rect 23891 43948 24308 43976
rect 23891 43945 23903 43948
rect 23845 43939 23903 43945
rect 24302 43936 24308 43948
rect 24360 43936 24366 43988
rect 24765 43979 24823 43985
rect 24765 43945 24777 43979
rect 24811 43976 24823 43979
rect 24854 43976 24860 43988
rect 24811 43948 24860 43976
rect 24811 43945 24823 43948
rect 24765 43939 24823 43945
rect 24854 43936 24860 43948
rect 24912 43936 24918 43988
rect 25958 43976 25964 43988
rect 25919 43948 25964 43976
rect 25958 43936 25964 43948
rect 26016 43936 26022 43988
rect 26326 43976 26332 43988
rect 26287 43948 26332 43976
rect 26326 43936 26332 43948
rect 26384 43936 26390 43988
rect 26602 43976 26608 43988
rect 26563 43948 26608 43976
rect 26602 43936 26608 43948
rect 26660 43936 26666 43988
rect 27982 43976 27988 43988
rect 27943 43948 27988 43976
rect 27982 43936 27988 43948
rect 28040 43936 28046 43988
rect 29362 43936 29368 43988
rect 29420 43976 29426 43988
rect 29641 43979 29699 43985
rect 29641 43976 29653 43979
rect 29420 43948 29653 43976
rect 29420 43936 29426 43948
rect 29641 43945 29653 43948
rect 29687 43945 29699 43979
rect 36078 43976 36084 43988
rect 36039 43948 36084 43976
rect 29641 43939 29699 43945
rect 36078 43936 36084 43948
rect 36136 43936 36142 43988
rect 28902 43868 28908 43920
rect 28960 43908 28966 43920
rect 30009 43911 30067 43917
rect 30009 43908 30021 43911
rect 28960 43880 30021 43908
rect 28960 43868 28966 43880
rect 30009 43877 30021 43880
rect 30055 43877 30067 43911
rect 30009 43871 30067 43877
rect 20898 43840 20904 43852
rect 20811 43812 20904 43840
rect 17957 43803 18015 43809
rect 20898 43800 20904 43812
rect 20956 43800 20962 43852
rect 23661 43843 23719 43849
rect 23661 43809 23673 43843
rect 23707 43840 23719 43843
rect 23842 43840 23848 43852
rect 23707 43812 23848 43840
rect 23707 43809 23719 43812
rect 23661 43803 23719 43809
rect 23842 43800 23848 43812
rect 23900 43800 23906 43852
rect 24210 43840 24216 43852
rect 24123 43812 24216 43840
rect 24210 43800 24216 43812
rect 24268 43840 24274 43852
rect 24857 43843 24915 43849
rect 24857 43840 24869 43843
rect 24268 43812 24869 43840
rect 24268 43800 24274 43812
rect 24857 43809 24869 43812
rect 24903 43809 24915 43843
rect 25222 43840 25228 43852
rect 25183 43812 25228 43840
rect 24857 43803 24915 43809
rect 25222 43800 25228 43812
rect 25280 43840 25286 43852
rect 25590 43840 25596 43852
rect 25280 43812 25596 43840
rect 25280 43800 25286 43812
rect 25590 43800 25596 43812
rect 25648 43800 25654 43852
rect 26510 43840 26516 43852
rect 26471 43812 26516 43840
rect 26510 43800 26516 43812
rect 26568 43800 26574 43852
rect 27065 43843 27123 43849
rect 27065 43809 27077 43843
rect 27111 43840 27123 43843
rect 27338 43840 27344 43852
rect 27111 43812 27344 43840
rect 27111 43809 27123 43812
rect 27065 43803 27123 43809
rect 27338 43800 27344 43812
rect 27396 43800 27402 43852
rect 27522 43800 27528 43852
rect 27580 43840 27586 43852
rect 27982 43840 27988 43852
rect 27580 43812 27988 43840
rect 27580 43800 27586 43812
rect 27982 43800 27988 43812
rect 28040 43800 28046 43852
rect 28350 43840 28356 43852
rect 28311 43812 28356 43840
rect 28350 43800 28356 43812
rect 28408 43800 28414 43852
rect 28994 43800 29000 43852
rect 29052 43840 29058 43852
rect 29181 43843 29239 43849
rect 29181 43840 29193 43843
rect 29052 43812 29193 43840
rect 29052 43800 29058 43812
rect 29181 43809 29193 43812
rect 29227 43840 29239 43843
rect 29454 43840 29460 43852
rect 29227 43812 29460 43840
rect 29227 43809 29239 43812
rect 29181 43803 29239 43809
rect 29454 43800 29460 43812
rect 29512 43800 29518 43852
rect 29914 43800 29920 43852
rect 29972 43840 29978 43852
rect 30193 43843 30251 43849
rect 30193 43840 30205 43843
rect 29972 43812 30205 43840
rect 29972 43800 29978 43812
rect 30193 43809 30205 43812
rect 30239 43809 30251 43843
rect 30193 43803 30251 43809
rect 11146 43732 11152 43784
rect 11204 43772 11210 43784
rect 11241 43775 11299 43781
rect 11241 43772 11253 43775
rect 11204 43744 11253 43772
rect 11204 43732 11210 43744
rect 11241 43741 11253 43744
rect 11287 43772 11299 43775
rect 12250 43772 12256 43784
rect 11287 43744 12256 43772
rect 11287 43741 11299 43744
rect 11241 43735 11299 43741
rect 12250 43732 12256 43744
rect 12308 43732 12314 43784
rect 15286 43772 15292 43784
rect 15247 43744 15292 43772
rect 15286 43732 15292 43744
rect 15344 43732 15350 43784
rect 21174 43772 21180 43784
rect 21135 43744 21180 43772
rect 21174 43732 21180 43744
rect 21232 43732 21238 43784
rect 28445 43775 28503 43781
rect 28445 43741 28457 43775
rect 28491 43772 28503 43775
rect 28626 43772 28632 43784
rect 28491 43744 28632 43772
rect 28491 43741 28503 43744
rect 28445 43735 28503 43741
rect 28626 43732 28632 43744
rect 28684 43732 28690 43784
rect 29270 43772 29276 43784
rect 29231 43744 29276 43772
rect 29270 43732 29276 43744
rect 29328 43732 29334 43784
rect 29546 43732 29552 43784
rect 29604 43772 29610 43784
rect 30653 43775 30711 43781
rect 30653 43772 30665 43775
rect 29604 43744 30665 43772
rect 29604 43732 29610 43744
rect 30653 43741 30665 43744
rect 30699 43741 30711 43775
rect 30653 43735 30711 43741
rect 23566 43704 23572 43716
rect 23479 43676 23572 43704
rect 23566 43664 23572 43676
rect 23624 43704 23630 43716
rect 25038 43704 25044 43716
rect 23624 43676 25044 43704
rect 23624 43664 23630 43676
rect 25038 43664 25044 43676
rect 25096 43664 25102 43716
rect 27430 43664 27436 43716
rect 27488 43704 27494 43716
rect 27617 43707 27675 43713
rect 27617 43704 27629 43707
rect 27488 43676 27629 43704
rect 27488 43664 27494 43676
rect 27617 43673 27629 43676
rect 27663 43704 27675 43707
rect 29914 43704 29920 43716
rect 27663 43676 29920 43704
rect 27663 43673 27675 43676
rect 27617 43667 27675 43673
rect 29914 43664 29920 43676
rect 29972 43664 29978 43716
rect 15102 43596 15108 43648
rect 15160 43636 15166 43648
rect 15565 43639 15623 43645
rect 15565 43636 15577 43639
rect 15160 43608 15577 43636
rect 15160 43596 15166 43608
rect 15565 43605 15577 43608
rect 15611 43605 15623 43639
rect 15565 43599 15623 43605
rect 22002 43596 22008 43648
rect 22060 43636 22066 43648
rect 22281 43639 22339 43645
rect 22281 43636 22293 43639
rect 22060 43608 22293 43636
rect 22060 43596 22066 43608
rect 22281 43605 22293 43608
rect 22327 43605 22339 43639
rect 30374 43636 30380 43648
rect 30335 43608 30380 43636
rect 22281 43599 22339 43605
rect 30374 43596 30380 43608
rect 30432 43596 30438 43648
rect 1104 43546 38824 43568
rect 1104 43494 4246 43546
rect 4298 43494 4310 43546
rect 4362 43494 4374 43546
rect 4426 43494 4438 43546
rect 4490 43494 34966 43546
rect 35018 43494 35030 43546
rect 35082 43494 35094 43546
rect 35146 43494 35158 43546
rect 35210 43494 38824 43546
rect 1104 43472 38824 43494
rect 11057 43435 11115 43441
rect 11057 43401 11069 43435
rect 11103 43432 11115 43435
rect 11146 43432 11152 43444
rect 11103 43404 11152 43432
rect 11103 43401 11115 43404
rect 11057 43395 11115 43401
rect 11146 43392 11152 43404
rect 11204 43392 11210 43444
rect 11330 43432 11336 43444
rect 11291 43404 11336 43432
rect 11330 43392 11336 43404
rect 11388 43392 11394 43444
rect 15286 43432 15292 43444
rect 15247 43404 15292 43432
rect 15286 43392 15292 43404
rect 15344 43392 15350 43444
rect 17770 43432 17776 43444
rect 17731 43404 17776 43432
rect 17770 43392 17776 43404
rect 17828 43392 17834 43444
rect 20993 43435 21051 43441
rect 20993 43401 21005 43435
rect 21039 43432 21051 43435
rect 21174 43432 21180 43444
rect 21039 43404 21180 43432
rect 21039 43401 21051 43404
rect 20993 43395 21051 43401
rect 21174 43392 21180 43404
rect 21232 43392 21238 43444
rect 27890 43432 27896 43444
rect 27851 43404 27896 43432
rect 27890 43392 27896 43404
rect 27948 43392 27954 43444
rect 28074 43392 28080 43444
rect 28132 43432 28138 43444
rect 28261 43435 28319 43441
rect 28261 43432 28273 43435
rect 28132 43404 28273 43432
rect 28132 43392 28138 43404
rect 28261 43401 28273 43404
rect 28307 43401 28319 43435
rect 28261 43395 28319 43401
rect 20898 43324 20904 43376
rect 20956 43364 20962 43376
rect 21269 43367 21327 43373
rect 21269 43364 21281 43367
rect 20956 43336 21281 43364
rect 20956 43324 20962 43336
rect 21269 43333 21281 43336
rect 21315 43364 21327 43367
rect 21358 43364 21364 43376
rect 21315 43336 21364 43364
rect 21315 43333 21327 43336
rect 21269 43327 21327 43333
rect 21358 43324 21364 43336
rect 21416 43324 21422 43376
rect 24397 43367 24455 43373
rect 24397 43333 24409 43367
rect 24443 43364 24455 43367
rect 28276 43364 28304 43395
rect 28350 43392 28356 43444
rect 28408 43432 28414 43444
rect 28629 43435 28687 43441
rect 28629 43432 28641 43435
rect 28408 43404 28641 43432
rect 28408 43392 28414 43404
rect 28629 43401 28641 43404
rect 28675 43432 28687 43435
rect 29178 43432 29184 43444
rect 28675 43404 29184 43432
rect 28675 43401 28687 43404
rect 28629 43395 28687 43401
rect 29178 43392 29184 43404
rect 29236 43392 29242 43444
rect 29914 43392 29920 43444
rect 29972 43432 29978 43444
rect 30653 43435 30711 43441
rect 30653 43432 30665 43435
rect 29972 43404 30665 43432
rect 29972 43392 29978 43404
rect 30653 43401 30665 43404
rect 30699 43401 30711 43435
rect 30653 43395 30711 43401
rect 28997 43367 29055 43373
rect 28997 43364 29009 43367
rect 24443 43336 25544 43364
rect 28276 43336 29009 43364
rect 24443 43333 24455 43336
rect 24397 43327 24455 43333
rect 25516 43308 25544 43336
rect 28997 43333 29009 43336
rect 29043 43364 29055 43367
rect 29270 43364 29276 43376
rect 29043 43336 29276 43364
rect 29043 43333 29055 43336
rect 28997 43327 29055 43333
rect 29270 43324 29276 43336
rect 29328 43364 29334 43376
rect 30374 43364 30380 43376
rect 29328 43336 30380 43364
rect 29328 43324 29334 43336
rect 13078 43296 13084 43308
rect 13039 43268 13084 43296
rect 13078 43256 13084 43268
rect 13136 43256 13142 43308
rect 14737 43299 14795 43305
rect 14737 43265 14749 43299
rect 14783 43296 14795 43299
rect 15378 43296 15384 43308
rect 14783 43268 15384 43296
rect 14783 43265 14795 43268
rect 14737 43259 14795 43265
rect 15378 43256 15384 43268
rect 15436 43296 15442 43308
rect 15657 43299 15715 43305
rect 15657 43296 15669 43299
rect 15436 43268 15669 43296
rect 15436 43256 15442 43268
rect 15657 43265 15669 43268
rect 15703 43265 15715 43299
rect 15657 43259 15715 43265
rect 24486 43256 24492 43308
rect 24544 43296 24550 43308
rect 24581 43299 24639 43305
rect 24581 43296 24593 43299
rect 24544 43268 24593 43296
rect 24544 43256 24550 43268
rect 24581 43265 24593 43268
rect 24627 43296 24639 43299
rect 24670 43296 24676 43308
rect 24627 43268 24676 43296
rect 24627 43265 24639 43268
rect 24581 43259 24639 43265
rect 24670 43256 24676 43268
rect 24728 43256 24734 43308
rect 25498 43296 25504 43308
rect 25459 43268 25504 43296
rect 25498 43256 25504 43268
rect 25556 43256 25562 43308
rect 25961 43299 26019 43305
rect 25961 43265 25973 43299
rect 26007 43296 26019 43299
rect 26694 43296 26700 43308
rect 26007 43268 26700 43296
rect 26007 43265 26019 43268
rect 25961 43259 26019 43265
rect 26694 43256 26700 43268
rect 26752 43296 26758 43308
rect 27430 43296 27436 43308
rect 26752 43268 27436 43296
rect 26752 43256 26758 43268
rect 27430 43256 27436 43268
rect 27488 43256 27494 43308
rect 29362 43296 29368 43308
rect 29323 43268 29368 43296
rect 29362 43256 29368 43268
rect 29420 43256 29426 43308
rect 30300 43305 30328 43336
rect 30374 43324 30380 43336
rect 30432 43324 30438 43376
rect 30285 43299 30343 43305
rect 30285 43265 30297 43299
rect 30331 43265 30343 43299
rect 30285 43259 30343 43265
rect 13357 43231 13415 43237
rect 13357 43228 13369 43231
rect 12912 43200 13369 43228
rect 12618 43052 12624 43104
rect 12676 43092 12682 43104
rect 12912 43101 12940 43200
rect 13357 43197 13369 43200
rect 13403 43228 13415 43231
rect 14090 43228 14096 43240
rect 13403 43200 14096 43228
rect 13403 43197 13415 43200
rect 13357 43191 13415 43197
rect 14090 43188 14096 43200
rect 14148 43188 14154 43240
rect 25130 43188 25136 43240
rect 25188 43228 25194 43240
rect 25409 43231 25467 43237
rect 25409 43228 25421 43231
rect 25188 43200 25421 43228
rect 25188 43188 25194 43200
rect 25409 43197 25421 43200
rect 25455 43197 25467 43231
rect 25409 43191 25467 43197
rect 26326 43188 26332 43240
rect 26384 43228 26390 43240
rect 26513 43231 26571 43237
rect 26513 43228 26525 43231
rect 26384 43200 26525 43228
rect 26384 43188 26390 43200
rect 26513 43197 26525 43200
rect 26559 43197 26571 43231
rect 26513 43191 26571 43197
rect 27154 43188 27160 43240
rect 27212 43228 27218 43240
rect 27341 43231 27399 43237
rect 27341 43228 27353 43231
rect 27212 43200 27353 43228
rect 27212 43188 27218 43200
rect 27341 43197 27353 43200
rect 27387 43197 27399 43231
rect 27341 43191 27399 43197
rect 29730 43188 29736 43240
rect 29788 43228 29794 43240
rect 30193 43231 30251 43237
rect 30193 43228 30205 43231
rect 29788 43200 30205 43228
rect 29788 43188 29794 43200
rect 30193 43197 30205 43200
rect 30239 43197 30251 43231
rect 30193 43191 30251 43197
rect 24670 43160 24676 43172
rect 24631 43132 24676 43160
rect 24670 43120 24676 43132
rect 24728 43120 24734 43172
rect 26605 43163 26663 43169
rect 26605 43129 26617 43163
rect 26651 43160 26663 43163
rect 27062 43160 27068 43172
rect 26651 43132 27068 43160
rect 26651 43129 26663 43132
rect 26605 43123 26663 43129
rect 27062 43120 27068 43132
rect 27120 43120 27126 43172
rect 29454 43160 29460 43172
rect 29415 43132 29460 43160
rect 29454 43120 29460 43132
rect 29512 43120 29518 43172
rect 12897 43095 12955 43101
rect 12897 43092 12909 43095
rect 12676 43064 12909 43092
rect 12676 43052 12682 43064
rect 12897 43061 12909 43064
rect 12943 43061 12955 43095
rect 23842 43092 23848 43104
rect 23803 43064 23848 43092
rect 12897 43055 12955 43061
rect 23842 43052 23848 43064
rect 23900 43052 23906 43104
rect 26329 43095 26387 43101
rect 26329 43061 26341 43095
rect 26375 43092 26387 43095
rect 26510 43092 26516 43104
rect 26375 43064 26516 43092
rect 26375 43061 26387 43064
rect 26329 43055 26387 43061
rect 26510 43052 26516 43064
rect 26568 43052 26574 43104
rect 1104 43002 38824 43024
rect 1104 42950 19606 43002
rect 19658 42950 19670 43002
rect 19722 42950 19734 43002
rect 19786 42950 19798 43002
rect 19850 42950 38824 43002
rect 1104 42928 38824 42950
rect 14090 42888 14096 42900
rect 14051 42860 14096 42888
rect 14090 42848 14096 42860
rect 14148 42888 14154 42900
rect 14734 42888 14740 42900
rect 14148 42860 14740 42888
rect 14148 42848 14154 42860
rect 14734 42848 14740 42860
rect 14792 42848 14798 42900
rect 24486 42888 24492 42900
rect 24447 42860 24492 42888
rect 24486 42848 24492 42860
rect 24544 42848 24550 42900
rect 24949 42891 25007 42897
rect 24949 42857 24961 42891
rect 24995 42888 25007 42891
rect 25130 42888 25136 42900
rect 24995 42860 25136 42888
rect 24995 42857 25007 42860
rect 24949 42851 25007 42857
rect 25130 42848 25136 42860
rect 25188 42848 25194 42900
rect 26329 42891 26387 42897
rect 26329 42857 26341 42891
rect 26375 42888 26387 42891
rect 27338 42888 27344 42900
rect 26375 42860 27344 42888
rect 26375 42857 26387 42860
rect 26329 42851 26387 42857
rect 27338 42848 27344 42860
rect 27396 42848 27402 42900
rect 28353 42891 28411 42897
rect 28353 42857 28365 42891
rect 28399 42888 28411 42891
rect 28994 42888 29000 42900
rect 28399 42860 29000 42888
rect 28399 42857 28411 42860
rect 28353 42851 28411 42857
rect 28994 42848 29000 42860
rect 29052 42848 29058 42900
rect 29086 42848 29092 42900
rect 29144 42888 29150 42900
rect 29730 42888 29736 42900
rect 29144 42860 29736 42888
rect 29144 42848 29150 42860
rect 29730 42848 29736 42860
rect 29788 42888 29794 42900
rect 29917 42891 29975 42897
rect 29917 42888 29929 42891
rect 29788 42860 29929 42888
rect 29788 42848 29794 42860
rect 29917 42857 29929 42860
rect 29963 42857 29975 42891
rect 29917 42851 29975 42857
rect 26602 42780 26608 42832
rect 26660 42820 26666 42832
rect 26660 42792 27752 42820
rect 26660 42780 26666 42792
rect 12894 42752 12900 42764
rect 12855 42724 12900 42752
rect 12894 42712 12900 42724
rect 12952 42712 12958 42764
rect 13078 42752 13084 42764
rect 13039 42724 13084 42752
rect 13078 42712 13084 42724
rect 13136 42712 13142 42764
rect 13265 42755 13323 42761
rect 13265 42721 13277 42755
rect 13311 42752 13323 42755
rect 13354 42752 13360 42764
rect 13311 42724 13360 42752
rect 13311 42721 13323 42724
rect 13265 42715 13323 42721
rect 13354 42712 13360 42724
rect 13412 42712 13418 42764
rect 14090 42712 14096 42764
rect 14148 42752 14154 42764
rect 14826 42752 14832 42764
rect 14148 42724 14832 42752
rect 14148 42712 14154 42724
rect 14826 42712 14832 42724
rect 14884 42712 14890 42764
rect 20898 42752 20904 42764
rect 20859 42724 20904 42752
rect 20898 42712 20904 42724
rect 20956 42712 20962 42764
rect 20990 42712 20996 42764
rect 21048 42752 21054 42764
rect 21177 42755 21235 42761
rect 21177 42752 21189 42755
rect 21048 42724 21189 42752
rect 21048 42712 21054 42724
rect 21177 42721 21189 42724
rect 21223 42752 21235 42755
rect 22002 42752 22008 42764
rect 21223 42724 22008 42752
rect 21223 42721 21235 42724
rect 21177 42715 21235 42721
rect 22002 42712 22008 42724
rect 22060 42712 22066 42764
rect 24118 42752 24124 42764
rect 24079 42724 24124 42752
rect 24118 42712 24124 42724
rect 24176 42712 24182 42764
rect 25774 42712 25780 42764
rect 25832 42752 25838 42764
rect 26789 42755 26847 42761
rect 26789 42752 26801 42755
rect 25832 42724 26801 42752
rect 25832 42712 25838 42724
rect 26789 42721 26801 42724
rect 26835 42752 26847 42755
rect 26970 42752 26976 42764
rect 26835 42724 26976 42752
rect 26835 42721 26847 42724
rect 26789 42715 26847 42721
rect 26970 42712 26976 42724
rect 27028 42712 27034 42764
rect 27246 42752 27252 42764
rect 27207 42724 27252 42752
rect 27246 42712 27252 42724
rect 27304 42712 27310 42764
rect 27614 42752 27620 42764
rect 27575 42724 27620 42752
rect 27614 42712 27620 42724
rect 27672 42712 27678 42764
rect 27724 42752 27752 42792
rect 28629 42755 28687 42761
rect 28629 42752 28641 42755
rect 27724 42724 28641 42752
rect 28629 42721 28641 42724
rect 28675 42752 28687 42755
rect 28994 42752 29000 42764
rect 28675 42724 29000 42752
rect 28675 42721 28687 42724
rect 28629 42715 28687 42721
rect 28994 42712 29000 42724
rect 29052 42712 29058 42764
rect 29454 42752 29460 42764
rect 29415 42724 29460 42752
rect 29454 42712 29460 42724
rect 29512 42712 29518 42764
rect 33781 42755 33839 42761
rect 33781 42721 33793 42755
rect 33827 42752 33839 42755
rect 34146 42752 34152 42764
rect 33827 42724 34152 42752
rect 33827 42721 33839 42724
rect 33781 42715 33839 42721
rect 34146 42712 34152 42724
rect 34204 42712 34210 42764
rect 26697 42687 26755 42693
rect 26697 42653 26709 42687
rect 26743 42684 26755 42687
rect 27522 42684 27528 42696
rect 26743 42656 27528 42684
rect 26743 42653 26755 42656
rect 26697 42647 26755 42653
rect 27522 42644 27528 42656
rect 27580 42644 27586 42696
rect 27985 42687 28043 42693
rect 27985 42653 27997 42687
rect 28031 42684 28043 42687
rect 28534 42684 28540 42696
rect 28031 42656 28540 42684
rect 28031 42653 28043 42656
rect 27985 42647 28043 42653
rect 28534 42644 28540 42656
rect 28592 42644 28598 42696
rect 28718 42644 28724 42696
rect 28776 42684 28782 42696
rect 28776 42656 28821 42684
rect 28776 42644 28782 42656
rect 29270 42644 29276 42696
rect 29328 42684 29334 42696
rect 29549 42687 29607 42693
rect 29549 42684 29561 42687
rect 29328 42656 29561 42684
rect 29328 42644 29334 42656
rect 29549 42653 29561 42656
rect 29595 42653 29607 42687
rect 34054 42684 34060 42696
rect 34015 42656 34060 42684
rect 29549 42647 29607 42653
rect 34054 42644 34060 42656
rect 34112 42644 34118 42696
rect 35158 42684 35164 42696
rect 35119 42656 35164 42684
rect 35158 42644 35164 42656
rect 35216 42644 35222 42696
rect 12710 42616 12716 42628
rect 12671 42588 12716 42616
rect 12710 42576 12716 42588
rect 12768 42576 12774 42628
rect 19613 42551 19671 42557
rect 19613 42517 19625 42551
rect 19659 42548 19671 42551
rect 19702 42548 19708 42560
rect 19659 42520 19708 42548
rect 19659 42517 19671 42520
rect 19613 42511 19671 42517
rect 19702 42508 19708 42520
rect 19760 42548 19766 42560
rect 22281 42551 22339 42557
rect 22281 42548 22293 42551
rect 19760 42520 22293 42548
rect 19760 42508 19766 42520
rect 22281 42517 22293 42520
rect 22327 42517 22339 42551
rect 25222 42548 25228 42560
rect 25183 42520 25228 42548
rect 22281 42511 22339 42517
rect 25222 42508 25228 42520
rect 25280 42508 25286 42560
rect 25685 42551 25743 42557
rect 25685 42517 25697 42551
rect 25731 42548 25743 42551
rect 25958 42548 25964 42560
rect 25731 42520 25964 42548
rect 25731 42517 25743 42520
rect 25685 42511 25743 42517
rect 25958 42508 25964 42520
rect 26016 42508 26022 42560
rect 1104 42458 38824 42480
rect 1104 42406 4246 42458
rect 4298 42406 4310 42458
rect 4362 42406 4374 42458
rect 4426 42406 4438 42458
rect 4490 42406 34966 42458
rect 35018 42406 35030 42458
rect 35082 42406 35094 42458
rect 35146 42406 35158 42458
rect 35210 42406 38824 42458
rect 1104 42384 38824 42406
rect 12621 42347 12679 42353
rect 12621 42313 12633 42347
rect 12667 42344 12679 42347
rect 12710 42344 12716 42356
rect 12667 42316 12716 42344
rect 12667 42313 12679 42316
rect 12621 42307 12679 42313
rect 12710 42304 12716 42316
rect 12768 42344 12774 42356
rect 12986 42344 12992 42356
rect 12768 42316 12992 42344
rect 12768 42304 12774 42316
rect 12986 42304 12992 42316
rect 13044 42304 13050 42356
rect 20990 42344 20996 42356
rect 20951 42316 20996 42344
rect 20990 42304 20996 42316
rect 21048 42304 21054 42356
rect 25501 42347 25559 42353
rect 25501 42313 25513 42347
rect 25547 42344 25559 42347
rect 26970 42344 26976 42356
rect 25547 42316 26648 42344
rect 26931 42316 26976 42344
rect 25547 42313 25559 42316
rect 25501 42307 25559 42313
rect 12158 42236 12164 42288
rect 12216 42276 12222 42288
rect 13265 42279 13323 42285
rect 13265 42276 13277 42279
rect 12216 42248 13277 42276
rect 12216 42236 12222 42248
rect 13265 42245 13277 42248
rect 13311 42276 13323 42279
rect 13354 42276 13360 42288
rect 13311 42248 13360 42276
rect 13311 42245 13323 42248
rect 13265 42239 13323 42245
rect 13354 42236 13360 42248
rect 13412 42236 13418 42288
rect 14366 42276 14372 42288
rect 14327 42248 14372 42276
rect 14366 42236 14372 42248
rect 14424 42236 14430 42288
rect 20898 42236 20904 42288
rect 20956 42276 20962 42288
rect 21269 42279 21327 42285
rect 21269 42276 21281 42279
rect 20956 42248 21281 42276
rect 20956 42236 20962 42248
rect 21269 42245 21281 42248
rect 21315 42245 21327 42279
rect 21269 42239 21327 42245
rect 25682 42236 25688 42288
rect 25740 42276 25746 42288
rect 25740 42248 25820 42276
rect 25740 42236 25746 42248
rect 12986 42208 12992 42220
rect 12452 42180 12992 42208
rect 12452 42149 12480 42180
rect 12986 42168 12992 42180
rect 13044 42208 13050 42220
rect 13722 42208 13728 42220
rect 13044 42180 13728 42208
rect 13044 42168 13050 42180
rect 13722 42168 13728 42180
rect 13780 42168 13786 42220
rect 15102 42208 15108 42220
rect 14568 42180 15108 42208
rect 12437 42143 12495 42149
rect 12437 42109 12449 42143
rect 12483 42109 12495 42143
rect 12437 42103 12495 42109
rect 14182 42100 14188 42152
rect 14240 42140 14246 42152
rect 14568 42149 14596 42180
rect 15102 42168 15108 42180
rect 15160 42168 15166 42220
rect 25792 42217 25820 42248
rect 26620 42217 26648 42316
rect 26970 42304 26976 42316
rect 27028 42304 27034 42356
rect 27433 42347 27491 42353
rect 27433 42313 27445 42347
rect 27479 42344 27491 42347
rect 27522 42344 27528 42356
rect 27479 42316 27528 42344
rect 27479 42313 27491 42316
rect 27433 42307 27491 42313
rect 27522 42304 27528 42316
rect 27580 42304 27586 42356
rect 28074 42344 28080 42356
rect 28035 42316 28080 42344
rect 28074 42304 28080 42316
rect 28132 42304 28138 42356
rect 28994 42344 29000 42356
rect 28955 42316 29000 42344
rect 28994 42304 29000 42316
rect 29052 42304 29058 42356
rect 29454 42344 29460 42356
rect 29415 42316 29460 42344
rect 29454 42304 29460 42316
rect 29512 42304 29518 42356
rect 34146 42344 34152 42356
rect 34107 42316 34152 42344
rect 34146 42304 34152 42316
rect 34204 42344 34210 42356
rect 34606 42344 34612 42356
rect 34204 42316 34612 42344
rect 34204 42304 34210 42316
rect 34606 42304 34612 42316
rect 34664 42304 34670 42356
rect 27709 42279 27767 42285
rect 27709 42245 27721 42279
rect 27755 42276 27767 42279
rect 27982 42276 27988 42288
rect 27755 42248 27988 42276
rect 27755 42245 27767 42248
rect 27709 42239 27767 42245
rect 27982 42236 27988 42248
rect 28040 42236 28046 42288
rect 28629 42279 28687 42285
rect 28629 42245 28641 42279
rect 28675 42276 28687 42279
rect 29270 42276 29276 42288
rect 28675 42248 29276 42276
rect 28675 42245 28687 42248
rect 28629 42239 28687 42245
rect 29270 42236 29276 42248
rect 29328 42236 29334 42288
rect 25777 42211 25835 42217
rect 25777 42177 25789 42211
rect 25823 42177 25835 42211
rect 25777 42171 25835 42177
rect 26605 42211 26663 42217
rect 26605 42177 26617 42211
rect 26651 42208 26663 42211
rect 26694 42208 26700 42220
rect 26651 42180 26700 42208
rect 26651 42177 26663 42180
rect 26605 42171 26663 42177
rect 26694 42168 26700 42180
rect 26752 42168 26758 42220
rect 14553 42143 14611 42149
rect 14553 42140 14565 42143
rect 14240 42112 14565 42140
rect 14240 42100 14246 42112
rect 14553 42109 14565 42112
rect 14599 42109 14611 42143
rect 14734 42140 14740 42152
rect 14695 42112 14740 42140
rect 14553 42103 14611 42109
rect 14734 42100 14740 42112
rect 14792 42100 14798 42152
rect 14921 42143 14979 42149
rect 14921 42109 14933 42143
rect 14967 42140 14979 42143
rect 15010 42140 15016 42152
rect 14967 42112 15016 42140
rect 14967 42109 14979 42112
rect 14921 42103 14979 42109
rect 12253 42007 12311 42013
rect 12253 41973 12265 42007
rect 12299 42004 12311 42007
rect 12894 42004 12900 42016
rect 12299 41976 12900 42004
rect 12299 41973 12311 41976
rect 12253 41967 12311 41973
rect 12894 41964 12900 41976
rect 12952 41964 12958 42016
rect 14001 42007 14059 42013
rect 14001 41973 14013 42007
rect 14047 42004 14059 42007
rect 14550 42004 14556 42016
rect 14047 41976 14556 42004
rect 14047 41973 14059 41976
rect 14001 41967 14059 41973
rect 14550 41964 14556 41976
rect 14608 42004 14614 42016
rect 14936 42004 14964 42103
rect 15010 42100 15016 42112
rect 15068 42100 15074 42152
rect 19521 42143 19579 42149
rect 19521 42140 19533 42143
rect 19076 42112 19533 42140
rect 19076 42016 19104 42112
rect 19521 42109 19533 42112
rect 19567 42109 19579 42143
rect 19702 42140 19708 42152
rect 19663 42112 19708 42140
rect 19521 42103 19579 42109
rect 19702 42100 19708 42112
rect 19760 42100 19766 42152
rect 19797 42143 19855 42149
rect 19797 42109 19809 42143
rect 19843 42109 19855 42143
rect 19797 42103 19855 42109
rect 24029 42143 24087 42149
rect 24029 42109 24041 42143
rect 24075 42109 24087 42143
rect 24029 42103 24087 42109
rect 19058 42004 19064 42016
rect 14608 41976 14964 42004
rect 19019 41976 19064 42004
rect 14608 41964 14614 41976
rect 19058 41964 19064 41976
rect 19116 41964 19122 42016
rect 19334 42004 19340 42016
rect 19295 41976 19340 42004
rect 19334 41964 19340 41976
rect 19392 42004 19398 42016
rect 19812 42004 19840 42103
rect 20257 42075 20315 42081
rect 20257 42041 20269 42075
rect 20303 42072 20315 42075
rect 20438 42072 20444 42084
rect 20303 42044 20444 42072
rect 20303 42041 20315 42044
rect 20257 42035 20315 42041
rect 20438 42032 20444 42044
rect 20496 42032 20502 42084
rect 23937 42075 23995 42081
rect 23937 42041 23949 42075
rect 23983 42072 23995 42075
rect 24044 42072 24072 42103
rect 24118 42100 24124 42152
rect 24176 42140 24182 42152
rect 24489 42143 24547 42149
rect 24489 42140 24501 42143
rect 24176 42112 24501 42140
rect 24176 42100 24182 42112
rect 24489 42109 24501 42112
rect 24535 42109 24547 42143
rect 25682 42140 25688 42152
rect 25643 42112 25688 42140
rect 24489 42103 24547 42109
rect 25682 42100 25688 42112
rect 25740 42100 25746 42152
rect 25958 42100 25964 42152
rect 26016 42140 26022 42152
rect 26513 42143 26571 42149
rect 26513 42140 26525 42143
rect 26016 42112 26525 42140
rect 26016 42100 26022 42112
rect 26513 42109 26525 42112
rect 26559 42109 26571 42143
rect 26513 42103 26571 42109
rect 27525 42143 27583 42149
rect 27525 42109 27537 42143
rect 27571 42140 27583 42143
rect 28074 42140 28080 42152
rect 27571 42112 28080 42140
rect 27571 42109 27583 42112
rect 27525 42103 27583 42109
rect 26528 42072 26556 42103
rect 28074 42100 28080 42112
rect 28132 42100 28138 42152
rect 28166 42072 28172 42084
rect 23983 42044 24440 42072
rect 26528 42044 28172 42072
rect 23983 42041 23995 42044
rect 23937 42035 23995 42041
rect 24302 42004 24308 42016
rect 19392 41976 19840 42004
rect 24263 41976 24308 42004
rect 19392 41964 19398 41976
rect 24302 41964 24308 41976
rect 24360 41964 24366 42016
rect 24412 42004 24440 42044
rect 28166 42032 28172 42044
rect 28224 42032 28230 42084
rect 26602 42004 26608 42016
rect 24412 41976 26608 42004
rect 26602 41964 26608 41976
rect 26660 41964 26666 42016
rect 28074 41964 28080 42016
rect 28132 42004 28138 42016
rect 28258 42004 28264 42016
rect 28132 41976 28264 42004
rect 28132 41964 28138 41976
rect 28258 41964 28264 41976
rect 28316 41964 28322 42016
rect 33873 42007 33931 42013
rect 33873 41973 33885 42007
rect 33919 42004 33931 42007
rect 34054 42004 34060 42016
rect 33919 41976 34060 42004
rect 33919 41973 33931 41976
rect 33873 41967 33931 41973
rect 34054 41964 34060 41976
rect 34112 41964 34118 42016
rect 1104 41914 38824 41936
rect 1104 41862 19606 41914
rect 19658 41862 19670 41914
rect 19722 41862 19734 41914
rect 19786 41862 19798 41914
rect 19850 41862 38824 41914
rect 1104 41840 38824 41862
rect 12434 41760 12440 41812
rect 12492 41800 12498 41812
rect 12529 41803 12587 41809
rect 12529 41800 12541 41803
rect 12492 41772 12541 41800
rect 12492 41760 12498 41772
rect 12529 41769 12541 41772
rect 12575 41800 12587 41803
rect 13078 41800 13084 41812
rect 12575 41772 13084 41800
rect 12575 41769 12587 41772
rect 12529 41763 12587 41769
rect 13078 41760 13084 41772
rect 13136 41760 13142 41812
rect 14182 41800 14188 41812
rect 14143 41772 14188 41800
rect 14182 41760 14188 41772
rect 14240 41760 14246 41812
rect 20898 41760 20904 41812
rect 20956 41800 20962 41812
rect 21085 41803 21143 41809
rect 21085 41800 21097 41803
rect 20956 41772 21097 41800
rect 20956 41760 20962 41772
rect 21085 41769 21097 41772
rect 21131 41769 21143 41803
rect 21085 41763 21143 41769
rect 24210 41760 24216 41812
rect 24268 41800 24274 41812
rect 25593 41803 25651 41809
rect 25593 41800 25605 41803
rect 24268 41772 25605 41800
rect 24268 41760 24274 41772
rect 25593 41769 25605 41772
rect 25639 41800 25651 41803
rect 25682 41800 25688 41812
rect 25639 41772 25688 41800
rect 25639 41769 25651 41772
rect 25593 41763 25651 41769
rect 25682 41760 25688 41772
rect 25740 41760 25746 41812
rect 26789 41803 26847 41809
rect 26789 41769 26801 41803
rect 26835 41800 26847 41803
rect 27154 41800 27160 41812
rect 26835 41772 27160 41800
rect 26835 41769 26847 41772
rect 26789 41763 26847 41769
rect 27154 41760 27160 41772
rect 27212 41760 27218 41812
rect 5718 41732 5724 41744
rect 5679 41704 5724 41732
rect 5718 41692 5724 41704
rect 5776 41692 5782 41744
rect 12894 41692 12900 41744
rect 12952 41732 12958 41744
rect 13633 41735 13691 41741
rect 13633 41732 13645 41735
rect 12952 41704 13645 41732
rect 12952 41692 12958 41704
rect 13633 41701 13645 41704
rect 13679 41701 13691 41735
rect 13633 41695 13691 41701
rect 4154 41624 4160 41676
rect 4212 41664 4218 41676
rect 4341 41667 4399 41673
rect 4341 41664 4353 41667
rect 4212 41636 4353 41664
rect 4212 41624 4218 41636
rect 4341 41633 4353 41636
rect 4387 41633 4399 41667
rect 4341 41627 4399 41633
rect 13173 41667 13231 41673
rect 13173 41633 13185 41667
rect 13219 41664 13231 41667
rect 13446 41664 13452 41676
rect 13219 41636 13452 41664
rect 13219 41633 13231 41636
rect 13173 41627 13231 41633
rect 13446 41624 13452 41636
rect 13504 41624 13510 41676
rect 19886 41664 19892 41676
rect 19847 41636 19892 41664
rect 19886 41624 19892 41636
rect 19944 41624 19950 41676
rect 23477 41667 23535 41673
rect 23477 41633 23489 41667
rect 23523 41664 23535 41667
rect 23566 41664 23572 41676
rect 23523 41636 23572 41664
rect 23523 41633 23535 41636
rect 23477 41627 23535 41633
rect 23566 41624 23572 41636
rect 23624 41624 23630 41676
rect 3970 41556 3976 41608
rect 4028 41596 4034 41608
rect 4065 41599 4123 41605
rect 4065 41596 4077 41599
rect 4028 41568 4077 41596
rect 4028 41556 4034 41568
rect 4065 41565 4077 41568
rect 4111 41565 4123 41599
rect 10318 41596 10324 41608
rect 10279 41568 10324 41596
rect 4065 41559 4123 41565
rect 10318 41556 10324 41568
rect 10376 41556 10382 41608
rect 10502 41556 10508 41608
rect 10560 41596 10566 41608
rect 10597 41599 10655 41605
rect 10597 41596 10609 41599
rect 10560 41568 10609 41596
rect 10560 41556 10566 41568
rect 10597 41565 10609 41568
rect 10643 41565 10655 41599
rect 10597 41559 10655 41565
rect 12618 41556 12624 41608
rect 12676 41596 12682 41608
rect 12894 41596 12900 41608
rect 12676 41568 12900 41596
rect 12676 41556 12682 41568
rect 12894 41556 12900 41568
rect 12952 41556 12958 41608
rect 13078 41596 13084 41608
rect 13039 41568 13084 41596
rect 13078 41556 13084 41568
rect 13136 41556 13142 41608
rect 19058 41556 19064 41608
rect 19116 41596 19122 41608
rect 19153 41599 19211 41605
rect 19153 41596 19165 41599
rect 19116 41568 19165 41596
rect 19116 41556 19122 41568
rect 19153 41565 19165 41568
rect 19199 41596 19211 41599
rect 19518 41596 19524 41608
rect 19199 41568 19524 41596
rect 19199 41565 19211 41568
rect 19153 41559 19211 41565
rect 19518 41556 19524 41568
rect 19576 41556 19582 41608
rect 23750 41596 23756 41608
rect 23711 41568 23756 41596
rect 23750 41556 23756 41568
rect 23808 41556 23814 41608
rect 27246 41596 27252 41608
rect 27207 41568 27252 41596
rect 27246 41556 27252 41568
rect 27304 41556 27310 41608
rect 27522 41596 27528 41608
rect 27483 41568 27528 41596
rect 27522 41556 27528 41568
rect 27580 41556 27586 41608
rect 28905 41599 28963 41605
rect 28905 41565 28917 41599
rect 28951 41596 28963 41599
rect 29273 41599 29331 41605
rect 29273 41596 29285 41599
rect 28951 41568 29285 41596
rect 28951 41565 28963 41568
rect 28905 41559 28963 41565
rect 29273 41565 29285 41568
rect 29319 41596 29331 41599
rect 30190 41596 30196 41608
rect 29319 41568 30196 41596
rect 29319 41565 29331 41568
rect 29273 41559 29331 41565
rect 30190 41556 30196 41568
rect 30248 41556 30254 41608
rect 11606 41420 11612 41472
rect 11664 41460 11670 41472
rect 11701 41463 11759 41469
rect 11701 41460 11713 41463
rect 11664 41432 11713 41460
rect 11664 41420 11670 41432
rect 11701 41429 11713 41432
rect 11747 41429 11759 41463
rect 11701 41423 11759 41429
rect 19426 41420 19432 41472
rect 19484 41460 19490 41472
rect 19521 41463 19579 41469
rect 19521 41460 19533 41463
rect 19484 41432 19533 41460
rect 19484 41420 19490 41432
rect 19521 41429 19533 41432
rect 19567 41429 19579 41463
rect 24854 41460 24860 41472
rect 24815 41432 24860 41460
rect 19521 41423 19579 41429
rect 24854 41420 24860 41432
rect 24912 41420 24918 41472
rect 29454 41420 29460 41472
rect 29512 41460 29518 41472
rect 30006 41460 30012 41472
rect 29512 41432 30012 41460
rect 29512 41420 29518 41432
rect 30006 41420 30012 41432
rect 30064 41420 30070 41472
rect 1104 41370 38824 41392
rect 1104 41318 4246 41370
rect 4298 41318 4310 41370
rect 4362 41318 4374 41370
rect 4426 41318 4438 41370
rect 4490 41318 34966 41370
rect 35018 41318 35030 41370
rect 35082 41318 35094 41370
rect 35146 41318 35158 41370
rect 35210 41318 38824 41370
rect 1104 41296 38824 41318
rect 10413 41259 10471 41265
rect 10413 41225 10425 41259
rect 10459 41256 10471 41259
rect 10502 41256 10508 41268
rect 10459 41228 10508 41256
rect 10459 41225 10471 41228
rect 10413 41219 10471 41225
rect 10502 41216 10508 41228
rect 10560 41216 10566 41268
rect 23750 41216 23756 41268
rect 23808 41256 23814 41268
rect 23845 41259 23903 41265
rect 23845 41256 23857 41259
rect 23808 41228 23857 41256
rect 23808 41216 23814 41228
rect 23845 41225 23857 41228
rect 23891 41225 23903 41259
rect 23845 41219 23903 41225
rect 27341 41259 27399 41265
rect 27341 41225 27353 41259
rect 27387 41256 27399 41259
rect 27522 41256 27528 41268
rect 27387 41228 27528 41256
rect 27387 41225 27399 41228
rect 27341 41219 27399 41225
rect 27522 41216 27528 41228
rect 27580 41216 27586 41268
rect 27706 41256 27712 41268
rect 27667 41228 27712 41256
rect 27706 41216 27712 41228
rect 27764 41216 27770 41268
rect 29089 41259 29147 41265
rect 29089 41225 29101 41259
rect 29135 41256 29147 41259
rect 29178 41256 29184 41268
rect 29135 41228 29184 41256
rect 29135 41225 29147 41228
rect 29089 41219 29147 41225
rect 29178 41216 29184 41228
rect 29236 41216 29242 41268
rect 34698 41216 34704 41268
rect 34756 41216 34762 41268
rect 19245 41191 19303 41197
rect 19245 41157 19257 41191
rect 19291 41188 19303 41191
rect 19886 41188 19892 41200
rect 19291 41160 19892 41188
rect 19291 41157 19303 41160
rect 19245 41151 19303 41157
rect 19886 41148 19892 41160
rect 19944 41148 19950 41200
rect 23566 41148 23572 41200
rect 23624 41188 23630 41200
rect 24213 41191 24271 41197
rect 24213 41188 24225 41191
rect 23624 41160 24225 41188
rect 23624 41148 23630 41160
rect 24213 41157 24225 41160
rect 24259 41157 24271 41191
rect 24213 41151 24271 41157
rect 18601 41123 18659 41129
rect 18601 41120 18613 41123
rect 18064 41092 18613 41120
rect 18064 41061 18092 41092
rect 18601 41089 18613 41092
rect 18647 41120 18659 41123
rect 19613 41123 19671 41129
rect 19613 41120 19625 41123
rect 18647 41092 19625 41120
rect 18647 41089 18659 41092
rect 18601 41083 18659 41089
rect 19613 41089 19625 41092
rect 19659 41089 19671 41123
rect 19613 41083 19671 41089
rect 20993 41123 21051 41129
rect 20993 41089 21005 41123
rect 21039 41120 21051 41123
rect 29196 41120 29224 41216
rect 34716 41188 34744 41216
rect 34882 41188 34888 41200
rect 34716 41160 34888 41188
rect 34882 41148 34888 41160
rect 34940 41148 34946 41200
rect 29365 41123 29423 41129
rect 29365 41120 29377 41123
rect 21039 41092 21404 41120
rect 29196 41092 29377 41120
rect 21039 41089 21051 41092
rect 20993 41083 21051 41089
rect 21376 41064 21404 41092
rect 29365 41089 29377 41092
rect 29411 41089 29423 41123
rect 29365 41083 29423 41089
rect 30006 41080 30012 41132
rect 30064 41120 30070 41132
rect 30285 41123 30343 41129
rect 30285 41120 30297 41123
rect 30064 41092 30297 41120
rect 30064 41080 30070 41092
rect 30285 41089 30297 41092
rect 30331 41089 30343 41123
rect 30285 41083 30343 41089
rect 18049 41055 18107 41061
rect 18049 41021 18061 41055
rect 18095 41021 18107 41055
rect 19153 41055 19211 41061
rect 19153 41052 19165 41055
rect 18049 41015 18107 41021
rect 18984 41024 19165 41052
rect 3970 40944 3976 40996
rect 4028 40984 4034 40996
rect 4433 40987 4491 40993
rect 4433 40984 4445 40987
rect 4028 40956 4445 40984
rect 4028 40944 4034 40956
rect 4433 40953 4445 40956
rect 4479 40953 4491 40987
rect 4433 40947 4491 40953
rect 13078 40944 13084 40996
rect 13136 40984 13142 40996
rect 13173 40987 13231 40993
rect 13173 40984 13185 40987
rect 13136 40956 13185 40984
rect 13136 40944 13142 40956
rect 13173 40953 13185 40956
rect 13219 40984 13231 40987
rect 13814 40984 13820 40996
rect 13219 40956 13820 40984
rect 13219 40953 13231 40956
rect 13173 40947 13231 40953
rect 13814 40944 13820 40956
rect 13872 40944 13878 40996
rect 18984 40928 19012 41024
rect 19153 41021 19165 41024
rect 19199 41052 19211 41055
rect 19334 41052 19340 41064
rect 19199 41024 19340 41052
rect 19199 41021 19211 41024
rect 19153 41015 19211 41021
rect 19334 41012 19340 41024
rect 19392 41012 19398 41064
rect 19429 41055 19487 41061
rect 19429 41021 19441 41055
rect 19475 41021 19487 41055
rect 19429 41015 19487 41021
rect 19444 40984 19472 41015
rect 19886 41012 19892 41064
rect 19944 41052 19950 41064
rect 20257 41055 20315 41061
rect 20257 41052 20269 41055
rect 19944 41024 20269 41052
rect 19944 41012 19950 41024
rect 20257 41021 20269 41024
rect 20303 41052 20315 41055
rect 20533 41055 20591 41061
rect 20533 41052 20545 41055
rect 20303 41024 20545 41052
rect 20303 41021 20315 41024
rect 20257 41015 20315 41021
rect 20533 41021 20545 41024
rect 20579 41021 20591 41055
rect 20533 41015 20591 41021
rect 20898 41012 20904 41064
rect 20956 41052 20962 41064
rect 21085 41055 21143 41061
rect 21085 41052 21097 41055
rect 20956 41024 21097 41052
rect 20956 41012 20962 41024
rect 21085 41021 21097 41024
rect 21131 41052 21143 41055
rect 21174 41052 21180 41064
rect 21131 41024 21180 41052
rect 21131 41021 21143 41024
rect 21085 41015 21143 41021
rect 21174 41012 21180 41024
rect 21232 41012 21238 41064
rect 21358 41052 21364 41064
rect 21319 41024 21364 41052
rect 21358 41012 21364 41024
rect 21416 41012 21422 41064
rect 30190 41052 30196 41064
rect 30151 41024 30196 41052
rect 30190 41012 30196 41024
rect 30248 41012 30254 41064
rect 19518 40984 19524 40996
rect 19431 40956 19524 40984
rect 19518 40944 19524 40956
rect 19576 40984 19582 40996
rect 29457 40987 29515 40993
rect 19576 40956 20300 40984
rect 19576 40944 19582 40956
rect 20272 40928 20300 40956
rect 29457 40953 29469 40987
rect 29503 40984 29515 40987
rect 29638 40984 29644 40996
rect 29503 40956 29644 40984
rect 29503 40953 29515 40956
rect 29457 40947 29515 40953
rect 29638 40944 29644 40956
rect 29696 40944 29702 40996
rect 4062 40916 4068 40928
rect 4023 40888 4068 40916
rect 4062 40876 4068 40888
rect 4120 40876 4126 40928
rect 10318 40876 10324 40928
rect 10376 40916 10382 40928
rect 10781 40919 10839 40925
rect 10781 40916 10793 40919
rect 10376 40888 10793 40916
rect 10376 40876 10382 40888
rect 10781 40885 10793 40888
rect 10827 40916 10839 40919
rect 11330 40916 11336 40928
rect 10827 40888 11336 40916
rect 10827 40885 10839 40888
rect 10781 40879 10839 40885
rect 11330 40876 11336 40888
rect 11388 40876 11394 40928
rect 13446 40916 13452 40928
rect 13407 40888 13452 40916
rect 13446 40876 13452 40888
rect 13504 40876 13510 40928
rect 18230 40916 18236 40928
rect 18191 40888 18236 40916
rect 18230 40876 18236 40888
rect 18288 40876 18294 40928
rect 18966 40916 18972 40928
rect 18927 40888 18972 40916
rect 18966 40876 18972 40888
rect 19024 40876 19030 40928
rect 20254 40876 20260 40928
rect 20312 40876 20318 40928
rect 22462 40916 22468 40928
rect 22423 40888 22468 40916
rect 22462 40876 22468 40888
rect 22520 40876 22526 40928
rect 1104 40826 38824 40848
rect 1104 40774 19606 40826
rect 19658 40774 19670 40826
rect 19722 40774 19734 40826
rect 19786 40774 19798 40826
rect 19850 40774 38824 40826
rect 1104 40752 38824 40774
rect 20714 40672 20720 40724
rect 20772 40712 20778 40724
rect 21085 40715 21143 40721
rect 21085 40712 21097 40715
rect 20772 40684 21097 40712
rect 20772 40672 20778 40684
rect 21085 40681 21097 40684
rect 21131 40681 21143 40715
rect 21085 40675 21143 40681
rect 21174 40672 21180 40724
rect 21232 40712 21238 40724
rect 21729 40715 21787 40721
rect 21729 40712 21741 40715
rect 21232 40684 21741 40712
rect 21232 40672 21238 40684
rect 21729 40681 21741 40684
rect 21775 40681 21787 40715
rect 23474 40712 23480 40724
rect 23435 40684 23480 40712
rect 21729 40675 21787 40681
rect 2406 40644 2412 40656
rect 2367 40616 2412 40644
rect 2406 40604 2412 40616
rect 2464 40604 2470 40656
rect 2961 40647 3019 40653
rect 2961 40613 2973 40647
rect 3007 40644 3019 40647
rect 4062 40644 4068 40656
rect 3007 40616 4068 40644
rect 3007 40613 3019 40616
rect 2961 40607 3019 40613
rect 4062 40604 4068 40616
rect 4120 40604 4126 40656
rect 12989 40647 13047 40653
rect 12989 40613 13001 40647
rect 13035 40644 13047 40647
rect 13446 40644 13452 40656
rect 13035 40616 13452 40644
rect 13035 40613 13047 40616
rect 12989 40607 13047 40613
rect 13446 40604 13452 40616
rect 13504 40604 13510 40656
rect 19352 40616 20116 40644
rect 19352 40588 19380 40616
rect 20088 40588 20116 40616
rect 2593 40579 2651 40585
rect 2593 40545 2605 40579
rect 2639 40545 2651 40579
rect 13814 40576 13820 40588
rect 13775 40548 13820 40576
rect 2593 40539 2651 40545
rect 2222 40468 2228 40520
rect 2280 40508 2286 40520
rect 2608 40508 2636 40539
rect 13814 40536 13820 40548
rect 13872 40536 13878 40588
rect 15930 40576 15936 40588
rect 15891 40548 15936 40576
rect 15930 40536 15936 40548
rect 15988 40536 15994 40588
rect 17681 40579 17739 40585
rect 17681 40545 17693 40579
rect 17727 40576 17739 40579
rect 17862 40576 17868 40588
rect 17727 40548 17868 40576
rect 17727 40545 17739 40548
rect 17681 40539 17739 40545
rect 17862 40536 17868 40548
rect 17920 40536 17926 40588
rect 18966 40576 18972 40588
rect 18879 40548 18972 40576
rect 18966 40536 18972 40548
rect 19024 40536 19030 40588
rect 19334 40576 19340 40588
rect 19295 40548 19340 40576
rect 19334 40536 19340 40548
rect 19392 40536 19398 40588
rect 19702 40576 19708 40588
rect 19663 40548 19708 40576
rect 19702 40536 19708 40548
rect 19760 40536 19766 40588
rect 19978 40576 19984 40588
rect 19939 40548 19984 40576
rect 19978 40536 19984 40548
rect 20036 40536 20042 40588
rect 20070 40536 20076 40588
rect 20128 40576 20134 40588
rect 20128 40548 20221 40576
rect 20128 40536 20134 40548
rect 20254 40536 20260 40588
rect 20312 40576 20318 40588
rect 20717 40579 20775 40585
rect 20312 40548 20357 40576
rect 20312 40536 20318 40548
rect 20717 40545 20729 40579
rect 20763 40576 20775 40579
rect 20901 40579 20959 40585
rect 20901 40576 20913 40579
rect 20763 40548 20913 40576
rect 20763 40545 20775 40548
rect 20717 40539 20775 40545
rect 20901 40545 20913 40548
rect 20947 40576 20959 40579
rect 21082 40576 21088 40588
rect 20947 40548 21088 40576
rect 20947 40545 20959 40548
rect 20901 40539 20959 40545
rect 21082 40536 21088 40548
rect 21140 40536 21146 40588
rect 21744 40576 21772 40675
rect 23474 40672 23480 40684
rect 23532 40672 23538 40724
rect 22097 40579 22155 40585
rect 22097 40576 22109 40579
rect 21744 40548 22109 40576
rect 22097 40545 22109 40548
rect 22143 40545 22155 40579
rect 22097 40539 22155 40545
rect 22373 40579 22431 40585
rect 22373 40545 22385 40579
rect 22419 40576 22431 40579
rect 23382 40576 23388 40588
rect 22419 40548 23388 40576
rect 22419 40545 22431 40548
rect 22373 40539 22431 40545
rect 23382 40536 23388 40548
rect 23440 40536 23446 40588
rect 34882 40536 34888 40588
rect 34940 40576 34946 40588
rect 35253 40579 35311 40585
rect 35253 40576 35265 40579
rect 34940 40548 35265 40576
rect 34940 40536 34946 40548
rect 35253 40545 35265 40548
rect 35299 40576 35311 40579
rect 35526 40576 35532 40588
rect 35299 40548 35532 40576
rect 35299 40545 35311 40548
rect 35253 40539 35311 40545
rect 35526 40536 35532 40548
rect 35584 40536 35590 40588
rect 11330 40508 11336 40520
rect 2280 40480 2636 40508
rect 11291 40480 11336 40508
rect 2280 40468 2286 40480
rect 11330 40468 11336 40480
rect 11388 40468 11394 40520
rect 11606 40508 11612 40520
rect 11567 40480 11612 40508
rect 11606 40468 11612 40480
rect 11664 40468 11670 40520
rect 17770 40508 17776 40520
rect 17731 40480 17776 40508
rect 17770 40468 17776 40480
rect 17828 40468 17834 40520
rect 18984 40508 19012 40536
rect 19996 40508 20024 40536
rect 18984 40480 20024 40508
rect 34606 40468 34612 40520
rect 34664 40508 34670 40520
rect 34977 40511 35035 40517
rect 34977 40508 34989 40511
rect 34664 40480 34989 40508
rect 34664 40468 34670 40480
rect 34977 40477 34989 40480
rect 35023 40508 35035 40511
rect 35434 40508 35440 40520
rect 35023 40480 35440 40508
rect 35023 40477 35035 40480
rect 34977 40471 35035 40477
rect 35434 40468 35440 40480
rect 35492 40468 35498 40520
rect 19702 40400 19708 40452
rect 19760 40440 19766 40452
rect 20254 40440 20260 40452
rect 19760 40412 20260 40440
rect 19760 40400 19766 40412
rect 20254 40400 20260 40412
rect 20312 40400 20318 40452
rect 1673 40375 1731 40381
rect 1673 40341 1685 40375
rect 1719 40372 1731 40375
rect 1946 40372 1952 40384
rect 1719 40344 1952 40372
rect 1719 40341 1731 40344
rect 1673 40335 1731 40341
rect 1946 40332 1952 40344
rect 2004 40332 2010 40384
rect 13998 40372 14004 40384
rect 13959 40344 14004 40372
rect 13998 40332 14004 40344
rect 14056 40332 14062 40384
rect 15194 40332 15200 40384
rect 15252 40372 15258 40384
rect 16117 40375 16175 40381
rect 16117 40372 16129 40375
rect 15252 40344 16129 40372
rect 15252 40332 15258 40344
rect 16117 40341 16129 40344
rect 16163 40341 16175 40375
rect 16117 40335 16175 40341
rect 18785 40375 18843 40381
rect 18785 40341 18797 40375
rect 18831 40372 18843 40375
rect 19334 40372 19340 40384
rect 18831 40344 19340 40372
rect 18831 40341 18843 40344
rect 18785 40335 18843 40341
rect 19334 40332 19340 40344
rect 19392 40332 19398 40384
rect 21358 40372 21364 40384
rect 21319 40344 21364 40372
rect 21358 40332 21364 40344
rect 21416 40332 21422 40384
rect 25682 40372 25688 40384
rect 25643 40344 25688 40372
rect 25682 40332 25688 40344
rect 25740 40332 25746 40384
rect 28442 40332 28448 40384
rect 28500 40372 28506 40384
rect 29273 40375 29331 40381
rect 29273 40372 29285 40375
rect 28500 40344 29285 40372
rect 28500 40332 28506 40344
rect 29273 40341 29285 40344
rect 29319 40372 29331 40375
rect 30006 40372 30012 40384
rect 29319 40344 30012 40372
rect 29319 40341 29331 40344
rect 29273 40335 29331 40341
rect 30006 40332 30012 40344
rect 30064 40332 30070 40384
rect 35710 40332 35716 40384
rect 35768 40372 35774 40384
rect 36357 40375 36415 40381
rect 36357 40372 36369 40375
rect 35768 40344 36369 40372
rect 35768 40332 35774 40344
rect 36357 40341 36369 40344
rect 36403 40341 36415 40375
rect 36357 40335 36415 40341
rect 1104 40282 38824 40304
rect 1104 40230 4246 40282
rect 4298 40230 4310 40282
rect 4362 40230 4374 40282
rect 4426 40230 4438 40282
rect 4490 40230 34966 40282
rect 35018 40230 35030 40282
rect 35082 40230 35094 40282
rect 35146 40230 35158 40282
rect 35210 40230 38824 40282
rect 1104 40208 38824 40230
rect 17126 40168 17132 40180
rect 17039 40140 17132 40168
rect 17126 40128 17132 40140
rect 17184 40168 17190 40180
rect 17862 40168 17868 40180
rect 17184 40140 17868 40168
rect 17184 40128 17190 40140
rect 17862 40128 17868 40140
rect 17920 40128 17926 40180
rect 23109 40171 23167 40177
rect 23109 40137 23121 40171
rect 23155 40168 23167 40171
rect 23382 40168 23388 40180
rect 23155 40140 23388 40168
rect 23155 40137 23167 40140
rect 23109 40131 23167 40137
rect 23382 40128 23388 40140
rect 23440 40128 23446 40180
rect 35434 40168 35440 40180
rect 35395 40140 35440 40168
rect 35434 40128 35440 40140
rect 35492 40128 35498 40180
rect 9674 40060 9680 40112
rect 9732 40100 9738 40112
rect 11330 40100 11336 40112
rect 9732 40072 11336 40100
rect 9732 40060 9738 40072
rect 11330 40060 11336 40072
rect 11388 40100 11394 40112
rect 11701 40103 11759 40109
rect 11701 40100 11713 40103
rect 11388 40072 11713 40100
rect 11388 40060 11394 40072
rect 11701 40069 11713 40072
rect 11747 40069 11759 40103
rect 11701 40063 11759 40069
rect 35161 40103 35219 40109
rect 35161 40069 35173 40103
rect 35207 40100 35219 40103
rect 35526 40100 35532 40112
rect 35207 40072 35532 40100
rect 35207 40069 35219 40072
rect 35161 40063 35219 40069
rect 35526 40060 35532 40072
rect 35584 40060 35590 40112
rect 1581 40035 1639 40041
rect 1581 40001 1593 40035
rect 1627 40032 1639 40035
rect 1946 40032 1952 40044
rect 1627 40004 1952 40032
rect 1627 40001 1639 40004
rect 1581 39995 1639 40001
rect 1946 39992 1952 40004
rect 2004 39992 2010 40044
rect 18325 40035 18383 40041
rect 18325 40001 18337 40035
rect 18371 40032 18383 40035
rect 20070 40032 20076 40044
rect 18371 40004 20076 40032
rect 18371 40001 18383 40004
rect 18325 39995 18383 40001
rect 20070 39992 20076 40004
rect 20128 40032 20134 40044
rect 20809 40035 20867 40041
rect 20809 40032 20821 40035
rect 20128 40004 20821 40032
rect 20128 39992 20134 40004
rect 20809 40001 20821 40004
rect 20855 40001 20867 40035
rect 21358 40032 21364 40044
rect 21319 40004 21364 40032
rect 20809 39995 20867 40001
rect 21358 39992 21364 40004
rect 21416 39992 21422 40044
rect 25682 39992 25688 40044
rect 25740 40032 25746 40044
rect 26145 40035 26203 40041
rect 26145 40032 26157 40035
rect 25740 40004 26157 40032
rect 25740 39992 25746 40004
rect 26145 40001 26157 40004
rect 26191 40032 26203 40035
rect 26510 40032 26516 40044
rect 26191 40004 26516 40032
rect 26191 40001 26203 40004
rect 26145 39995 26203 40001
rect 26510 39992 26516 40004
rect 26568 39992 26574 40044
rect 1670 39924 1676 39976
rect 1728 39964 1734 39976
rect 1857 39967 1915 39973
rect 1857 39964 1869 39967
rect 1728 39936 1869 39964
rect 1728 39924 1734 39936
rect 1857 39933 1869 39936
rect 1903 39933 1915 39967
rect 13078 39964 13084 39976
rect 13039 39936 13084 39964
rect 1857 39927 1915 39933
rect 13078 39924 13084 39936
rect 13136 39964 13142 39976
rect 13541 39967 13599 39973
rect 13541 39964 13553 39967
rect 13136 39936 13553 39964
rect 13136 39924 13142 39936
rect 13541 39933 13553 39936
rect 13587 39933 13599 39967
rect 13541 39927 13599 39933
rect 15565 39967 15623 39973
rect 15565 39933 15577 39967
rect 15611 39964 15623 39967
rect 15930 39964 15936 39976
rect 15611 39936 15936 39964
rect 15611 39933 15623 39936
rect 15565 39927 15623 39933
rect 15930 39924 15936 39936
rect 15988 39964 15994 39976
rect 16482 39964 16488 39976
rect 15988 39936 16488 39964
rect 15988 39924 15994 39936
rect 16482 39924 16488 39936
rect 16540 39924 16546 39976
rect 17862 39964 17868 39976
rect 17823 39936 17868 39964
rect 17862 39924 17868 39936
rect 17920 39924 17926 39976
rect 21085 39967 21143 39973
rect 21085 39933 21097 39967
rect 21131 39964 21143 39967
rect 21174 39964 21180 39976
rect 21131 39936 21180 39964
rect 21131 39933 21143 39936
rect 21085 39927 21143 39933
rect 21174 39924 21180 39936
rect 21232 39964 21238 39976
rect 23385 39967 23443 39973
rect 23385 39964 23397 39967
rect 21232 39936 23397 39964
rect 21232 39924 21238 39936
rect 23385 39933 23397 39936
rect 23431 39964 23443 39967
rect 23566 39964 23572 39976
rect 23431 39936 23572 39964
rect 23431 39933 23443 39936
rect 23385 39927 23443 39933
rect 23566 39924 23572 39936
rect 23624 39924 23630 39976
rect 25130 39964 25136 39976
rect 25043 39936 25136 39964
rect 25130 39924 25136 39936
rect 25188 39964 25194 39976
rect 26283 39967 26341 39973
rect 26283 39964 26295 39967
rect 25188 39936 26295 39964
rect 25188 39924 25194 39936
rect 26283 39933 26295 39936
rect 26329 39933 26341 39967
rect 26283 39927 26341 39933
rect 26421 39967 26479 39973
rect 26421 39933 26433 39967
rect 26467 39964 26479 39967
rect 26878 39964 26884 39976
rect 26467 39936 26884 39964
rect 26467 39933 26479 39936
rect 26421 39927 26479 39933
rect 3237 39899 3295 39905
rect 3237 39865 3249 39899
rect 3283 39896 3295 39899
rect 4062 39896 4068 39908
rect 3283 39868 4068 39896
rect 3283 39865 3295 39868
rect 3237 39859 3295 39865
rect 4062 39856 4068 39868
rect 4120 39856 4126 39908
rect 16025 39899 16083 39905
rect 16025 39865 16037 39899
rect 16071 39865 16083 39899
rect 16025 39859 16083 39865
rect 18785 39899 18843 39905
rect 18785 39865 18797 39899
rect 18831 39865 18843 39899
rect 18785 39859 18843 39865
rect 11425 39831 11483 39837
rect 11425 39797 11437 39831
rect 11471 39828 11483 39831
rect 11606 39828 11612 39840
rect 11471 39800 11612 39828
rect 11471 39797 11483 39800
rect 11425 39791 11483 39797
rect 11606 39788 11612 39800
rect 11664 39828 11670 39840
rect 12434 39828 12440 39840
rect 11664 39800 12440 39828
rect 11664 39788 11670 39800
rect 12434 39788 12440 39800
rect 12492 39788 12498 39840
rect 13265 39831 13323 39837
rect 13265 39797 13277 39831
rect 13311 39828 13323 39831
rect 13446 39828 13452 39840
rect 13311 39800 13452 39828
rect 13311 39797 13323 39800
rect 13265 39791 13323 39797
rect 13446 39788 13452 39800
rect 13504 39828 13510 39840
rect 13814 39828 13820 39840
rect 13504 39800 13820 39828
rect 13504 39788 13510 39800
rect 13814 39788 13820 39800
rect 13872 39828 13878 39840
rect 13909 39831 13967 39837
rect 13909 39828 13921 39831
rect 13872 39800 13921 39828
rect 13872 39788 13878 39800
rect 13909 39797 13921 39800
rect 13955 39797 13967 39831
rect 13909 39791 13967 39797
rect 15197 39831 15255 39837
rect 15197 39797 15209 39831
rect 15243 39828 15255 39831
rect 15470 39828 15476 39840
rect 15243 39800 15476 39828
rect 15243 39797 15255 39800
rect 15197 39791 15255 39797
rect 15470 39788 15476 39800
rect 15528 39788 15534 39840
rect 15930 39788 15936 39840
rect 15988 39828 15994 39840
rect 16040 39828 16068 39859
rect 18598 39828 18604 39840
rect 15988 39800 16068 39828
rect 18559 39800 18604 39828
rect 15988 39788 15994 39800
rect 18598 39788 18604 39800
rect 18656 39828 18662 39840
rect 18800 39828 18828 39859
rect 20346 39856 20352 39908
rect 20404 39896 20410 39908
rect 20530 39896 20536 39908
rect 20404 39868 20536 39896
rect 20404 39856 20410 39868
rect 20530 39856 20536 39868
rect 20588 39856 20594 39908
rect 25593 39899 25651 39905
rect 25593 39865 25605 39899
rect 25639 39896 25651 39899
rect 25774 39896 25780 39908
rect 25639 39868 25780 39896
rect 25639 39865 25651 39868
rect 25593 39859 25651 39865
rect 25774 39856 25780 39868
rect 25832 39856 25838 39908
rect 18656 39800 18828 39828
rect 18656 39788 18662 39800
rect 20990 39788 20996 39840
rect 21048 39828 21054 39840
rect 22465 39831 22523 39837
rect 22465 39828 22477 39831
rect 21048 39800 22477 39828
rect 21048 39788 21054 39800
rect 22465 39797 22477 39800
rect 22511 39797 22523 39831
rect 22465 39791 22523 39797
rect 25501 39831 25559 39837
rect 25501 39797 25513 39831
rect 25547 39828 25559 39831
rect 26436 39828 26464 39927
rect 26878 39924 26884 39936
rect 26936 39924 26942 39976
rect 25547 39800 26464 39828
rect 25547 39797 25559 39800
rect 25501 39791 25559 39797
rect 1104 39738 38824 39760
rect 1104 39686 19606 39738
rect 19658 39686 19670 39738
rect 19722 39686 19734 39738
rect 19786 39686 19798 39738
rect 19850 39686 38824 39738
rect 1104 39664 38824 39686
rect 2406 39584 2412 39636
rect 2464 39624 2470 39636
rect 2777 39627 2835 39633
rect 2777 39624 2789 39627
rect 2464 39596 2789 39624
rect 2464 39584 2470 39596
rect 2777 39593 2789 39596
rect 2823 39593 2835 39627
rect 19058 39624 19064 39636
rect 19019 39596 19064 39624
rect 2777 39587 2835 39593
rect 19058 39584 19064 39596
rect 19116 39584 19122 39636
rect 21082 39624 21088 39636
rect 21043 39596 21088 39624
rect 21082 39584 21088 39596
rect 21140 39584 21146 39636
rect 21358 39584 21364 39636
rect 21416 39624 21422 39636
rect 22741 39627 22799 39633
rect 22741 39624 22753 39627
rect 21416 39596 22753 39624
rect 21416 39584 21422 39596
rect 22741 39593 22753 39596
rect 22787 39593 22799 39627
rect 25130 39624 25136 39636
rect 25091 39596 25136 39624
rect 22741 39587 22799 39593
rect 25130 39584 25136 39596
rect 25188 39584 25194 39636
rect 1578 39556 1584 39568
rect 1539 39528 1584 39556
rect 1578 39516 1584 39528
rect 1636 39516 1642 39568
rect 18785 39559 18843 39565
rect 18785 39525 18797 39559
rect 18831 39556 18843 39559
rect 19978 39556 19984 39568
rect 18831 39528 19984 39556
rect 18831 39525 18843 39528
rect 18785 39519 18843 39525
rect 19978 39516 19984 39528
rect 20036 39556 20042 39568
rect 20257 39559 20315 39565
rect 20257 39556 20269 39559
rect 20036 39528 20269 39556
rect 20036 39516 20042 39528
rect 20257 39525 20269 39528
rect 20303 39525 20315 39559
rect 26510 39556 26516 39568
rect 26471 39528 26516 39556
rect 20257 39519 20315 39525
rect 26510 39516 26516 39528
rect 26568 39516 26574 39568
rect 15562 39488 15568 39500
rect 15523 39460 15568 39488
rect 15562 39448 15568 39460
rect 15620 39448 15626 39500
rect 16574 39448 16580 39500
rect 16632 39488 16638 39500
rect 17865 39491 17923 39497
rect 17865 39488 17877 39491
rect 16632 39460 17877 39488
rect 16632 39448 16638 39460
rect 17865 39457 17877 39460
rect 17911 39457 17923 39491
rect 18230 39488 18236 39500
rect 18191 39460 18236 39488
rect 17865 39451 17923 39457
rect 18230 39448 18236 39460
rect 18288 39448 18294 39500
rect 19886 39488 19892 39500
rect 19847 39460 19892 39488
rect 19886 39448 19892 39460
rect 19944 39448 19950 39500
rect 21174 39448 21180 39500
rect 21232 39488 21238 39500
rect 21361 39491 21419 39497
rect 21361 39488 21373 39491
rect 21232 39460 21373 39488
rect 21232 39448 21238 39460
rect 21361 39457 21373 39460
rect 21407 39457 21419 39491
rect 25038 39488 25044 39500
rect 24999 39460 25044 39488
rect 21361 39451 21419 39457
rect 25038 39448 25044 39460
rect 25096 39448 25102 39500
rect 26602 39488 26608 39500
rect 26563 39460 26608 39488
rect 26602 39448 26608 39460
rect 26660 39448 26666 39500
rect 35345 39491 35403 39497
rect 35345 39457 35357 39491
rect 35391 39488 35403 39491
rect 35710 39488 35716 39500
rect 35391 39460 35716 39488
rect 35391 39457 35403 39460
rect 35345 39451 35403 39457
rect 35710 39448 35716 39460
rect 35768 39448 35774 39500
rect 14182 39380 14188 39432
rect 14240 39420 14246 39432
rect 14461 39423 14519 39429
rect 14461 39420 14473 39423
rect 14240 39392 14473 39420
rect 14240 39380 14246 39392
rect 14461 39389 14473 39392
rect 14507 39389 14519 39423
rect 14461 39383 14519 39389
rect 15473 39423 15531 39429
rect 15473 39389 15485 39423
rect 15519 39389 15531 39423
rect 16022 39420 16028 39432
rect 15983 39392 16028 39420
rect 15473 39383 15531 39389
rect 13817 39355 13875 39361
rect 13817 39321 13829 39355
rect 13863 39352 13875 39355
rect 15102 39352 15108 39364
rect 13863 39324 15108 39352
rect 13863 39321 13875 39324
rect 13817 39315 13875 39321
rect 15102 39312 15108 39324
rect 15160 39312 15166 39364
rect 15488 39352 15516 39383
rect 16022 39380 16028 39392
rect 16080 39380 16086 39432
rect 16114 39380 16120 39432
rect 16172 39420 16178 39432
rect 17221 39423 17279 39429
rect 17221 39420 17233 39423
rect 16172 39392 17233 39420
rect 16172 39380 16178 39392
rect 17221 39389 17233 39392
rect 17267 39389 17279 39423
rect 17770 39420 17776 39432
rect 17731 39392 17776 39420
rect 17221 39383 17279 39389
rect 17770 39380 17776 39392
rect 17828 39380 17834 39432
rect 18325 39423 18383 39429
rect 18325 39389 18337 39423
rect 18371 39389 18383 39423
rect 18325 39383 18383 39389
rect 21637 39423 21695 39429
rect 21637 39389 21649 39423
rect 21683 39420 21695 39423
rect 21726 39420 21732 39432
rect 21683 39392 21732 39420
rect 21683 39389 21695 39392
rect 21637 39383 21695 39389
rect 16206 39352 16212 39364
rect 15488 39324 16212 39352
rect 16206 39312 16212 39324
rect 16264 39312 16270 39364
rect 17129 39355 17187 39361
rect 17129 39321 17141 39355
rect 17175 39352 17187 39355
rect 18046 39352 18052 39364
rect 17175 39324 18052 39352
rect 17175 39321 17187 39324
rect 17129 39315 17187 39321
rect 18046 39312 18052 39324
rect 18104 39352 18110 39364
rect 18340 39352 18368 39383
rect 21726 39380 21732 39392
rect 21784 39380 21790 39432
rect 34698 39420 34704 39432
rect 34659 39392 34704 39420
rect 34698 39380 34704 39392
rect 34756 39380 34762 39432
rect 18104 39324 18368 39352
rect 18104 39312 18110 39324
rect 2222 39244 2228 39296
rect 2280 39284 2286 39296
rect 2409 39287 2467 39293
rect 2409 39284 2421 39287
rect 2280 39256 2421 39284
rect 2280 39244 2286 39256
rect 2409 39253 2421 39256
rect 2455 39253 2467 39287
rect 2409 39247 2467 39253
rect 14185 39287 14243 39293
rect 14185 39253 14197 39287
rect 14231 39284 14243 39287
rect 14274 39284 14280 39296
rect 14231 39256 14280 39284
rect 14231 39253 14243 39256
rect 14185 39247 14243 39253
rect 14274 39244 14280 39256
rect 14332 39244 14338 39296
rect 15010 39284 15016 39296
rect 14971 39256 15016 39284
rect 15010 39244 15016 39256
rect 15068 39244 15074 39296
rect 16298 39284 16304 39296
rect 16259 39256 16304 39284
rect 16298 39244 16304 39256
rect 16356 39244 16362 39296
rect 16574 39244 16580 39296
rect 16632 39284 16638 39296
rect 16669 39287 16727 39293
rect 16669 39284 16681 39287
rect 16632 39256 16681 39284
rect 16632 39244 16638 39256
rect 16669 39253 16681 39256
rect 16715 39253 16727 39287
rect 16669 39247 16727 39253
rect 20254 39244 20260 39296
rect 20312 39284 20318 39296
rect 20717 39287 20775 39293
rect 20717 39284 20729 39287
rect 20312 39256 20729 39284
rect 20312 39244 20318 39256
rect 20717 39253 20729 39256
rect 20763 39284 20775 39287
rect 22462 39284 22468 39296
rect 20763 39256 22468 39284
rect 20763 39253 20775 39256
rect 20717 39247 20775 39253
rect 22462 39244 22468 39256
rect 22520 39244 22526 39296
rect 1104 39194 38824 39216
rect 1104 39142 4246 39194
rect 4298 39142 4310 39194
rect 4362 39142 4374 39194
rect 4426 39142 4438 39194
rect 4490 39142 34966 39194
rect 35018 39142 35030 39194
rect 35082 39142 35094 39194
rect 35146 39142 35158 39194
rect 35210 39142 38824 39194
rect 1104 39120 38824 39142
rect 9398 39080 9404 39092
rect 9359 39052 9404 39080
rect 9398 39040 9404 39052
rect 9456 39040 9462 39092
rect 15562 39040 15568 39092
rect 15620 39080 15626 39092
rect 16301 39083 16359 39089
rect 16301 39080 16313 39083
rect 15620 39052 16313 39080
rect 15620 39040 15626 39052
rect 16301 39049 16313 39052
rect 16347 39049 16359 39083
rect 16758 39080 16764 39092
rect 16719 39052 16764 39080
rect 16301 39043 16359 39049
rect 1670 38944 1676 38956
rect 1583 38916 1676 38944
rect 1670 38904 1676 38916
rect 1728 38944 1734 38956
rect 2406 38944 2412 38956
rect 1728 38916 2412 38944
rect 1728 38904 1734 38916
rect 2406 38904 2412 38916
rect 2464 38904 2470 38956
rect 9416 38944 9444 39040
rect 9861 38947 9919 38953
rect 9861 38944 9873 38947
rect 9416 38916 9873 38944
rect 9861 38913 9873 38916
rect 9907 38913 9919 38947
rect 9861 38907 9919 38913
rect 13265 38947 13323 38953
rect 13265 38913 13277 38947
rect 13311 38944 13323 38947
rect 16316 38944 16344 39043
rect 16758 39040 16764 39052
rect 16816 39040 16822 39092
rect 17770 39080 17776 39092
rect 17731 39052 17776 39080
rect 17770 39040 17776 39052
rect 17828 39040 17834 39092
rect 19334 39080 19340 39092
rect 19295 39052 19340 39080
rect 19334 39040 19340 39052
rect 19392 39040 19398 39092
rect 20990 39080 20996 39092
rect 20951 39052 20996 39080
rect 20990 39040 20996 39052
rect 21048 39040 21054 39092
rect 22373 39083 22431 39089
rect 22373 39049 22385 39083
rect 22419 39080 22431 39083
rect 22462 39080 22468 39092
rect 22419 39052 22468 39080
rect 22419 39049 22431 39052
rect 22373 39043 22431 39049
rect 22462 39040 22468 39052
rect 22520 39040 22526 39092
rect 26329 39083 26387 39089
rect 26329 39049 26341 39083
rect 26375 39080 26387 39083
rect 26602 39080 26608 39092
rect 26375 39052 26608 39080
rect 26375 39049 26387 39052
rect 26329 39043 26387 39049
rect 26602 39040 26608 39052
rect 26660 39040 26666 39092
rect 29454 39040 29460 39092
rect 29512 39080 29518 39092
rect 29733 39083 29791 39089
rect 29733 39080 29745 39083
rect 29512 39052 29745 39080
rect 29512 39040 29518 39052
rect 29733 39049 29745 39052
rect 29779 39049 29791 39083
rect 29733 39043 29791 39049
rect 35161 39083 35219 39089
rect 35161 39049 35173 39083
rect 35207 39080 35219 39083
rect 35710 39080 35716 39092
rect 35207 39052 35716 39080
rect 35207 39049 35219 39052
rect 35161 39043 35219 39049
rect 19352 39012 19380 39040
rect 18616 38984 19380 39012
rect 18046 38944 18052 38956
rect 13311 38916 15700 38944
rect 16316 38916 16620 38944
rect 18007 38916 18052 38944
rect 13311 38913 13323 38916
rect 13265 38907 13323 38913
rect 1397 38879 1455 38885
rect 1397 38845 1409 38879
rect 1443 38876 1455 38879
rect 1946 38876 1952 38888
rect 1443 38848 1952 38876
rect 1443 38845 1455 38848
rect 1397 38839 1455 38845
rect 1946 38836 1952 38848
rect 2004 38836 2010 38888
rect 9125 38879 9183 38885
rect 9125 38845 9137 38879
rect 9171 38876 9183 38879
rect 9398 38876 9404 38888
rect 9171 38848 9404 38876
rect 9171 38845 9183 38848
rect 9125 38839 9183 38845
rect 9398 38836 9404 38848
rect 9456 38876 9462 38888
rect 9585 38879 9643 38885
rect 9585 38876 9597 38879
rect 9456 38848 9597 38876
rect 9456 38836 9462 38848
rect 9585 38845 9597 38848
rect 9631 38876 9643 38879
rect 9674 38876 9680 38888
rect 9631 38848 9680 38876
rect 9631 38845 9643 38848
rect 9585 38839 9643 38845
rect 9674 38836 9680 38848
rect 9732 38836 9738 38888
rect 13725 38879 13783 38885
rect 13725 38876 13737 38879
rect 13096 38848 13737 38876
rect 13096 38752 13124 38848
rect 13725 38845 13737 38848
rect 13771 38845 13783 38879
rect 13725 38839 13783 38845
rect 13906 38836 13912 38888
rect 13964 38876 13970 38888
rect 14093 38879 14151 38885
rect 14093 38876 14105 38879
rect 13964 38848 14105 38876
rect 13964 38836 13970 38848
rect 14093 38845 14105 38848
rect 14139 38845 14151 38879
rect 14274 38876 14280 38888
rect 14235 38848 14280 38876
rect 14093 38839 14151 38845
rect 14274 38836 14280 38848
rect 14332 38836 14338 38888
rect 14737 38879 14795 38885
rect 14737 38845 14749 38879
rect 14783 38876 14795 38879
rect 14918 38876 14924 38888
rect 14783 38848 14924 38876
rect 14783 38845 14795 38848
rect 14737 38839 14795 38845
rect 13633 38811 13691 38817
rect 13633 38777 13645 38811
rect 13679 38808 13691 38811
rect 14752 38808 14780 38839
rect 14918 38836 14924 38848
rect 14976 38836 14982 38888
rect 15102 38876 15108 38888
rect 15063 38848 15108 38876
rect 15102 38836 15108 38848
rect 15160 38836 15166 38888
rect 15672 38885 15700 38916
rect 16592 38888 16620 38916
rect 18046 38904 18052 38916
rect 18104 38904 18110 38956
rect 18414 38904 18420 38956
rect 18472 38944 18478 38956
rect 18616 38953 18644 38984
rect 19978 38972 19984 39024
rect 20036 39021 20042 39024
rect 20036 39015 20085 39021
rect 20036 38981 20039 39015
rect 20073 38981 20085 39015
rect 20036 38975 20085 38981
rect 20165 39015 20223 39021
rect 20165 38981 20177 39015
rect 20211 38981 20223 39015
rect 20165 38975 20223 38981
rect 26697 39015 26755 39021
rect 26697 38981 26709 39015
rect 26743 39012 26755 39015
rect 27246 39012 27252 39024
rect 26743 38984 27252 39012
rect 26743 38981 26755 38984
rect 26697 38975 26755 38981
rect 20036 38972 20042 38975
rect 18601 38947 18659 38953
rect 18601 38944 18613 38947
rect 18472 38916 18613 38944
rect 18472 38904 18478 38916
rect 18601 38913 18613 38916
rect 18647 38913 18659 38947
rect 19058 38944 19064 38956
rect 19019 38916 19064 38944
rect 18601 38907 18659 38913
rect 19058 38904 19064 38916
rect 19116 38904 19122 38956
rect 15657 38879 15715 38885
rect 15657 38845 15669 38879
rect 15703 38876 15715 38879
rect 16114 38876 16120 38888
rect 15703 38848 16120 38876
rect 15703 38845 15715 38848
rect 15657 38839 15715 38845
rect 16114 38836 16120 38848
rect 16172 38836 16178 38888
rect 16298 38836 16304 38888
rect 16356 38876 16362 38888
rect 16482 38876 16488 38888
rect 16356 38848 16488 38876
rect 16356 38836 16362 38848
rect 16482 38836 16488 38848
rect 16540 38836 16546 38888
rect 16574 38836 16580 38888
rect 16632 38876 16638 38888
rect 17313 38879 17371 38885
rect 17313 38876 17325 38879
rect 16632 38848 17325 38876
rect 16632 38836 16638 38848
rect 17313 38845 17325 38848
rect 17359 38845 17371 38879
rect 17313 38839 17371 38845
rect 18877 38879 18935 38885
rect 18877 38845 18889 38879
rect 18923 38876 18935 38879
rect 19150 38876 19156 38888
rect 18923 38848 19156 38876
rect 18923 38845 18935 38848
rect 18877 38839 18935 38845
rect 19150 38836 19156 38848
rect 19208 38836 19214 38888
rect 19797 38879 19855 38885
rect 19797 38845 19809 38879
rect 19843 38876 19855 38879
rect 20070 38876 20076 38888
rect 19843 38848 20076 38876
rect 19843 38845 19855 38848
rect 19797 38839 19855 38845
rect 20070 38836 20076 38848
rect 20128 38876 20134 38888
rect 20180 38876 20208 38975
rect 27246 38972 27252 38984
rect 27304 39012 27310 39024
rect 27304 38984 27844 39012
rect 27304 38972 27310 38984
rect 20254 38904 20260 38956
rect 20312 38944 20318 38956
rect 24397 38947 24455 38953
rect 20312 38916 20357 38944
rect 20312 38904 20318 38916
rect 24397 38913 24409 38947
rect 24443 38944 24455 38947
rect 25041 38947 25099 38953
rect 25041 38944 25053 38947
rect 24443 38916 25053 38944
rect 24443 38913 24455 38916
rect 24397 38907 24455 38913
rect 25041 38913 25053 38916
rect 25087 38944 25099 38947
rect 25130 38944 25136 38956
rect 25087 38916 25136 38944
rect 25087 38913 25099 38916
rect 25041 38907 25099 38913
rect 25130 38904 25136 38916
rect 25188 38904 25194 38956
rect 25961 38947 26019 38953
rect 25961 38913 25973 38947
rect 26007 38944 26019 38947
rect 26050 38944 26056 38956
rect 26007 38916 26056 38944
rect 26007 38913 26019 38916
rect 25961 38907 26019 38913
rect 26050 38904 26056 38916
rect 26108 38904 26114 38956
rect 26510 38904 26516 38956
rect 26568 38944 26574 38956
rect 27154 38944 27160 38956
rect 26568 38916 27160 38944
rect 26568 38904 26574 38916
rect 27154 38904 27160 38916
rect 27212 38944 27218 38956
rect 27816 38953 27844 38984
rect 27341 38947 27399 38953
rect 27341 38944 27353 38947
rect 27212 38916 27353 38944
rect 27212 38904 27218 38916
rect 27341 38913 27353 38916
rect 27387 38913 27399 38947
rect 27341 38907 27399 38913
rect 27801 38947 27859 38953
rect 27801 38913 27813 38947
rect 27847 38913 27859 38947
rect 29748 38944 29776 39043
rect 35710 39040 35716 39052
rect 35768 39040 35774 39092
rect 30193 38947 30251 38953
rect 30193 38944 30205 38947
rect 29748 38916 30205 38944
rect 27801 38907 27859 38913
rect 30193 38913 30205 38916
rect 30239 38913 30251 38947
rect 30193 38907 30251 38913
rect 20128 38848 20208 38876
rect 20625 38879 20683 38885
rect 20128 38836 20134 38848
rect 20625 38845 20637 38879
rect 20671 38876 20683 38879
rect 21453 38879 21511 38885
rect 21453 38876 21465 38879
rect 20671 38848 21465 38876
rect 20671 38845 20683 38848
rect 20625 38839 20683 38845
rect 21453 38845 21465 38848
rect 21499 38876 21511 38879
rect 21913 38879 21971 38885
rect 21913 38876 21925 38879
rect 21499 38848 21925 38876
rect 21499 38845 21511 38848
rect 21453 38839 21511 38845
rect 21913 38845 21925 38848
rect 21959 38845 21971 38879
rect 21913 38839 21971 38845
rect 24765 38879 24823 38885
rect 24765 38845 24777 38879
rect 24811 38876 24823 38879
rect 25406 38876 25412 38888
rect 24811 38848 25412 38876
rect 24811 38845 24823 38848
rect 24765 38839 24823 38845
rect 25406 38836 25412 38848
rect 25464 38836 25470 38888
rect 25774 38876 25780 38888
rect 25735 38848 25780 38876
rect 25774 38836 25780 38848
rect 25832 38836 25838 38888
rect 26878 38836 26884 38888
rect 26936 38876 26942 38888
rect 27617 38879 27675 38885
rect 27617 38876 27629 38879
rect 26936 38848 27629 38876
rect 26936 38836 26942 38848
rect 27617 38845 27629 38848
rect 27663 38876 27675 38879
rect 28074 38876 28080 38888
rect 27663 38848 28080 38876
rect 27663 38845 27675 38848
rect 27617 38839 27675 38845
rect 28074 38836 28080 38848
rect 28132 38836 28138 38888
rect 29546 38836 29552 38888
rect 29604 38876 29610 38888
rect 29914 38876 29920 38888
rect 29604 38848 29920 38876
rect 29604 38836 29610 38848
rect 29914 38836 29920 38848
rect 29972 38836 29978 38888
rect 19886 38808 19892 38820
rect 13679 38780 14780 38808
rect 19799 38780 19892 38808
rect 13679 38777 13691 38780
rect 13633 38771 13691 38777
rect 19886 38768 19892 38780
rect 19944 38808 19950 38820
rect 20990 38808 20996 38820
rect 19944 38780 20996 38808
rect 19944 38768 19950 38780
rect 20990 38768 20996 38780
rect 21048 38768 21054 38820
rect 21361 38811 21419 38817
rect 21361 38777 21373 38811
rect 21407 38808 21419 38811
rect 21726 38808 21732 38820
rect 21407 38780 21732 38808
rect 21407 38777 21419 38780
rect 21361 38771 21419 38777
rect 21726 38768 21732 38780
rect 21784 38808 21790 38820
rect 22462 38808 22468 38820
rect 21784 38780 22468 38808
rect 21784 38768 21790 38780
rect 22462 38768 22468 38780
rect 22520 38768 22526 38820
rect 24029 38811 24087 38817
rect 24029 38777 24041 38811
rect 24075 38808 24087 38811
rect 25792 38808 25820 38836
rect 26786 38808 26792 38820
rect 24075 38780 25820 38808
rect 26747 38780 26792 38808
rect 24075 38777 24087 38780
rect 24029 38771 24087 38777
rect 26786 38768 26792 38780
rect 26844 38768 26850 38820
rect 2774 38700 2780 38752
rect 2832 38740 2838 38752
rect 11146 38740 11152 38752
rect 2832 38712 2877 38740
rect 11107 38712 11152 38740
rect 2832 38700 2838 38712
rect 11146 38700 11152 38712
rect 11204 38700 11210 38752
rect 12897 38743 12955 38749
rect 12897 38709 12909 38743
rect 12943 38740 12955 38743
rect 13078 38740 13084 38752
rect 12943 38712 13084 38740
rect 12943 38709 12955 38712
rect 12897 38703 12955 38709
rect 13078 38700 13084 38712
rect 13136 38700 13142 38752
rect 16025 38743 16083 38749
rect 16025 38709 16037 38743
rect 16071 38740 16083 38743
rect 16206 38740 16212 38752
rect 16071 38712 16212 38740
rect 16071 38709 16083 38712
rect 16025 38703 16083 38709
rect 16206 38700 16212 38712
rect 16264 38700 16270 38752
rect 21634 38740 21640 38752
rect 21595 38712 21640 38740
rect 21634 38700 21640 38712
rect 21692 38700 21698 38752
rect 30466 38700 30472 38752
rect 30524 38740 30530 38752
rect 31297 38743 31355 38749
rect 31297 38740 31309 38743
rect 30524 38712 31309 38740
rect 30524 38700 30530 38712
rect 31297 38709 31309 38712
rect 31343 38709 31355 38743
rect 31297 38703 31355 38709
rect 1104 38650 38824 38672
rect 1104 38598 19606 38650
rect 19658 38598 19670 38650
rect 19722 38598 19734 38650
rect 19786 38598 19798 38650
rect 19850 38598 38824 38650
rect 1104 38576 38824 38598
rect 1670 38536 1676 38548
rect 1631 38508 1676 38536
rect 1670 38496 1676 38508
rect 1728 38496 1734 38548
rect 1946 38536 1952 38548
rect 1907 38508 1952 38536
rect 1946 38496 1952 38508
rect 2004 38496 2010 38548
rect 13722 38496 13728 38548
rect 13780 38536 13786 38548
rect 13906 38536 13912 38548
rect 13780 38508 13912 38536
rect 13780 38496 13786 38508
rect 13906 38496 13912 38508
rect 13964 38496 13970 38548
rect 15930 38536 15936 38548
rect 15891 38508 15936 38536
rect 15930 38496 15936 38508
rect 15988 38496 15994 38548
rect 19334 38496 19340 38548
rect 19392 38536 19398 38548
rect 19978 38536 19984 38548
rect 19392 38508 19984 38536
rect 19392 38496 19398 38508
rect 19978 38496 19984 38508
rect 20036 38496 20042 38548
rect 20717 38539 20775 38545
rect 20717 38505 20729 38539
rect 20763 38536 20775 38539
rect 20990 38536 20996 38548
rect 20763 38508 20996 38536
rect 20763 38505 20775 38508
rect 20717 38499 20775 38505
rect 20990 38496 20996 38508
rect 21048 38496 21054 38548
rect 21174 38496 21180 38548
rect 21232 38536 21238 38548
rect 21729 38539 21787 38545
rect 21729 38536 21741 38539
rect 21232 38508 21741 38536
rect 21232 38496 21238 38508
rect 21729 38505 21741 38508
rect 21775 38505 21787 38539
rect 21729 38499 21787 38505
rect 25038 38496 25044 38548
rect 25096 38536 25102 38548
rect 25685 38539 25743 38545
rect 25685 38536 25697 38539
rect 25096 38508 25697 38536
rect 25096 38496 25102 38508
rect 25685 38505 25697 38508
rect 25731 38505 25743 38539
rect 26878 38536 26884 38548
rect 26839 38508 26884 38536
rect 25685 38499 25743 38505
rect 26878 38496 26884 38508
rect 26936 38496 26942 38548
rect 27154 38536 27160 38548
rect 27115 38508 27160 38536
rect 27154 38496 27160 38508
rect 27212 38496 27218 38548
rect 29914 38536 29920 38548
rect 29875 38508 29920 38536
rect 29914 38496 29920 38508
rect 29972 38496 29978 38548
rect 12158 38468 12164 38480
rect 11808 38440 12164 38468
rect 11808 38412 11836 38440
rect 12158 38428 12164 38440
rect 12216 38428 12222 38480
rect 13265 38471 13323 38477
rect 13265 38437 13277 38471
rect 13311 38468 13323 38471
rect 13311 38440 14412 38468
rect 13311 38437 13323 38440
rect 13265 38431 13323 38437
rect 14384 38412 14412 38440
rect 18046 38428 18052 38480
rect 18104 38468 18110 38480
rect 18141 38471 18199 38477
rect 18141 38468 18153 38471
rect 18104 38440 18153 38468
rect 18104 38428 18110 38440
rect 18141 38437 18153 38440
rect 18187 38468 18199 38471
rect 18187 38440 19196 38468
rect 18187 38437 18199 38440
rect 18141 38431 18199 38437
rect 19168 38412 19196 38440
rect 25314 38428 25320 38480
rect 25372 38428 25378 38480
rect 11790 38400 11796 38412
rect 11703 38372 11796 38400
rect 11790 38360 11796 38372
rect 11848 38360 11854 38412
rect 11974 38400 11980 38412
rect 11935 38372 11980 38400
rect 11974 38360 11980 38372
rect 12032 38360 12038 38412
rect 12250 38360 12256 38412
rect 12308 38400 12314 38412
rect 12345 38403 12403 38409
rect 12345 38400 12357 38403
rect 12308 38372 12357 38400
rect 12308 38360 12314 38372
rect 12345 38369 12357 38372
rect 12391 38369 12403 38403
rect 12345 38363 12403 38369
rect 12529 38403 12587 38409
rect 12529 38369 12541 38403
rect 12575 38400 12587 38403
rect 12618 38400 12624 38412
rect 12575 38372 12624 38400
rect 12575 38369 12587 38372
rect 12529 38363 12587 38369
rect 12618 38360 12624 38372
rect 12676 38360 12682 38412
rect 14090 38360 14096 38412
rect 14148 38400 14154 38412
rect 14185 38403 14243 38409
rect 14185 38400 14197 38403
rect 14148 38372 14197 38400
rect 14148 38360 14154 38372
rect 14185 38369 14197 38372
rect 14231 38369 14243 38403
rect 14366 38400 14372 38412
rect 14327 38372 14372 38400
rect 14185 38363 14243 38369
rect 14366 38360 14372 38372
rect 14424 38360 14430 38412
rect 16022 38400 16028 38412
rect 15983 38372 16028 38400
rect 16022 38360 16028 38372
rect 16080 38360 16086 38412
rect 16114 38360 16120 38412
rect 16172 38400 16178 38412
rect 16393 38403 16451 38409
rect 16393 38400 16405 38403
rect 16172 38372 16405 38400
rect 16172 38360 16178 38372
rect 16393 38369 16405 38372
rect 16439 38369 16451 38403
rect 16393 38363 16451 38369
rect 16853 38403 16911 38409
rect 16853 38369 16865 38403
rect 16899 38369 16911 38403
rect 19058 38400 19064 38412
rect 19019 38372 19064 38400
rect 16853 38363 16911 38369
rect 11330 38332 11336 38344
rect 11291 38304 11336 38332
rect 11330 38292 11336 38304
rect 11388 38292 11394 38344
rect 13354 38332 13360 38344
rect 13315 38304 13360 38332
rect 13354 38292 13360 38304
rect 13412 38292 13418 38344
rect 13906 38332 13912 38344
rect 13867 38304 13912 38332
rect 13906 38292 13912 38304
rect 13964 38332 13970 38344
rect 16868 38332 16896 38363
rect 19058 38360 19064 38372
rect 19116 38360 19122 38412
rect 19150 38360 19156 38412
rect 19208 38400 19214 38412
rect 19429 38403 19487 38409
rect 19429 38400 19441 38403
rect 19208 38372 19441 38400
rect 19208 38360 19214 38372
rect 19429 38369 19441 38372
rect 19475 38400 19487 38403
rect 20438 38400 20444 38412
rect 19475 38372 20444 38400
rect 19475 38369 19487 38372
rect 19429 38363 19487 38369
rect 20438 38360 20444 38372
rect 20496 38360 20502 38412
rect 20990 38400 20996 38412
rect 20951 38372 20996 38400
rect 20990 38360 20996 38372
rect 21048 38360 21054 38412
rect 24302 38360 24308 38412
rect 24360 38400 24366 38412
rect 24397 38403 24455 38409
rect 24397 38400 24409 38403
rect 24360 38372 24409 38400
rect 24360 38360 24366 38372
rect 24397 38369 24409 38372
rect 24443 38369 24455 38403
rect 24397 38363 24455 38369
rect 25225 38403 25283 38409
rect 25225 38369 25237 38403
rect 25271 38400 25283 38403
rect 25332 38400 25360 38428
rect 25271 38372 25360 38400
rect 27985 38403 28043 38409
rect 25271 38369 25283 38372
rect 25225 38363 25283 38369
rect 27985 38369 27997 38403
rect 28031 38400 28043 38403
rect 28074 38400 28080 38412
rect 28031 38372 28080 38400
rect 28031 38369 28043 38372
rect 27985 38363 28043 38369
rect 17402 38332 17408 38344
rect 13964 38304 17408 38332
rect 13964 38292 13970 38304
rect 17402 38292 17408 38304
rect 17460 38292 17466 38344
rect 17862 38292 17868 38344
rect 17920 38332 17926 38344
rect 18693 38335 18751 38341
rect 18693 38332 18705 38335
rect 17920 38304 18705 38332
rect 17920 38292 17926 38304
rect 18693 38301 18705 38304
rect 18739 38332 18751 38335
rect 20901 38335 20959 38341
rect 18739 38304 20760 38332
rect 18739 38301 18751 38304
rect 18693 38295 18751 38301
rect 16850 38264 16856 38276
rect 16811 38236 16856 38264
rect 16850 38224 16856 38236
rect 16908 38224 16914 38276
rect 17497 38267 17555 38273
rect 17497 38233 17509 38267
rect 17543 38264 17555 38267
rect 18230 38264 18236 38276
rect 17543 38236 18236 38264
rect 17543 38233 17555 38236
rect 17497 38227 17555 38233
rect 18230 38224 18236 38236
rect 18288 38264 18294 38276
rect 19337 38267 19395 38273
rect 19337 38264 19349 38267
rect 18288 38236 19349 38264
rect 18288 38224 18294 38236
rect 19337 38233 19349 38236
rect 19383 38233 19395 38267
rect 20732 38264 20760 38304
rect 20901 38301 20913 38335
rect 20947 38332 20959 38335
rect 21082 38332 21088 38344
rect 20947 38304 21088 38332
rect 20947 38301 20959 38304
rect 20901 38295 20959 38301
rect 21082 38292 21088 38304
rect 21140 38292 21146 38344
rect 24486 38332 24492 38344
rect 24447 38304 24492 38332
rect 24486 38292 24492 38304
rect 24544 38292 24550 38344
rect 25240 38264 25268 38363
rect 28074 38360 28080 38372
rect 28132 38360 28138 38412
rect 25317 38335 25375 38341
rect 25317 38301 25329 38335
rect 25363 38332 25375 38335
rect 25498 38332 25504 38344
rect 25363 38304 25504 38332
rect 25363 38301 25375 38304
rect 25317 38295 25375 38301
rect 25498 38292 25504 38304
rect 25556 38292 25562 38344
rect 27709 38335 27767 38341
rect 27709 38301 27721 38335
rect 27755 38332 27767 38335
rect 28350 38332 28356 38344
rect 27755 38304 28356 38332
rect 27755 38301 27767 38304
rect 27709 38295 27767 38301
rect 28350 38292 28356 38304
rect 28408 38292 28414 38344
rect 20732 38236 21220 38264
rect 19337 38227 19395 38233
rect 11054 38156 11060 38208
rect 11112 38196 11118 38208
rect 11149 38199 11207 38205
rect 11149 38196 11161 38199
rect 11112 38168 11161 38196
rect 11112 38156 11118 38168
rect 11149 38165 11161 38168
rect 11195 38196 11207 38199
rect 12250 38196 12256 38208
rect 11195 38168 12256 38196
rect 11195 38165 11207 38168
rect 11149 38159 11207 38165
rect 12250 38156 12256 38168
rect 12308 38156 12314 38208
rect 12526 38156 12532 38208
rect 12584 38196 12590 38208
rect 12805 38199 12863 38205
rect 12805 38196 12817 38199
rect 12584 38168 12817 38196
rect 12584 38156 12590 38168
rect 12805 38165 12817 38168
rect 12851 38165 12863 38199
rect 14734 38196 14740 38208
rect 14695 38168 14740 38196
rect 12805 38159 12863 38165
rect 14734 38156 14740 38168
rect 14792 38156 14798 38208
rect 15102 38196 15108 38208
rect 15063 38168 15108 38196
rect 15102 38156 15108 38168
rect 15160 38156 15166 38208
rect 15286 38156 15292 38208
rect 15344 38196 15350 38208
rect 15473 38199 15531 38205
rect 15473 38196 15485 38199
rect 15344 38168 15485 38196
rect 15344 38156 15350 38168
rect 15473 38165 15485 38168
rect 15519 38165 15531 38199
rect 15473 38159 15531 38165
rect 18782 38156 18788 38208
rect 18840 38196 18846 38208
rect 21192 38205 21220 38236
rect 24136 38236 25268 38264
rect 24136 38208 24164 38236
rect 20257 38199 20315 38205
rect 20257 38196 20269 38199
rect 18840 38168 20269 38196
rect 18840 38156 18846 38168
rect 20257 38165 20269 38168
rect 20303 38165 20315 38199
rect 20257 38159 20315 38165
rect 21177 38199 21235 38205
rect 21177 38165 21189 38199
rect 21223 38165 21235 38199
rect 24118 38196 24124 38208
rect 24079 38168 24124 38196
rect 21177 38159 21235 38165
rect 24118 38156 24124 38168
rect 24176 38156 24182 38208
rect 27617 38199 27675 38205
rect 27617 38165 27629 38199
rect 27663 38196 27675 38199
rect 27706 38196 27712 38208
rect 27663 38168 27712 38196
rect 27663 38165 27675 38168
rect 27617 38159 27675 38165
rect 27706 38156 27712 38168
rect 27764 38196 27770 38208
rect 29089 38199 29147 38205
rect 29089 38196 29101 38199
rect 27764 38168 29101 38196
rect 27764 38156 27770 38168
rect 29089 38165 29101 38168
rect 29135 38165 29147 38199
rect 29089 38159 29147 38165
rect 1104 38106 38824 38128
rect 1104 38054 4246 38106
rect 4298 38054 4310 38106
rect 4362 38054 4374 38106
rect 4426 38054 4438 38106
rect 4490 38054 34966 38106
rect 35018 38054 35030 38106
rect 35082 38054 35094 38106
rect 35146 38054 35158 38106
rect 35210 38054 38824 38106
rect 1104 38032 38824 38054
rect 11057 37995 11115 38001
rect 11057 37961 11069 37995
rect 11103 37992 11115 37995
rect 12618 37992 12624 38004
rect 11103 37964 12624 37992
rect 11103 37961 11115 37964
rect 11057 37955 11115 37961
rect 12618 37952 12624 37964
rect 12676 37952 12682 38004
rect 13630 37992 13636 38004
rect 13591 37964 13636 37992
rect 13630 37952 13636 37964
rect 13688 37952 13694 38004
rect 13906 37952 13912 38004
rect 13964 37992 13970 38004
rect 14093 37995 14151 38001
rect 14093 37992 14105 37995
rect 13964 37964 14105 37992
rect 13964 37952 13970 37964
rect 14093 37961 14105 37964
rect 14139 37961 14151 37995
rect 14093 37955 14151 37961
rect 15841 37995 15899 38001
rect 15841 37961 15853 37995
rect 15887 37992 15899 37995
rect 16022 37992 16028 38004
rect 15887 37964 16028 37992
rect 15887 37961 15899 37964
rect 15841 37955 15899 37961
rect 16022 37952 16028 37964
rect 16080 37952 16086 38004
rect 17402 37992 17408 38004
rect 17363 37964 17408 37992
rect 17402 37952 17408 37964
rect 17460 37952 17466 38004
rect 17862 37992 17868 38004
rect 17823 37964 17868 37992
rect 17862 37952 17868 37964
rect 17920 37952 17926 38004
rect 19794 37992 19800 38004
rect 19755 37964 19800 37992
rect 19794 37952 19800 37964
rect 19852 37952 19858 38004
rect 23477 37995 23535 38001
rect 23477 37961 23489 37995
rect 23523 37992 23535 37995
rect 24302 37992 24308 38004
rect 23523 37964 24308 37992
rect 23523 37961 23535 37964
rect 23477 37955 23535 37961
rect 24302 37952 24308 37964
rect 24360 37952 24366 38004
rect 25498 37952 25504 38004
rect 25556 37992 25562 38004
rect 26237 37995 26295 38001
rect 26237 37992 26249 37995
rect 25556 37964 26249 37992
rect 25556 37952 25562 37964
rect 26237 37961 26249 37964
rect 26283 37961 26295 37995
rect 26237 37955 26295 37961
rect 11425 37927 11483 37933
rect 11425 37893 11437 37927
rect 11471 37924 11483 37927
rect 11790 37924 11796 37936
rect 11471 37896 11796 37924
rect 11471 37893 11483 37896
rect 11425 37887 11483 37893
rect 11790 37884 11796 37896
rect 11848 37884 11854 37936
rect 15473 37927 15531 37933
rect 15473 37893 15485 37927
rect 15519 37924 15531 37927
rect 17126 37924 17132 37936
rect 15519 37896 17132 37924
rect 15519 37893 15531 37896
rect 15473 37887 15531 37893
rect 17126 37884 17132 37896
rect 17184 37884 17190 37936
rect 19812 37924 19840 37952
rect 24029 37927 24087 37933
rect 19812 37896 20484 37924
rect 12526 37856 12532 37868
rect 12487 37828 12532 37856
rect 12526 37816 12532 37828
rect 12584 37816 12590 37868
rect 14274 37816 14280 37868
rect 14332 37856 14338 37868
rect 14829 37859 14887 37865
rect 14829 37856 14841 37859
rect 14332 37828 14841 37856
rect 14332 37816 14338 37828
rect 14829 37825 14841 37828
rect 14875 37856 14887 37859
rect 15930 37856 15936 37868
rect 14875 37828 15936 37856
rect 14875 37825 14887 37828
rect 14829 37819 14887 37825
rect 12621 37791 12679 37797
rect 12621 37757 12633 37791
rect 12667 37757 12679 37791
rect 12621 37751 12679 37757
rect 13173 37791 13231 37797
rect 13173 37757 13185 37791
rect 13219 37757 13231 37791
rect 13173 37751 13231 37757
rect 13357 37791 13415 37797
rect 13357 37757 13369 37791
rect 13403 37788 13415 37791
rect 13538 37788 13544 37800
rect 13403 37760 13544 37788
rect 13403 37757 13415 37760
rect 13357 37751 13415 37757
rect 10689 37723 10747 37729
rect 10689 37689 10701 37723
rect 10735 37720 10747 37723
rect 11974 37720 11980 37732
rect 10735 37692 11980 37720
rect 10735 37689 10747 37692
rect 10689 37683 10747 37689
rect 11974 37680 11980 37692
rect 12032 37680 12038 37732
rect 12636 37720 12664 37751
rect 13188 37720 13216 37751
rect 13538 37748 13544 37760
rect 13596 37748 13602 37800
rect 14936 37797 14964 37828
rect 15930 37816 15936 37828
rect 15988 37856 15994 37868
rect 16485 37859 16543 37865
rect 16485 37856 16497 37859
rect 15988 37828 16497 37856
rect 15988 37816 15994 37828
rect 16485 37825 16497 37828
rect 16531 37825 16543 37859
rect 16485 37819 16543 37825
rect 14921 37791 14979 37797
rect 14921 37757 14933 37791
rect 14967 37757 14979 37791
rect 16574 37788 16580 37800
rect 16535 37760 16580 37788
rect 14921 37751 14979 37757
rect 16574 37748 16580 37760
rect 16632 37748 16638 37800
rect 16942 37788 16948 37800
rect 16903 37760 16948 37788
rect 16942 37748 16948 37760
rect 17000 37748 17006 37800
rect 17126 37788 17132 37800
rect 17087 37760 17132 37788
rect 17126 37748 17132 37760
rect 17184 37748 17190 37800
rect 18230 37788 18236 37800
rect 18143 37760 18236 37788
rect 18230 37748 18236 37760
rect 18288 37788 18294 37800
rect 18414 37788 18420 37800
rect 18288 37760 18420 37788
rect 18288 37748 18294 37760
rect 18414 37748 18420 37760
rect 18472 37748 18478 37800
rect 18782 37788 18788 37800
rect 18743 37760 18788 37788
rect 18782 37748 18788 37760
rect 18840 37748 18846 37800
rect 18874 37748 18880 37800
rect 18932 37788 18938 37800
rect 18932 37760 18977 37788
rect 18932 37748 18938 37760
rect 19058 37748 19064 37800
rect 19116 37788 19122 37800
rect 19521 37791 19579 37797
rect 19521 37788 19533 37791
rect 19116 37760 19533 37788
rect 19116 37748 19122 37760
rect 19521 37757 19533 37760
rect 19567 37788 19579 37791
rect 20070 37788 20076 37800
rect 19567 37760 20076 37788
rect 19567 37757 19579 37760
rect 19521 37751 19579 37757
rect 20070 37748 20076 37760
rect 20128 37748 20134 37800
rect 20456 37797 20484 37896
rect 24029 37893 24041 37927
rect 24075 37924 24087 37927
rect 25516 37924 25544 37952
rect 24075 37896 25544 37924
rect 26252 37924 26280 37955
rect 28074 37952 28080 38004
rect 28132 37992 28138 38004
rect 28169 37995 28227 38001
rect 28169 37992 28181 37995
rect 28132 37964 28181 37992
rect 28132 37952 28138 37964
rect 28169 37961 28181 37964
rect 28215 37961 28227 37995
rect 28169 37955 28227 37961
rect 28350 37952 28356 38004
rect 28408 37992 28414 38004
rect 28629 37995 28687 38001
rect 28629 37992 28641 37995
rect 28408 37964 28641 37992
rect 28408 37952 28414 37964
rect 28629 37961 28641 37964
rect 28675 37992 28687 37995
rect 29546 37992 29552 38004
rect 28675 37964 29552 37992
rect 28675 37961 28687 37964
rect 28629 37955 28687 37961
rect 29546 37952 29552 37964
rect 29604 37952 29610 38004
rect 26252 37896 27844 37924
rect 24075 37893 24087 37896
rect 24029 37887 24087 37893
rect 21542 37816 21548 37868
rect 21600 37856 21606 37868
rect 21637 37859 21695 37865
rect 21637 37856 21649 37859
rect 21600 37828 21649 37856
rect 21600 37816 21606 37828
rect 21637 37825 21649 37828
rect 21683 37825 21695 37859
rect 21637 37819 21695 37825
rect 24765 37859 24823 37865
rect 24765 37825 24777 37859
rect 24811 37856 24823 37859
rect 25041 37859 25099 37865
rect 25041 37856 25053 37859
rect 24811 37828 25053 37856
rect 24811 37825 24823 37828
rect 24765 37819 24823 37825
rect 25041 37825 25053 37828
rect 25087 37856 25099 37859
rect 27246 37856 27252 37868
rect 25087 37828 27252 37856
rect 25087 37825 25099 37828
rect 25041 37819 25099 37825
rect 27246 37816 27252 37828
rect 27304 37816 27310 37868
rect 27816 37865 27844 37896
rect 27801 37859 27859 37865
rect 27801 37825 27813 37859
rect 27847 37825 27859 37859
rect 27801 37819 27859 37825
rect 20441 37791 20499 37797
rect 20441 37757 20453 37791
rect 20487 37757 20499 37791
rect 20441 37751 20499 37757
rect 20625 37791 20683 37797
rect 20625 37757 20637 37791
rect 20671 37757 20683 37791
rect 20806 37788 20812 37800
rect 20767 37760 20812 37788
rect 20625 37751 20683 37757
rect 15930 37720 15936 37732
rect 12636 37692 13216 37720
rect 15891 37692 15936 37720
rect 11885 37655 11943 37661
rect 11885 37621 11897 37655
rect 11931 37652 11943 37655
rect 12161 37655 12219 37661
rect 12161 37652 12173 37655
rect 11931 37624 12173 37652
rect 11931 37621 11943 37624
rect 11885 37615 11943 37621
rect 12161 37621 12173 37624
rect 12207 37652 12219 37655
rect 12636 37652 12664 37692
rect 15930 37680 15936 37692
rect 15988 37680 15994 37732
rect 19978 37720 19984 37732
rect 19939 37692 19984 37720
rect 19978 37680 19984 37692
rect 20036 37680 20042 37732
rect 20346 37680 20352 37732
rect 20404 37720 20410 37732
rect 20640 37720 20668 37751
rect 20806 37748 20812 37760
rect 20864 37748 20870 37800
rect 24397 37791 24455 37797
rect 24397 37757 24409 37791
rect 24443 37788 24455 37791
rect 25406 37788 25412 37800
rect 24443 37760 25412 37788
rect 24443 37757 24455 37760
rect 24397 37751 24455 37757
rect 25406 37748 25412 37760
rect 25464 37748 25470 37800
rect 25682 37788 25688 37800
rect 25643 37760 25688 37788
rect 25682 37748 25688 37760
rect 25740 37788 25746 37800
rect 26605 37791 26663 37797
rect 26605 37788 26617 37791
rect 25740 37760 26617 37788
rect 25740 37748 25746 37760
rect 26605 37757 26617 37760
rect 26651 37788 26663 37791
rect 26786 37788 26792 37800
rect 26651 37760 26792 37788
rect 26651 37757 26663 37760
rect 26605 37751 26663 37757
rect 26786 37748 26792 37760
rect 26844 37788 26850 37800
rect 26881 37791 26939 37797
rect 26881 37788 26893 37791
rect 26844 37760 26893 37788
rect 26844 37748 26850 37760
rect 26881 37757 26893 37760
rect 26927 37757 26939 37791
rect 27706 37788 27712 37800
rect 27667 37760 27712 37788
rect 26881 37751 26939 37757
rect 27706 37748 27712 37760
rect 27764 37748 27770 37800
rect 25958 37720 25964 37732
rect 20404 37692 20668 37720
rect 25919 37692 25964 37720
rect 20404 37680 20410 37692
rect 25958 37680 25964 37692
rect 26016 37680 26022 37732
rect 26973 37723 27031 37729
rect 26973 37720 26985 37723
rect 26896 37692 26985 37720
rect 26896 37664 26924 37692
rect 26973 37689 26985 37692
rect 27019 37689 27031 37723
rect 26973 37683 27031 37689
rect 12802 37652 12808 37664
rect 12207 37624 12808 37652
rect 12207 37621 12219 37624
rect 12161 37615 12219 37621
rect 12802 37612 12808 37624
rect 12860 37612 12866 37664
rect 13262 37612 13268 37664
rect 13320 37652 13326 37664
rect 15105 37655 15163 37661
rect 15105 37652 15117 37655
rect 13320 37624 15117 37652
rect 13320 37612 13326 37624
rect 15105 37621 15117 37624
rect 15151 37652 15163 37655
rect 16850 37652 16856 37664
rect 15151 37624 16856 37652
rect 15151 37621 15163 37624
rect 15105 37615 15163 37621
rect 16850 37612 16856 37624
rect 16908 37612 16914 37664
rect 17954 37612 17960 37664
rect 18012 37652 18018 37664
rect 18141 37655 18199 37661
rect 18141 37652 18153 37655
rect 18012 37624 18153 37652
rect 18012 37612 18018 37624
rect 18141 37621 18153 37624
rect 18187 37652 18199 37655
rect 19150 37652 19156 37664
rect 18187 37624 19156 37652
rect 18187 37621 18199 37624
rect 18141 37615 18199 37621
rect 19150 37612 19156 37624
rect 19208 37612 19214 37664
rect 20438 37612 20444 37664
rect 20496 37652 20502 37664
rect 21082 37652 21088 37664
rect 20496 37624 21088 37652
rect 20496 37612 20502 37624
rect 21082 37612 21088 37624
rect 21140 37652 21146 37664
rect 21269 37655 21327 37661
rect 21269 37652 21281 37655
rect 21140 37624 21281 37652
rect 21140 37612 21146 37624
rect 21269 37621 21281 37624
rect 21315 37621 21327 37655
rect 21269 37615 21327 37621
rect 26878 37612 26884 37664
rect 26936 37612 26942 37664
rect 1104 37562 38824 37584
rect 1104 37510 19606 37562
rect 19658 37510 19670 37562
rect 19722 37510 19734 37562
rect 19786 37510 19798 37562
rect 19850 37510 38824 37562
rect 1104 37488 38824 37510
rect 11974 37408 11980 37460
rect 12032 37448 12038 37460
rect 12161 37451 12219 37457
rect 12161 37448 12173 37451
rect 12032 37420 12173 37448
rect 12032 37408 12038 37420
rect 12161 37417 12173 37420
rect 12207 37417 12219 37451
rect 12161 37411 12219 37417
rect 12529 37451 12587 37457
rect 12529 37417 12541 37451
rect 12575 37448 12587 37451
rect 13173 37451 13231 37457
rect 13173 37448 13185 37451
rect 12575 37420 13185 37448
rect 12575 37417 12587 37420
rect 12529 37411 12587 37417
rect 13173 37417 13185 37420
rect 13219 37448 13231 37451
rect 13538 37448 13544 37460
rect 13219 37420 13544 37448
rect 13219 37417 13231 37420
rect 13173 37411 13231 37417
rect 13538 37408 13544 37420
rect 13596 37408 13602 37460
rect 15473 37451 15531 37457
rect 15473 37448 15485 37451
rect 14292 37420 15485 37448
rect 14292 37324 14320 37420
rect 15473 37417 15485 37420
rect 15519 37417 15531 37451
rect 15473 37411 15531 37417
rect 18046 37408 18052 37460
rect 18104 37448 18110 37460
rect 18141 37451 18199 37457
rect 18141 37448 18153 37451
rect 18104 37420 18153 37448
rect 18104 37408 18110 37420
rect 18141 37417 18153 37420
rect 18187 37417 18199 37451
rect 18414 37448 18420 37460
rect 18375 37420 18420 37448
rect 18141 37411 18199 37417
rect 18414 37408 18420 37420
rect 18472 37408 18478 37460
rect 18506 37408 18512 37460
rect 18564 37448 18570 37460
rect 20073 37451 20131 37457
rect 20073 37448 20085 37451
rect 18564 37420 20085 37448
rect 18564 37408 18570 37420
rect 20073 37417 20085 37420
rect 20119 37448 20131 37451
rect 20346 37448 20352 37460
rect 20119 37420 20352 37448
rect 20119 37417 20131 37420
rect 20073 37411 20131 37417
rect 20346 37408 20352 37420
rect 20404 37408 20410 37460
rect 20441 37451 20499 37457
rect 20441 37417 20453 37451
rect 20487 37448 20499 37451
rect 20806 37448 20812 37460
rect 20487 37420 20812 37448
rect 20487 37417 20499 37420
rect 20441 37411 20499 37417
rect 20806 37408 20812 37420
rect 20864 37408 20870 37460
rect 25133 37451 25191 37457
rect 25133 37417 25145 37451
rect 25179 37448 25191 37451
rect 25682 37448 25688 37460
rect 25179 37420 25688 37448
rect 25179 37417 25191 37420
rect 25133 37411 25191 37417
rect 25682 37408 25688 37420
rect 25740 37408 25746 37460
rect 27157 37451 27215 37457
rect 27157 37417 27169 37451
rect 27203 37448 27215 37451
rect 27246 37448 27252 37460
rect 27203 37420 27252 37448
rect 27203 37417 27215 37420
rect 27157 37411 27215 37417
rect 27246 37408 27252 37420
rect 27304 37408 27310 37460
rect 33502 37448 33508 37460
rect 33463 37420 33508 37448
rect 33502 37408 33508 37420
rect 33560 37408 33566 37460
rect 14734 37340 14740 37392
rect 14792 37380 14798 37392
rect 15746 37380 15752 37392
rect 14792 37352 15752 37380
rect 14792 37340 14798 37352
rect 15746 37340 15752 37352
rect 15804 37380 15810 37392
rect 16301 37383 16359 37389
rect 16301 37380 16313 37383
rect 15804 37352 16313 37380
rect 15804 37340 15810 37352
rect 16301 37349 16313 37352
rect 16347 37349 16359 37383
rect 17954 37380 17960 37392
rect 16301 37343 16359 37349
rect 16960 37352 17960 37380
rect 16960 37324 16988 37352
rect 17954 37340 17960 37352
rect 18012 37340 18018 37392
rect 19978 37380 19984 37392
rect 18524 37352 19984 37380
rect 9398 37272 9404 37324
rect 9456 37312 9462 37324
rect 10597 37315 10655 37321
rect 10597 37312 10609 37315
rect 9456 37284 10609 37312
rect 9456 37272 9462 37284
rect 10597 37281 10609 37284
rect 10643 37312 10655 37315
rect 10781 37315 10839 37321
rect 10781 37312 10793 37315
rect 10643 37284 10793 37312
rect 10643 37281 10655 37284
rect 10597 37275 10655 37281
rect 10781 37281 10793 37284
rect 10827 37281 10839 37315
rect 11054 37312 11060 37324
rect 11015 37284 11060 37312
rect 10781 37275 10839 37281
rect 11054 37272 11060 37284
rect 11112 37272 11118 37324
rect 13722 37312 13728 37324
rect 12360 37284 13728 37312
rect 11882 37204 11888 37256
rect 11940 37244 11946 37256
rect 12360 37244 12388 37284
rect 13722 37272 13728 37284
rect 13780 37272 13786 37324
rect 14185 37315 14243 37321
rect 14185 37281 14197 37315
rect 14231 37312 14243 37315
rect 14274 37312 14280 37324
rect 14231 37284 14280 37312
rect 14231 37281 14243 37284
rect 14185 37275 14243 37281
rect 14274 37272 14280 37284
rect 14332 37272 14338 37324
rect 15289 37315 15347 37321
rect 15289 37281 15301 37315
rect 15335 37312 15347 37315
rect 15378 37312 15384 37324
rect 15335 37284 15384 37312
rect 15335 37281 15347 37284
rect 15289 37275 15347 37281
rect 15378 37272 15384 37284
rect 15436 37272 15442 37324
rect 16114 37312 16120 37324
rect 16075 37284 16120 37312
rect 16114 37272 16120 37284
rect 16172 37272 16178 37324
rect 16942 37312 16948 37324
rect 16903 37284 16948 37312
rect 16942 37272 16948 37284
rect 17000 37272 17006 37324
rect 17310 37312 17316 37324
rect 17271 37284 17316 37312
rect 17310 37272 17316 37284
rect 17368 37272 17374 37324
rect 17865 37315 17923 37321
rect 17865 37281 17877 37315
rect 17911 37312 17923 37315
rect 18230 37312 18236 37324
rect 17911 37284 18236 37312
rect 17911 37281 17923 37284
rect 17865 37275 17923 37281
rect 18230 37272 18236 37284
rect 18288 37272 18294 37324
rect 18524 37321 18552 37352
rect 19978 37340 19984 37352
rect 20036 37340 20042 37392
rect 18509 37315 18567 37321
rect 18509 37281 18521 37315
rect 18555 37281 18567 37315
rect 18966 37312 18972 37324
rect 18927 37284 18972 37312
rect 18509 37275 18567 37281
rect 18966 37272 18972 37284
rect 19024 37272 19030 37324
rect 19150 37312 19156 37324
rect 19111 37284 19156 37312
rect 19150 37272 19156 37284
rect 19208 37272 19214 37324
rect 23842 37272 23848 37324
rect 23900 37312 23906 37324
rect 24946 37312 24952 37324
rect 23900 37284 24952 37312
rect 23900 37272 23906 37284
rect 24946 37272 24952 37284
rect 25004 37272 25010 37324
rect 27430 37312 27436 37324
rect 27391 37284 27436 37312
rect 27430 37272 27436 37284
rect 27488 37272 27494 37324
rect 32214 37272 32220 37324
rect 32272 37312 32278 37324
rect 32401 37315 32459 37321
rect 32401 37312 32413 37315
rect 32272 37284 32413 37312
rect 32272 37272 32278 37284
rect 32401 37281 32413 37284
rect 32447 37281 32459 37315
rect 32401 37275 32459 37281
rect 11940 37216 12388 37244
rect 11940 37204 11946 37216
rect 13354 37204 13360 37256
rect 13412 37244 13418 37256
rect 13449 37247 13507 37253
rect 13449 37244 13461 37247
rect 13412 37216 13461 37244
rect 13412 37204 13418 37216
rect 13449 37213 13461 37216
rect 13495 37244 13507 37247
rect 14826 37244 14832 37256
rect 13495 37216 14832 37244
rect 13495 37213 13507 37216
rect 13449 37207 13507 37213
rect 14826 37204 14832 37216
rect 14884 37204 14890 37256
rect 16850 37244 16856 37256
rect 16811 37216 16856 37244
rect 16850 37204 16856 37216
rect 16908 37204 16914 37256
rect 17126 37204 17132 37256
rect 17184 37244 17190 37256
rect 17405 37247 17463 37253
rect 17405 37244 17417 37247
rect 17184 37216 17417 37244
rect 17184 37204 17190 37216
rect 17405 37213 17417 37216
rect 17451 37213 17463 37247
rect 23106 37244 23112 37256
rect 23067 37216 23112 37244
rect 17405 37207 17463 37213
rect 23106 37204 23112 37216
rect 23164 37204 23170 37256
rect 23290 37204 23296 37256
rect 23348 37244 23354 37256
rect 23385 37247 23443 37253
rect 23385 37244 23397 37247
rect 23348 37216 23397 37244
rect 23348 37204 23354 37216
rect 23385 37213 23397 37216
rect 23431 37213 23443 37247
rect 23385 37207 23443 37213
rect 32125 37247 32183 37253
rect 32125 37213 32137 37247
rect 32171 37244 32183 37247
rect 32490 37244 32496 37256
rect 32171 37216 32496 37244
rect 32171 37213 32183 37216
rect 32125 37207 32183 37213
rect 32490 37204 32496 37216
rect 32548 37204 32554 37256
rect 11790 37136 11796 37188
rect 11848 37176 11854 37188
rect 12529 37179 12587 37185
rect 12529 37176 12541 37179
rect 11848 37148 12541 37176
rect 11848 37136 11854 37148
rect 12529 37145 12541 37148
rect 12575 37145 12587 37179
rect 12529 37139 12587 37145
rect 14185 37179 14243 37185
rect 14185 37145 14197 37179
rect 14231 37176 14243 37179
rect 14366 37176 14372 37188
rect 14231 37148 14372 37176
rect 14231 37145 14243 37148
rect 14185 37139 14243 37145
rect 14366 37136 14372 37148
rect 14424 37136 14430 37188
rect 16206 37136 16212 37188
rect 16264 37176 16270 37188
rect 17586 37176 17592 37188
rect 16264 37148 17592 37176
rect 16264 37136 16270 37148
rect 17586 37136 17592 37148
rect 17644 37136 17650 37188
rect 12802 37108 12808 37120
rect 12763 37080 12808 37108
rect 12802 37068 12808 37080
rect 12860 37068 12866 37120
rect 14734 37108 14740 37120
rect 14695 37080 14740 37108
rect 14734 37068 14740 37080
rect 14792 37068 14798 37120
rect 15105 37111 15163 37117
rect 15105 37077 15117 37111
rect 15151 37108 15163 37111
rect 15654 37108 15660 37120
rect 15151 37080 15660 37108
rect 15151 37077 15163 37080
rect 15105 37071 15163 37077
rect 15654 37068 15660 37080
rect 15712 37068 15718 37120
rect 24210 37068 24216 37120
rect 24268 37108 24274 37120
rect 24489 37111 24547 37117
rect 24489 37108 24501 37111
rect 24268 37080 24501 37108
rect 24268 37068 24274 37080
rect 24489 37077 24501 37080
rect 24535 37077 24547 37111
rect 24489 37071 24547 37077
rect 1104 37018 38824 37040
rect 1104 36966 4246 37018
rect 4298 36966 4310 37018
rect 4362 36966 4374 37018
rect 4426 36966 4438 37018
rect 4490 36966 34966 37018
rect 35018 36966 35030 37018
rect 35082 36966 35094 37018
rect 35146 36966 35158 37018
rect 35210 36966 38824 37018
rect 1104 36944 38824 36966
rect 9953 36907 10011 36913
rect 9953 36873 9965 36907
rect 9999 36904 10011 36907
rect 11054 36904 11060 36916
rect 9999 36876 11060 36904
rect 9999 36873 10011 36876
rect 9953 36867 10011 36873
rect 11054 36864 11060 36876
rect 11112 36864 11118 36916
rect 12710 36864 12716 36916
rect 12768 36904 12774 36916
rect 13170 36904 13176 36916
rect 12768 36876 13176 36904
rect 12768 36864 12774 36876
rect 13170 36864 13176 36876
rect 13228 36864 13234 36916
rect 14458 36864 14464 36916
rect 14516 36904 14522 36916
rect 14734 36904 14740 36916
rect 14516 36876 14740 36904
rect 14516 36864 14522 36876
rect 14734 36864 14740 36876
rect 14792 36864 14798 36916
rect 15378 36864 15384 36916
rect 15436 36904 15442 36916
rect 16022 36904 16028 36916
rect 15436 36876 16028 36904
rect 15436 36864 15442 36876
rect 16022 36864 16028 36876
rect 16080 36904 16086 36916
rect 16209 36907 16267 36913
rect 16209 36904 16221 36907
rect 16080 36876 16221 36904
rect 16080 36864 16086 36876
rect 16209 36873 16221 36876
rect 16255 36873 16267 36907
rect 16209 36867 16267 36873
rect 16669 36907 16727 36913
rect 16669 36873 16681 36907
rect 16715 36904 16727 36907
rect 17126 36904 17132 36916
rect 16715 36876 17132 36904
rect 16715 36873 16727 36876
rect 16669 36867 16727 36873
rect 17126 36864 17132 36876
rect 17184 36864 17190 36916
rect 17497 36907 17555 36913
rect 17497 36873 17509 36907
rect 17543 36904 17555 36907
rect 17770 36904 17776 36916
rect 17543 36876 17776 36904
rect 17543 36873 17555 36876
rect 17497 36867 17555 36873
rect 11422 36796 11428 36848
rect 11480 36836 11486 36848
rect 14369 36839 14427 36845
rect 14369 36836 14381 36839
rect 11480 36808 14381 36836
rect 11480 36796 11486 36808
rect 14369 36805 14381 36808
rect 14415 36836 14427 36839
rect 15102 36836 15108 36848
rect 14415 36808 15108 36836
rect 14415 36805 14427 36808
rect 14369 36799 14427 36805
rect 15102 36796 15108 36808
rect 15160 36836 15166 36848
rect 15160 36808 15884 36836
rect 15160 36796 15166 36808
rect 11517 36771 11575 36777
rect 11517 36737 11529 36771
rect 11563 36768 11575 36771
rect 11790 36768 11796 36780
rect 11563 36740 11796 36768
rect 11563 36737 11575 36740
rect 11517 36731 11575 36737
rect 11790 36728 11796 36740
rect 11848 36728 11854 36780
rect 12253 36771 12311 36777
rect 12253 36737 12265 36771
rect 12299 36768 12311 36771
rect 12299 36740 12756 36768
rect 12299 36737 12311 36740
rect 12253 36731 12311 36737
rect 10873 36703 10931 36709
rect 10873 36700 10885 36703
rect 10244 36672 10885 36700
rect 10134 36524 10140 36576
rect 10192 36564 10198 36576
rect 10244 36573 10272 36672
rect 10873 36669 10885 36672
rect 10919 36669 10931 36703
rect 10873 36663 10931 36669
rect 11885 36703 11943 36709
rect 11885 36669 11897 36703
rect 11931 36700 11943 36703
rect 12618 36700 12624 36712
rect 11931 36672 12624 36700
rect 11931 36669 11943 36672
rect 11885 36663 11943 36669
rect 12618 36660 12624 36672
rect 12676 36660 12682 36712
rect 12728 36700 12756 36740
rect 12802 36728 12808 36780
rect 12860 36768 12866 36780
rect 13541 36771 13599 36777
rect 13541 36768 13553 36771
rect 12860 36740 13553 36768
rect 12860 36728 12866 36740
rect 13541 36737 13553 36740
rect 13587 36737 13599 36771
rect 13541 36731 13599 36737
rect 14461 36771 14519 36777
rect 14461 36737 14473 36771
rect 14507 36768 14519 36771
rect 14642 36768 14648 36780
rect 14507 36740 14648 36768
rect 14507 36737 14519 36740
rect 14461 36731 14519 36737
rect 14642 36728 14648 36740
rect 14700 36728 14706 36780
rect 15856 36777 15884 36808
rect 15841 36771 15899 36777
rect 15841 36737 15853 36771
rect 15887 36737 15899 36771
rect 15841 36731 15899 36737
rect 13354 36700 13360 36712
rect 12728 36672 13360 36700
rect 13354 36660 13360 36672
rect 13412 36700 13418 36712
rect 13449 36703 13507 36709
rect 13449 36700 13461 36703
rect 13412 36672 13461 36700
rect 13412 36660 13418 36672
rect 13449 36669 13461 36672
rect 13495 36669 13507 36703
rect 14918 36700 14924 36712
rect 14879 36672 14924 36700
rect 13449 36663 13507 36669
rect 14918 36660 14924 36672
rect 14976 36660 14982 36712
rect 15194 36700 15200 36712
rect 15155 36672 15200 36700
rect 15194 36660 15200 36672
rect 15252 36660 15258 36712
rect 15289 36703 15347 36709
rect 15289 36669 15301 36703
rect 15335 36669 15347 36703
rect 15654 36700 15660 36712
rect 15615 36672 15660 36700
rect 15289 36663 15347 36669
rect 12713 36635 12771 36641
rect 12713 36601 12725 36635
rect 12759 36632 12771 36635
rect 13630 36632 13636 36644
rect 12759 36604 13636 36632
rect 12759 36601 12771 36604
rect 12713 36595 12771 36601
rect 13630 36592 13636 36604
rect 13688 36592 13694 36644
rect 14001 36635 14059 36641
rect 14001 36601 14013 36635
rect 14047 36632 14059 36635
rect 14458 36632 14464 36644
rect 14047 36604 14464 36632
rect 14047 36601 14059 36604
rect 14001 36595 14059 36601
rect 14458 36592 14464 36604
rect 14516 36592 14522 36644
rect 15010 36592 15016 36644
rect 15068 36632 15074 36644
rect 15304 36632 15332 36663
rect 15654 36660 15660 36672
rect 15712 36660 15718 36712
rect 16945 36703 17003 36709
rect 16945 36669 16957 36703
rect 16991 36700 17003 36703
rect 17512 36700 17540 36867
rect 17770 36864 17776 36876
rect 17828 36864 17834 36916
rect 19978 36864 19984 36916
rect 20036 36904 20042 36916
rect 20165 36907 20223 36913
rect 20165 36904 20177 36907
rect 20036 36876 20177 36904
rect 20036 36864 20042 36876
rect 20165 36873 20177 36876
rect 20211 36873 20223 36907
rect 20165 36867 20223 36873
rect 20254 36864 20260 36916
rect 20312 36904 20318 36916
rect 20533 36907 20591 36913
rect 20533 36904 20545 36907
rect 20312 36876 20545 36904
rect 20312 36864 20318 36876
rect 20533 36873 20545 36876
rect 20579 36873 20591 36907
rect 21634 36904 21640 36916
rect 21595 36876 21640 36904
rect 20533 36867 20591 36873
rect 21634 36864 21640 36876
rect 21692 36864 21698 36916
rect 23201 36907 23259 36913
rect 23201 36873 23213 36907
rect 23247 36904 23259 36907
rect 23290 36904 23296 36916
rect 23247 36876 23296 36904
rect 23247 36873 23259 36876
rect 23201 36867 23259 36873
rect 23290 36864 23296 36876
rect 23348 36864 23354 36916
rect 26786 36904 26792 36916
rect 26747 36876 26792 36904
rect 26786 36864 26792 36876
rect 26844 36864 26850 36916
rect 27430 36904 27436 36916
rect 27391 36876 27436 36904
rect 27430 36864 27436 36876
rect 27488 36864 27494 36916
rect 32490 36904 32496 36916
rect 32451 36876 32496 36904
rect 32490 36864 32496 36876
rect 32548 36864 32554 36916
rect 25317 36771 25375 36777
rect 25317 36737 25329 36771
rect 25363 36768 25375 36771
rect 25363 36740 25728 36768
rect 25363 36737 25375 36740
rect 25317 36731 25375 36737
rect 25700 36712 25728 36740
rect 18230 36700 18236 36712
rect 16991 36672 17540 36700
rect 18191 36672 18236 36700
rect 16991 36669 17003 36672
rect 16945 36663 17003 36669
rect 18230 36660 18236 36672
rect 18288 36660 18294 36712
rect 18785 36703 18843 36709
rect 18785 36669 18797 36703
rect 18831 36669 18843 36703
rect 18785 36663 18843 36669
rect 17402 36632 17408 36644
rect 15068 36604 15332 36632
rect 17144 36604 17408 36632
rect 15068 36592 15074 36604
rect 10229 36567 10287 36573
rect 10229 36564 10241 36567
rect 10192 36536 10241 36564
rect 10192 36524 10198 36536
rect 10229 36533 10241 36536
rect 10275 36533 10287 36567
rect 10594 36564 10600 36576
rect 10555 36536 10600 36564
rect 10229 36527 10287 36533
rect 10594 36524 10600 36536
rect 10652 36524 10658 36576
rect 17144 36573 17172 36604
rect 17402 36592 17408 36604
rect 17460 36592 17466 36644
rect 17586 36592 17592 36644
rect 17644 36632 17650 36644
rect 17865 36635 17923 36641
rect 17865 36632 17877 36635
rect 17644 36604 17877 36632
rect 17644 36592 17650 36604
rect 17865 36601 17877 36604
rect 17911 36632 17923 36635
rect 18800 36632 18828 36663
rect 18874 36660 18880 36712
rect 18932 36700 18938 36712
rect 19061 36703 19119 36709
rect 19061 36700 19073 36703
rect 18932 36672 19073 36700
rect 18932 36660 18938 36672
rect 19061 36669 19073 36672
rect 19107 36700 19119 36703
rect 25406 36700 25412 36712
rect 19107 36672 19564 36700
rect 25367 36672 25412 36700
rect 19107 36669 19119 36672
rect 19061 36663 19119 36669
rect 17911 36604 19104 36632
rect 17911 36601 17923 36604
rect 17865 36595 17923 36601
rect 19076 36576 19104 36604
rect 17129 36567 17187 36573
rect 17129 36533 17141 36567
rect 17175 36533 17187 36567
rect 17129 36527 17187 36533
rect 18141 36567 18199 36573
rect 18141 36533 18153 36567
rect 18187 36564 18199 36567
rect 18506 36564 18512 36576
rect 18187 36536 18512 36564
rect 18187 36533 18199 36536
rect 18141 36527 18199 36533
rect 18506 36524 18512 36536
rect 18564 36524 18570 36576
rect 19058 36524 19064 36576
rect 19116 36524 19122 36576
rect 19536 36573 19564 36672
rect 25406 36660 25412 36672
rect 25464 36660 25470 36712
rect 25682 36700 25688 36712
rect 25643 36672 25688 36700
rect 25682 36660 25688 36672
rect 25740 36660 25746 36712
rect 19521 36567 19579 36573
rect 19521 36533 19533 36567
rect 19567 36564 19579 36567
rect 19889 36567 19947 36573
rect 19889 36564 19901 36567
rect 19567 36536 19901 36564
rect 19567 36533 19579 36536
rect 19521 36527 19579 36533
rect 19889 36533 19901 36536
rect 19935 36564 19947 36567
rect 19978 36564 19984 36576
rect 19935 36536 19984 36564
rect 19935 36533 19947 36536
rect 19889 36527 19947 36533
rect 19978 36524 19984 36536
rect 20036 36524 20042 36576
rect 20898 36564 20904 36576
rect 20859 36536 20904 36564
rect 20898 36524 20904 36536
rect 20956 36524 20962 36576
rect 21174 36524 21180 36576
rect 21232 36564 21238 36576
rect 21269 36567 21327 36573
rect 21269 36564 21281 36567
rect 21232 36536 21281 36564
rect 21232 36524 21238 36536
rect 21269 36533 21281 36536
rect 21315 36533 21327 36567
rect 21269 36527 21327 36533
rect 23106 36524 23112 36576
rect 23164 36564 23170 36576
rect 23290 36564 23296 36576
rect 23164 36536 23296 36564
rect 23164 36524 23170 36536
rect 23290 36524 23296 36536
rect 23348 36564 23354 36576
rect 23845 36567 23903 36573
rect 23845 36564 23857 36567
rect 23348 36536 23857 36564
rect 23348 36524 23354 36536
rect 23845 36533 23857 36536
rect 23891 36533 23903 36567
rect 32122 36564 32128 36576
rect 32083 36536 32128 36564
rect 23845 36527 23903 36533
rect 32122 36524 32128 36536
rect 32180 36524 32186 36576
rect 1104 36474 38824 36496
rect 1104 36422 19606 36474
rect 19658 36422 19670 36474
rect 19722 36422 19734 36474
rect 19786 36422 19798 36474
rect 19850 36422 38824 36474
rect 1104 36400 38824 36422
rect 10962 36360 10968 36372
rect 10923 36332 10968 36360
rect 10962 36320 10968 36332
rect 11020 36320 11026 36372
rect 11609 36363 11667 36369
rect 11609 36329 11621 36363
rect 11655 36360 11667 36363
rect 11882 36360 11888 36372
rect 11655 36332 11888 36360
rect 11655 36329 11667 36332
rect 11609 36323 11667 36329
rect 11882 36320 11888 36332
rect 11940 36320 11946 36372
rect 12250 36320 12256 36372
rect 12308 36360 12314 36372
rect 13265 36363 13323 36369
rect 13265 36360 13277 36363
rect 12308 36332 13277 36360
rect 12308 36320 12314 36332
rect 13265 36329 13277 36332
rect 13311 36329 13323 36363
rect 14826 36360 14832 36372
rect 14787 36332 14832 36360
rect 13265 36323 13323 36329
rect 14826 36320 14832 36332
rect 14884 36320 14890 36372
rect 15378 36320 15384 36372
rect 15436 36360 15442 36372
rect 16666 36360 16672 36372
rect 15436 36332 16672 36360
rect 15436 36320 15442 36332
rect 16666 36320 16672 36332
rect 16724 36320 16730 36372
rect 17497 36363 17555 36369
rect 17497 36329 17509 36363
rect 17543 36360 17555 36363
rect 17862 36360 17868 36372
rect 17543 36332 17868 36360
rect 17543 36329 17555 36332
rect 17497 36323 17555 36329
rect 17862 36320 17868 36332
rect 17920 36320 17926 36372
rect 18230 36320 18236 36372
rect 18288 36360 18294 36372
rect 18601 36363 18659 36369
rect 18601 36360 18613 36363
rect 18288 36332 18613 36360
rect 18288 36320 18294 36332
rect 18601 36329 18613 36332
rect 18647 36329 18659 36363
rect 18966 36360 18972 36372
rect 18927 36332 18972 36360
rect 18601 36323 18659 36329
rect 18966 36320 18972 36332
rect 19024 36320 19030 36372
rect 23842 36320 23848 36372
rect 23900 36360 23906 36372
rect 24489 36363 24547 36369
rect 24489 36360 24501 36363
rect 23900 36332 24501 36360
rect 23900 36320 23906 36332
rect 24489 36329 24501 36332
rect 24535 36329 24547 36363
rect 29546 36360 29552 36372
rect 29507 36332 29552 36360
rect 24489 36323 24547 36329
rect 29546 36320 29552 36332
rect 29604 36320 29610 36372
rect 15289 36295 15347 36301
rect 15289 36261 15301 36295
rect 15335 36292 15347 36295
rect 15838 36292 15844 36304
rect 15335 36264 15844 36292
rect 15335 36261 15347 36264
rect 15289 36255 15347 36261
rect 15838 36252 15844 36264
rect 15896 36252 15902 36304
rect 17218 36252 17224 36304
rect 17276 36292 17282 36304
rect 17678 36292 17684 36304
rect 17276 36264 17684 36292
rect 17276 36252 17282 36264
rect 17678 36252 17684 36264
rect 17736 36252 17742 36304
rect 18322 36292 18328 36304
rect 18283 36264 18328 36292
rect 18322 36252 18328 36264
rect 18380 36252 18386 36304
rect 21729 36295 21787 36301
rect 21729 36292 21741 36295
rect 20088 36264 21741 36292
rect 11054 36224 11060 36236
rect 10967 36196 11060 36224
rect 11054 36184 11060 36196
rect 11112 36224 11118 36236
rect 11422 36224 11428 36236
rect 11112 36196 11428 36224
rect 11112 36184 11118 36196
rect 11422 36184 11428 36196
rect 11480 36184 11486 36236
rect 12158 36184 12164 36236
rect 12216 36224 12222 36236
rect 12253 36227 12311 36233
rect 12253 36224 12265 36227
rect 12216 36196 12265 36224
rect 12216 36184 12222 36196
rect 12253 36193 12265 36196
rect 12299 36224 12311 36227
rect 12802 36224 12808 36236
rect 12299 36196 12808 36224
rect 12299 36193 12311 36196
rect 12253 36187 12311 36193
rect 12802 36184 12808 36196
rect 12860 36184 12866 36236
rect 12986 36224 12992 36236
rect 12947 36196 12992 36224
rect 12986 36184 12992 36196
rect 13044 36184 13050 36236
rect 15746 36224 15752 36236
rect 15707 36196 15752 36224
rect 15746 36184 15752 36196
rect 15804 36184 15810 36236
rect 15930 36224 15936 36236
rect 15891 36196 15936 36224
rect 15930 36184 15936 36196
rect 15988 36184 15994 36236
rect 16117 36227 16175 36233
rect 16117 36193 16129 36227
rect 16163 36193 16175 36227
rect 16666 36224 16672 36236
rect 16627 36196 16672 36224
rect 16117 36187 16175 36193
rect 12069 36159 12127 36165
rect 12069 36156 12081 36159
rect 11992 36128 12081 36156
rect 11992 36088 12020 36128
rect 12069 36125 12081 36128
rect 12115 36125 12127 36159
rect 12069 36119 12127 36125
rect 14918 36116 14924 36168
rect 14976 36156 14982 36168
rect 16132 36156 16160 36187
rect 16666 36184 16672 36196
rect 16724 36184 16730 36236
rect 17402 36184 17408 36236
rect 17460 36224 17466 36236
rect 17589 36227 17647 36233
rect 17589 36224 17601 36227
rect 17460 36196 17601 36224
rect 17460 36184 17466 36196
rect 17589 36193 17601 36196
rect 17635 36193 17647 36227
rect 17589 36187 17647 36193
rect 17773 36227 17831 36233
rect 17773 36193 17785 36227
rect 17819 36193 17831 36227
rect 17773 36187 17831 36193
rect 14976 36128 16160 36156
rect 14976 36116 14982 36128
rect 16298 36116 16304 36168
rect 16356 36156 16362 36168
rect 16393 36159 16451 36165
rect 16393 36156 16405 36159
rect 16356 36128 16405 36156
rect 16356 36116 16362 36128
rect 16393 36125 16405 36128
rect 16439 36125 16451 36159
rect 17788 36156 17816 36187
rect 17862 36184 17868 36236
rect 17920 36224 17926 36236
rect 17920 36196 17965 36224
rect 17920 36184 17926 36196
rect 18874 36184 18880 36236
rect 18932 36224 18938 36236
rect 19153 36227 19211 36233
rect 19153 36224 19165 36227
rect 18932 36196 19165 36224
rect 18932 36184 18938 36196
rect 19153 36193 19165 36196
rect 19199 36193 19211 36227
rect 19153 36187 19211 36193
rect 19334 36184 19340 36236
rect 19392 36224 19398 36236
rect 20088 36224 20116 36264
rect 21729 36261 21741 36264
rect 21775 36261 21787 36295
rect 21729 36255 21787 36261
rect 19392 36196 20116 36224
rect 20901 36227 20959 36233
rect 19392 36184 19398 36196
rect 20901 36193 20913 36227
rect 20947 36224 20959 36227
rect 21174 36224 21180 36236
rect 20947 36196 21180 36224
rect 20947 36193 20959 36196
rect 20901 36187 20959 36193
rect 21174 36184 21180 36196
rect 21232 36184 21238 36236
rect 23382 36224 23388 36236
rect 23343 36196 23388 36224
rect 23382 36184 23388 36196
rect 23440 36184 23446 36236
rect 28169 36227 28227 36233
rect 28169 36193 28181 36227
rect 28215 36224 28227 36227
rect 28258 36224 28264 36236
rect 28215 36196 28264 36224
rect 28215 36193 28227 36196
rect 28169 36187 28227 36193
rect 28258 36184 28264 36196
rect 28316 36184 28322 36236
rect 19705 36159 19763 36165
rect 19705 36156 19717 36159
rect 17788 36128 19717 36156
rect 16393 36119 16451 36125
rect 19705 36125 19717 36128
rect 19751 36156 19763 36159
rect 21361 36159 21419 36165
rect 21361 36156 21373 36159
rect 19751 36128 21373 36156
rect 19751 36125 19763 36128
rect 19705 36119 19763 36125
rect 21361 36125 21373 36128
rect 21407 36125 21419 36159
rect 21361 36119 21419 36125
rect 22557 36159 22615 36165
rect 22557 36125 22569 36159
rect 22603 36156 22615 36159
rect 23109 36159 23167 36165
rect 23109 36156 23121 36159
rect 22603 36128 23121 36156
rect 22603 36125 22615 36128
rect 22557 36119 22615 36125
rect 23109 36125 23121 36128
rect 23155 36156 23167 36159
rect 23290 36156 23296 36168
rect 23155 36128 23296 36156
rect 23155 36125 23167 36128
rect 23109 36119 23167 36125
rect 23290 36116 23296 36128
rect 23348 36156 23354 36168
rect 25406 36156 25412 36168
rect 23348 36128 25412 36156
rect 23348 36116 23354 36128
rect 25406 36116 25412 36128
rect 25464 36116 25470 36168
rect 28442 36156 28448 36168
rect 28403 36128 28448 36156
rect 28442 36116 28448 36128
rect 28500 36116 28506 36168
rect 16758 36088 16764 36100
rect 11992 36060 16764 36088
rect 11992 36032 12020 36060
rect 16758 36048 16764 36060
rect 16816 36088 16822 36100
rect 17678 36088 17684 36100
rect 16816 36060 17684 36088
rect 16816 36048 16822 36060
rect 17678 36048 17684 36060
rect 17736 36048 17742 36100
rect 19242 36048 19248 36100
rect 19300 36088 19306 36100
rect 20349 36091 20407 36097
rect 20349 36088 20361 36091
rect 19300 36060 20361 36088
rect 19300 36048 19306 36060
rect 20349 36057 20361 36060
rect 20395 36057 20407 36091
rect 20349 36051 20407 36057
rect 11241 36023 11299 36029
rect 11241 35989 11253 36023
rect 11287 36020 11299 36023
rect 11422 36020 11428 36032
rect 11287 35992 11428 36020
rect 11287 35989 11299 35992
rect 11241 35983 11299 35989
rect 11422 35980 11428 35992
rect 11480 35980 11486 36032
rect 11974 36020 11980 36032
rect 11935 35992 11980 36020
rect 11974 35980 11980 35992
rect 12032 35980 12038 36032
rect 14001 36023 14059 36029
rect 14001 35989 14013 36023
rect 14047 36020 14059 36023
rect 14553 36023 14611 36029
rect 14553 36020 14565 36023
rect 14047 35992 14565 36020
rect 14047 35989 14059 35992
rect 14001 35983 14059 35989
rect 14553 35989 14565 35992
rect 14599 36020 14611 36023
rect 14918 36020 14924 36032
rect 14599 35992 14924 36020
rect 14599 35989 14611 35992
rect 14553 35983 14611 35989
rect 14918 35980 14924 35992
rect 14976 35980 14982 36032
rect 16942 35980 16948 36032
rect 17000 36020 17006 36032
rect 17037 36023 17095 36029
rect 17037 36020 17049 36023
rect 17000 35992 17049 36020
rect 17000 35980 17006 35992
rect 17037 35989 17049 35992
rect 17083 35989 17095 36023
rect 17037 35983 17095 35989
rect 18230 35980 18236 36032
rect 18288 36020 18294 36032
rect 19150 36020 19156 36032
rect 18288 35992 19156 36020
rect 18288 35980 18294 35992
rect 19150 35980 19156 35992
rect 19208 35980 19214 36032
rect 19426 35980 19432 36032
rect 19484 36020 19490 36032
rect 19981 36023 20039 36029
rect 19981 36020 19993 36023
rect 19484 35992 19993 36020
rect 19484 35980 19490 35992
rect 19981 35989 19993 35992
rect 20027 35989 20039 36023
rect 21082 36020 21088 36032
rect 21043 35992 21088 36020
rect 19981 35983 20039 35989
rect 21082 35980 21088 35992
rect 21140 35980 21146 36032
rect 21174 35980 21180 36032
rect 21232 36020 21238 36032
rect 22097 36023 22155 36029
rect 22097 36020 22109 36023
rect 21232 35992 22109 36020
rect 21232 35980 21238 35992
rect 22097 35989 22109 35992
rect 22143 36020 22155 36023
rect 24210 36020 24216 36032
rect 22143 35992 24216 36020
rect 22143 35989 22155 35992
rect 22097 35983 22155 35989
rect 24210 35980 24216 35992
rect 24268 35980 24274 36032
rect 1104 35930 38824 35952
rect 1104 35878 4246 35930
rect 4298 35878 4310 35930
rect 4362 35878 4374 35930
rect 4426 35878 4438 35930
rect 4490 35878 34966 35930
rect 35018 35878 35030 35930
rect 35082 35878 35094 35930
rect 35146 35878 35158 35930
rect 35210 35878 38824 35930
rect 1104 35856 38824 35878
rect 10778 35816 10784 35828
rect 10739 35788 10784 35816
rect 10778 35776 10784 35788
rect 10836 35776 10842 35828
rect 11054 35816 11060 35828
rect 11015 35788 11060 35816
rect 11054 35776 11060 35788
rect 11112 35776 11118 35828
rect 11422 35776 11428 35828
rect 11480 35816 11486 35828
rect 11701 35819 11759 35825
rect 11701 35816 11713 35819
rect 11480 35788 11713 35816
rect 11480 35776 11486 35788
rect 11701 35785 11713 35788
rect 11747 35816 11759 35819
rect 12069 35819 12127 35825
rect 12069 35816 12081 35819
rect 11747 35788 12081 35816
rect 11747 35785 11759 35788
rect 11701 35779 11759 35785
rect 12069 35785 12081 35788
rect 12115 35816 12127 35819
rect 12158 35816 12164 35828
rect 12115 35788 12164 35816
rect 12115 35785 12127 35788
rect 12069 35779 12127 35785
rect 12158 35776 12164 35788
rect 12216 35776 12222 35828
rect 12618 35776 12624 35828
rect 12676 35816 12682 35828
rect 12805 35819 12863 35825
rect 12805 35816 12817 35819
rect 12676 35788 12817 35816
rect 12676 35776 12682 35788
rect 12805 35785 12817 35788
rect 12851 35785 12863 35819
rect 12805 35779 12863 35785
rect 13354 35776 13360 35828
rect 13412 35816 13418 35828
rect 13725 35819 13783 35825
rect 13725 35816 13737 35819
rect 13412 35788 13737 35816
rect 13412 35776 13418 35788
rect 13725 35785 13737 35788
rect 13771 35816 13783 35819
rect 14090 35816 14096 35828
rect 13771 35788 14096 35816
rect 13771 35785 13783 35788
rect 13725 35779 13783 35785
rect 14090 35776 14096 35788
rect 14148 35776 14154 35828
rect 16022 35816 16028 35828
rect 15983 35788 16028 35816
rect 16022 35776 16028 35788
rect 16080 35816 16086 35828
rect 16347 35819 16405 35825
rect 16347 35816 16359 35819
rect 16080 35788 16359 35816
rect 16080 35776 16086 35788
rect 16347 35785 16359 35788
rect 16393 35785 16405 35819
rect 16482 35816 16488 35828
rect 16443 35788 16488 35816
rect 16347 35779 16405 35785
rect 16482 35776 16488 35788
rect 16540 35776 16546 35828
rect 16666 35816 16672 35828
rect 16627 35788 16672 35816
rect 16666 35776 16672 35788
rect 16724 35776 16730 35828
rect 16758 35776 16764 35828
rect 16816 35816 16822 35828
rect 17313 35819 17371 35825
rect 17313 35816 17325 35819
rect 16816 35788 17325 35816
rect 16816 35776 16822 35788
rect 17313 35785 17325 35788
rect 17359 35785 17371 35819
rect 17313 35779 17371 35785
rect 17402 35776 17408 35828
rect 17460 35816 17466 35828
rect 17681 35819 17739 35825
rect 17681 35816 17693 35819
rect 17460 35788 17693 35816
rect 17460 35776 17466 35788
rect 17681 35785 17693 35788
rect 17727 35816 17739 35819
rect 17865 35819 17923 35825
rect 17865 35816 17877 35819
rect 17727 35788 17877 35816
rect 17727 35785 17739 35788
rect 17681 35779 17739 35785
rect 17865 35785 17877 35788
rect 17911 35785 17923 35819
rect 17865 35779 17923 35785
rect 17954 35776 17960 35828
rect 18012 35816 18018 35828
rect 18509 35819 18567 35825
rect 18509 35816 18521 35819
rect 18012 35788 18521 35816
rect 18012 35776 18018 35788
rect 18509 35785 18521 35788
rect 18555 35785 18567 35819
rect 18509 35779 18567 35785
rect 23201 35819 23259 35825
rect 23201 35785 23213 35819
rect 23247 35816 23259 35819
rect 23382 35816 23388 35828
rect 23247 35788 23388 35816
rect 23247 35785 23259 35788
rect 23201 35779 23259 35785
rect 23382 35776 23388 35788
rect 23440 35776 23446 35828
rect 28258 35776 28264 35828
rect 28316 35816 28322 35828
rect 28537 35819 28595 35825
rect 28537 35816 28549 35819
rect 28316 35788 28549 35816
rect 28316 35776 28322 35788
rect 28537 35785 28549 35788
rect 28583 35785 28595 35819
rect 28537 35779 28595 35785
rect 13262 35708 13268 35760
rect 13320 35708 13326 35760
rect 13906 35708 13912 35760
rect 13964 35748 13970 35760
rect 15838 35748 15844 35760
rect 13964 35720 15844 35748
rect 13964 35708 13970 35720
rect 15838 35708 15844 35720
rect 15896 35708 15902 35760
rect 20441 35751 20499 35757
rect 20441 35748 20453 35751
rect 16500 35720 20453 35748
rect 10413 35683 10471 35689
rect 10413 35649 10425 35683
rect 10459 35680 10471 35683
rect 10962 35680 10968 35692
rect 10459 35652 10968 35680
rect 10459 35649 10471 35652
rect 10413 35643 10471 35649
rect 10962 35640 10968 35652
rect 11020 35640 11026 35692
rect 11054 35640 11060 35692
rect 11112 35680 11118 35692
rect 13280 35680 13308 35708
rect 11112 35652 13308 35680
rect 11112 35640 11118 35652
rect 14090 35640 14096 35692
rect 14148 35680 14154 35692
rect 15013 35683 15071 35689
rect 15013 35680 15025 35683
rect 14148 35652 15025 35680
rect 14148 35640 14154 35652
rect 15013 35649 15025 35652
rect 15059 35649 15071 35683
rect 15286 35680 15292 35692
rect 15247 35652 15292 35680
rect 15013 35643 15071 35649
rect 15286 35640 15292 35652
rect 15344 35640 15350 35692
rect 16500 35680 16528 35720
rect 20441 35717 20453 35720
rect 20487 35717 20499 35751
rect 20441 35711 20499 35717
rect 16224 35652 16528 35680
rect 16577 35683 16635 35689
rect 12713 35615 12771 35621
rect 12713 35581 12725 35615
rect 12759 35612 12771 35615
rect 13262 35612 13268 35624
rect 12759 35584 13268 35612
rect 12759 35581 12771 35584
rect 12713 35575 12771 35581
rect 13262 35572 13268 35584
rect 13320 35612 13326 35624
rect 13357 35615 13415 35621
rect 13357 35612 13369 35615
rect 13320 35584 13369 35612
rect 13320 35572 13326 35584
rect 13357 35581 13369 35584
rect 13403 35581 13415 35615
rect 14366 35612 14372 35624
rect 14327 35584 14372 35612
rect 13357 35575 13415 35581
rect 14366 35572 14372 35584
rect 14424 35572 14430 35624
rect 14458 35572 14464 35624
rect 14516 35612 14522 35624
rect 14553 35615 14611 35621
rect 14553 35612 14565 35615
rect 14516 35584 14565 35612
rect 14516 35572 14522 35584
rect 14553 35581 14565 35584
rect 14599 35581 14611 35615
rect 14553 35575 14611 35581
rect 14829 35615 14887 35621
rect 14829 35581 14841 35615
rect 14875 35612 14887 35615
rect 14918 35612 14924 35624
rect 14875 35584 14924 35612
rect 14875 35581 14887 35584
rect 14829 35575 14887 35581
rect 14918 35572 14924 35584
rect 14976 35572 14982 35624
rect 12526 35544 12532 35556
rect 12487 35516 12532 35544
rect 12526 35504 12532 35516
rect 12584 35504 12590 35556
rect 13906 35544 13912 35556
rect 13867 35516 13912 35544
rect 13906 35504 13912 35516
rect 13964 35504 13970 35556
rect 15194 35504 15200 35556
rect 15252 35544 15258 35556
rect 16224 35553 16252 35652
rect 16577 35649 16589 35683
rect 16623 35649 16635 35683
rect 16577 35643 16635 35649
rect 17865 35683 17923 35689
rect 17865 35649 17877 35683
rect 17911 35680 17923 35683
rect 17954 35680 17960 35692
rect 17911 35652 17960 35680
rect 17911 35649 17923 35652
rect 17865 35643 17923 35649
rect 16209 35547 16267 35553
rect 16209 35544 16221 35547
rect 15252 35516 16221 35544
rect 15252 35504 15258 35516
rect 16209 35513 16221 35516
rect 16255 35513 16267 35547
rect 16209 35507 16267 35513
rect 16592 35544 16620 35643
rect 17954 35640 17960 35652
rect 18012 35680 18018 35692
rect 18049 35683 18107 35689
rect 18049 35680 18061 35683
rect 18012 35652 18061 35680
rect 18012 35640 18018 35652
rect 18049 35649 18061 35652
rect 18095 35649 18107 35683
rect 19426 35680 19432 35692
rect 18049 35643 18107 35649
rect 18248 35652 19432 35680
rect 18248 35621 18276 35652
rect 19426 35640 19432 35652
rect 19484 35640 19490 35692
rect 20901 35683 20959 35689
rect 20901 35649 20913 35683
rect 20947 35680 20959 35683
rect 23290 35680 23296 35692
rect 20947 35652 23296 35680
rect 20947 35649 20959 35652
rect 20901 35643 20959 35649
rect 23290 35640 23296 35652
rect 23348 35640 23354 35692
rect 18233 35615 18291 35621
rect 18233 35581 18245 35615
rect 18279 35581 18291 35615
rect 18233 35575 18291 35581
rect 18322 35572 18328 35624
rect 18380 35612 18386 35624
rect 19242 35612 19248 35624
rect 18380 35584 19248 35612
rect 18380 35572 18386 35584
rect 19242 35572 19248 35584
rect 19300 35572 19306 35624
rect 19613 35615 19671 35621
rect 19613 35581 19625 35615
rect 19659 35612 19671 35615
rect 21174 35612 21180 35624
rect 19659 35584 20208 35612
rect 21135 35584 21180 35612
rect 19659 35581 19671 35584
rect 19613 35575 19671 35581
rect 19886 35544 19892 35556
rect 16592 35516 19892 35544
rect 10045 35479 10103 35485
rect 10045 35445 10057 35479
rect 10091 35476 10103 35479
rect 10134 35476 10140 35488
rect 10091 35448 10140 35476
rect 10091 35445 10103 35448
rect 10045 35439 10103 35445
rect 10134 35436 10140 35448
rect 10192 35436 10198 35488
rect 15749 35479 15807 35485
rect 15749 35445 15761 35479
rect 15795 35476 15807 35479
rect 16592 35476 16620 35516
rect 19886 35504 19892 35516
rect 19944 35504 19950 35556
rect 20180 35553 20208 35584
rect 21174 35572 21180 35584
rect 21232 35572 21238 35624
rect 20165 35547 20223 35553
rect 20165 35513 20177 35547
rect 20211 35544 20223 35547
rect 20622 35544 20628 35556
rect 20211 35516 20628 35544
rect 20211 35513 20223 35516
rect 20165 35507 20223 35513
rect 20622 35504 20628 35516
rect 20680 35504 20686 35556
rect 22554 35544 22560 35556
rect 22515 35516 22560 35544
rect 22554 35504 22560 35516
rect 22612 35504 22618 35556
rect 28261 35547 28319 35553
rect 28261 35513 28273 35547
rect 28307 35544 28319 35547
rect 28442 35544 28448 35556
rect 28307 35516 28448 35544
rect 28307 35513 28319 35516
rect 28261 35507 28319 35513
rect 28442 35504 28448 35516
rect 28500 35544 28506 35556
rect 28810 35544 28816 35556
rect 28500 35516 28816 35544
rect 28500 35504 28506 35516
rect 28810 35504 28816 35516
rect 28868 35504 28874 35556
rect 15795 35448 16620 35476
rect 15795 35445 15807 35448
rect 15749 35439 15807 35445
rect 18874 35436 18880 35488
rect 18932 35476 18938 35488
rect 19153 35479 19211 35485
rect 19153 35476 19165 35479
rect 18932 35448 19165 35476
rect 18932 35436 18938 35448
rect 19153 35445 19165 35448
rect 19199 35476 19211 35479
rect 19797 35479 19855 35485
rect 19797 35476 19809 35479
rect 19199 35448 19809 35476
rect 19199 35445 19211 35448
rect 19153 35439 19211 35445
rect 19797 35445 19809 35448
rect 19843 35445 19855 35479
rect 23934 35476 23940 35488
rect 23895 35448 23940 35476
rect 19797 35439 19855 35445
rect 23934 35436 23940 35448
rect 23992 35436 23998 35488
rect 1104 35386 38824 35408
rect 1104 35334 19606 35386
rect 19658 35334 19670 35386
rect 19722 35334 19734 35386
rect 19786 35334 19798 35386
rect 19850 35334 38824 35386
rect 1104 35312 38824 35334
rect 1670 35232 1676 35284
rect 1728 35272 1734 35284
rect 1765 35275 1823 35281
rect 1765 35272 1777 35275
rect 1728 35244 1777 35272
rect 1728 35232 1734 35244
rect 1765 35241 1777 35244
rect 1811 35272 1823 35275
rect 1946 35272 1952 35284
rect 1811 35244 1952 35272
rect 1811 35241 1823 35244
rect 1765 35235 1823 35241
rect 1946 35232 1952 35244
rect 2004 35232 2010 35284
rect 11330 35272 11336 35284
rect 11291 35244 11336 35272
rect 11330 35232 11336 35244
rect 11388 35232 11394 35284
rect 11698 35272 11704 35284
rect 11659 35244 11704 35272
rect 11698 35232 11704 35244
rect 11756 35232 11762 35284
rect 12526 35232 12532 35284
rect 12584 35272 12590 35284
rect 13081 35275 13139 35281
rect 13081 35272 13093 35275
rect 12584 35244 13093 35272
rect 12584 35232 12590 35244
rect 13081 35241 13093 35244
rect 13127 35272 13139 35275
rect 13722 35272 13728 35284
rect 13127 35244 13728 35272
rect 13127 35241 13139 35244
rect 13081 35235 13139 35241
rect 13722 35232 13728 35244
rect 13780 35232 13786 35284
rect 17497 35275 17555 35281
rect 17497 35241 17509 35275
rect 17543 35272 17555 35275
rect 17586 35272 17592 35284
rect 17543 35244 17592 35272
rect 17543 35241 17555 35244
rect 17497 35235 17555 35241
rect 17586 35232 17592 35244
rect 17644 35232 17650 35284
rect 17954 35232 17960 35284
rect 18012 35272 18018 35284
rect 18325 35275 18383 35281
rect 18325 35272 18337 35275
rect 18012 35244 18337 35272
rect 18012 35232 18018 35244
rect 18325 35241 18337 35244
rect 18371 35241 18383 35275
rect 18325 35235 18383 35241
rect 19334 35232 19340 35284
rect 19392 35272 19398 35284
rect 19705 35275 19763 35281
rect 19705 35272 19717 35275
rect 19392 35244 19717 35272
rect 19392 35232 19398 35244
rect 19705 35241 19717 35244
rect 19751 35241 19763 35275
rect 19705 35235 19763 35241
rect 21177 35275 21235 35281
rect 21177 35241 21189 35275
rect 21223 35272 21235 35275
rect 21266 35272 21272 35284
rect 21223 35244 21272 35272
rect 21223 35241 21235 35244
rect 21177 35235 21235 35241
rect 21266 35232 21272 35244
rect 21324 35232 21330 35284
rect 22646 35232 22652 35284
rect 22704 35272 22710 35284
rect 22741 35275 22799 35281
rect 22741 35272 22753 35275
rect 22704 35244 22753 35272
rect 22704 35232 22710 35244
rect 22741 35241 22753 35244
rect 22787 35272 22799 35275
rect 23382 35272 23388 35284
rect 22787 35244 23388 35272
rect 22787 35241 22799 35244
rect 22741 35235 22799 35241
rect 23382 35232 23388 35244
rect 23440 35232 23446 35284
rect 10597 35207 10655 35213
rect 10597 35173 10609 35207
rect 10643 35204 10655 35207
rect 10643 35176 12112 35204
rect 10643 35173 10655 35176
rect 10597 35167 10655 35173
rect 10229 35139 10287 35145
rect 10229 35105 10241 35139
rect 10275 35136 10287 35139
rect 11882 35136 11888 35148
rect 10275 35108 11888 35136
rect 10275 35105 10287 35108
rect 10229 35099 10287 35105
rect 11882 35096 11888 35108
rect 11940 35096 11946 35148
rect 12084 35136 12112 35176
rect 12250 35164 12256 35216
rect 12308 35204 12314 35216
rect 12345 35207 12403 35213
rect 12345 35204 12357 35207
rect 12308 35176 12357 35204
rect 12308 35164 12314 35176
rect 12345 35173 12357 35176
rect 12391 35173 12403 35207
rect 12345 35167 12403 35173
rect 12437 35207 12495 35213
rect 12437 35173 12449 35207
rect 12483 35204 12495 35207
rect 12713 35207 12771 35213
rect 12713 35204 12725 35207
rect 12483 35176 12725 35204
rect 12483 35173 12495 35176
rect 12437 35167 12495 35173
rect 12713 35173 12725 35176
rect 12759 35204 12771 35207
rect 12986 35204 12992 35216
rect 12759 35176 12992 35204
rect 12759 35173 12771 35176
rect 12713 35167 12771 35173
rect 12986 35164 12992 35176
rect 13044 35164 13050 35216
rect 13173 35207 13231 35213
rect 13173 35173 13185 35207
rect 13219 35204 13231 35207
rect 13538 35204 13544 35216
rect 13219 35176 13544 35204
rect 13219 35173 13231 35176
rect 13173 35167 13231 35173
rect 13538 35164 13544 35176
rect 13596 35164 13602 35216
rect 14458 35164 14464 35216
rect 14516 35204 14522 35216
rect 15289 35207 15347 35213
rect 15289 35204 15301 35207
rect 14516 35176 15301 35204
rect 14516 35164 14522 35176
rect 15289 35173 15301 35176
rect 15335 35173 15347 35207
rect 16761 35207 16819 35213
rect 16761 35204 16773 35207
rect 15289 35167 15347 35173
rect 15948 35176 16773 35204
rect 15948 35148 15976 35176
rect 16761 35173 16773 35176
rect 16807 35173 16819 35207
rect 17678 35204 17684 35216
rect 17639 35176 17684 35204
rect 16761 35167 16819 35173
rect 17678 35164 17684 35176
rect 17736 35164 17742 35216
rect 18046 35204 18052 35216
rect 18007 35176 18052 35204
rect 18046 35164 18052 35176
rect 18104 35164 18110 35216
rect 19426 35204 19432 35216
rect 19387 35176 19432 35204
rect 19426 35164 19432 35176
rect 19484 35164 19490 35216
rect 22465 35207 22523 35213
rect 22465 35204 22477 35207
rect 21560 35176 22477 35204
rect 13814 35136 13820 35148
rect 12084 35108 13820 35136
rect 13814 35096 13820 35108
rect 13872 35096 13878 35148
rect 14182 35136 14188 35148
rect 14143 35108 14188 35136
rect 14182 35096 14188 35108
rect 14240 35136 14246 35148
rect 15930 35136 15936 35148
rect 14240 35108 15608 35136
rect 15891 35108 15936 35136
rect 14240 35096 14246 35108
rect 11606 35028 11612 35080
rect 11664 35068 11670 35080
rect 11793 35071 11851 35077
rect 11793 35068 11805 35071
rect 11664 35040 11805 35068
rect 11664 35028 11670 35040
rect 11793 35037 11805 35040
rect 11839 35037 11851 35071
rect 11793 35031 11851 35037
rect 13725 35071 13783 35077
rect 13725 35037 13737 35071
rect 13771 35037 13783 35071
rect 13725 35031 13783 35037
rect 14277 35071 14335 35077
rect 14277 35037 14289 35071
rect 14323 35068 14335 35071
rect 14642 35068 14648 35080
rect 14323 35040 14648 35068
rect 14323 35037 14335 35040
rect 14277 35031 14335 35037
rect 10965 35003 11023 35009
rect 10965 34969 10977 35003
rect 11011 35000 11023 35003
rect 11011 34972 13308 35000
rect 11011 34969 11023 34972
rect 10965 34963 11023 34969
rect 9398 34932 9404 34944
rect 9359 34904 9404 34932
rect 9398 34892 9404 34904
rect 9456 34892 9462 34944
rect 12250 34892 12256 34944
rect 12308 34932 12314 34944
rect 12437 34935 12495 34941
rect 12437 34932 12449 34935
rect 12308 34904 12449 34932
rect 12308 34892 12314 34904
rect 12437 34901 12449 34904
rect 12483 34901 12495 34935
rect 13280 34932 13308 34972
rect 13354 34960 13360 35012
rect 13412 35000 13418 35012
rect 13740 35000 13768 35031
rect 14642 35028 14648 35040
rect 14700 35028 14706 35080
rect 15580 35068 15608 35108
rect 15930 35096 15936 35108
rect 15988 35096 15994 35148
rect 16022 35096 16028 35148
rect 16080 35136 16086 35148
rect 16301 35139 16359 35145
rect 16301 35136 16313 35139
rect 16080 35108 16125 35136
rect 16224 35108 16313 35136
rect 16080 35096 16086 35108
rect 16224 35068 16252 35108
rect 16301 35105 16313 35108
rect 16347 35105 16359 35139
rect 16301 35099 16359 35105
rect 17589 35139 17647 35145
rect 17589 35105 17601 35139
rect 17635 35105 17647 35139
rect 18874 35136 18880 35148
rect 18835 35108 18880 35136
rect 17589 35099 17647 35105
rect 16390 35068 16396 35080
rect 15580 35040 16252 35068
rect 16351 35040 16396 35068
rect 16390 35028 16396 35040
rect 16448 35028 16454 35080
rect 17313 35071 17371 35077
rect 17313 35037 17325 35071
rect 17359 35068 17371 35071
rect 17402 35068 17408 35080
rect 17359 35040 17408 35068
rect 17359 35037 17371 35040
rect 17313 35031 17371 35037
rect 17402 35028 17408 35040
rect 17460 35028 17466 35080
rect 16022 35000 16028 35012
rect 13412 34972 16028 35000
rect 13412 34960 13418 34972
rect 16022 34960 16028 34972
rect 16080 34960 16086 35012
rect 13722 34932 13728 34944
rect 13280 34904 13728 34932
rect 12437 34895 12495 34901
rect 13722 34892 13728 34904
rect 13780 34892 13786 34944
rect 14458 34892 14464 34944
rect 14516 34932 14522 34944
rect 14645 34935 14703 34941
rect 14645 34932 14657 34935
rect 14516 34904 14657 34932
rect 14516 34892 14522 34904
rect 14645 34901 14657 34904
rect 14691 34901 14703 34935
rect 14645 34895 14703 34901
rect 14918 34892 14924 34944
rect 14976 34932 14982 34944
rect 15013 34935 15071 34941
rect 15013 34932 15025 34935
rect 14976 34904 15025 34932
rect 14976 34892 14982 34904
rect 15013 34901 15025 34904
rect 15059 34901 15071 34935
rect 17126 34932 17132 34944
rect 17087 34904 17132 34932
rect 15013 34895 15071 34901
rect 17126 34892 17132 34904
rect 17184 34932 17190 34944
rect 17604 34932 17632 35099
rect 18874 35096 18880 35108
rect 18932 35096 18938 35148
rect 19061 35139 19119 35145
rect 19061 35105 19073 35139
rect 19107 35136 19119 35139
rect 19150 35136 19156 35148
rect 19107 35108 19156 35136
rect 19107 35105 19119 35108
rect 19061 35099 19119 35105
rect 17954 35028 17960 35080
rect 18012 35068 18018 35080
rect 19076 35068 19104 35099
rect 19150 35096 19156 35108
rect 19208 35096 19214 35148
rect 19334 35096 19340 35148
rect 19392 35136 19398 35148
rect 20441 35139 20499 35145
rect 20441 35136 20453 35139
rect 19392 35108 20453 35136
rect 19392 35096 19398 35108
rect 20441 35105 20453 35108
rect 20487 35105 20499 35139
rect 20441 35099 20499 35105
rect 21082 35096 21088 35148
rect 21140 35136 21146 35148
rect 21560 35145 21588 35176
rect 22465 35173 22477 35176
rect 22511 35204 22523 35207
rect 23474 35204 23480 35216
rect 22511 35176 23480 35204
rect 22511 35173 22523 35176
rect 22465 35167 22523 35173
rect 23474 35164 23480 35176
rect 23532 35164 23538 35216
rect 21361 35139 21419 35145
rect 21361 35136 21373 35139
rect 21140 35108 21373 35136
rect 21140 35096 21146 35108
rect 21361 35105 21373 35108
rect 21407 35105 21419 35139
rect 21361 35099 21419 35105
rect 21545 35139 21603 35145
rect 21545 35105 21557 35139
rect 21591 35105 21603 35139
rect 21545 35099 21603 35105
rect 21913 35139 21971 35145
rect 21913 35105 21925 35139
rect 21959 35136 21971 35139
rect 22554 35136 22560 35148
rect 21959 35108 22560 35136
rect 21959 35105 21971 35108
rect 21913 35099 21971 35105
rect 22554 35096 22560 35108
rect 22612 35096 22618 35148
rect 21821 35071 21879 35077
rect 21821 35068 21833 35071
rect 18012 35040 19104 35068
rect 19352 35040 21833 35068
rect 18012 35028 18018 35040
rect 19352 35012 19380 35040
rect 21821 35037 21833 35040
rect 21867 35068 21879 35071
rect 22646 35068 22652 35080
rect 21867 35040 22652 35068
rect 21867 35037 21879 35040
rect 21821 35031 21879 35037
rect 22646 35028 22652 35040
rect 22704 35028 22710 35080
rect 23569 35071 23627 35077
rect 23569 35068 23581 35071
rect 22756 35040 23581 35068
rect 19334 34960 19340 35012
rect 19392 34960 19398 35012
rect 20070 35000 20076 35012
rect 20031 34972 20076 35000
rect 20070 34960 20076 34972
rect 20128 34960 20134 35012
rect 20346 34960 20352 35012
rect 20404 35000 20410 35012
rect 22756 35000 22784 35040
rect 23569 35037 23581 35040
rect 23615 35068 23627 35071
rect 27890 35068 27896 35080
rect 23615 35040 27896 35068
rect 23615 35037 23627 35040
rect 23569 35031 23627 35037
rect 27890 35028 27896 35040
rect 27948 35028 27954 35080
rect 20404 34972 22784 35000
rect 20404 34960 20410 34972
rect 23290 34960 23296 35012
rect 23348 35000 23354 35012
rect 23934 35000 23940 35012
rect 23348 34972 23940 35000
rect 23348 34960 23354 34972
rect 23934 34960 23940 34972
rect 23992 35000 23998 35012
rect 24213 35003 24271 35009
rect 24213 35000 24225 35003
rect 23992 34972 24225 35000
rect 23992 34960 23998 34972
rect 24213 34969 24225 34972
rect 24259 34969 24271 35003
rect 24213 34963 24271 34969
rect 18690 34932 18696 34944
rect 17184 34904 17632 34932
rect 18651 34904 18696 34932
rect 17184 34892 17190 34904
rect 18690 34892 18696 34904
rect 18748 34892 18754 34944
rect 19610 34892 19616 34944
rect 19668 34932 19674 34944
rect 22830 34932 22836 34944
rect 19668 34904 22836 34932
rect 19668 34892 19674 34904
rect 22830 34892 22836 34904
rect 22888 34932 22894 34944
rect 23109 34935 23167 34941
rect 23109 34932 23121 34935
rect 22888 34904 23121 34932
rect 22888 34892 22894 34904
rect 23109 34901 23121 34904
rect 23155 34901 23167 34935
rect 23842 34932 23848 34944
rect 23803 34904 23848 34932
rect 23109 34895 23167 34901
rect 23842 34892 23848 34904
rect 23900 34892 23906 34944
rect 1104 34842 38824 34864
rect 1104 34790 4246 34842
rect 4298 34790 4310 34842
rect 4362 34790 4374 34842
rect 4426 34790 4438 34842
rect 4490 34790 34966 34842
rect 35018 34790 35030 34842
rect 35082 34790 35094 34842
rect 35146 34790 35158 34842
rect 35210 34790 38824 34842
rect 1104 34768 38824 34790
rect 3050 34728 3056 34740
rect 3011 34700 3056 34728
rect 3050 34688 3056 34700
rect 3108 34688 3114 34740
rect 8938 34728 8944 34740
rect 8899 34700 8944 34728
rect 8938 34688 8944 34700
rect 8996 34688 9002 34740
rect 9214 34728 9220 34740
rect 9175 34700 9220 34728
rect 9214 34688 9220 34700
rect 9272 34688 9278 34740
rect 11517 34731 11575 34737
rect 11517 34697 11529 34731
rect 11563 34728 11575 34731
rect 11606 34728 11612 34740
rect 11563 34700 11612 34728
rect 11563 34697 11575 34700
rect 11517 34691 11575 34697
rect 11606 34688 11612 34700
rect 11664 34688 11670 34740
rect 13354 34728 13360 34740
rect 13315 34700 13360 34728
rect 13354 34688 13360 34700
rect 13412 34688 13418 34740
rect 13725 34731 13783 34737
rect 13725 34697 13737 34731
rect 13771 34728 13783 34731
rect 14090 34728 14096 34740
rect 13771 34700 14096 34728
rect 13771 34697 13783 34700
rect 13725 34691 13783 34697
rect 14090 34688 14096 34700
rect 14148 34728 14154 34740
rect 14826 34728 14832 34740
rect 14148 34700 14832 34728
rect 14148 34688 14154 34700
rect 14826 34688 14832 34700
rect 14884 34688 14890 34740
rect 15565 34731 15623 34737
rect 15565 34697 15577 34731
rect 15611 34728 15623 34731
rect 16022 34728 16028 34740
rect 15611 34700 16028 34728
rect 15611 34697 15623 34700
rect 15565 34691 15623 34697
rect 16022 34688 16028 34700
rect 16080 34688 16086 34740
rect 16282 34731 16340 34737
rect 16282 34697 16294 34731
rect 16328 34728 16340 34731
rect 16574 34728 16580 34740
rect 16328 34700 16580 34728
rect 16328 34697 16340 34700
rect 16282 34691 16340 34697
rect 16574 34688 16580 34700
rect 16632 34688 16638 34740
rect 16761 34731 16819 34737
rect 16761 34697 16773 34731
rect 16807 34728 16819 34731
rect 18322 34728 18328 34740
rect 16807 34700 18328 34728
rect 16807 34697 16819 34700
rect 16761 34691 16819 34697
rect 18322 34688 18328 34700
rect 18380 34688 18386 34740
rect 19886 34728 19892 34740
rect 19847 34700 19892 34728
rect 19886 34688 19892 34700
rect 19944 34688 19950 34740
rect 21082 34688 21088 34740
rect 21140 34728 21146 34740
rect 21453 34731 21511 34737
rect 21453 34728 21465 34731
rect 21140 34700 21465 34728
rect 21140 34688 21146 34700
rect 21453 34697 21465 34700
rect 21499 34697 21511 34731
rect 21453 34691 21511 34697
rect 22554 34688 22560 34740
rect 22612 34728 22618 34740
rect 23201 34731 23259 34737
rect 23201 34728 23213 34731
rect 22612 34700 23213 34728
rect 22612 34688 22618 34700
rect 23201 34697 23213 34700
rect 23247 34697 23259 34731
rect 23201 34691 23259 34697
rect 24210 34688 24216 34740
rect 24268 34728 24274 34740
rect 24670 34728 24676 34740
rect 24268 34700 24676 34728
rect 24268 34688 24274 34700
rect 24670 34688 24676 34700
rect 24728 34688 24734 34740
rect 27801 34731 27859 34737
rect 27801 34697 27813 34731
rect 27847 34728 27859 34731
rect 28166 34728 28172 34740
rect 27847 34700 28172 34728
rect 27847 34697 27859 34700
rect 27801 34691 27859 34697
rect 28166 34688 28172 34700
rect 28224 34688 28230 34740
rect 1670 34592 1676 34604
rect 1631 34564 1676 34592
rect 1670 34552 1676 34564
rect 1728 34552 1734 34604
rect 9232 34592 9260 34688
rect 14918 34620 14924 34672
rect 14976 34660 14982 34672
rect 16390 34660 16396 34672
rect 14976 34632 16160 34660
rect 16351 34632 16396 34660
rect 14976 34620 14982 34632
rect 9677 34595 9735 34601
rect 9677 34592 9689 34595
rect 9232 34564 9689 34592
rect 9677 34561 9689 34564
rect 9723 34561 9735 34595
rect 9677 34555 9735 34561
rect 11885 34595 11943 34601
rect 11885 34561 11897 34595
rect 11931 34592 11943 34595
rect 11974 34592 11980 34604
rect 11931 34564 11980 34592
rect 11931 34561 11943 34564
rect 11885 34555 11943 34561
rect 11974 34552 11980 34564
rect 12032 34592 12038 34604
rect 12437 34595 12495 34601
rect 12437 34592 12449 34595
rect 12032 34564 12449 34592
rect 12032 34552 12038 34564
rect 12437 34561 12449 34564
rect 12483 34592 12495 34595
rect 12802 34592 12808 34604
rect 12483 34564 12808 34592
rect 12483 34561 12495 34564
rect 12437 34555 12495 34561
rect 12802 34552 12808 34564
rect 12860 34552 12866 34604
rect 13817 34595 13875 34601
rect 13817 34561 13829 34595
rect 13863 34592 13875 34595
rect 15930 34592 15936 34604
rect 13863 34564 15936 34592
rect 13863 34561 13875 34564
rect 13817 34555 13875 34561
rect 15930 34552 15936 34564
rect 15988 34552 15994 34604
rect 16132 34592 16160 34632
rect 16390 34620 16396 34632
rect 16448 34620 16454 34672
rect 18690 34620 18696 34672
rect 18748 34660 18754 34672
rect 19429 34663 19487 34669
rect 19429 34660 19441 34663
rect 18748 34632 19441 34660
rect 18748 34620 18754 34632
rect 19429 34629 19441 34632
rect 19475 34629 19487 34663
rect 20806 34660 20812 34672
rect 20767 34632 20812 34660
rect 19429 34623 19487 34629
rect 20806 34620 20812 34632
rect 20864 34620 20870 34672
rect 20990 34620 20996 34672
rect 21048 34660 21054 34672
rect 21177 34663 21235 34669
rect 21177 34660 21189 34663
rect 21048 34632 21189 34660
rect 21048 34620 21054 34632
rect 21177 34629 21189 34632
rect 21223 34629 21235 34663
rect 21177 34623 21235 34629
rect 16485 34595 16543 34601
rect 16485 34592 16497 34595
rect 16132 34564 16497 34592
rect 16224 34536 16252 34564
rect 16485 34561 16497 34564
rect 16531 34561 16543 34595
rect 16485 34555 16543 34561
rect 18785 34595 18843 34601
rect 18785 34561 18797 34595
rect 18831 34592 18843 34595
rect 26145 34595 26203 34601
rect 18831 34564 21036 34592
rect 18831 34561 18843 34564
rect 18785 34555 18843 34561
rect 1946 34524 1952 34536
rect 1907 34496 1952 34524
rect 1946 34484 1952 34496
rect 2004 34484 2010 34536
rect 9214 34484 9220 34536
rect 9272 34524 9278 34536
rect 9398 34524 9404 34536
rect 9272 34496 9404 34524
rect 9272 34484 9278 34496
rect 9398 34484 9404 34496
rect 9456 34484 9462 34536
rect 12529 34527 12587 34533
rect 12529 34493 12541 34527
rect 12575 34493 12587 34527
rect 12986 34524 12992 34536
rect 12947 34496 12992 34524
rect 12529 34487 12587 34493
rect 10870 34416 10876 34468
rect 10928 34456 10934 34468
rect 12161 34459 12219 34465
rect 12161 34456 12173 34459
rect 10928 34428 12173 34456
rect 10928 34416 10934 34428
rect 12161 34425 12173 34428
rect 12207 34456 12219 34459
rect 12544 34456 12572 34487
rect 12986 34484 12992 34496
rect 13044 34484 13050 34536
rect 14277 34527 14335 34533
rect 14277 34524 14289 34527
rect 13096 34496 14289 34524
rect 12207 34428 12572 34456
rect 12207 34425 12219 34428
rect 12161 34419 12219 34425
rect 12618 34416 12624 34468
rect 12676 34456 12682 34468
rect 13096 34456 13124 34496
rect 14277 34493 14289 34496
rect 14323 34493 14335 34527
rect 14458 34524 14464 34536
rect 14419 34496 14464 34524
rect 14277 34487 14335 34493
rect 14458 34484 14464 34496
rect 14516 34484 14522 34536
rect 14645 34527 14703 34533
rect 14645 34493 14657 34527
rect 14691 34493 14703 34527
rect 14645 34487 14703 34493
rect 12676 34428 13124 34456
rect 12676 34416 12682 34428
rect 14090 34416 14096 34468
rect 14148 34456 14154 34468
rect 14660 34456 14688 34487
rect 14826 34484 14832 34536
rect 14884 34524 14890 34536
rect 14921 34527 14979 34533
rect 14921 34524 14933 34527
rect 14884 34496 14933 34524
rect 14884 34484 14890 34496
rect 14921 34493 14933 34496
rect 14967 34493 14979 34527
rect 15194 34524 15200 34536
rect 15155 34496 15200 34524
rect 14921 34487 14979 34493
rect 15194 34484 15200 34496
rect 15252 34524 15258 34536
rect 16025 34527 16083 34533
rect 16025 34524 16037 34527
rect 15252 34496 16037 34524
rect 15252 34484 15258 34496
rect 16025 34493 16037 34496
rect 16071 34493 16083 34527
rect 16025 34487 16083 34493
rect 16206 34484 16212 34536
rect 16264 34484 16270 34536
rect 17405 34527 17463 34533
rect 17405 34493 17417 34527
rect 17451 34524 17463 34527
rect 17586 34524 17592 34536
rect 17451 34496 17592 34524
rect 17451 34493 17463 34496
rect 17405 34487 17463 34493
rect 17586 34484 17592 34496
rect 17644 34484 17650 34536
rect 17865 34527 17923 34533
rect 17865 34493 17877 34527
rect 17911 34524 17923 34527
rect 18141 34527 18199 34533
rect 18141 34524 18153 34527
rect 17911 34496 18153 34524
rect 17911 34493 17923 34496
rect 17865 34487 17923 34493
rect 18141 34493 18153 34496
rect 18187 34524 18199 34527
rect 18874 34524 18880 34536
rect 18187 34496 18880 34524
rect 18187 34493 18199 34496
rect 18141 34487 18199 34493
rect 18874 34484 18880 34496
rect 18932 34524 18938 34536
rect 19061 34527 19119 34533
rect 19061 34524 19073 34527
rect 18932 34496 19073 34524
rect 18932 34484 18938 34496
rect 19061 34493 19073 34496
rect 19107 34493 19119 34527
rect 19610 34524 19616 34536
rect 19571 34496 19616 34524
rect 19061 34487 19119 34493
rect 19610 34484 19616 34496
rect 19668 34484 19674 34536
rect 19705 34527 19763 34533
rect 19705 34493 19717 34527
rect 19751 34524 19763 34527
rect 20346 34524 20352 34536
rect 19751 34496 20352 34524
rect 19751 34493 19763 34496
rect 19705 34487 19763 34493
rect 20346 34484 20352 34496
rect 20404 34484 20410 34536
rect 21008 34533 21036 34564
rect 26145 34561 26157 34595
rect 26191 34592 26203 34595
rect 26513 34595 26571 34601
rect 26513 34592 26525 34595
rect 26191 34564 26525 34592
rect 26191 34561 26203 34564
rect 26145 34555 26203 34561
rect 26513 34561 26525 34564
rect 26559 34592 26571 34595
rect 26694 34592 26700 34604
rect 26559 34564 26700 34592
rect 26559 34561 26571 34564
rect 26513 34555 26571 34561
rect 26694 34552 26700 34564
rect 26752 34552 26758 34604
rect 29089 34595 29147 34601
rect 29089 34561 29101 34595
rect 29135 34592 29147 34595
rect 30650 34592 30656 34604
rect 29135 34564 29592 34592
rect 30611 34564 30656 34592
rect 29135 34561 29147 34564
rect 29089 34555 29147 34561
rect 20993 34527 21051 34533
rect 20993 34493 21005 34527
rect 21039 34524 21051 34527
rect 21082 34524 21088 34536
rect 21039 34496 21088 34524
rect 21039 34493 21051 34496
rect 20993 34487 21051 34493
rect 21082 34484 21088 34496
rect 21140 34524 21146 34536
rect 21821 34527 21879 34533
rect 21821 34524 21833 34527
rect 21140 34496 21833 34524
rect 21140 34484 21146 34496
rect 21821 34493 21833 34496
rect 21867 34493 21879 34527
rect 21821 34487 21879 34493
rect 22005 34527 22063 34533
rect 22005 34493 22017 34527
rect 22051 34524 22063 34527
rect 22554 34524 22560 34536
rect 22051 34496 22560 34524
rect 22051 34493 22063 34496
rect 22005 34487 22063 34493
rect 22554 34484 22560 34496
rect 22612 34484 22618 34536
rect 23474 34484 23480 34536
rect 23532 34524 23538 34536
rect 23937 34527 23995 34533
rect 23937 34524 23949 34527
rect 23532 34496 23949 34524
rect 23532 34484 23538 34496
rect 23937 34493 23949 34496
rect 23983 34524 23995 34527
rect 24486 34524 24492 34536
rect 23983 34496 24492 34524
rect 23983 34493 23995 34496
rect 23937 34487 23995 34493
rect 24486 34484 24492 34496
rect 24544 34484 24550 34536
rect 26234 34524 26240 34536
rect 26195 34496 26240 34524
rect 26234 34484 26240 34496
rect 26292 34484 26298 34536
rect 28258 34484 28264 34536
rect 28316 34524 28322 34536
rect 29270 34524 29276 34536
rect 28316 34496 29276 34524
rect 28316 34484 28322 34496
rect 29270 34484 29276 34496
rect 29328 34484 29334 34536
rect 29564 34533 29592 34564
rect 30650 34552 30656 34564
rect 30708 34552 30714 34604
rect 29549 34527 29607 34533
rect 29549 34493 29561 34527
rect 29595 34524 29607 34527
rect 29822 34524 29828 34536
rect 29595 34496 29828 34524
rect 29595 34493 29607 34496
rect 29549 34487 29607 34493
rect 29822 34484 29828 34496
rect 29880 34484 29886 34536
rect 14148 34428 14688 34456
rect 16117 34459 16175 34465
rect 14148 34416 14154 34428
rect 16117 34425 16129 34459
rect 16163 34456 16175 34459
rect 16298 34456 16304 34468
rect 16163 34428 16304 34456
rect 16163 34425 16175 34428
rect 16117 34419 16175 34425
rect 8478 34348 8484 34400
rect 8536 34388 8542 34400
rect 10965 34391 11023 34397
rect 10965 34388 10977 34391
rect 8536 34360 10977 34388
rect 8536 34348 8542 34360
rect 10965 34357 10977 34360
rect 11011 34388 11023 34391
rect 12066 34388 12072 34400
rect 11011 34360 12072 34388
rect 11011 34357 11023 34360
rect 10965 34351 11023 34357
rect 12066 34348 12072 34360
rect 12124 34348 12130 34400
rect 13722 34348 13728 34400
rect 13780 34388 13786 34400
rect 16132 34388 16160 34419
rect 16298 34416 16304 34428
rect 16356 34416 16362 34468
rect 19426 34416 19432 34468
rect 19484 34456 19490 34468
rect 21358 34456 21364 34468
rect 19484 34428 21364 34456
rect 19484 34416 19490 34428
rect 21358 34416 21364 34428
rect 21416 34416 21422 34468
rect 22646 34416 22652 34468
rect 22704 34456 22710 34468
rect 22925 34459 22983 34465
rect 22925 34456 22937 34459
rect 22704 34428 22937 34456
rect 22704 34416 22710 34428
rect 22925 34425 22937 34428
rect 22971 34456 22983 34459
rect 24854 34456 24860 34468
rect 22971 34428 24860 34456
rect 22971 34425 22983 34428
rect 22925 34419 22983 34425
rect 24854 34416 24860 34428
rect 24912 34416 24918 34468
rect 13780 34360 16160 34388
rect 13780 34348 13786 34360
rect 20346 34348 20352 34400
rect 20404 34388 20410 34400
rect 20441 34391 20499 34397
rect 20441 34388 20453 34391
rect 20404 34360 20453 34388
rect 20404 34348 20410 34360
rect 20441 34357 20453 34360
rect 20487 34357 20499 34391
rect 20441 34351 20499 34357
rect 22094 34348 22100 34400
rect 22152 34388 22158 34400
rect 22189 34391 22247 34397
rect 22189 34388 22201 34391
rect 22152 34360 22201 34388
rect 22152 34348 22158 34360
rect 22189 34357 22201 34360
rect 22235 34357 22247 34391
rect 22189 34351 22247 34357
rect 24026 34348 24032 34400
rect 24084 34388 24090 34400
rect 24213 34391 24271 34397
rect 24213 34388 24225 34391
rect 24084 34360 24225 34388
rect 24084 34348 24090 34360
rect 24213 34357 24225 34360
rect 24259 34357 24271 34391
rect 24213 34351 24271 34357
rect 1104 34298 38824 34320
rect 1104 34246 19606 34298
rect 19658 34246 19670 34298
rect 19722 34246 19734 34298
rect 19786 34246 19798 34298
rect 19850 34246 38824 34298
rect 1104 34224 38824 34246
rect 10594 34184 10600 34196
rect 10555 34156 10600 34184
rect 10594 34144 10600 34156
rect 10652 34144 10658 34196
rect 10962 34144 10968 34196
rect 11020 34184 11026 34196
rect 11020 34156 12388 34184
rect 11020 34144 11026 34156
rect 10321 34119 10379 34125
rect 10321 34085 10333 34119
rect 10367 34116 10379 34119
rect 11054 34116 11060 34128
rect 10367 34088 11060 34116
rect 10367 34085 10379 34088
rect 10321 34079 10379 34085
rect 11054 34076 11060 34088
rect 11112 34076 11118 34128
rect 11517 34119 11575 34125
rect 11517 34085 11529 34119
rect 11563 34116 11575 34119
rect 12250 34116 12256 34128
rect 11563 34088 12256 34116
rect 11563 34085 11575 34088
rect 11517 34079 11575 34085
rect 12250 34076 12256 34088
rect 12308 34076 12314 34128
rect 12360 34116 12388 34156
rect 12434 34144 12440 34196
rect 12492 34184 12498 34196
rect 16301 34187 16359 34193
rect 12492 34156 12537 34184
rect 12492 34144 12498 34156
rect 16301 34153 16313 34187
rect 16347 34184 16359 34187
rect 16942 34184 16948 34196
rect 16347 34156 16948 34184
rect 16347 34153 16359 34156
rect 16301 34147 16359 34153
rect 16942 34144 16948 34156
rect 17000 34184 17006 34196
rect 17865 34187 17923 34193
rect 17865 34184 17877 34187
rect 17000 34156 17877 34184
rect 17000 34144 17006 34156
rect 17865 34153 17877 34156
rect 17911 34184 17923 34187
rect 18690 34184 18696 34196
rect 17911 34156 18696 34184
rect 17911 34153 17923 34156
rect 17865 34147 17923 34153
rect 18690 34144 18696 34156
rect 18748 34144 18754 34196
rect 18785 34187 18843 34193
rect 18785 34153 18797 34187
rect 18831 34184 18843 34187
rect 19429 34187 19487 34193
rect 19429 34184 19441 34187
rect 18831 34156 19441 34184
rect 18831 34153 18843 34156
rect 18785 34147 18843 34153
rect 19429 34153 19441 34156
rect 19475 34184 19487 34187
rect 19475 34156 20668 34184
rect 19475 34153 19487 34156
rect 19429 34147 19487 34153
rect 16393 34119 16451 34125
rect 16393 34116 16405 34119
rect 12360 34088 16405 34116
rect 7558 34008 7564 34060
rect 7616 34048 7622 34060
rect 8849 34051 8907 34057
rect 8849 34048 8861 34051
rect 7616 34020 8861 34048
rect 7616 34008 7622 34020
rect 8849 34017 8861 34020
rect 8895 34017 8907 34051
rect 11146 34048 11152 34060
rect 11107 34020 11152 34048
rect 8849 34011 8907 34017
rect 11146 34008 11152 34020
rect 11204 34008 11210 34060
rect 12989 34051 13047 34057
rect 12989 34048 13001 34051
rect 12544 34020 13001 34048
rect 12544 33992 12572 34020
rect 12989 34017 13001 34020
rect 13035 34017 13047 34051
rect 13354 34048 13360 34060
rect 13315 34020 13360 34048
rect 12989 34011 13047 34017
rect 13354 34008 13360 34020
rect 13412 34008 13418 34060
rect 13556 34057 13584 34088
rect 16393 34085 16405 34088
rect 16439 34116 16451 34119
rect 16850 34116 16856 34128
rect 16439 34088 16856 34116
rect 16439 34085 16451 34088
rect 16393 34079 16451 34085
rect 13541 34051 13599 34057
rect 13541 34017 13553 34051
rect 13587 34017 13599 34051
rect 13541 34011 13599 34017
rect 14182 34008 14188 34060
rect 14240 34008 14246 34060
rect 16206 34048 16212 34060
rect 16167 34020 16212 34048
rect 16206 34008 16212 34020
rect 16264 34008 16270 34060
rect 11882 33980 11888 33992
rect 11843 33952 11888 33980
rect 11882 33940 11888 33952
rect 11940 33940 11946 33992
rect 12526 33940 12532 33992
rect 12584 33940 12590 33992
rect 12802 33980 12808 33992
rect 12763 33952 12808 33980
rect 12802 33940 12808 33952
rect 12860 33940 12866 33992
rect 13906 33940 13912 33992
rect 13964 33980 13970 33992
rect 14200 33980 14228 34008
rect 16592 33992 16620 34088
rect 16850 34076 16856 34088
rect 16908 34076 16914 34128
rect 17954 34116 17960 34128
rect 17915 34088 17960 34116
rect 17954 34076 17960 34088
rect 18012 34076 18018 34128
rect 18322 34116 18328 34128
rect 18283 34088 18328 34116
rect 18322 34076 18328 34088
rect 18380 34076 18386 34128
rect 19242 34076 19248 34128
rect 19300 34116 19306 34128
rect 19613 34119 19671 34125
rect 19613 34116 19625 34119
rect 19300 34088 19625 34116
rect 19300 34076 19306 34088
rect 19613 34085 19625 34088
rect 19659 34116 19671 34119
rect 20254 34116 20260 34128
rect 19659 34088 20260 34116
rect 19659 34085 19671 34088
rect 19613 34079 19671 34085
rect 20254 34076 20260 34088
rect 20312 34076 20318 34128
rect 20640 34116 20668 34156
rect 20714 34144 20720 34196
rect 20772 34184 20778 34196
rect 21177 34187 21235 34193
rect 21177 34184 21189 34187
rect 20772 34156 21189 34184
rect 20772 34144 20778 34156
rect 21177 34153 21189 34156
rect 21223 34153 21235 34187
rect 24118 34184 24124 34196
rect 24079 34156 24124 34184
rect 21177 34147 21235 34153
rect 24118 34144 24124 34156
rect 24176 34144 24182 34196
rect 25038 34184 25044 34196
rect 24999 34156 25044 34184
rect 25038 34144 25044 34156
rect 25096 34144 25102 34196
rect 29270 34184 29276 34196
rect 29231 34156 29276 34184
rect 29270 34144 29276 34156
rect 29328 34144 29334 34196
rect 22094 34116 22100 34128
rect 20640 34088 22100 34116
rect 22094 34076 22100 34088
rect 22152 34076 22158 34128
rect 17773 34051 17831 34057
rect 17773 34017 17785 34051
rect 17819 34048 17831 34051
rect 18230 34048 18236 34060
rect 17819 34020 18236 34048
rect 17819 34017 17831 34020
rect 17773 34011 17831 34017
rect 18230 34008 18236 34020
rect 18288 34008 18294 34060
rect 19521 34051 19579 34057
rect 19521 34017 19533 34051
rect 19567 34048 19579 34051
rect 20346 34048 20352 34060
rect 19567 34020 20352 34048
rect 19567 34017 19579 34020
rect 19521 34011 19579 34017
rect 20346 34008 20352 34020
rect 20404 34008 20410 34060
rect 20898 34048 20904 34060
rect 20859 34020 20904 34048
rect 20898 34008 20904 34020
rect 20956 34008 20962 34060
rect 20990 34008 20996 34060
rect 21048 34048 21054 34060
rect 21085 34051 21143 34057
rect 21085 34048 21097 34051
rect 21048 34020 21097 34048
rect 21048 34008 21054 34020
rect 21085 34017 21097 34020
rect 21131 34017 21143 34051
rect 21085 34011 21143 34017
rect 22741 34051 22799 34057
rect 22741 34017 22753 34051
rect 22787 34048 22799 34051
rect 23290 34048 23296 34060
rect 22787 34020 23296 34048
rect 22787 34017 22799 34020
rect 22741 34011 22799 34017
rect 23290 34008 23296 34020
rect 23348 34008 23354 34060
rect 27614 34048 27620 34060
rect 27575 34020 27620 34048
rect 27614 34008 27620 34020
rect 27672 34008 27678 34060
rect 32398 34048 32404 34060
rect 32359 34020 32404 34048
rect 32398 34008 32404 34020
rect 32456 34008 32462 34060
rect 15013 33983 15071 33989
rect 15013 33980 15025 33983
rect 13964 33952 15025 33980
rect 13964 33940 13970 33952
rect 15013 33949 15025 33952
rect 15059 33949 15071 33983
rect 16025 33983 16083 33989
rect 16025 33980 16037 33983
rect 15013 33943 15071 33949
rect 15580 33952 16037 33980
rect 15580 33856 15608 33952
rect 16025 33949 16037 33952
rect 16071 33949 16083 33983
rect 16025 33943 16083 33949
rect 16574 33940 16580 33992
rect 16632 33940 16638 33992
rect 16761 33983 16819 33989
rect 16761 33949 16773 33983
rect 16807 33949 16819 33983
rect 16761 33943 16819 33949
rect 17589 33983 17647 33989
rect 17589 33949 17601 33983
rect 17635 33980 17647 33983
rect 17678 33980 17684 33992
rect 17635 33952 17684 33980
rect 17635 33949 17647 33952
rect 17589 33943 17647 33949
rect 16776 33912 16804 33943
rect 17678 33940 17684 33952
rect 17736 33940 17742 33992
rect 19245 33983 19303 33989
rect 19245 33949 19257 33983
rect 19291 33949 19303 33983
rect 19245 33943 19303 33949
rect 19981 33983 20039 33989
rect 19981 33949 19993 33983
rect 20027 33980 20039 33983
rect 20622 33980 20628 33992
rect 20027 33952 20628 33980
rect 20027 33949 20039 33952
rect 19981 33943 20039 33949
rect 17862 33912 17868 33924
rect 16776 33884 17868 33912
rect 17862 33872 17868 33884
rect 17920 33872 17926 33924
rect 1765 33847 1823 33853
rect 1765 33813 1777 33847
rect 1811 33844 1823 33847
rect 1946 33844 1952 33856
rect 1811 33816 1952 33844
rect 1811 33813 1823 33816
rect 1765 33807 1823 33813
rect 1946 33804 1952 33816
rect 2004 33804 2010 33856
rect 8110 33844 8116 33856
rect 8071 33816 8116 33844
rect 8110 33804 8116 33816
rect 8168 33804 8174 33856
rect 8478 33844 8484 33856
rect 8439 33816 8484 33844
rect 8478 33804 8484 33816
rect 8536 33804 8542 33856
rect 8665 33847 8723 33853
rect 8665 33813 8677 33847
rect 8711 33844 8723 33847
rect 9214 33844 9220 33856
rect 8711 33816 9220 33844
rect 8711 33813 8723 33816
rect 8665 33807 8723 33813
rect 9214 33804 9220 33816
rect 9272 33804 9278 33856
rect 9493 33847 9551 33853
rect 9493 33813 9505 33847
rect 9539 33844 9551 33847
rect 9582 33844 9588 33856
rect 9539 33816 9588 33844
rect 9539 33813 9551 33816
rect 9493 33807 9551 33813
rect 9582 33804 9588 33816
rect 9640 33804 9646 33856
rect 9950 33844 9956 33856
rect 9911 33816 9956 33844
rect 9950 33804 9956 33816
rect 10008 33804 10014 33856
rect 12253 33847 12311 33853
rect 12253 33813 12265 33847
rect 12299 33844 12311 33847
rect 12618 33844 12624 33856
rect 12299 33816 12624 33844
rect 12299 33813 12311 33816
rect 12253 33807 12311 33813
rect 12618 33804 12624 33816
rect 12676 33804 12682 33856
rect 13909 33847 13967 33853
rect 13909 33813 13921 33847
rect 13955 33844 13967 33847
rect 14090 33844 14096 33856
rect 13955 33816 14096 33844
rect 13955 33813 13967 33816
rect 13909 33807 13967 33813
rect 14090 33804 14096 33816
rect 14148 33804 14154 33856
rect 14274 33844 14280 33856
rect 14235 33816 14280 33844
rect 14274 33804 14280 33816
rect 14332 33844 14338 33856
rect 14645 33847 14703 33853
rect 14645 33844 14657 33847
rect 14332 33816 14657 33844
rect 14332 33804 14338 33816
rect 14645 33813 14657 33816
rect 14691 33813 14703 33847
rect 15562 33844 15568 33856
rect 15523 33816 15568 33844
rect 14645 33807 14703 33813
rect 15562 33804 15568 33816
rect 15620 33804 15626 33856
rect 15930 33844 15936 33856
rect 15891 33816 15936 33844
rect 15930 33804 15936 33816
rect 15988 33804 15994 33856
rect 17402 33844 17408 33856
rect 17315 33816 17408 33844
rect 17402 33804 17408 33816
rect 17460 33844 17466 33856
rect 18046 33844 18052 33856
rect 17460 33816 18052 33844
rect 17460 33804 17466 33816
rect 18046 33804 18052 33816
rect 18104 33804 18110 33856
rect 19150 33844 19156 33856
rect 19111 33816 19156 33844
rect 19150 33804 19156 33816
rect 19208 33844 19214 33856
rect 19260 33844 19288 33943
rect 20622 33940 20628 33952
rect 20680 33940 20686 33992
rect 23014 33980 23020 33992
rect 22975 33952 23020 33980
rect 23014 33940 23020 33952
rect 23072 33940 23078 33992
rect 27341 33983 27399 33989
rect 27341 33949 27353 33983
rect 27387 33980 27399 33983
rect 28258 33980 28264 33992
rect 27387 33952 28264 33980
rect 27387 33949 27399 33952
rect 27341 33943 27399 33949
rect 28258 33940 28264 33952
rect 28316 33940 28322 33992
rect 32125 33983 32183 33989
rect 32125 33949 32137 33983
rect 32171 33980 32183 33983
rect 32490 33980 32496 33992
rect 32171 33952 32496 33980
rect 32171 33949 32183 33952
rect 32125 33943 32183 33949
rect 32490 33940 32496 33952
rect 32548 33940 32554 33992
rect 21542 33872 21548 33924
rect 21600 33912 21606 33924
rect 22097 33915 22155 33921
rect 22097 33912 22109 33915
rect 21600 33884 22109 33912
rect 21600 33872 21606 33884
rect 22097 33881 22109 33884
rect 22143 33881 22155 33915
rect 22097 33875 22155 33881
rect 23750 33872 23756 33924
rect 23808 33912 23814 33924
rect 25409 33915 25467 33921
rect 25409 33912 25421 33915
rect 23808 33884 25421 33912
rect 23808 33872 23814 33884
rect 25409 33881 25421 33884
rect 25455 33912 25467 33915
rect 26326 33912 26332 33924
rect 25455 33884 26332 33912
rect 25455 33881 25467 33884
rect 25409 33875 25467 33881
rect 26326 33872 26332 33884
rect 26384 33872 26390 33924
rect 19208 33816 19288 33844
rect 19208 33804 19214 33816
rect 19334 33804 19340 33856
rect 19392 33844 19398 33856
rect 20257 33847 20315 33853
rect 20257 33844 20269 33847
rect 19392 33816 20269 33844
rect 19392 33804 19398 33816
rect 20257 33813 20269 33816
rect 20303 33813 20315 33847
rect 20714 33844 20720 33856
rect 20675 33816 20720 33844
rect 20257 33807 20315 33813
rect 20714 33804 20720 33816
rect 20772 33804 20778 33856
rect 21266 33804 21272 33856
rect 21324 33844 21330 33856
rect 21729 33847 21787 33853
rect 21729 33844 21741 33847
rect 21324 33816 21741 33844
rect 21324 33804 21330 33816
rect 21729 33813 21741 33816
rect 21775 33813 21787 33847
rect 22462 33844 22468 33856
rect 22423 33816 22468 33844
rect 21729 33807 21787 33813
rect 22462 33804 22468 33816
rect 22520 33804 22526 33856
rect 24670 33844 24676 33856
rect 24631 33816 24676 33844
rect 24670 33804 24676 33816
rect 24728 33804 24734 33856
rect 26234 33844 26240 33856
rect 26195 33816 26240 33844
rect 26234 33804 26240 33816
rect 26292 33804 26298 33856
rect 27706 33804 27712 33856
rect 27764 33844 27770 33856
rect 28721 33847 28779 33853
rect 28721 33844 28733 33847
rect 27764 33816 28733 33844
rect 27764 33804 27770 33816
rect 28721 33813 28733 33816
rect 28767 33813 28779 33847
rect 33502 33844 33508 33856
rect 33463 33816 33508 33844
rect 28721 33807 28779 33813
rect 33502 33804 33508 33816
rect 33560 33804 33566 33856
rect 1104 33754 38824 33776
rect 1104 33702 4246 33754
rect 4298 33702 4310 33754
rect 4362 33702 4374 33754
rect 4426 33702 4438 33754
rect 4490 33702 34966 33754
rect 35018 33702 35030 33754
rect 35082 33702 35094 33754
rect 35146 33702 35158 33754
rect 35210 33702 38824 33754
rect 1104 33680 38824 33702
rect 5442 33600 5448 33652
rect 5500 33640 5506 33652
rect 6457 33643 6515 33649
rect 6457 33640 6469 33643
rect 5500 33612 6469 33640
rect 5500 33600 5506 33612
rect 6457 33609 6469 33612
rect 6503 33640 6515 33643
rect 7558 33640 7564 33652
rect 6503 33612 7564 33640
rect 6503 33609 6515 33612
rect 6457 33603 6515 33609
rect 7558 33600 7564 33612
rect 7616 33600 7622 33652
rect 9398 33640 9404 33652
rect 9359 33612 9404 33640
rect 9398 33600 9404 33612
rect 9456 33600 9462 33652
rect 10042 33640 10048 33652
rect 10003 33612 10048 33640
rect 10042 33600 10048 33612
rect 10100 33600 10106 33652
rect 14182 33600 14188 33652
rect 14240 33640 14246 33652
rect 15010 33640 15016 33652
rect 14240 33612 15016 33640
rect 14240 33600 14246 33612
rect 15010 33600 15016 33612
rect 15068 33600 15074 33652
rect 15654 33600 15660 33652
rect 15712 33600 15718 33652
rect 16850 33640 16856 33652
rect 16811 33612 16856 33640
rect 16850 33600 16856 33612
rect 16908 33600 16914 33652
rect 17497 33643 17555 33649
rect 17497 33609 17509 33643
rect 17543 33640 17555 33643
rect 17865 33643 17923 33649
rect 17865 33640 17877 33643
rect 17543 33612 17877 33640
rect 17543 33609 17555 33612
rect 17497 33603 17555 33609
rect 17865 33609 17877 33612
rect 17911 33640 17923 33643
rect 18230 33640 18236 33652
rect 17911 33612 18236 33640
rect 17911 33609 17923 33612
rect 17865 33603 17923 33609
rect 18230 33600 18236 33612
rect 18288 33600 18294 33652
rect 19337 33643 19395 33649
rect 19337 33609 19349 33643
rect 19383 33640 19395 33643
rect 19426 33640 19432 33652
rect 19383 33612 19432 33640
rect 19383 33609 19395 33612
rect 19337 33603 19395 33609
rect 19426 33600 19432 33612
rect 19484 33600 19490 33652
rect 20898 33600 20904 33652
rect 20956 33640 20962 33652
rect 22002 33640 22008 33652
rect 20956 33612 22008 33640
rect 20956 33600 20962 33612
rect 22002 33600 22008 33612
rect 22060 33640 22066 33652
rect 22189 33643 22247 33649
rect 22189 33640 22201 33643
rect 22060 33612 22201 33640
rect 22060 33600 22066 33612
rect 22189 33609 22201 33612
rect 22235 33609 22247 33643
rect 22189 33603 22247 33609
rect 23937 33643 23995 33649
rect 23937 33609 23949 33643
rect 23983 33640 23995 33643
rect 24762 33640 24768 33652
rect 23983 33612 24768 33640
rect 23983 33609 23995 33612
rect 23937 33603 23995 33609
rect 24762 33600 24768 33612
rect 24820 33600 24826 33652
rect 25590 33640 25596 33652
rect 25551 33612 25596 33640
rect 25590 33600 25596 33612
rect 25648 33600 25654 33652
rect 27433 33643 27491 33649
rect 27433 33609 27445 33643
rect 27479 33640 27491 33643
rect 27614 33640 27620 33652
rect 27479 33612 27620 33640
rect 27479 33609 27491 33612
rect 27433 33603 27491 33609
rect 27614 33600 27620 33612
rect 27672 33600 27678 33652
rect 27801 33643 27859 33649
rect 27801 33609 27813 33643
rect 27847 33640 27859 33643
rect 28258 33640 28264 33652
rect 27847 33612 28264 33640
rect 27847 33609 27859 33612
rect 27801 33603 27859 33609
rect 28258 33600 28264 33612
rect 28316 33600 28322 33652
rect 32217 33643 32275 33649
rect 32217 33609 32229 33643
rect 32263 33640 32275 33643
rect 32398 33640 32404 33652
rect 32263 33612 32404 33640
rect 32263 33609 32275 33612
rect 32217 33603 32275 33609
rect 32398 33600 32404 33612
rect 32456 33600 32462 33652
rect 32490 33600 32496 33652
rect 32548 33640 32554 33652
rect 32548 33612 32593 33640
rect 32548 33600 32554 33612
rect 10413 33575 10471 33581
rect 10413 33541 10425 33575
rect 10459 33572 10471 33575
rect 15672 33572 15700 33600
rect 10459 33544 15700 33572
rect 10459 33541 10471 33544
rect 10413 33535 10471 33541
rect 20070 33532 20076 33584
rect 20128 33572 20134 33584
rect 20128 33544 22032 33572
rect 20128 33532 20134 33544
rect 9033 33507 9091 33513
rect 9033 33473 9045 33507
rect 9079 33504 9091 33507
rect 11514 33504 11520 33516
rect 9079 33476 11376 33504
rect 11475 33476 11520 33504
rect 9079 33473 9091 33476
rect 9033 33467 9091 33473
rect 6641 33439 6699 33445
rect 6641 33405 6653 33439
rect 6687 33436 6699 33439
rect 9493 33439 9551 33445
rect 6687 33408 7144 33436
rect 6687 33405 6699 33408
rect 6641 33399 6699 33405
rect 7116 33377 7144 33408
rect 9493 33405 9505 33439
rect 9539 33405 9551 33439
rect 9493 33399 9551 33405
rect 7101 33371 7159 33377
rect 7101 33337 7113 33371
rect 7147 33368 7159 33371
rect 7926 33368 7932 33380
rect 7147 33340 7932 33368
rect 7147 33337 7159 33340
rect 7101 33331 7159 33337
rect 7926 33328 7932 33340
rect 7984 33328 7990 33380
rect 9508 33368 9536 33399
rect 9582 33396 9588 33448
rect 9640 33436 9646 33448
rect 10502 33436 10508 33448
rect 9640 33408 10508 33436
rect 9640 33396 9646 33408
rect 10502 33396 10508 33408
rect 10560 33396 10566 33448
rect 10778 33396 10784 33448
rect 10836 33436 10842 33448
rect 11054 33436 11060 33448
rect 10836 33408 11060 33436
rect 10836 33396 10842 33408
rect 11054 33396 11060 33408
rect 11112 33396 11118 33448
rect 11348 33445 11376 33476
rect 11514 33464 11520 33476
rect 11572 33464 11578 33516
rect 12437 33507 12495 33513
rect 12437 33473 12449 33507
rect 12483 33504 12495 33507
rect 12526 33504 12532 33516
rect 12483 33476 12532 33504
rect 12483 33473 12495 33476
rect 12437 33467 12495 33473
rect 12526 33464 12532 33476
rect 12584 33464 12590 33516
rect 12912 33476 13308 33504
rect 11333 33439 11391 33445
rect 11333 33405 11345 33439
rect 11379 33405 11391 33439
rect 11333 33399 11391 33405
rect 10042 33368 10048 33380
rect 9508 33340 10048 33368
rect 10042 33328 10048 33340
rect 10100 33328 10106 33380
rect 11348 33368 11376 33399
rect 11606 33396 11612 33448
rect 11664 33436 11670 33448
rect 12253 33439 12311 33445
rect 12253 33436 12265 33439
rect 11664 33408 12265 33436
rect 11664 33396 11670 33408
rect 12253 33405 12265 33408
rect 12299 33436 12311 33439
rect 12912 33436 12940 33476
rect 13280 33448 13308 33476
rect 13814 33464 13820 33516
rect 13872 33504 13878 33516
rect 14277 33507 14335 33513
rect 14277 33504 14289 33507
rect 13872 33476 14289 33504
rect 13872 33464 13878 33476
rect 14277 33473 14289 33476
rect 14323 33473 14335 33507
rect 14277 33467 14335 33473
rect 14366 33464 14372 33516
rect 14424 33504 14430 33516
rect 15194 33504 15200 33516
rect 14424 33476 15200 33504
rect 14424 33464 14430 33476
rect 15194 33464 15200 33476
rect 15252 33504 15258 33516
rect 15657 33507 15715 33513
rect 15657 33504 15669 33507
rect 15252 33476 15669 33504
rect 15252 33464 15258 33476
rect 15657 33473 15669 33476
rect 15703 33504 15715 33507
rect 19610 33504 19616 33516
rect 15703 33476 16712 33504
rect 19571 33476 19616 33504
rect 15703 33473 15715 33476
rect 15657 33467 15715 33473
rect 12299 33408 12940 33436
rect 12989 33439 13047 33445
rect 12299 33405 12311 33408
rect 12253 33399 12311 33405
rect 12989 33405 13001 33439
rect 13035 33405 13047 33439
rect 13262 33436 13268 33448
rect 13223 33408 13268 33436
rect 12989 33399 13047 33405
rect 12434 33368 12440 33380
rect 11348 33340 12440 33368
rect 12434 33328 12440 33340
rect 12492 33328 12498 33380
rect 13004 33368 13032 33399
rect 13262 33396 13268 33408
rect 13320 33396 13326 33448
rect 13449 33439 13507 33445
rect 13449 33405 13461 33439
rect 13495 33436 13507 33439
rect 14642 33436 14648 33448
rect 13495 33408 14648 33436
rect 13495 33405 13507 33408
rect 13449 33399 13507 33405
rect 13538 33368 13544 33380
rect 13004 33340 13544 33368
rect 13538 33328 13544 33340
rect 13596 33328 13602 33380
rect 7837 33303 7895 33309
rect 7837 33269 7849 33303
rect 7883 33300 7895 33303
rect 8297 33303 8355 33309
rect 8297 33300 8309 33303
rect 7883 33272 8309 33300
rect 7883 33269 7895 33272
rect 7837 33263 7895 33269
rect 8297 33269 8309 33272
rect 8343 33300 8355 33303
rect 8478 33300 8484 33312
rect 8343 33272 8484 33300
rect 8343 33269 8355 33272
rect 8297 33263 8355 33269
rect 8478 33260 8484 33272
rect 8536 33300 8542 33312
rect 8573 33303 8631 33309
rect 8573 33300 8585 33303
rect 8536 33272 8585 33300
rect 8536 33260 8542 33272
rect 8573 33269 8585 33272
rect 8619 33269 8631 33303
rect 8573 33263 8631 33269
rect 9677 33303 9735 33309
rect 9677 33269 9689 33303
rect 9723 33300 9735 33303
rect 9950 33300 9956 33312
rect 9723 33272 9956 33300
rect 9723 33269 9735 33272
rect 9677 33263 9735 33269
rect 9950 33260 9956 33272
rect 10008 33260 10014 33312
rect 11885 33303 11943 33309
rect 11885 33269 11897 33303
rect 11931 33300 11943 33303
rect 11974 33300 11980 33312
rect 11931 33272 11980 33300
rect 11931 33269 11943 33272
rect 11885 33263 11943 33269
rect 11974 33260 11980 33272
rect 12032 33260 12038 33312
rect 12066 33260 12072 33312
rect 12124 33300 12130 33312
rect 13648 33300 13676 33408
rect 14642 33396 14648 33408
rect 14700 33396 14706 33448
rect 14826 33436 14832 33448
rect 14787 33408 14832 33436
rect 14826 33396 14832 33408
rect 14884 33396 14890 33448
rect 15010 33436 15016 33448
rect 14971 33408 15016 33436
rect 15010 33396 15016 33408
rect 15068 33396 15074 33448
rect 15105 33439 15163 33445
rect 15105 33405 15117 33439
rect 15151 33405 15163 33439
rect 15105 33399 15163 33405
rect 15565 33439 15623 33445
rect 15565 33405 15577 33439
rect 15611 33405 15623 33439
rect 16574 33436 16580 33448
rect 16535 33408 16580 33436
rect 15565 33399 15623 33405
rect 15120 33368 15148 33399
rect 15470 33368 15476 33380
rect 14384 33340 15476 33368
rect 14384 33312 14412 33340
rect 15470 33328 15476 33340
rect 15528 33328 15534 33380
rect 15580 33368 15608 33399
rect 16574 33396 16580 33408
rect 16632 33396 16638 33448
rect 16684 33445 16712 33476
rect 19610 33464 19616 33476
rect 19668 33464 19674 33516
rect 19978 33464 19984 33516
rect 20036 33504 20042 33516
rect 20349 33507 20407 33513
rect 20349 33504 20361 33507
rect 20036 33476 20361 33504
rect 20036 33464 20042 33476
rect 20349 33473 20361 33476
rect 20395 33473 20407 33507
rect 20349 33467 20407 33473
rect 20809 33507 20867 33513
rect 20809 33473 20821 33507
rect 20855 33504 20867 33507
rect 21177 33507 21235 33513
rect 21177 33504 21189 33507
rect 20855 33476 21189 33504
rect 20855 33473 20867 33476
rect 20809 33467 20867 33473
rect 21177 33473 21189 33476
rect 21223 33504 21235 33507
rect 21726 33504 21732 33516
rect 21223 33476 21732 33504
rect 21223 33473 21235 33476
rect 21177 33467 21235 33473
rect 21726 33464 21732 33476
rect 21784 33464 21790 33516
rect 16669 33439 16727 33445
rect 16669 33405 16681 33439
rect 16715 33405 16727 33439
rect 16669 33399 16727 33405
rect 16942 33396 16948 33448
rect 17000 33436 17006 33448
rect 18325 33439 18383 33445
rect 18325 33436 18337 33439
rect 17000 33408 18337 33436
rect 17000 33396 17006 33408
rect 18325 33405 18337 33408
rect 18371 33405 18383 33439
rect 18690 33436 18696 33448
rect 18325 33399 18383 33405
rect 18432 33408 18696 33436
rect 15654 33368 15660 33380
rect 15567 33340 15660 33368
rect 15654 33328 15660 33340
rect 15712 33368 15718 33380
rect 16850 33368 16856 33380
rect 15712 33340 16856 33368
rect 15712 33328 15718 33340
rect 16850 33328 16856 33340
rect 16908 33328 16914 33380
rect 17678 33328 17684 33380
rect 17736 33368 17742 33380
rect 18432 33377 18460 33408
rect 18690 33396 18696 33408
rect 18748 33396 18754 33448
rect 19426 33396 19432 33448
rect 19484 33436 19490 33448
rect 19521 33439 19579 33445
rect 19521 33436 19533 33439
rect 19484 33408 19533 33436
rect 19484 33396 19490 33408
rect 19521 33405 19533 33408
rect 19567 33436 19579 33439
rect 19797 33439 19855 33445
rect 19797 33436 19809 33439
rect 19567 33408 19809 33436
rect 19567 33405 19579 33408
rect 19521 33399 19579 33405
rect 19797 33405 19809 33408
rect 19843 33436 19855 33439
rect 20898 33436 20904 33448
rect 19843 33408 20904 33436
rect 19843 33405 19855 33408
rect 19797 33399 19855 33405
rect 20898 33396 20904 33408
rect 20956 33396 20962 33448
rect 21358 33396 21364 33448
rect 21416 33436 21422 33448
rect 21913 33439 21971 33445
rect 21913 33436 21925 33439
rect 21416 33408 21925 33436
rect 21416 33396 21422 33408
rect 21913 33405 21925 33408
rect 21959 33405 21971 33439
rect 21913 33399 21971 33405
rect 18049 33371 18107 33377
rect 18049 33368 18061 33371
rect 17736 33340 18061 33368
rect 17736 33328 17742 33340
rect 18049 33337 18061 33340
rect 18095 33368 18107 33371
rect 18417 33371 18475 33377
rect 18095 33340 18368 33368
rect 18095 33337 18107 33340
rect 18049 33331 18107 33337
rect 12124 33272 13676 33300
rect 13817 33303 13875 33309
rect 12124 33260 12130 33272
rect 13817 33269 13829 33303
rect 13863 33300 13875 33303
rect 13906 33300 13912 33312
rect 13863 33272 13912 33300
rect 13863 33269 13875 33272
rect 13817 33263 13875 33269
rect 13906 33260 13912 33272
rect 13964 33260 13970 33312
rect 14090 33260 14096 33312
rect 14148 33300 14154 33312
rect 14185 33303 14243 33309
rect 14185 33300 14197 33303
rect 14148 33272 14197 33300
rect 14148 33260 14154 33272
rect 14185 33269 14197 33272
rect 14231 33300 14243 33303
rect 14366 33300 14372 33312
rect 14231 33272 14372 33300
rect 14231 33269 14243 33272
rect 14185 33263 14243 33269
rect 14366 33260 14372 33272
rect 14424 33260 14430 33312
rect 15194 33260 15200 33312
rect 15252 33300 15258 33312
rect 16025 33303 16083 33309
rect 16025 33300 16037 33303
rect 15252 33272 16037 33300
rect 15252 33260 15258 33272
rect 16025 33269 16037 33272
rect 16071 33300 16083 33303
rect 16206 33300 16212 33312
rect 16071 33272 16212 33300
rect 16071 33269 16083 33272
rect 16025 33263 16083 33269
rect 16206 33260 16212 33272
rect 16264 33260 16270 33312
rect 16390 33300 16396 33312
rect 16351 33272 16396 33300
rect 16390 33260 16396 33272
rect 16448 33260 16454 33312
rect 16574 33260 16580 33312
rect 16632 33300 16638 33312
rect 18230 33300 18236 33312
rect 16632 33272 18236 33300
rect 16632 33260 16638 33272
rect 18230 33260 18236 33272
rect 18288 33260 18294 33312
rect 18340 33300 18368 33340
rect 18417 33337 18429 33371
rect 18463 33337 18475 33371
rect 18782 33368 18788 33380
rect 18743 33340 18788 33368
rect 18417 33331 18475 33337
rect 18782 33328 18788 33340
rect 18840 33328 18846 33380
rect 19150 33328 19156 33380
rect 19208 33368 19214 33380
rect 19981 33371 20039 33377
rect 19981 33368 19993 33371
rect 19208 33340 19993 33368
rect 19208 33328 19214 33340
rect 19981 33337 19993 33340
rect 20027 33368 20039 33371
rect 20254 33368 20260 33380
rect 20027 33340 20260 33368
rect 20027 33337 20039 33340
rect 19981 33331 20039 33337
rect 20254 33328 20260 33340
rect 20312 33368 20318 33380
rect 20809 33371 20867 33377
rect 20809 33368 20821 33371
rect 20312 33340 20821 33368
rect 20312 33328 20318 33340
rect 20809 33337 20821 33340
rect 20855 33337 20867 33371
rect 20809 33331 20867 33337
rect 21545 33371 21603 33377
rect 21545 33337 21557 33371
rect 21591 33368 21603 33371
rect 21634 33368 21640 33380
rect 21591 33340 21640 33368
rect 21591 33337 21603 33340
rect 21545 33331 21603 33337
rect 21634 33328 21640 33340
rect 21692 33328 21698 33380
rect 22004 33312 22032 33544
rect 23477 33439 23535 33445
rect 23477 33405 23489 33439
rect 23523 33436 23535 33439
rect 23750 33436 23756 33448
rect 23523 33408 23756 33436
rect 23523 33405 23535 33408
rect 23477 33399 23535 33405
rect 23750 33396 23756 33408
rect 23808 33396 23814 33448
rect 24118 33436 24124 33448
rect 24079 33408 24124 33436
rect 24118 33396 24124 33408
rect 24176 33396 24182 33448
rect 24305 33439 24363 33445
rect 24305 33405 24317 33439
rect 24351 33436 24363 33439
rect 24486 33436 24492 33448
rect 24351 33408 24492 33436
rect 24351 33405 24363 33408
rect 24305 33399 24363 33405
rect 24486 33396 24492 33408
rect 24544 33396 24550 33448
rect 24670 33436 24676 33448
rect 24631 33408 24676 33436
rect 24670 33396 24676 33408
rect 24728 33396 24734 33448
rect 24854 33436 24860 33448
rect 24767 33408 24860 33436
rect 24854 33396 24860 33408
rect 24912 33436 24918 33448
rect 25225 33439 25283 33445
rect 25225 33436 25237 33439
rect 24912 33408 25237 33436
rect 24912 33396 24918 33408
rect 25225 33405 25237 33408
rect 25271 33436 25283 33439
rect 25498 33436 25504 33448
rect 25271 33408 25504 33436
rect 25271 33405 25283 33408
rect 25225 33399 25283 33405
rect 25498 33396 25504 33408
rect 25556 33396 25562 33448
rect 22833 33371 22891 33377
rect 22833 33337 22845 33371
rect 22879 33368 22891 33371
rect 23014 33368 23020 33380
rect 22879 33340 23020 33368
rect 22879 33337 22891 33340
rect 22833 33331 22891 33337
rect 23014 33328 23020 33340
rect 23072 33328 23078 33380
rect 25314 33328 25320 33380
rect 25372 33368 25378 33380
rect 25869 33371 25927 33377
rect 25869 33368 25881 33371
rect 25372 33340 25881 33368
rect 25372 33328 25378 33340
rect 25869 33337 25881 33340
rect 25915 33337 25927 33371
rect 25869 33331 25927 33337
rect 19061 33303 19119 33309
rect 19061 33300 19073 33303
rect 18340 33272 19073 33300
rect 19061 33269 19073 33272
rect 19107 33269 19119 33303
rect 19061 33263 19119 33269
rect 19337 33303 19395 33309
rect 19337 33269 19349 33303
rect 19383 33300 19395 33303
rect 19889 33303 19947 33309
rect 19889 33300 19901 33303
rect 19383 33272 19901 33300
rect 19383 33269 19395 33272
rect 19337 33263 19395 33269
rect 19889 33269 19901 33272
rect 19935 33269 19947 33303
rect 19889 33263 19947 33269
rect 20346 33260 20352 33312
rect 20404 33300 20410 33312
rect 21266 33300 21272 33312
rect 20404 33272 21272 33300
rect 20404 33260 20410 33272
rect 21266 33260 21272 33272
rect 21324 33300 21330 33312
rect 21361 33303 21419 33309
rect 21361 33300 21373 33303
rect 21324 33272 21373 33300
rect 21324 33260 21330 33272
rect 21361 33269 21373 33272
rect 21407 33269 21419 33303
rect 21361 33263 21419 33269
rect 21450 33260 21456 33312
rect 21508 33300 21514 33312
rect 21508 33272 21553 33300
rect 21508 33260 21514 33272
rect 22002 33260 22008 33312
rect 22060 33260 22066 33312
rect 23106 33300 23112 33312
rect 23067 33272 23112 33300
rect 23106 33260 23112 33272
rect 23164 33260 23170 33312
rect 23290 33300 23296 33312
rect 23203 33272 23296 33300
rect 23290 33260 23296 33272
rect 23348 33300 23354 33312
rect 23750 33300 23756 33312
rect 23348 33272 23756 33300
rect 23348 33260 23354 33272
rect 23750 33260 23756 33272
rect 23808 33300 23814 33312
rect 26234 33300 26240 33312
rect 23808 33272 26240 33300
rect 23808 33260 23814 33272
rect 26234 33260 26240 33272
rect 26292 33260 26298 33312
rect 29270 33260 29276 33312
rect 29328 33300 29334 33312
rect 32490 33300 32496 33312
rect 29328 33272 32496 33300
rect 29328 33260 29334 33272
rect 32490 33260 32496 33272
rect 32548 33260 32554 33312
rect 1104 33210 38824 33232
rect 1104 33158 19606 33210
rect 19658 33158 19670 33210
rect 19722 33158 19734 33210
rect 19786 33158 19798 33210
rect 19850 33158 38824 33210
rect 1104 33136 38824 33158
rect 8110 33096 8116 33108
rect 8071 33068 8116 33096
rect 8110 33056 8116 33068
rect 8168 33056 8174 33108
rect 8754 33096 8760 33108
rect 8715 33068 8760 33096
rect 8754 33056 8760 33068
rect 8812 33056 8818 33108
rect 9493 33099 9551 33105
rect 9493 33065 9505 33099
rect 9539 33096 9551 33099
rect 9582 33096 9588 33108
rect 9539 33068 9588 33096
rect 9539 33065 9551 33068
rect 9493 33059 9551 33065
rect 9582 33056 9588 33068
rect 9640 33056 9646 33108
rect 11054 33096 11060 33108
rect 11015 33068 11060 33096
rect 11054 33056 11060 33068
rect 11112 33096 11118 33108
rect 15470 33096 15476 33108
rect 11112 33068 14320 33096
rect 15431 33068 15476 33096
rect 11112 33056 11118 33068
rect 8481 33031 8539 33037
rect 8481 32997 8493 33031
rect 8527 33028 8539 33031
rect 9030 33028 9036 33040
rect 8527 33000 9036 33028
rect 8527 32997 8539 33000
rect 8481 32991 8539 32997
rect 9030 32988 9036 33000
rect 9088 32988 9094 33040
rect 13078 32988 13084 33040
rect 13136 33028 13142 33040
rect 13173 33031 13231 33037
rect 13173 33028 13185 33031
rect 13136 33000 13185 33028
rect 13136 32988 13142 33000
rect 13173 32997 13185 33000
rect 13219 32997 13231 33031
rect 13173 32991 13231 32997
rect 13538 32988 13544 33040
rect 13596 33028 13602 33040
rect 13906 33028 13912 33040
rect 13596 33000 13912 33028
rect 13596 32988 13602 33000
rect 13906 32988 13912 33000
rect 13964 32988 13970 33040
rect 8570 32960 8576 32972
rect 8531 32932 8576 32960
rect 8570 32920 8576 32932
rect 8628 32920 8634 32972
rect 9125 32963 9183 32969
rect 9125 32929 9137 32963
rect 9171 32960 9183 32963
rect 10962 32960 10968 32972
rect 9171 32932 10968 32960
rect 9171 32929 9183 32932
rect 9125 32923 9183 32929
rect 10962 32920 10968 32932
rect 11020 32920 11026 32972
rect 12158 32960 12164 32972
rect 12119 32932 12164 32960
rect 12158 32920 12164 32932
rect 12216 32920 12222 32972
rect 12986 32920 12992 32972
rect 13044 32960 13050 32972
rect 14292 32969 14320 33068
rect 15470 33056 15476 33068
rect 15528 33056 15534 33108
rect 17589 33099 17647 33105
rect 17589 33096 17601 33099
rect 16408 33068 17601 33096
rect 16408 33028 16436 33068
rect 17589 33065 17601 33068
rect 17635 33096 17647 33099
rect 17678 33096 17684 33108
rect 17635 33068 17684 33096
rect 17635 33065 17647 33068
rect 17589 33059 17647 33065
rect 17678 33056 17684 33068
rect 17736 33056 17742 33108
rect 18598 33096 18604 33108
rect 18559 33068 18604 33096
rect 18598 33056 18604 33068
rect 18656 33056 18662 33108
rect 20073 33099 20131 33105
rect 20073 33065 20085 33099
rect 20119 33096 20131 33099
rect 20254 33096 20260 33108
rect 20119 33068 20260 33096
rect 20119 33065 20131 33068
rect 20073 33059 20131 33065
rect 20254 33056 20260 33068
rect 20312 33056 20318 33108
rect 21284 33068 21496 33096
rect 16574 33028 16580 33040
rect 15396 33000 16436 33028
rect 16535 33000 16580 33028
rect 13817 32963 13875 32969
rect 13817 32960 13829 32963
rect 13044 32932 13829 32960
rect 13044 32920 13050 32932
rect 13817 32929 13829 32932
rect 13863 32929 13875 32963
rect 13817 32923 13875 32929
rect 14185 32963 14243 32969
rect 14185 32929 14197 32963
rect 14231 32929 14243 32963
rect 14185 32923 14243 32929
rect 14277 32963 14335 32969
rect 14277 32929 14289 32963
rect 14323 32929 14335 32963
rect 14277 32923 14335 32929
rect 15289 32963 15347 32969
rect 15289 32929 15301 32963
rect 15335 32960 15347 32963
rect 15396 32960 15424 33000
rect 16574 32988 16580 33000
rect 16632 32988 16638 33040
rect 16758 33028 16764 33040
rect 16719 33000 16764 33028
rect 16758 32988 16764 33000
rect 16816 32988 16822 33040
rect 17770 33028 17776 33040
rect 17604 33000 17776 33028
rect 15335 32932 15424 32960
rect 15335 32929 15347 32932
rect 15289 32923 15347 32929
rect 9214 32852 9220 32904
rect 9272 32892 9278 32904
rect 9674 32892 9680 32904
rect 9272 32864 9680 32892
rect 9272 32852 9278 32864
rect 9674 32852 9680 32864
rect 9732 32852 9738 32904
rect 9858 32852 9864 32904
rect 9916 32892 9922 32904
rect 9953 32895 10011 32901
rect 9953 32892 9965 32895
rect 9916 32864 9965 32892
rect 9916 32852 9922 32864
rect 9953 32861 9965 32864
rect 9999 32861 10011 32895
rect 9953 32855 10011 32861
rect 11514 32852 11520 32904
rect 11572 32892 11578 32904
rect 13081 32895 13139 32901
rect 13081 32892 13093 32895
rect 11572 32864 13093 32892
rect 11572 32852 11578 32864
rect 13081 32861 13093 32864
rect 13127 32892 13139 32895
rect 13725 32895 13783 32901
rect 13725 32892 13737 32895
rect 13127 32864 13737 32892
rect 13127 32861 13139 32864
rect 13081 32855 13139 32861
rect 13725 32861 13737 32864
rect 13771 32861 13783 32895
rect 13725 32855 13783 32861
rect 12618 32824 12624 32836
rect 11348 32796 12624 32824
rect 11348 32768 11376 32796
rect 12618 32784 12624 32796
rect 12676 32784 12682 32836
rect 12710 32784 12716 32836
rect 12768 32824 12774 32836
rect 14200 32824 14228 32923
rect 15396 32904 15424 32932
rect 15654 32920 15660 32972
rect 15712 32960 15718 32972
rect 16390 32960 16396 32972
rect 15712 32932 16396 32960
rect 15712 32920 15718 32932
rect 16390 32920 16396 32932
rect 16448 32920 16454 32972
rect 16669 32963 16727 32969
rect 16669 32929 16681 32963
rect 16715 32960 16727 32963
rect 16942 32960 16948 32972
rect 16715 32932 16948 32960
rect 16715 32929 16727 32932
rect 16669 32923 16727 32929
rect 16942 32920 16948 32932
rect 17000 32920 17006 32972
rect 17604 32904 17632 33000
rect 17770 32988 17776 33000
rect 17828 32988 17834 33040
rect 21284 33037 21312 33068
rect 21269 33031 21327 33037
rect 21269 32997 21281 33031
rect 21315 32997 21327 33031
rect 21468 33028 21496 33068
rect 21726 33056 21732 33108
rect 21784 33096 21790 33108
rect 21913 33099 21971 33105
rect 21913 33096 21925 33099
rect 21784 33068 21925 33096
rect 21784 33056 21790 33068
rect 21913 33065 21925 33068
rect 21959 33065 21971 33099
rect 25869 33099 25927 33105
rect 25869 33096 25881 33099
rect 21913 33059 21971 33065
rect 22020 33068 25881 33096
rect 22020 33040 22048 33068
rect 25869 33065 25881 33068
rect 25915 33065 25927 33099
rect 25869 33059 25927 33065
rect 26234 33056 26240 33108
rect 26292 33096 26298 33108
rect 26697 33099 26755 33105
rect 26697 33096 26709 33099
rect 26292 33068 26709 33096
rect 26292 33056 26298 33068
rect 26697 33065 26709 33068
rect 26743 33065 26755 33099
rect 26697 33059 26755 33065
rect 22002 33028 22008 33040
rect 21468 33000 22008 33028
rect 21269 32991 21327 32997
rect 22002 32988 22008 33000
rect 22060 32988 22066 33040
rect 17954 32960 17960 32972
rect 17915 32932 17960 32960
rect 17954 32920 17960 32932
rect 18012 32920 18018 32972
rect 19426 32920 19432 32972
rect 19484 32960 19490 32972
rect 19521 32963 19579 32969
rect 19521 32960 19533 32963
rect 19484 32932 19533 32960
rect 19484 32920 19490 32932
rect 19521 32929 19533 32932
rect 19567 32929 19579 32963
rect 19521 32923 19579 32929
rect 21085 32963 21143 32969
rect 21085 32929 21097 32963
rect 21131 32929 21143 32963
rect 21085 32923 21143 32929
rect 21177 32963 21235 32969
rect 21177 32929 21189 32963
rect 21223 32929 21235 32963
rect 21177 32923 21235 32929
rect 22557 32963 22615 32969
rect 22557 32929 22569 32963
rect 22603 32960 22615 32963
rect 22922 32960 22928 32972
rect 22603 32932 22928 32960
rect 22603 32929 22615 32932
rect 22557 32923 22615 32929
rect 15378 32852 15384 32904
rect 15436 32852 15442 32904
rect 17129 32895 17187 32901
rect 17129 32861 17141 32895
rect 17175 32861 17187 32895
rect 17129 32855 17187 32861
rect 12768 32796 14228 32824
rect 12768 32784 12774 32796
rect 16022 32784 16028 32836
rect 16080 32824 16086 32836
rect 17144 32824 17172 32855
rect 17586 32852 17592 32904
rect 17644 32852 17650 32904
rect 17770 32852 17776 32904
rect 17828 32892 17834 32904
rect 18322 32892 18328 32904
rect 17828 32864 18328 32892
rect 17828 32852 17834 32864
rect 18322 32852 18328 32864
rect 18380 32852 18386 32904
rect 19337 32895 19395 32901
rect 19337 32861 19349 32895
rect 19383 32892 19395 32895
rect 20346 32892 20352 32904
rect 19383 32864 20352 32892
rect 19383 32861 19395 32864
rect 19337 32855 19395 32861
rect 20346 32852 20352 32864
rect 20404 32852 20410 32904
rect 20806 32852 20812 32904
rect 20864 32892 20870 32904
rect 20901 32895 20959 32901
rect 20901 32892 20913 32895
rect 20864 32864 20913 32892
rect 20864 32852 20870 32864
rect 20901 32861 20913 32864
rect 20947 32861 20959 32895
rect 20901 32855 20959 32861
rect 16080 32796 17172 32824
rect 18233 32827 18291 32833
rect 16080 32784 16086 32796
rect 18233 32793 18245 32827
rect 18279 32824 18291 32827
rect 18782 32824 18788 32836
rect 18279 32796 18788 32824
rect 18279 32793 18291 32796
rect 18233 32787 18291 32793
rect 18782 32784 18788 32796
rect 18840 32784 18846 32836
rect 19610 32784 19616 32836
rect 19668 32824 19674 32836
rect 20530 32824 20536 32836
rect 19668 32796 20536 32824
rect 19668 32784 19674 32796
rect 20530 32784 20536 32796
rect 20588 32784 20594 32836
rect 11330 32716 11336 32768
rect 11388 32716 11394 32768
rect 11698 32756 11704 32768
rect 11659 32728 11704 32756
rect 11698 32716 11704 32728
rect 11756 32716 11762 32768
rect 12066 32756 12072 32768
rect 12027 32728 12072 32756
rect 12066 32716 12072 32728
rect 12124 32716 12130 32768
rect 12250 32716 12256 32768
rect 12308 32756 12314 32768
rect 12345 32759 12403 32765
rect 12345 32756 12357 32759
rect 12308 32728 12357 32756
rect 12308 32716 12314 32728
rect 12345 32725 12357 32728
rect 12391 32725 12403 32759
rect 12345 32719 12403 32725
rect 12802 32716 12808 32768
rect 12860 32756 12866 32768
rect 13354 32756 13360 32768
rect 12860 32728 13360 32756
rect 12860 32716 12866 32728
rect 13354 32716 13360 32728
rect 13412 32716 13418 32768
rect 13814 32716 13820 32768
rect 13872 32756 13878 32768
rect 14458 32756 14464 32768
rect 13872 32728 14464 32756
rect 13872 32716 13878 32728
rect 14458 32716 14464 32728
rect 14516 32756 14522 32768
rect 14645 32759 14703 32765
rect 14645 32756 14657 32759
rect 14516 32728 14657 32756
rect 14516 32716 14522 32728
rect 14645 32725 14657 32728
rect 14691 32756 14703 32759
rect 15010 32756 15016 32768
rect 14691 32728 15016 32756
rect 14691 32725 14703 32728
rect 14645 32719 14703 32725
rect 15010 32716 15016 32728
rect 15068 32716 15074 32768
rect 15746 32716 15752 32768
rect 15804 32756 15810 32768
rect 15933 32759 15991 32765
rect 15933 32756 15945 32759
rect 15804 32728 15945 32756
rect 15804 32716 15810 32728
rect 15933 32725 15945 32728
rect 15979 32756 15991 32759
rect 16298 32756 16304 32768
rect 15979 32728 16304 32756
rect 15979 32725 15991 32728
rect 15933 32719 15991 32725
rect 16298 32716 16304 32728
rect 16356 32756 16362 32768
rect 16666 32756 16672 32768
rect 16356 32728 16672 32756
rect 16356 32716 16362 32728
rect 16666 32716 16672 32728
rect 16724 32716 16730 32768
rect 17862 32716 17868 32768
rect 17920 32756 17926 32768
rect 18122 32759 18180 32765
rect 18122 32756 18134 32759
rect 17920 32728 18134 32756
rect 17920 32716 17926 32728
rect 18122 32725 18134 32728
rect 18168 32756 18180 32759
rect 18322 32756 18328 32768
rect 18168 32728 18328 32756
rect 18168 32725 18180 32728
rect 18122 32719 18180 32725
rect 18322 32716 18328 32728
rect 18380 32716 18386 32768
rect 18874 32716 18880 32768
rect 18932 32756 18938 32768
rect 18969 32759 19027 32765
rect 18969 32756 18981 32759
rect 18932 32728 18981 32756
rect 18932 32716 18938 32728
rect 18969 32725 18981 32728
rect 19015 32756 19027 32759
rect 19058 32756 19064 32768
rect 19015 32728 19064 32756
rect 19015 32725 19027 32728
rect 18969 32719 19027 32725
rect 19058 32716 19064 32728
rect 19116 32716 19122 32768
rect 19426 32716 19432 32768
rect 19484 32756 19490 32768
rect 19705 32759 19763 32765
rect 19705 32756 19717 32759
rect 19484 32728 19717 32756
rect 19484 32716 19490 32728
rect 19705 32725 19717 32728
rect 19751 32725 19763 32759
rect 20714 32756 20720 32768
rect 20675 32728 20720 32756
rect 19705 32719 19763 32725
rect 20714 32716 20720 32728
rect 20772 32756 20778 32768
rect 21100 32756 21128 32923
rect 21192 32824 21220 32923
rect 22922 32920 22928 32932
rect 22980 32920 22986 32972
rect 24210 32960 24216 32972
rect 24171 32932 24216 32960
rect 24210 32920 24216 32932
rect 24268 32920 24274 32972
rect 27157 32963 27215 32969
rect 27157 32929 27169 32963
rect 27203 32960 27215 32963
rect 27338 32960 27344 32972
rect 27203 32932 27344 32960
rect 27203 32929 27215 32932
rect 27157 32923 27215 32929
rect 27338 32920 27344 32932
rect 27396 32960 27402 32972
rect 28258 32960 28264 32972
rect 27396 32932 28264 32960
rect 27396 32920 27402 32932
rect 28258 32920 28264 32932
rect 28316 32960 28322 32972
rect 28442 32960 28448 32972
rect 28316 32932 28448 32960
rect 28316 32920 28322 32932
rect 28442 32920 28448 32932
rect 28500 32960 28506 32972
rect 28629 32963 28687 32969
rect 28629 32960 28641 32963
rect 28500 32932 28641 32960
rect 28500 32920 28506 32932
rect 28629 32929 28641 32932
rect 28675 32929 28687 32963
rect 28902 32960 28908 32972
rect 28863 32932 28908 32960
rect 28629 32923 28687 32929
rect 28902 32920 28908 32932
rect 28960 32920 28966 32972
rect 21634 32852 21640 32904
rect 21692 32892 21698 32904
rect 21692 32864 21737 32892
rect 21692 32852 21698 32864
rect 22094 32852 22100 32904
rect 22152 32892 22158 32904
rect 22462 32892 22468 32904
rect 22152 32864 22468 32892
rect 22152 32852 22158 32864
rect 22462 32852 22468 32864
rect 22520 32852 22526 32904
rect 23658 32892 23664 32904
rect 23619 32864 23664 32892
rect 23658 32852 23664 32864
rect 23716 32852 23722 32904
rect 23750 32852 23756 32904
rect 23808 32892 23814 32904
rect 23937 32895 23995 32901
rect 23937 32892 23949 32895
rect 23808 32864 23949 32892
rect 23808 32852 23814 32864
rect 23937 32861 23949 32864
rect 23983 32861 23995 32895
rect 25314 32892 25320 32904
rect 25275 32864 25320 32892
rect 23937 32855 23995 32861
rect 25314 32852 25320 32864
rect 25372 32852 25378 32904
rect 22373 32827 22431 32833
rect 22373 32824 22385 32827
rect 21192 32796 22385 32824
rect 22373 32793 22385 32796
rect 22419 32824 22431 32827
rect 22646 32824 22652 32836
rect 22419 32796 22652 32824
rect 22419 32793 22431 32796
rect 22373 32787 22431 32793
rect 22646 32784 22652 32796
rect 22704 32784 22710 32836
rect 24946 32784 24952 32836
rect 25004 32824 25010 32836
rect 26329 32827 26387 32833
rect 26329 32824 26341 32827
rect 25004 32796 26341 32824
rect 25004 32784 25010 32796
rect 26329 32793 26341 32796
rect 26375 32824 26387 32827
rect 28166 32824 28172 32836
rect 26375 32796 28172 32824
rect 26375 32793 26387 32796
rect 26329 32787 26387 32793
rect 28166 32784 28172 32796
rect 28224 32784 28230 32836
rect 20772 32728 21128 32756
rect 20772 32716 20778 32728
rect 22554 32716 22560 32768
rect 22612 32756 22618 32768
rect 22741 32759 22799 32765
rect 22741 32756 22753 32759
rect 22612 32728 22753 32756
rect 22612 32716 22618 32728
rect 22741 32725 22753 32728
rect 22787 32725 22799 32759
rect 23290 32756 23296 32768
rect 23251 32728 23296 32756
rect 22741 32719 22799 32725
rect 23290 32716 23296 32728
rect 23348 32716 23354 32768
rect 30006 32756 30012 32768
rect 29967 32728 30012 32756
rect 30006 32716 30012 32728
rect 30064 32716 30070 32768
rect 1104 32666 38824 32688
rect 1104 32614 4246 32666
rect 4298 32614 4310 32666
rect 4362 32614 4374 32666
rect 4426 32614 4438 32666
rect 4490 32614 34966 32666
rect 35018 32614 35030 32666
rect 35082 32614 35094 32666
rect 35146 32614 35158 32666
rect 35210 32614 38824 32666
rect 1104 32592 38824 32614
rect 1670 32512 1676 32564
rect 1728 32552 1734 32564
rect 4893 32555 4951 32561
rect 4893 32552 4905 32555
rect 1728 32524 4905 32552
rect 1728 32512 1734 32524
rect 4893 32521 4905 32524
rect 4939 32521 4951 32555
rect 5442 32552 5448 32564
rect 5403 32524 5448 32552
rect 4893 32515 4951 32521
rect 5442 32512 5448 32524
rect 5500 32512 5506 32564
rect 7742 32552 7748 32564
rect 7703 32524 7748 32552
rect 7742 32512 7748 32524
rect 7800 32512 7806 32564
rect 9125 32555 9183 32561
rect 9125 32552 9137 32555
rect 8312 32524 9137 32552
rect 5077 32351 5135 32357
rect 5077 32317 5089 32351
rect 5123 32348 5135 32351
rect 5442 32348 5448 32360
rect 5123 32320 5448 32348
rect 5123 32317 5135 32320
rect 5077 32311 5135 32317
rect 5442 32308 5448 32320
rect 5500 32308 5506 32360
rect 8312 32357 8340 32524
rect 9125 32521 9137 32524
rect 9171 32552 9183 32555
rect 9214 32552 9220 32564
rect 9171 32524 9220 32552
rect 9171 32521 9183 32524
rect 9125 32515 9183 32521
rect 9214 32512 9220 32524
rect 9272 32512 9278 32564
rect 9858 32512 9864 32564
rect 9916 32552 9922 32564
rect 10413 32555 10471 32561
rect 10413 32552 10425 32555
rect 9916 32524 10425 32552
rect 9916 32512 9922 32524
rect 10413 32521 10425 32524
rect 10459 32521 10471 32555
rect 11882 32552 11888 32564
rect 11843 32524 11888 32552
rect 10413 32515 10471 32521
rect 11882 32512 11888 32524
rect 11940 32512 11946 32564
rect 12158 32552 12164 32564
rect 12119 32524 12164 32552
rect 12158 32512 12164 32524
rect 12216 32512 12222 32564
rect 12713 32555 12771 32561
rect 12713 32521 12725 32555
rect 12759 32552 12771 32555
rect 15378 32552 15384 32564
rect 12759 32524 15384 32552
rect 12759 32521 12771 32524
rect 12713 32515 12771 32521
rect 15378 32512 15384 32524
rect 15436 32512 15442 32564
rect 16022 32512 16028 32564
rect 16080 32561 16086 32564
rect 16080 32555 16129 32561
rect 16080 32521 16083 32555
rect 16117 32521 16129 32555
rect 16080 32515 16129 32521
rect 16080 32512 16086 32515
rect 16758 32512 16764 32564
rect 16816 32552 16822 32564
rect 16945 32555 17003 32561
rect 16945 32552 16957 32555
rect 16816 32524 16957 32552
rect 16816 32512 16822 32524
rect 16945 32521 16957 32524
rect 16991 32521 17003 32555
rect 17310 32552 17316 32564
rect 16945 32515 17003 32521
rect 17236 32524 17316 32552
rect 13078 32484 13084 32496
rect 12452 32456 13084 32484
rect 8757 32419 8815 32425
rect 8757 32385 8769 32419
rect 8803 32416 8815 32419
rect 9306 32416 9312 32428
rect 8803 32388 9312 32416
rect 8803 32385 8815 32388
rect 8757 32379 8815 32385
rect 9306 32376 9312 32388
rect 9364 32376 9370 32428
rect 9493 32419 9551 32425
rect 9493 32385 9505 32419
rect 9539 32416 9551 32419
rect 9539 32388 9720 32416
rect 9539 32385 9551 32388
rect 9493 32379 9551 32385
rect 9692 32360 9720 32388
rect 10962 32376 10968 32428
rect 11020 32425 11026 32428
rect 11020 32419 11033 32425
rect 11021 32416 11033 32419
rect 11514 32416 11520 32428
rect 11021 32388 11065 32416
rect 11475 32388 11520 32416
rect 11021 32385 11033 32388
rect 11020 32379 11033 32385
rect 11020 32376 11026 32379
rect 11514 32376 11520 32388
rect 11572 32376 11578 32428
rect 8205 32351 8263 32357
rect 8205 32348 8217 32351
rect 8128 32320 8217 32348
rect 8128 32224 8156 32320
rect 8205 32317 8217 32320
rect 8251 32317 8263 32351
rect 8205 32311 8263 32317
rect 8297 32351 8355 32357
rect 8297 32317 8309 32351
rect 8343 32317 8355 32351
rect 8297 32311 8355 32317
rect 9030 32308 9036 32360
rect 9088 32348 9094 32360
rect 9585 32351 9643 32357
rect 9585 32348 9597 32351
rect 9088 32320 9597 32348
rect 9088 32308 9094 32320
rect 9585 32317 9597 32320
rect 9631 32317 9643 32351
rect 9585 32311 9643 32317
rect 9674 32308 9680 32360
rect 9732 32348 9738 32360
rect 11054 32348 11060 32360
rect 9732 32320 9777 32348
rect 10967 32320 11060 32348
rect 9732 32308 9738 32320
rect 11054 32308 11060 32320
rect 11112 32348 11118 32360
rect 11882 32348 11888 32360
rect 11112 32320 11888 32348
rect 11112 32308 11118 32320
rect 11882 32308 11888 32320
rect 11940 32308 11946 32360
rect 12452 32348 12480 32456
rect 13078 32444 13084 32456
rect 13136 32444 13142 32496
rect 14366 32484 14372 32496
rect 13556 32456 14372 32484
rect 13556 32428 13584 32456
rect 14366 32444 14372 32456
rect 14424 32444 14430 32496
rect 15286 32444 15292 32496
rect 15344 32484 15350 32496
rect 16206 32484 16212 32496
rect 15344 32456 16212 32484
rect 15344 32444 15350 32456
rect 16206 32444 16212 32456
rect 16264 32444 16270 32496
rect 13449 32419 13507 32425
rect 13449 32385 13461 32419
rect 13495 32416 13507 32419
rect 13538 32416 13544 32428
rect 13495 32388 13544 32416
rect 13495 32385 13507 32388
rect 13449 32379 13507 32385
rect 13538 32376 13544 32388
rect 13596 32376 13602 32428
rect 15838 32416 15844 32428
rect 14108 32388 15844 32416
rect 12529 32351 12587 32357
rect 12529 32348 12541 32351
rect 12452 32320 12541 32348
rect 12529 32317 12541 32320
rect 12575 32317 12587 32351
rect 12529 32311 12587 32317
rect 12618 32308 12624 32360
rect 12676 32348 12682 32360
rect 13814 32348 13820 32360
rect 12676 32320 13820 32348
rect 12676 32308 12682 32320
rect 13814 32308 13820 32320
rect 13872 32308 13878 32360
rect 14001 32351 14059 32357
rect 14001 32317 14013 32351
rect 14047 32348 14059 32351
rect 14108 32348 14136 32388
rect 15838 32376 15844 32388
rect 15896 32376 15902 32428
rect 16298 32416 16304 32428
rect 16259 32388 16304 32416
rect 16298 32376 16304 32388
rect 16356 32376 16362 32428
rect 14047 32320 14136 32348
rect 14277 32351 14335 32357
rect 14047 32317 14059 32320
rect 14001 32311 14059 32317
rect 14277 32317 14289 32351
rect 14323 32317 14335 32351
rect 14277 32311 14335 32317
rect 10134 32280 10140 32292
rect 10095 32252 10140 32280
rect 10134 32240 10140 32252
rect 10192 32240 10198 32292
rect 10870 32280 10876 32292
rect 10831 32252 10876 32280
rect 10870 32240 10876 32252
rect 10928 32240 10934 32292
rect 12434 32240 12440 32292
rect 12492 32280 12498 32292
rect 13541 32283 13599 32289
rect 13541 32280 13553 32283
rect 12492 32252 13553 32280
rect 12492 32240 12498 32252
rect 13541 32249 13553 32252
rect 13587 32249 13599 32283
rect 13832 32280 13860 32308
rect 14292 32280 14320 32311
rect 14366 32308 14372 32360
rect 14424 32348 14430 32360
rect 14642 32348 14648 32360
rect 14424 32320 14469 32348
rect 14603 32320 14648 32348
rect 14424 32308 14430 32320
rect 14642 32308 14648 32320
rect 14700 32308 14706 32360
rect 14826 32308 14832 32360
rect 14884 32348 14890 32360
rect 14921 32351 14979 32357
rect 14921 32348 14933 32351
rect 14884 32320 14933 32348
rect 14884 32308 14890 32320
rect 14921 32317 14933 32320
rect 14967 32317 14979 32351
rect 14921 32311 14979 32317
rect 15749 32351 15807 32357
rect 15749 32317 15761 32351
rect 15795 32348 15807 32351
rect 16574 32348 16580 32360
rect 15795 32320 16580 32348
rect 15795 32317 15807 32320
rect 15749 32311 15807 32317
rect 13832 32252 14320 32280
rect 13541 32243 13599 32249
rect 7377 32215 7435 32221
rect 7377 32181 7389 32215
rect 7423 32212 7435 32215
rect 7558 32212 7564 32224
rect 7423 32184 7564 32212
rect 7423 32181 7435 32184
rect 7377 32175 7435 32181
rect 7558 32172 7564 32184
rect 7616 32172 7622 32224
rect 8110 32212 8116 32224
rect 8071 32184 8116 32212
rect 8110 32172 8116 32184
rect 8168 32172 8174 32224
rect 13078 32172 13084 32224
rect 13136 32212 13142 32224
rect 13446 32212 13452 32224
rect 13136 32184 13452 32212
rect 13136 32172 13142 32184
rect 13446 32172 13452 32184
rect 13504 32172 13510 32224
rect 13814 32172 13820 32224
rect 13872 32212 13878 32224
rect 15764 32212 15792 32311
rect 16574 32308 16580 32320
rect 16632 32308 16638 32360
rect 15838 32240 15844 32292
rect 15896 32280 15902 32292
rect 15933 32283 15991 32289
rect 15933 32280 15945 32283
rect 15896 32252 15945 32280
rect 15896 32240 15902 32252
rect 15933 32249 15945 32252
rect 15979 32249 15991 32283
rect 17236 32280 17264 32524
rect 17310 32512 17316 32524
rect 17368 32512 17374 32564
rect 17405 32555 17463 32561
rect 17405 32521 17417 32555
rect 17451 32552 17463 32555
rect 17451 32524 19012 32552
rect 17451 32521 17463 32524
rect 17405 32515 17463 32521
rect 17310 32376 17316 32428
rect 17368 32416 17374 32428
rect 17420 32416 17448 32515
rect 18874 32484 18880 32496
rect 17368 32388 17448 32416
rect 18800 32456 18880 32484
rect 17368 32376 17374 32388
rect 17586 32308 17592 32360
rect 17644 32348 17650 32360
rect 17681 32351 17739 32357
rect 17681 32348 17693 32351
rect 17644 32320 17693 32348
rect 17644 32308 17650 32320
rect 17681 32317 17693 32320
rect 17727 32317 17739 32351
rect 17681 32311 17739 32317
rect 18325 32351 18383 32357
rect 18325 32317 18337 32351
rect 18371 32348 18383 32351
rect 18414 32348 18420 32360
rect 18371 32320 18420 32348
rect 18371 32317 18383 32320
rect 18325 32311 18383 32317
rect 18414 32308 18420 32320
rect 18472 32308 18478 32360
rect 18800 32357 18828 32456
rect 18874 32444 18880 32456
rect 18932 32444 18938 32496
rect 18984 32416 19012 32524
rect 19886 32512 19892 32564
rect 19944 32552 19950 32564
rect 20070 32552 20076 32564
rect 19944 32524 20076 32552
rect 19944 32512 19950 32524
rect 20070 32512 20076 32524
rect 20128 32512 20134 32564
rect 20533 32555 20591 32561
rect 20533 32521 20545 32555
rect 20579 32552 20591 32555
rect 21082 32552 21088 32564
rect 20579 32524 21088 32552
rect 20579 32521 20591 32524
rect 20533 32515 20591 32521
rect 21082 32512 21088 32524
rect 21140 32512 21146 32564
rect 22094 32512 22100 32564
rect 22152 32552 22158 32564
rect 22465 32555 22523 32561
rect 22465 32552 22477 32555
rect 22152 32524 22477 32552
rect 22152 32512 22158 32524
rect 22465 32521 22477 32524
rect 22511 32521 22523 32555
rect 22465 32515 22523 32521
rect 23400 32524 24624 32552
rect 20790 32487 20848 32493
rect 20790 32453 20802 32487
rect 20836 32484 20848 32487
rect 20901 32487 20959 32493
rect 20836 32453 20852 32484
rect 20790 32447 20852 32453
rect 20901 32453 20913 32487
rect 20947 32484 20959 32487
rect 21726 32484 21732 32496
rect 20947 32456 21732 32484
rect 20947 32453 20959 32456
rect 20901 32447 20959 32453
rect 19613 32419 19671 32425
rect 18984 32388 19196 32416
rect 19168 32357 19196 32388
rect 19613 32385 19625 32419
rect 19659 32416 19671 32419
rect 19886 32416 19892 32428
rect 19659 32388 19892 32416
rect 19659 32385 19671 32388
rect 19613 32379 19671 32385
rect 19886 32376 19892 32388
rect 19944 32376 19950 32428
rect 20824 32416 20852 32447
rect 21726 32444 21732 32456
rect 21784 32484 21790 32496
rect 23290 32484 23296 32496
rect 21784 32456 23296 32484
rect 21784 32444 21790 32456
rect 23290 32444 23296 32456
rect 23348 32444 23354 32496
rect 20993 32419 21051 32425
rect 20088 32388 20668 32416
rect 20824 32388 20944 32416
rect 18785 32351 18843 32357
rect 18785 32317 18797 32351
rect 18831 32317 18843 32351
rect 18785 32311 18843 32317
rect 18969 32351 19027 32357
rect 18969 32317 18981 32351
rect 19015 32317 19027 32351
rect 18969 32311 19027 32317
rect 19153 32351 19211 32357
rect 19153 32317 19165 32351
rect 19199 32317 19211 32351
rect 19153 32311 19211 32317
rect 17236 32252 17632 32280
rect 15933 32243 15991 32249
rect 17604 32224 17632 32252
rect 17954 32240 17960 32292
rect 18012 32280 18018 32292
rect 18984 32280 19012 32311
rect 19242 32308 19248 32360
rect 19300 32348 19306 32360
rect 19797 32351 19855 32357
rect 19797 32348 19809 32351
rect 19300 32320 19809 32348
rect 19300 32308 19306 32320
rect 19797 32317 19809 32320
rect 19843 32348 19855 32351
rect 20088 32348 20116 32388
rect 19843 32320 20116 32348
rect 20640 32348 20668 32388
rect 20806 32348 20812 32360
rect 20640 32320 20812 32348
rect 19843 32317 19855 32320
rect 19797 32311 19855 32317
rect 20806 32308 20812 32320
rect 20864 32308 20870 32360
rect 20916 32348 20944 32388
rect 20993 32385 21005 32419
rect 21039 32416 21051 32419
rect 21082 32416 21088 32428
rect 21039 32388 21088 32416
rect 21039 32385 21051 32388
rect 20993 32379 21051 32385
rect 21082 32376 21088 32388
rect 21140 32376 21146 32428
rect 21450 32376 21456 32428
rect 21508 32416 21514 32428
rect 22002 32416 22008 32428
rect 21508 32388 22008 32416
rect 21508 32376 21514 32388
rect 21652 32348 21680 32388
rect 22002 32376 22008 32388
rect 22060 32376 22066 32428
rect 22189 32419 22247 32425
rect 22189 32385 22201 32419
rect 22235 32416 22247 32419
rect 23400 32416 23428 32524
rect 24596 32484 24624 32524
rect 24854 32512 24860 32564
rect 24912 32552 24918 32564
rect 25041 32555 25099 32561
rect 25041 32552 25053 32555
rect 24912 32524 25053 32552
rect 24912 32512 24918 32524
rect 25041 32521 25053 32524
rect 25087 32521 25099 32555
rect 25590 32552 25596 32564
rect 25551 32524 25596 32552
rect 25041 32515 25099 32521
rect 25590 32512 25596 32524
rect 25648 32512 25654 32564
rect 26326 32512 26332 32564
rect 26384 32552 26390 32564
rect 27157 32555 27215 32561
rect 27157 32552 27169 32555
rect 26384 32524 27169 32552
rect 26384 32512 26390 32524
rect 27157 32521 27169 32524
rect 27203 32552 27215 32555
rect 28261 32555 28319 32561
rect 28261 32552 28273 32555
rect 27203 32524 28273 32552
rect 27203 32521 27215 32524
rect 27157 32515 27215 32521
rect 28261 32521 28273 32524
rect 28307 32521 28319 32555
rect 28442 32552 28448 32564
rect 28403 32524 28448 32552
rect 28261 32515 28319 32521
rect 25774 32484 25780 32496
rect 24596 32456 25780 32484
rect 25774 32444 25780 32456
rect 25832 32444 25838 32496
rect 24118 32416 24124 32428
rect 22235 32388 23428 32416
rect 23952 32388 24124 32416
rect 22235 32385 22247 32388
rect 22189 32379 22247 32385
rect 22204 32348 22232 32379
rect 23952 32360 23980 32388
rect 24118 32376 24124 32388
rect 24176 32416 24182 32428
rect 25961 32419 26019 32425
rect 25961 32416 25973 32419
rect 24176 32388 25973 32416
rect 24176 32376 24182 32388
rect 25961 32385 25973 32388
rect 26007 32385 26019 32419
rect 25961 32379 26019 32385
rect 20916 32320 21680 32348
rect 21744 32320 22232 32348
rect 22281 32351 22339 32357
rect 18012 32252 19012 32280
rect 18012 32240 18018 32252
rect 18432 32224 18460 32252
rect 19058 32240 19064 32292
rect 19116 32280 19122 32292
rect 19610 32280 19616 32292
rect 19116 32252 19616 32280
rect 19116 32240 19122 32252
rect 19610 32240 19616 32252
rect 19668 32280 19674 32292
rect 20625 32283 20683 32289
rect 20625 32280 20637 32283
rect 19668 32252 20637 32280
rect 19668 32240 19674 32252
rect 20625 32249 20637 32252
rect 20671 32249 20683 32283
rect 20625 32243 20683 32249
rect 20990 32240 20996 32292
rect 21048 32240 21054 32292
rect 21174 32240 21180 32292
rect 21232 32280 21238 32292
rect 21637 32283 21695 32289
rect 21637 32280 21649 32283
rect 21232 32252 21649 32280
rect 21232 32240 21238 32252
rect 21637 32249 21649 32252
rect 21683 32249 21695 32283
rect 21637 32243 21695 32249
rect 16574 32212 16580 32224
rect 13872 32184 15792 32212
rect 16535 32184 16580 32212
rect 13872 32172 13878 32184
rect 16574 32172 16580 32184
rect 16632 32172 16638 32224
rect 17402 32172 17408 32224
rect 17460 32212 17466 32224
rect 17497 32215 17555 32221
rect 17497 32212 17509 32215
rect 17460 32184 17509 32212
rect 17460 32172 17466 32184
rect 17497 32181 17509 32184
rect 17543 32181 17555 32215
rect 17497 32175 17555 32181
rect 17586 32172 17592 32224
rect 17644 32172 17650 32224
rect 18414 32172 18420 32224
rect 18472 32172 18478 32224
rect 20165 32215 20223 32221
rect 20165 32181 20177 32215
rect 20211 32212 20223 32215
rect 20898 32212 20904 32224
rect 20211 32184 20904 32212
rect 20211 32181 20223 32184
rect 20165 32175 20223 32181
rect 20898 32172 20904 32184
rect 20956 32172 20962 32224
rect 21008 32212 21036 32240
rect 21269 32215 21327 32221
rect 21269 32212 21281 32215
rect 21008 32184 21281 32212
rect 21269 32181 21281 32184
rect 21315 32181 21327 32215
rect 21269 32175 21327 32181
rect 21542 32172 21548 32224
rect 21600 32212 21606 32224
rect 21744 32212 21772 32320
rect 22281 32317 22293 32351
rect 22327 32348 22339 32351
rect 22554 32348 22560 32360
rect 22327 32320 22560 32348
rect 22327 32317 22339 32320
rect 22281 32311 22339 32317
rect 22554 32308 22560 32320
rect 22612 32348 22618 32360
rect 23385 32351 23443 32357
rect 23385 32348 23397 32351
rect 22612 32320 23397 32348
rect 22612 32308 22618 32320
rect 23385 32317 23397 32320
rect 23431 32317 23443 32351
rect 23658 32348 23664 32360
rect 23619 32320 23664 32348
rect 23385 32311 23443 32317
rect 23658 32308 23664 32320
rect 23716 32308 23722 32360
rect 23934 32348 23940 32360
rect 23895 32320 23940 32348
rect 23934 32308 23940 32320
rect 23992 32308 23998 32360
rect 26145 32351 26203 32357
rect 26145 32317 26157 32351
rect 26191 32348 26203 32351
rect 26418 32348 26424 32360
rect 26191 32320 26424 32348
rect 26191 32317 26203 32320
rect 26145 32311 26203 32317
rect 26418 32308 26424 32320
rect 26476 32308 26482 32360
rect 27154 32308 27160 32360
rect 27212 32348 27218 32360
rect 27341 32351 27399 32357
rect 27341 32348 27353 32351
rect 27212 32320 27353 32348
rect 27212 32308 27218 32320
rect 27341 32317 27353 32320
rect 27387 32348 27399 32351
rect 27617 32351 27675 32357
rect 27617 32348 27629 32351
rect 27387 32320 27629 32348
rect 27387 32317 27399 32320
rect 27341 32311 27399 32317
rect 27617 32317 27629 32320
rect 27663 32317 27675 32351
rect 28276 32348 28304 32515
rect 28442 32512 28448 32524
rect 28500 32512 28506 32564
rect 28902 32552 28908 32564
rect 28863 32524 28908 32552
rect 28902 32512 28908 32524
rect 28960 32512 28966 32564
rect 28460 32484 28488 32512
rect 29178 32484 29184 32496
rect 28460 32456 29184 32484
rect 29178 32444 29184 32456
rect 29236 32484 29242 32496
rect 29457 32487 29515 32493
rect 29457 32484 29469 32487
rect 29236 32456 29469 32484
rect 29236 32444 29242 32456
rect 29457 32453 29469 32456
rect 29503 32453 29515 32487
rect 29457 32447 29515 32453
rect 28629 32351 28687 32357
rect 28629 32348 28641 32351
rect 28276 32320 28641 32348
rect 27617 32311 27675 32317
rect 28629 32317 28641 32320
rect 28675 32317 28687 32351
rect 28629 32311 28687 32317
rect 22097 32283 22155 32289
rect 22097 32249 22109 32283
rect 22143 32280 22155 32283
rect 22462 32280 22468 32292
rect 22143 32252 22468 32280
rect 22143 32249 22155 32252
rect 22097 32243 22155 32249
rect 22462 32240 22468 32252
rect 22520 32280 22526 32292
rect 22520 32252 23152 32280
rect 22520 32240 22526 32252
rect 21600 32184 21772 32212
rect 21600 32172 21606 32184
rect 22922 32172 22928 32224
rect 22980 32212 22986 32224
rect 23017 32215 23075 32221
rect 23017 32212 23029 32215
rect 22980 32184 23029 32212
rect 22980 32172 22986 32184
rect 23017 32181 23029 32184
rect 23063 32181 23075 32215
rect 23124 32212 23152 32252
rect 26234 32240 26240 32292
rect 26292 32280 26298 32292
rect 26973 32283 27031 32289
rect 26973 32280 26985 32283
rect 26292 32252 26985 32280
rect 26292 32240 26298 32252
rect 26973 32249 26985 32252
rect 27019 32249 27031 32283
rect 26973 32243 27031 32249
rect 25682 32212 25688 32224
rect 23124 32184 25688 32212
rect 23017 32175 23075 32181
rect 25682 32172 25688 32184
rect 25740 32172 25746 32224
rect 26326 32212 26332 32224
rect 26287 32184 26332 32212
rect 26326 32172 26332 32184
rect 26384 32172 26390 32224
rect 26418 32172 26424 32224
rect 26476 32212 26482 32224
rect 26605 32215 26663 32221
rect 26605 32212 26617 32215
rect 26476 32184 26617 32212
rect 26476 32172 26482 32184
rect 26605 32181 26617 32184
rect 26651 32181 26663 32215
rect 26605 32175 26663 32181
rect 1104 32122 38824 32144
rect 1104 32070 19606 32122
rect 19658 32070 19670 32122
rect 19722 32070 19734 32122
rect 19786 32070 19798 32122
rect 19850 32070 38824 32122
rect 1104 32048 38824 32070
rect 6914 31968 6920 32020
rect 6972 32008 6978 32020
rect 7377 32011 7435 32017
rect 7377 32008 7389 32011
rect 6972 31980 7389 32008
rect 6972 31968 6978 31980
rect 7377 31977 7389 31980
rect 7423 32008 7435 32011
rect 7834 32008 7840 32020
rect 7423 31980 7840 32008
rect 7423 31977 7435 31980
rect 7377 31971 7435 31977
rect 7834 31968 7840 31980
rect 7892 31968 7898 32020
rect 8481 32011 8539 32017
rect 8481 31977 8493 32011
rect 8527 32008 8539 32011
rect 9030 32008 9036 32020
rect 8527 31980 9036 32008
rect 8527 31977 8539 31980
rect 8481 31971 8539 31977
rect 9030 31968 9036 31980
rect 9088 31968 9094 32020
rect 10134 31968 10140 32020
rect 10192 32008 10198 32020
rect 10321 32011 10379 32017
rect 10321 32008 10333 32011
rect 10192 31980 10333 32008
rect 10192 31968 10198 31980
rect 10321 31977 10333 31980
rect 10367 32008 10379 32011
rect 10594 32008 10600 32020
rect 10367 31980 10600 32008
rect 10367 31977 10379 31980
rect 10321 31971 10379 31977
rect 10594 31968 10600 31980
rect 10652 31968 10658 32020
rect 12805 32011 12863 32017
rect 12805 31977 12817 32011
rect 12851 32008 12863 32011
rect 12986 32008 12992 32020
rect 12851 31980 12992 32008
rect 12851 31977 12863 31980
rect 12805 31971 12863 31977
rect 12986 31968 12992 31980
rect 13044 31968 13050 32020
rect 13262 32008 13268 32020
rect 13223 31980 13268 32008
rect 13262 31968 13268 31980
rect 13320 31968 13326 32020
rect 14458 32008 14464 32020
rect 13464 31980 14464 32008
rect 7282 31900 7288 31952
rect 7340 31940 7346 31952
rect 8021 31943 8079 31949
rect 8021 31940 8033 31943
rect 7340 31912 8033 31940
rect 7340 31900 7346 31912
rect 8021 31909 8033 31912
rect 8067 31909 8079 31943
rect 10226 31940 10232 31952
rect 8021 31903 8079 31909
rect 9876 31912 10232 31940
rect 7561 31875 7619 31881
rect 7561 31841 7573 31875
rect 7607 31872 7619 31875
rect 8570 31872 8576 31884
rect 7607 31844 8064 31872
rect 8531 31844 8576 31872
rect 7607 31841 7619 31844
rect 7561 31835 7619 31841
rect 8036 31816 8064 31844
rect 8570 31832 8576 31844
rect 8628 31832 8634 31884
rect 9876 31872 9904 31912
rect 10226 31900 10232 31912
rect 10284 31900 10290 31952
rect 12710 31900 12716 31952
rect 12768 31940 12774 31952
rect 13464 31949 13492 31980
rect 14458 31968 14464 31980
rect 14516 32008 14522 32020
rect 14642 32008 14648 32020
rect 14516 31980 14648 32008
rect 14516 31968 14522 31980
rect 14642 31968 14648 31980
rect 14700 31968 14706 32020
rect 15746 31968 15752 32020
rect 15804 32008 15810 32020
rect 16022 32008 16028 32020
rect 15804 31980 16028 32008
rect 15804 31968 15810 31980
rect 16022 31968 16028 31980
rect 16080 31968 16086 32020
rect 16114 31968 16120 32020
rect 16172 32008 16178 32020
rect 16485 32011 16543 32017
rect 16485 32008 16497 32011
rect 16172 31980 16497 32008
rect 16172 31968 16178 31980
rect 16485 31977 16497 31980
rect 16531 31977 16543 32011
rect 16485 31971 16543 31977
rect 16666 31968 16672 32020
rect 16724 32008 16730 32020
rect 18966 32008 18972 32020
rect 16724 31980 18552 32008
rect 18927 31980 18972 32008
rect 16724 31968 16730 31980
rect 13081 31943 13139 31949
rect 13081 31940 13093 31943
rect 12768 31912 13093 31940
rect 12768 31900 12774 31912
rect 13081 31909 13093 31912
rect 13127 31940 13139 31943
rect 13449 31943 13507 31949
rect 13449 31940 13461 31943
rect 13127 31912 13461 31940
rect 13127 31909 13139 31912
rect 13081 31903 13139 31909
rect 13449 31909 13461 31912
rect 13495 31909 13507 31943
rect 13814 31940 13820 31952
rect 13775 31912 13820 31940
rect 13449 31903 13507 31909
rect 13814 31900 13820 31912
rect 13872 31900 13878 31952
rect 14001 31943 14059 31949
rect 14001 31909 14013 31943
rect 14047 31940 14059 31943
rect 15764 31940 15792 31968
rect 14047 31912 14136 31940
rect 14047 31909 14059 31912
rect 14001 31903 14059 31909
rect 9784 31844 9904 31872
rect 10045 31875 10103 31881
rect 9784 31816 9812 31844
rect 10045 31841 10057 31875
rect 10091 31872 10103 31875
rect 11146 31872 11152 31884
rect 10091 31844 11152 31872
rect 10091 31841 10103 31844
rect 10045 31835 10103 31841
rect 11146 31832 11152 31844
rect 11204 31832 11210 31884
rect 13906 31832 13912 31884
rect 13964 31872 13970 31884
rect 13964 31844 14009 31872
rect 13964 31832 13970 31844
rect 7650 31764 7656 31816
rect 7708 31764 7714 31816
rect 8018 31764 8024 31816
rect 8076 31764 8082 31816
rect 8938 31764 8944 31816
rect 8996 31804 9002 31816
rect 9125 31807 9183 31813
rect 9125 31804 9137 31807
rect 8996 31776 9137 31804
rect 8996 31764 9002 31776
rect 9125 31773 9137 31776
rect 9171 31804 9183 31807
rect 9171 31776 9536 31804
rect 9171 31773 9183 31776
rect 9125 31767 9183 31773
rect 7668 31736 7696 31764
rect 9508 31748 9536 31776
rect 9766 31764 9772 31816
rect 9824 31764 9830 31816
rect 9858 31764 9864 31816
rect 9916 31804 9922 31816
rect 10505 31807 10563 31813
rect 10505 31804 10517 31807
rect 9916 31776 10517 31804
rect 9916 31764 9922 31776
rect 10505 31773 10517 31776
rect 10551 31773 10563 31807
rect 10778 31804 10784 31816
rect 10739 31776 10784 31804
rect 10505 31767 10563 31773
rect 10778 31764 10784 31776
rect 10836 31764 10842 31816
rect 10962 31764 10968 31816
rect 11020 31804 11026 31816
rect 13538 31804 13544 31816
rect 11020 31776 13544 31804
rect 11020 31764 11026 31776
rect 13538 31764 13544 31776
rect 13596 31804 13602 31816
rect 13633 31807 13691 31813
rect 13633 31804 13645 31807
rect 13596 31776 13645 31804
rect 13596 31764 13602 31776
rect 13633 31773 13645 31776
rect 13679 31773 13691 31807
rect 13633 31767 13691 31773
rect 7745 31739 7803 31745
rect 7745 31736 7757 31739
rect 7668 31708 7757 31736
rect 7745 31705 7757 31708
rect 7791 31705 7803 31739
rect 8754 31736 8760 31748
rect 8715 31708 8760 31736
rect 7745 31699 7803 31705
rect 8754 31696 8760 31708
rect 8812 31696 8818 31748
rect 9490 31736 9496 31748
rect 9403 31708 9496 31736
rect 9490 31696 9496 31708
rect 9548 31696 9554 31748
rect 12250 31696 12256 31748
rect 12308 31736 12314 31748
rect 12434 31736 12440 31748
rect 12308 31708 12440 31736
rect 12308 31696 12314 31708
rect 12434 31696 12440 31708
rect 12492 31696 12498 31748
rect 12526 31696 12532 31748
rect 12584 31736 12590 31748
rect 12802 31736 12808 31748
rect 12584 31708 12808 31736
rect 12584 31696 12590 31708
rect 12802 31696 12808 31708
rect 12860 31736 12866 31748
rect 14108 31736 14136 31912
rect 15580 31912 15792 31940
rect 14366 31872 14372 31884
rect 14327 31844 14372 31872
rect 14366 31832 14372 31844
rect 14424 31832 14430 31884
rect 14642 31832 14648 31884
rect 14700 31872 14706 31884
rect 14918 31872 14924 31884
rect 14700 31844 14924 31872
rect 14700 31832 14706 31844
rect 14918 31832 14924 31844
rect 14976 31832 14982 31884
rect 15580 31881 15608 31912
rect 15838 31900 15844 31952
rect 15896 31940 15902 31952
rect 15896 31912 16344 31940
rect 15896 31900 15902 31912
rect 15565 31875 15623 31881
rect 15565 31841 15577 31875
rect 15611 31841 15623 31875
rect 15746 31872 15752 31884
rect 15707 31844 15752 31872
rect 15565 31835 15623 31841
rect 15746 31832 15752 31844
rect 15804 31832 15810 31884
rect 16114 31872 16120 31884
rect 16075 31844 16120 31872
rect 16114 31832 16120 31844
rect 16172 31832 16178 31884
rect 15105 31807 15163 31813
rect 15105 31773 15117 31807
rect 15151 31804 15163 31807
rect 16132 31804 16160 31832
rect 15151 31776 16160 31804
rect 16316 31804 16344 31912
rect 16390 31900 16396 31952
rect 16448 31940 16454 31952
rect 16448 31912 17632 31940
rect 16448 31900 16454 31912
rect 16669 31875 16727 31881
rect 16669 31841 16681 31875
rect 16715 31872 16727 31875
rect 16758 31872 16764 31884
rect 16715 31844 16764 31872
rect 16715 31841 16727 31844
rect 16669 31835 16727 31841
rect 16758 31832 16764 31844
rect 16816 31832 16822 31884
rect 17604 31881 17632 31912
rect 17589 31875 17647 31881
rect 17589 31841 17601 31875
rect 17635 31841 17647 31875
rect 18322 31872 18328 31884
rect 18283 31844 18328 31872
rect 17589 31835 17647 31841
rect 18322 31832 18328 31844
rect 18380 31832 18386 31884
rect 18417 31875 18475 31881
rect 18417 31841 18429 31875
rect 18463 31841 18475 31875
rect 18524 31872 18552 31980
rect 18966 31968 18972 31980
rect 19024 31968 19030 32020
rect 20254 32008 20260 32020
rect 19628 31980 20260 32008
rect 19628 31952 19656 31980
rect 20254 31968 20260 31980
rect 20312 31968 20318 32020
rect 20806 31968 20812 32020
rect 20864 32008 20870 32020
rect 21177 32011 21235 32017
rect 21177 32008 21189 32011
rect 20864 31980 21189 32008
rect 20864 31968 20870 31980
rect 21177 31977 21189 31980
rect 21223 31977 21235 32011
rect 21177 31971 21235 31977
rect 21266 31968 21272 32020
rect 21324 32008 21330 32020
rect 21542 32008 21548 32020
rect 21324 31980 21548 32008
rect 21324 31968 21330 31980
rect 21542 31968 21548 31980
rect 21600 31968 21606 32020
rect 23290 32008 23296 32020
rect 23251 31980 23296 32008
rect 23290 31968 23296 31980
rect 23348 31968 23354 32020
rect 24210 32008 24216 32020
rect 23768 31980 24216 32008
rect 19610 31900 19616 31952
rect 19668 31900 19674 31952
rect 19886 31900 19892 31952
rect 19944 31940 19950 31952
rect 19981 31943 20039 31949
rect 19981 31940 19993 31943
rect 19944 31912 19993 31940
rect 19944 31900 19950 31912
rect 19981 31909 19993 31912
rect 20027 31940 20039 31943
rect 20530 31940 20536 31952
rect 20027 31912 20536 31940
rect 20027 31909 20039 31912
rect 19981 31903 20039 31909
rect 20530 31900 20536 31912
rect 20588 31900 20594 31952
rect 22830 31940 22836 31952
rect 22791 31912 22836 31940
rect 22830 31900 22836 31912
rect 22888 31900 22894 31952
rect 23768 31949 23796 31980
rect 24210 31968 24216 31980
rect 24268 31968 24274 32020
rect 24854 32008 24860 32020
rect 24815 31980 24860 32008
rect 24854 31968 24860 31980
rect 24912 31968 24918 32020
rect 25038 31968 25044 32020
rect 25096 32008 25102 32020
rect 25133 32011 25191 32017
rect 25133 32008 25145 32011
rect 25096 31980 25145 32008
rect 25096 31968 25102 31980
rect 25133 31977 25145 31980
rect 25179 31977 25191 32011
rect 25133 31971 25191 31977
rect 27706 31968 27712 32020
rect 27764 31968 27770 32020
rect 23753 31943 23811 31949
rect 23753 31909 23765 31943
rect 23799 31909 23811 31943
rect 23753 31903 23811 31909
rect 24118 31900 24124 31952
rect 24176 31940 24182 31952
rect 24397 31943 24455 31949
rect 24397 31940 24409 31943
rect 24176 31912 24409 31940
rect 24176 31900 24182 31912
rect 24397 31909 24409 31912
rect 24443 31909 24455 31943
rect 24397 31903 24455 31909
rect 25590 31900 25596 31952
rect 25648 31940 25654 31952
rect 26145 31943 26203 31949
rect 26145 31940 26157 31943
rect 25648 31912 26157 31940
rect 25648 31900 25654 31912
rect 26145 31909 26157 31912
rect 26191 31909 26203 31943
rect 26145 31903 26203 31909
rect 18785 31875 18843 31881
rect 18785 31872 18797 31875
rect 18524 31844 18797 31872
rect 18417 31835 18475 31841
rect 18785 31841 18797 31844
rect 18831 31841 18843 31875
rect 18785 31835 18843 31841
rect 16574 31804 16580 31816
rect 16316 31776 16580 31804
rect 15151 31773 15163 31776
rect 15105 31767 15163 31773
rect 16574 31764 16580 31776
rect 16632 31764 16638 31816
rect 17497 31807 17555 31813
rect 17497 31773 17509 31807
rect 17543 31804 17555 31807
rect 17954 31804 17960 31816
rect 17543 31776 17960 31804
rect 17543 31773 17555 31776
rect 17497 31767 17555 31773
rect 17954 31764 17960 31776
rect 18012 31764 18018 31816
rect 18432 31804 18460 31835
rect 20254 31832 20260 31884
rect 20312 31872 20318 31884
rect 20438 31872 20444 31884
rect 20312 31844 20444 31872
rect 20312 31832 20318 31844
rect 20438 31832 20444 31844
rect 20496 31832 20502 31884
rect 21358 31872 21364 31884
rect 21319 31844 21364 31872
rect 21358 31832 21364 31844
rect 21416 31832 21422 31884
rect 21450 31832 21456 31884
rect 21508 31872 21514 31884
rect 21545 31875 21603 31881
rect 21545 31872 21557 31875
rect 21508 31844 21557 31872
rect 21508 31832 21514 31844
rect 21545 31841 21557 31844
rect 21591 31841 21603 31875
rect 21545 31835 21603 31841
rect 21913 31875 21971 31881
rect 21913 31841 21925 31875
rect 21959 31841 21971 31875
rect 22462 31872 22468 31884
rect 22423 31844 22468 31872
rect 21913 31835 21971 31841
rect 18874 31804 18880 31816
rect 18432 31776 18880 31804
rect 18874 31764 18880 31776
rect 18932 31804 18938 31816
rect 19334 31804 19340 31816
rect 18932 31776 19340 31804
rect 18932 31764 18938 31776
rect 19334 31764 19340 31776
rect 19392 31764 19398 31816
rect 20714 31764 20720 31816
rect 20772 31804 20778 31816
rect 21634 31804 21640 31816
rect 20772 31776 21640 31804
rect 20772 31764 20778 31776
rect 21634 31764 21640 31776
rect 21692 31804 21698 31816
rect 21928 31804 21956 31835
rect 22462 31832 22468 31844
rect 22520 31832 22526 31884
rect 23106 31832 23112 31884
rect 23164 31872 23170 31884
rect 23569 31875 23627 31881
rect 23569 31872 23581 31875
rect 23164 31844 23581 31872
rect 23164 31832 23170 31844
rect 23569 31841 23581 31844
rect 23615 31841 23627 31875
rect 23569 31835 23627 31841
rect 23661 31875 23719 31881
rect 23661 31841 23673 31875
rect 23707 31872 23719 31875
rect 24762 31872 24768 31884
rect 23707 31844 24768 31872
rect 23707 31841 23719 31844
rect 23661 31835 23719 31841
rect 24762 31832 24768 31844
rect 24820 31832 24826 31884
rect 24946 31872 24952 31884
rect 24907 31844 24952 31872
rect 24946 31832 24952 31844
rect 25004 31832 25010 31884
rect 26786 31832 26792 31884
rect 26844 31872 26850 31884
rect 26973 31875 27031 31881
rect 26973 31872 26985 31875
rect 26844 31844 26985 31872
rect 26844 31832 26850 31844
rect 26973 31841 26985 31844
rect 27019 31872 27031 31875
rect 27724 31872 27752 31968
rect 28074 31900 28080 31952
rect 28132 31940 28138 31952
rect 28718 31940 28724 31952
rect 28132 31912 28724 31940
rect 28132 31900 28138 31912
rect 28718 31900 28724 31912
rect 28776 31900 28782 31952
rect 29178 31872 29184 31884
rect 27019 31844 27752 31872
rect 29139 31844 29184 31872
rect 27019 31841 27031 31844
rect 26973 31835 27031 31841
rect 29178 31832 29184 31844
rect 29236 31832 29242 31884
rect 29454 31872 29460 31884
rect 29415 31844 29460 31872
rect 29454 31832 29460 31844
rect 29512 31832 29518 31884
rect 23290 31804 23296 31816
rect 21692 31776 21956 31804
rect 22112 31776 23296 31804
rect 21692 31764 21698 31776
rect 12860 31708 14136 31736
rect 12860 31696 12866 31708
rect 19886 31696 19892 31748
rect 19944 31736 19950 31748
rect 22112 31736 22140 31776
rect 23290 31764 23296 31776
rect 23348 31764 23354 31816
rect 23385 31807 23443 31813
rect 23385 31773 23397 31807
rect 23431 31773 23443 31807
rect 23385 31767 23443 31773
rect 24121 31807 24179 31813
rect 24121 31773 24133 31807
rect 24167 31804 24179 31807
rect 24302 31804 24308 31816
rect 24167 31776 24308 31804
rect 24167 31773 24179 31776
rect 24121 31767 24179 31773
rect 19944 31708 22140 31736
rect 23400 31736 23428 31767
rect 24302 31764 24308 31776
rect 24360 31764 24366 31816
rect 25130 31804 25136 31816
rect 24872 31776 25136 31804
rect 23934 31736 23940 31748
rect 23400 31708 23940 31736
rect 19944 31696 19950 31708
rect 23934 31696 23940 31708
rect 23992 31696 23998 31748
rect 7101 31671 7159 31677
rect 7101 31637 7113 31671
rect 7147 31668 7159 31671
rect 7558 31668 7564 31680
rect 7147 31640 7564 31668
rect 7147 31637 7159 31640
rect 7101 31631 7159 31637
rect 7558 31628 7564 31640
rect 7616 31628 7622 31680
rect 11146 31628 11152 31680
rect 11204 31668 11210 31680
rect 11514 31668 11520 31680
rect 11204 31640 11520 31668
rect 11204 31628 11210 31640
rect 11514 31628 11520 31640
rect 11572 31628 11578 31680
rect 11790 31628 11796 31680
rect 11848 31668 11854 31680
rect 11885 31671 11943 31677
rect 11885 31668 11897 31671
rect 11848 31640 11897 31668
rect 11848 31628 11854 31640
rect 11885 31637 11897 31640
rect 11931 31637 11943 31671
rect 11885 31631 11943 31637
rect 13265 31671 13323 31677
rect 13265 31637 13277 31671
rect 13311 31668 13323 31671
rect 13446 31668 13452 31680
rect 13311 31640 13452 31668
rect 13311 31637 13323 31640
rect 13265 31631 13323 31637
rect 13446 31628 13452 31640
rect 13504 31628 13510 31680
rect 16666 31628 16672 31680
rect 16724 31668 16730 31680
rect 17037 31671 17095 31677
rect 17037 31668 17049 31671
rect 16724 31640 17049 31668
rect 16724 31628 16730 31640
rect 17037 31637 17049 31640
rect 17083 31637 17095 31671
rect 17037 31631 17095 31637
rect 19334 31628 19340 31680
rect 19392 31668 19398 31680
rect 19613 31671 19671 31677
rect 19613 31668 19625 31671
rect 19392 31640 19625 31668
rect 19392 31628 19398 31640
rect 19613 31637 19625 31640
rect 19659 31637 19671 31671
rect 19613 31631 19671 31637
rect 20717 31671 20775 31677
rect 20717 31637 20729 31671
rect 20763 31668 20775 31671
rect 20806 31668 20812 31680
rect 20763 31640 20812 31668
rect 20763 31637 20775 31640
rect 20717 31631 20775 31637
rect 20806 31628 20812 31640
rect 20864 31628 20870 31680
rect 21266 31628 21272 31680
rect 21324 31668 21330 31680
rect 24872 31668 24900 31776
rect 25130 31764 25136 31776
rect 25188 31804 25194 31816
rect 25409 31807 25467 31813
rect 25409 31804 25421 31807
rect 25188 31776 25421 31804
rect 25188 31764 25194 31776
rect 25409 31773 25421 31776
rect 25455 31773 25467 31807
rect 25409 31767 25467 31773
rect 26697 31807 26755 31813
rect 26697 31773 26709 31807
rect 26743 31804 26755 31807
rect 27338 31804 27344 31816
rect 26743 31776 27344 31804
rect 26743 31773 26755 31776
rect 26697 31767 26755 31773
rect 27338 31764 27344 31776
rect 27396 31764 27402 31816
rect 27614 31764 27620 31816
rect 27672 31804 27678 31816
rect 28077 31807 28135 31813
rect 28077 31804 28089 31807
rect 27672 31776 28089 31804
rect 27672 31764 27678 31776
rect 28077 31773 28089 31776
rect 28123 31773 28135 31807
rect 30558 31804 30564 31816
rect 30519 31776 30564 31804
rect 28077 31767 28135 31773
rect 30558 31764 30564 31776
rect 30616 31764 30622 31816
rect 25774 31736 25780 31748
rect 25687 31708 25780 31736
rect 25774 31696 25780 31708
rect 25832 31736 25838 31748
rect 25832 31708 26556 31736
rect 25832 31696 25838 31708
rect 21324 31640 24900 31668
rect 26528 31668 26556 31708
rect 27706 31668 27712 31680
rect 26528 31640 27712 31668
rect 21324 31628 21330 31640
rect 27706 31628 27712 31640
rect 27764 31628 27770 31680
rect 1104 31578 38824 31600
rect 1104 31526 4246 31578
rect 4298 31526 4310 31578
rect 4362 31526 4374 31578
rect 4426 31526 4438 31578
rect 4490 31526 34966 31578
rect 35018 31526 35030 31578
rect 35082 31526 35094 31578
rect 35146 31526 35158 31578
rect 35210 31526 38824 31578
rect 1104 31504 38824 31526
rect 8478 31424 8484 31476
rect 8536 31464 8542 31476
rect 8754 31464 8760 31476
rect 8536 31436 8760 31464
rect 8536 31424 8542 31436
rect 8754 31424 8760 31436
rect 8812 31424 8818 31476
rect 11882 31464 11888 31476
rect 11843 31436 11888 31464
rect 11882 31424 11888 31436
rect 11940 31424 11946 31476
rect 12434 31424 12440 31476
rect 12492 31464 12498 31476
rect 13262 31464 13268 31476
rect 12492 31436 13268 31464
rect 12492 31424 12498 31436
rect 13262 31424 13268 31436
rect 13320 31424 13326 31476
rect 13814 31464 13820 31476
rect 13775 31436 13820 31464
rect 13814 31424 13820 31436
rect 13872 31424 13878 31476
rect 15838 31464 15844 31476
rect 15799 31436 15844 31464
rect 15838 31424 15844 31436
rect 15896 31424 15902 31476
rect 19334 31424 19340 31476
rect 19392 31464 19398 31476
rect 19392 31436 21220 31464
rect 19392 31424 19398 31436
rect 10870 31356 10876 31408
rect 10928 31396 10934 31408
rect 10928 31368 13492 31396
rect 10928 31356 10934 31368
rect 6641 31331 6699 31337
rect 6641 31297 6653 31331
rect 6687 31328 6699 31331
rect 7558 31328 7564 31340
rect 6687 31300 7564 31328
rect 6687 31297 6699 31300
rect 6641 31291 6699 31297
rect 7558 31288 7564 31300
rect 7616 31288 7622 31340
rect 7834 31328 7840 31340
rect 7795 31300 7840 31328
rect 7834 31288 7840 31300
rect 7892 31288 7898 31340
rect 10689 31331 10747 31337
rect 10689 31297 10701 31331
rect 10735 31328 10747 31331
rect 10781 31331 10839 31337
rect 10781 31328 10793 31331
rect 10735 31300 10793 31328
rect 10735 31297 10747 31300
rect 10689 31291 10747 31297
rect 10781 31297 10793 31300
rect 10827 31328 10839 31331
rect 10962 31328 10968 31340
rect 10827 31300 10968 31328
rect 10827 31297 10839 31300
rect 10781 31291 10839 31297
rect 10962 31288 10968 31300
rect 11020 31288 11026 31340
rect 11054 31288 11060 31340
rect 11112 31328 11118 31340
rect 11112 31300 11192 31328
rect 11112 31288 11118 31300
rect 11164 31260 11192 31300
rect 11514 31288 11520 31340
rect 11572 31288 11578 31340
rect 13464 31328 13492 31368
rect 13538 31356 13544 31408
rect 13596 31396 13602 31408
rect 14093 31399 14151 31405
rect 14093 31396 14105 31399
rect 13596 31368 14105 31396
rect 13596 31356 13602 31368
rect 14093 31365 14105 31368
rect 14139 31365 14151 31399
rect 14093 31359 14151 31365
rect 15286 31356 15292 31408
rect 15344 31396 15350 31408
rect 16209 31399 16267 31405
rect 16209 31396 16221 31399
rect 15344 31368 16221 31396
rect 15344 31356 15350 31368
rect 16209 31365 16221 31368
rect 16255 31396 16267 31399
rect 16298 31396 16304 31408
rect 16255 31368 16304 31396
rect 16255 31365 16267 31368
rect 16209 31359 16267 31365
rect 16298 31356 16304 31368
rect 16356 31396 16362 31408
rect 16356 31368 16436 31396
rect 16356 31356 16362 31368
rect 13464 31300 14412 31328
rect 11532 31260 11560 31288
rect 14384 31272 14412 31300
rect 14458 31288 14464 31340
rect 14516 31328 14522 31340
rect 14737 31331 14795 31337
rect 14737 31328 14749 31331
rect 14516 31300 14749 31328
rect 14516 31288 14522 31300
rect 14737 31297 14749 31300
rect 14783 31297 14795 31331
rect 15470 31328 15476 31340
rect 15431 31300 15476 31328
rect 14737 31291 14795 31297
rect 15470 31288 15476 31300
rect 15528 31288 15534 31340
rect 16408 31337 16436 31368
rect 17678 31356 17684 31408
rect 17736 31396 17742 31408
rect 19521 31399 19579 31405
rect 19521 31396 19533 31399
rect 17736 31368 19533 31396
rect 17736 31356 17742 31368
rect 19521 31365 19533 31368
rect 19567 31396 19579 31399
rect 19567 31368 21128 31396
rect 19567 31365 19579 31368
rect 19521 31359 19579 31365
rect 16393 31331 16451 31337
rect 16393 31297 16405 31331
rect 16439 31297 16451 31331
rect 16393 31291 16451 31297
rect 16574 31288 16580 31340
rect 16632 31328 16638 31340
rect 17129 31331 17187 31337
rect 17129 31328 17141 31331
rect 16632 31300 17141 31328
rect 16632 31288 16638 31300
rect 17129 31297 17141 31300
rect 17175 31297 17187 31331
rect 17129 31291 17187 31297
rect 18785 31331 18843 31337
rect 18785 31297 18797 31331
rect 18831 31328 18843 31331
rect 19058 31328 19064 31340
rect 18831 31300 19064 31328
rect 18831 31297 18843 31300
rect 18785 31291 18843 31297
rect 19058 31288 19064 31300
rect 19116 31288 19122 31340
rect 19334 31288 19340 31340
rect 19392 31328 19398 31340
rect 19613 31331 19671 31337
rect 19613 31328 19625 31331
rect 19392 31300 19625 31328
rect 19392 31288 19398 31300
rect 19613 31297 19625 31300
rect 19659 31297 19671 31331
rect 19613 31291 19671 31297
rect 11164 31232 11560 31260
rect 10321 31195 10379 31201
rect 10321 31161 10333 31195
rect 10367 31192 10379 31195
rect 10502 31192 10508 31204
rect 10367 31164 10508 31192
rect 10367 31161 10379 31164
rect 10321 31155 10379 31161
rect 10502 31152 10508 31164
rect 10560 31192 10566 31204
rect 11164 31201 11192 31232
rect 11974 31220 11980 31272
rect 12032 31260 12038 31272
rect 12437 31263 12495 31269
rect 12437 31260 12449 31263
rect 12032 31232 12449 31260
rect 12032 31220 12038 31232
rect 12437 31229 12449 31232
rect 12483 31229 12495 31263
rect 12894 31260 12900 31272
rect 12855 31232 12900 31260
rect 12437 31223 12495 31229
rect 12894 31220 12900 31232
rect 12952 31220 12958 31272
rect 13262 31260 13268 31272
rect 13223 31232 13268 31260
rect 13262 31220 13268 31232
rect 13320 31220 13326 31272
rect 13357 31263 13415 31269
rect 13357 31229 13369 31263
rect 13403 31260 13415 31263
rect 13446 31260 13452 31272
rect 13403 31232 13452 31260
rect 13403 31229 13415 31232
rect 13357 31223 13415 31229
rect 13446 31220 13452 31232
rect 13504 31220 13510 31272
rect 14366 31220 14372 31272
rect 14424 31220 14430 31272
rect 14921 31263 14979 31269
rect 14921 31229 14933 31263
rect 14967 31260 14979 31263
rect 15010 31260 15016 31272
rect 14967 31232 15016 31260
rect 14967 31229 14979 31232
rect 14921 31223 14979 31229
rect 15010 31220 15016 31232
rect 15068 31220 15074 31272
rect 17310 31260 17316 31272
rect 16684 31232 17316 31260
rect 11057 31195 11115 31201
rect 11057 31192 11069 31195
rect 10560 31164 11069 31192
rect 10560 31152 10566 31164
rect 11057 31161 11069 31164
rect 11103 31161 11115 31195
rect 11057 31155 11115 31161
rect 11149 31195 11207 31201
rect 11149 31161 11161 31195
rect 11195 31161 11207 31195
rect 11149 31155 11207 31161
rect 11517 31195 11575 31201
rect 11517 31161 11529 31195
rect 11563 31192 11575 31195
rect 11882 31192 11888 31204
rect 11563 31164 11888 31192
rect 11563 31161 11575 31164
rect 11517 31155 11575 31161
rect 7006 31124 7012 31136
rect 6967 31096 7012 31124
rect 7006 31084 7012 31096
rect 7064 31084 7070 31136
rect 7466 31124 7472 31136
rect 7427 31096 7472 31124
rect 7466 31084 7472 31096
rect 7524 31084 7530 31136
rect 8941 31127 8999 31133
rect 8941 31093 8953 31127
rect 8987 31124 8999 31127
rect 9030 31124 9036 31136
rect 8987 31096 9036 31124
rect 8987 31093 8999 31096
rect 8941 31087 8999 31093
rect 9030 31084 9036 31096
rect 9088 31084 9094 31136
rect 9582 31124 9588 31136
rect 9543 31096 9588 31124
rect 9582 31084 9588 31096
rect 9640 31084 9646 31136
rect 9950 31124 9956 31136
rect 9863 31096 9956 31124
rect 9950 31084 9956 31096
rect 10008 31124 10014 31136
rect 10226 31124 10232 31136
rect 10008 31096 10232 31124
rect 10008 31084 10014 31096
rect 10226 31084 10232 31096
rect 10284 31084 10290 31136
rect 10962 31124 10968 31136
rect 10923 31096 10968 31124
rect 10962 31084 10968 31096
rect 11020 31084 11026 31136
rect 11072 31124 11100 31155
rect 11882 31152 11888 31164
rect 11940 31152 11946 31204
rect 15105 31195 15163 31201
rect 12084 31164 13308 31192
rect 12084 31124 12112 31164
rect 13280 31136 13308 31164
rect 15105 31161 15117 31195
rect 15151 31192 15163 31195
rect 15286 31192 15292 31204
rect 15151 31164 15292 31192
rect 15151 31161 15163 31164
rect 15105 31155 15163 31161
rect 15286 31152 15292 31164
rect 15344 31152 15350 31204
rect 15838 31152 15844 31204
rect 15896 31192 15902 31204
rect 16684 31201 16712 31232
rect 17310 31220 17316 31232
rect 17368 31220 17374 31272
rect 17586 31220 17592 31272
rect 17644 31260 17650 31272
rect 19812 31269 19840 31368
rect 19886 31288 19892 31340
rect 19944 31328 19950 31340
rect 19944 31300 20024 31328
rect 19944 31288 19950 31300
rect 18325 31263 18383 31269
rect 18325 31260 18337 31263
rect 17644 31232 18337 31260
rect 17644 31220 17650 31232
rect 18325 31229 18337 31232
rect 18371 31229 18383 31263
rect 18325 31223 18383 31229
rect 19797 31263 19855 31269
rect 19797 31229 19809 31263
rect 19843 31229 19855 31263
rect 19797 31223 19855 31229
rect 16669 31195 16727 31201
rect 16669 31192 16681 31195
rect 15896 31164 16681 31192
rect 15896 31152 15902 31164
rect 16669 31161 16681 31164
rect 16715 31161 16727 31195
rect 16669 31155 16727 31161
rect 16758 31152 16764 31204
rect 16816 31192 16822 31204
rect 17218 31192 17224 31204
rect 16816 31164 17224 31192
rect 16816 31152 16822 31164
rect 17218 31152 17224 31164
rect 17276 31152 17282 31204
rect 17865 31195 17923 31201
rect 17865 31161 17877 31195
rect 17911 31192 17923 31195
rect 18046 31192 18052 31204
rect 17911 31164 18052 31192
rect 17911 31161 17923 31164
rect 17865 31155 17923 31161
rect 18046 31152 18052 31164
rect 18104 31152 18110 31204
rect 18417 31195 18475 31201
rect 18417 31161 18429 31195
rect 18463 31192 18475 31195
rect 18598 31192 18604 31204
rect 18463 31164 18604 31192
rect 18463 31161 18475 31164
rect 18417 31155 18475 31161
rect 18598 31152 18604 31164
rect 18656 31192 18662 31204
rect 19996 31201 20024 31300
rect 21100 31269 21128 31368
rect 21192 31337 21220 31436
rect 21450 31424 21456 31476
rect 21508 31464 21514 31476
rect 22557 31467 22615 31473
rect 22557 31464 22569 31467
rect 21508 31436 22569 31464
rect 21508 31424 21514 31436
rect 22557 31433 22569 31436
rect 22603 31433 22615 31467
rect 23106 31464 23112 31476
rect 23067 31436 23112 31464
rect 22557 31427 22615 31433
rect 23106 31424 23112 31436
rect 23164 31424 23170 31476
rect 24486 31424 24492 31476
rect 24544 31464 24550 31476
rect 24946 31464 24952 31476
rect 24544 31436 24952 31464
rect 24544 31424 24550 31436
rect 24946 31424 24952 31436
rect 25004 31424 25010 31476
rect 26050 31464 26056 31476
rect 26011 31436 26056 31464
rect 26050 31424 26056 31436
rect 26108 31424 26114 31476
rect 26786 31464 26792 31476
rect 26747 31436 26792 31464
rect 26786 31424 26792 31436
rect 26844 31424 26850 31476
rect 26970 31424 26976 31476
rect 27028 31464 27034 31476
rect 27065 31467 27123 31473
rect 27065 31464 27077 31467
rect 27028 31436 27077 31464
rect 27028 31424 27034 31436
rect 27065 31433 27077 31436
rect 27111 31433 27123 31467
rect 27430 31464 27436 31476
rect 27391 31436 27436 31464
rect 27065 31427 27123 31433
rect 27430 31424 27436 31436
rect 27488 31424 27494 31476
rect 28074 31464 28080 31476
rect 28035 31436 28080 31464
rect 28074 31424 28080 31436
rect 28132 31424 28138 31476
rect 29454 31464 29460 31476
rect 29415 31436 29460 31464
rect 29454 31424 29460 31436
rect 29512 31424 29518 31476
rect 23477 31399 23535 31405
rect 23477 31365 23489 31399
rect 23523 31396 23535 31399
rect 24026 31396 24032 31408
rect 23523 31368 24032 31396
rect 23523 31365 23535 31368
rect 23477 31359 23535 31365
rect 24026 31356 24032 31368
rect 24084 31356 24090 31408
rect 21177 31331 21235 31337
rect 21177 31297 21189 31331
rect 21223 31328 21235 31331
rect 21634 31328 21640 31340
rect 21223 31300 21640 31328
rect 21223 31297 21235 31300
rect 21177 31291 21235 31297
rect 21634 31288 21640 31300
rect 21692 31288 21698 31340
rect 21913 31331 21971 31337
rect 21913 31297 21925 31331
rect 21959 31328 21971 31331
rect 22002 31328 22008 31340
rect 21959 31300 22008 31328
rect 21959 31297 21971 31300
rect 21913 31291 21971 31297
rect 22002 31288 22008 31300
rect 22060 31288 22066 31340
rect 23661 31331 23719 31337
rect 23661 31297 23673 31331
rect 23707 31328 23719 31331
rect 23934 31328 23940 31340
rect 23707 31300 23940 31328
rect 23707 31297 23719 31300
rect 23661 31291 23719 31297
rect 23934 31288 23940 31300
rect 23992 31288 23998 31340
rect 25685 31331 25743 31337
rect 25685 31328 25697 31331
rect 24044 31300 25697 31328
rect 21085 31263 21143 31269
rect 21085 31229 21097 31263
rect 21131 31260 21143 31263
rect 21361 31263 21419 31269
rect 21361 31260 21373 31263
rect 21131 31232 21373 31260
rect 21131 31229 21143 31232
rect 21085 31223 21143 31229
rect 21361 31229 21373 31232
rect 21407 31260 21419 31263
rect 21450 31260 21456 31272
rect 21407 31232 21456 31260
rect 21407 31229 21419 31232
rect 21361 31223 21419 31229
rect 21450 31220 21456 31232
rect 21508 31220 21514 31272
rect 23474 31220 23480 31272
rect 23532 31260 23538 31272
rect 24044 31260 24072 31300
rect 25685 31297 25697 31300
rect 25731 31328 25743 31331
rect 25774 31328 25780 31340
rect 25731 31300 25780 31328
rect 25731 31297 25743 31300
rect 25685 31291 25743 31297
rect 25774 31288 25780 31300
rect 25832 31288 25838 31340
rect 28442 31328 28448 31340
rect 25884 31300 28448 31328
rect 23532 31232 24072 31260
rect 23532 31220 23538 31232
rect 19061 31195 19119 31201
rect 19061 31192 19073 31195
rect 18656 31164 19073 31192
rect 18656 31152 18662 31164
rect 19061 31161 19073 31164
rect 19107 31192 19119 31195
rect 19889 31195 19947 31201
rect 19889 31192 19901 31195
rect 19107 31164 19656 31192
rect 19107 31161 19119 31164
rect 19061 31155 19119 31161
rect 12250 31124 12256 31136
rect 11072 31096 12112 31124
rect 12211 31096 12256 31124
rect 12250 31084 12256 31096
rect 12308 31084 12314 31136
rect 13262 31084 13268 31136
rect 13320 31124 13326 31136
rect 14553 31127 14611 31133
rect 14553 31124 14565 31127
rect 13320 31096 14565 31124
rect 13320 31084 13326 31096
rect 14553 31093 14565 31096
rect 14599 31124 14611 31127
rect 15013 31127 15071 31133
rect 15013 31124 15025 31127
rect 14599 31096 15025 31124
rect 14599 31093 14611 31096
rect 14553 31087 14611 31093
rect 15013 31093 15025 31096
rect 15059 31093 15071 31127
rect 16574 31124 16580 31136
rect 16535 31096 16580 31124
rect 15013 31087 15071 31093
rect 16574 31084 16580 31096
rect 16632 31084 16638 31136
rect 17497 31127 17555 31133
rect 17497 31093 17509 31127
rect 17543 31124 17555 31127
rect 17954 31124 17960 31136
rect 17543 31096 17960 31124
rect 17543 31093 17555 31096
rect 17497 31087 17555 31093
rect 17954 31084 17960 31096
rect 18012 31124 18018 31136
rect 18233 31127 18291 31133
rect 18233 31124 18245 31127
rect 18012 31096 18245 31124
rect 18012 31084 18018 31096
rect 18233 31093 18245 31096
rect 18279 31124 18291 31127
rect 19426 31124 19432 31136
rect 18279 31096 19432 31124
rect 18279 31093 18291 31096
rect 18233 31087 18291 31093
rect 19426 31084 19432 31096
rect 19484 31084 19490 31136
rect 19628 31124 19656 31164
rect 19812 31164 19901 31192
rect 19812 31124 19840 31164
rect 19889 31161 19901 31164
rect 19935 31161 19947 31195
rect 19889 31155 19947 31161
rect 19981 31195 20039 31201
rect 19981 31161 19993 31195
rect 20027 31161 20039 31195
rect 20346 31192 20352 31204
rect 20307 31164 20352 31192
rect 19981 31155 20039 31161
rect 19628 31096 19840 31124
rect 19904 31124 19932 31155
rect 20346 31152 20352 31164
rect 20404 31152 20410 31204
rect 21545 31195 21603 31201
rect 21545 31161 21557 31195
rect 21591 31192 21603 31195
rect 22646 31192 22652 31204
rect 21591 31164 22652 31192
rect 21591 31161 21603 31164
rect 21545 31155 21603 31161
rect 22646 31152 22652 31164
rect 22704 31192 22710 31204
rect 22830 31192 22836 31204
rect 22704 31164 22836 31192
rect 22704 31152 22710 31164
rect 22830 31152 22836 31164
rect 22888 31152 22894 31204
rect 23750 31152 23756 31204
rect 23808 31192 23814 31204
rect 24044 31201 24072 31232
rect 25225 31263 25283 31269
rect 25225 31229 25237 31263
rect 25271 31260 25283 31263
rect 25314 31260 25320 31272
rect 25271 31232 25320 31260
rect 25271 31229 25283 31232
rect 25225 31223 25283 31229
rect 25314 31220 25320 31232
rect 25372 31260 25378 31272
rect 25884 31260 25912 31300
rect 28442 31288 28448 31300
rect 28500 31288 28506 31340
rect 26234 31260 26240 31272
rect 25372 31232 25912 31260
rect 26195 31232 26240 31260
rect 25372 31220 25378 31232
rect 26234 31220 26240 31232
rect 26292 31220 26298 31272
rect 27246 31260 27252 31272
rect 27207 31232 27252 31260
rect 27246 31220 27252 31232
rect 27304 31260 27310 31272
rect 27709 31263 27767 31269
rect 27709 31260 27721 31263
rect 27304 31232 27721 31260
rect 27304 31220 27310 31232
rect 27709 31229 27721 31232
rect 27755 31229 27767 31263
rect 27709 31223 27767 31229
rect 23845 31195 23903 31201
rect 23845 31192 23857 31195
rect 23808 31164 23857 31192
rect 23808 31152 23814 31164
rect 23845 31161 23857 31164
rect 23891 31161 23903 31195
rect 23845 31155 23903 31161
rect 24029 31195 24087 31201
rect 24029 31161 24041 31195
rect 24075 31161 24087 31195
rect 24029 31155 24087 31161
rect 24397 31195 24455 31201
rect 24397 31161 24409 31195
rect 24443 31192 24455 31195
rect 24486 31192 24492 31204
rect 24443 31164 24492 31192
rect 24443 31161 24455 31164
rect 24397 31155 24455 31161
rect 24486 31152 24492 31164
rect 24544 31152 24550 31204
rect 24762 31152 24768 31204
rect 24820 31192 24826 31204
rect 25133 31195 25191 31201
rect 25133 31192 25145 31195
rect 24820 31164 25145 31192
rect 24820 31152 24826 31164
rect 25133 31161 25145 31164
rect 25179 31192 25191 31195
rect 26326 31192 26332 31204
rect 25179 31164 26332 31192
rect 25179 31161 25191 31164
rect 25133 31155 25191 31161
rect 26326 31152 26332 31164
rect 26384 31152 26390 31204
rect 20625 31127 20683 31133
rect 20625 31124 20637 31127
rect 19904 31096 20637 31124
rect 20625 31093 20637 31096
rect 20671 31124 20683 31127
rect 21450 31124 21456 31136
rect 20671 31096 21456 31124
rect 20671 31093 20683 31096
rect 20625 31087 20683 31093
rect 21450 31084 21456 31096
rect 21508 31084 21514 31136
rect 21634 31084 21640 31136
rect 21692 31124 21698 31136
rect 22189 31127 22247 31133
rect 22189 31124 22201 31127
rect 21692 31096 22201 31124
rect 21692 31084 21698 31096
rect 22189 31093 22201 31096
rect 22235 31093 22247 31127
rect 22189 31087 22247 31093
rect 22462 31084 22468 31136
rect 22520 31124 22526 31136
rect 23106 31124 23112 31136
rect 22520 31096 23112 31124
rect 22520 31084 22526 31096
rect 23106 31084 23112 31096
rect 23164 31084 23170 31136
rect 23382 31084 23388 31136
rect 23440 31124 23446 31136
rect 23768 31124 23796 31152
rect 23440 31096 23796 31124
rect 23937 31127 23995 31133
rect 23440 31084 23446 31096
rect 23937 31093 23949 31127
rect 23983 31124 23995 31127
rect 24673 31127 24731 31133
rect 24673 31124 24685 31127
rect 23983 31096 24685 31124
rect 23983 31093 23995 31096
rect 23937 31087 23995 31093
rect 24673 31093 24685 31096
rect 24719 31124 24731 31127
rect 24946 31124 24952 31136
rect 24719 31096 24952 31124
rect 24719 31093 24731 31096
rect 24673 31087 24731 31093
rect 24946 31084 24952 31096
rect 25004 31084 25010 31136
rect 25406 31124 25412 31136
rect 25367 31096 25412 31124
rect 25406 31084 25412 31096
rect 25464 31084 25470 31136
rect 26421 31127 26479 31133
rect 26421 31093 26433 31127
rect 26467 31124 26479 31127
rect 26786 31124 26792 31136
rect 26467 31096 26792 31124
rect 26467 31093 26479 31096
rect 26421 31087 26479 31093
rect 26786 31084 26792 31096
rect 26844 31084 26850 31136
rect 28718 31084 28724 31136
rect 28776 31124 28782 31136
rect 28813 31127 28871 31133
rect 28813 31124 28825 31127
rect 28776 31096 28825 31124
rect 28776 31084 28782 31096
rect 28813 31093 28825 31096
rect 28859 31093 28871 31127
rect 28813 31087 28871 31093
rect 29178 31084 29184 31136
rect 29236 31124 29242 31136
rect 29454 31124 29460 31136
rect 29236 31096 29460 31124
rect 29236 31084 29242 31096
rect 29454 31084 29460 31096
rect 29512 31124 29518 31136
rect 29825 31127 29883 31133
rect 29825 31124 29837 31127
rect 29512 31096 29837 31124
rect 29512 31084 29518 31096
rect 29825 31093 29837 31096
rect 29871 31093 29883 31127
rect 29825 31087 29883 31093
rect 1104 31034 38824 31056
rect 1104 30982 19606 31034
rect 19658 30982 19670 31034
rect 19722 30982 19734 31034
rect 19786 30982 19798 31034
rect 19850 30982 38824 31034
rect 1104 30960 38824 30982
rect 6733 30923 6791 30929
rect 6733 30889 6745 30923
rect 6779 30920 6791 30923
rect 7006 30920 7012 30932
rect 6779 30892 7012 30920
rect 6779 30889 6791 30892
rect 6733 30883 6791 30889
rect 7006 30880 7012 30892
rect 7064 30880 7070 30932
rect 7742 30920 7748 30932
rect 7703 30892 7748 30920
rect 7742 30880 7748 30892
rect 7800 30880 7806 30932
rect 8570 30880 8576 30932
rect 8628 30920 8634 30932
rect 8757 30923 8815 30929
rect 8757 30920 8769 30923
rect 8628 30892 8769 30920
rect 8628 30880 8634 30892
rect 8757 30889 8769 30892
rect 8803 30920 8815 30923
rect 9582 30920 9588 30932
rect 8803 30892 9588 30920
rect 8803 30889 8815 30892
rect 8757 30883 8815 30889
rect 9582 30880 9588 30892
rect 9640 30880 9646 30932
rect 10321 30923 10379 30929
rect 10321 30889 10333 30923
rect 10367 30920 10379 30923
rect 10778 30920 10784 30932
rect 10367 30892 10784 30920
rect 10367 30889 10379 30892
rect 10321 30883 10379 30889
rect 10336 30852 10364 30883
rect 10778 30880 10784 30892
rect 10836 30880 10842 30932
rect 11238 30920 11244 30932
rect 11199 30892 11244 30920
rect 11238 30880 11244 30892
rect 11296 30880 11302 30932
rect 11514 30880 11520 30932
rect 11572 30920 11578 30932
rect 11698 30920 11704 30932
rect 11572 30892 11704 30920
rect 11572 30880 11578 30892
rect 11698 30880 11704 30892
rect 11756 30880 11762 30932
rect 12434 30880 12440 30932
rect 12492 30920 12498 30932
rect 13541 30923 13599 30929
rect 13541 30920 13553 30923
rect 12492 30892 13553 30920
rect 12492 30880 12498 30892
rect 13541 30889 13553 30892
rect 13587 30920 13599 30923
rect 13722 30920 13728 30932
rect 13587 30892 13728 30920
rect 13587 30889 13599 30892
rect 13541 30883 13599 30889
rect 13722 30880 13728 30892
rect 13780 30880 13786 30932
rect 15194 30920 15200 30932
rect 13924 30892 15200 30920
rect 12526 30852 12532 30864
rect 9968 30824 10364 30852
rect 11624 30824 12532 30852
rect 7558 30784 7564 30796
rect 7519 30756 7564 30784
rect 7558 30744 7564 30756
rect 7616 30744 7622 30796
rect 8573 30787 8631 30793
rect 8573 30753 8585 30787
rect 8619 30784 8631 30787
rect 9122 30784 9128 30796
rect 8619 30756 9128 30784
rect 8619 30753 8631 30756
rect 8573 30747 8631 30753
rect 9122 30744 9128 30756
rect 9180 30744 9186 30796
rect 7469 30719 7527 30725
rect 7469 30685 7481 30719
rect 7515 30716 7527 30719
rect 8110 30716 8116 30728
rect 7515 30688 8116 30716
rect 7515 30685 7527 30688
rect 7469 30679 7527 30685
rect 8110 30676 8116 30688
rect 8168 30716 8174 30728
rect 9033 30719 9091 30725
rect 9033 30716 9045 30719
rect 8168 30688 9045 30716
rect 8168 30676 8174 30688
rect 9033 30685 9045 30688
rect 9079 30685 9091 30719
rect 9033 30679 9091 30685
rect 7101 30651 7159 30657
rect 7101 30617 7113 30651
rect 7147 30648 7159 30651
rect 8202 30648 8208 30660
rect 7147 30620 8208 30648
rect 7147 30617 7159 30620
rect 7101 30611 7159 30617
rect 8202 30608 8208 30620
rect 8260 30608 8266 30660
rect 9122 30608 9128 30660
rect 9180 30648 9186 30660
rect 9968 30648 9996 30824
rect 10137 30787 10195 30793
rect 10137 30753 10149 30787
rect 10183 30784 10195 30787
rect 10870 30784 10876 30796
rect 10183 30756 10876 30784
rect 10183 30753 10195 30756
rect 10137 30747 10195 30753
rect 10870 30744 10876 30756
rect 10928 30744 10934 30796
rect 11624 30725 11652 30824
rect 12526 30812 12532 30824
rect 12584 30812 12590 30864
rect 13817 30855 13875 30861
rect 13817 30821 13829 30855
rect 13863 30852 13875 30855
rect 13924 30852 13952 30892
rect 14200 30864 14228 30892
rect 15194 30880 15200 30892
rect 15252 30920 15258 30932
rect 15473 30923 15531 30929
rect 15473 30920 15485 30923
rect 15252 30892 15485 30920
rect 15252 30880 15258 30892
rect 15473 30889 15485 30892
rect 15519 30889 15531 30923
rect 15473 30883 15531 30889
rect 16206 30880 16212 30932
rect 16264 30920 16270 30932
rect 18049 30923 18107 30929
rect 16264 30892 17080 30920
rect 16264 30880 16270 30892
rect 13863 30824 13952 30852
rect 14001 30855 14059 30861
rect 13863 30821 13875 30824
rect 13817 30815 13875 30821
rect 14001 30821 14013 30855
rect 14047 30821 14059 30855
rect 14001 30815 14059 30821
rect 11790 30784 11796 30796
rect 11751 30756 11796 30784
rect 11790 30744 11796 30756
rect 11848 30744 11854 30796
rect 11974 30744 11980 30796
rect 12032 30784 12038 30796
rect 12161 30787 12219 30793
rect 12161 30784 12173 30787
rect 12032 30756 12173 30784
rect 12032 30744 12038 30756
rect 12161 30753 12173 30756
rect 12207 30753 12219 30787
rect 12161 30747 12219 30753
rect 12618 30744 12624 30796
rect 12676 30784 12682 30796
rect 13909 30787 13967 30793
rect 13909 30784 13921 30787
rect 12676 30756 13921 30784
rect 12676 30744 12682 30756
rect 13909 30753 13921 30756
rect 13955 30753 13967 30787
rect 14016 30784 14044 30815
rect 14182 30812 14188 30864
rect 14240 30812 14246 30864
rect 14369 30855 14427 30861
rect 14369 30821 14381 30855
rect 14415 30852 14427 30855
rect 14918 30852 14924 30864
rect 14415 30824 14924 30852
rect 14415 30821 14427 30824
rect 14369 30815 14427 30821
rect 14918 30812 14924 30824
rect 14976 30812 14982 30864
rect 16298 30852 16304 30864
rect 16259 30824 16304 30852
rect 16298 30812 16304 30824
rect 16356 30812 16362 30864
rect 16669 30855 16727 30861
rect 16669 30821 16681 30855
rect 16715 30852 16727 30855
rect 16850 30852 16856 30864
rect 16715 30824 16856 30852
rect 16715 30821 16727 30824
rect 16669 30815 16727 30821
rect 16850 30812 16856 30824
rect 16908 30812 16914 30864
rect 17052 30861 17080 30892
rect 18049 30889 18061 30923
rect 18095 30920 18107 30923
rect 18322 30920 18328 30932
rect 18095 30892 18328 30920
rect 18095 30889 18107 30892
rect 18049 30883 18107 30889
rect 18322 30880 18328 30892
rect 18380 30880 18386 30932
rect 18690 30880 18696 30932
rect 18748 30920 18754 30932
rect 18785 30923 18843 30929
rect 18785 30920 18797 30923
rect 18748 30892 18797 30920
rect 18748 30880 18754 30892
rect 18785 30889 18797 30892
rect 18831 30889 18843 30923
rect 19242 30920 19248 30932
rect 19203 30892 19248 30920
rect 18785 30883 18843 30889
rect 19242 30880 19248 30892
rect 19300 30880 19306 30932
rect 20714 30920 20720 30932
rect 20675 30892 20720 30920
rect 20714 30880 20720 30892
rect 20772 30880 20778 30932
rect 21082 30880 21088 30932
rect 21140 30920 21146 30932
rect 21177 30923 21235 30929
rect 21177 30920 21189 30923
rect 21140 30892 21189 30920
rect 21140 30880 21146 30892
rect 21177 30889 21189 30892
rect 21223 30889 21235 30923
rect 21177 30883 21235 30889
rect 21358 30880 21364 30932
rect 21416 30920 21422 30932
rect 21913 30923 21971 30929
rect 21913 30920 21925 30923
rect 21416 30892 21925 30920
rect 21416 30880 21422 30892
rect 21913 30889 21925 30892
rect 21959 30889 21971 30923
rect 22922 30920 22928 30932
rect 22883 30892 22928 30920
rect 21913 30883 21971 30889
rect 22922 30880 22928 30892
rect 22980 30880 22986 30932
rect 23658 30880 23664 30932
rect 23716 30920 23722 30932
rect 23753 30923 23811 30929
rect 23753 30920 23765 30923
rect 23716 30892 23765 30920
rect 23716 30880 23722 30892
rect 23753 30889 23765 30892
rect 23799 30920 23811 30923
rect 23934 30920 23940 30932
rect 23799 30892 23940 30920
rect 23799 30889 23811 30892
rect 23753 30883 23811 30889
rect 23934 30880 23940 30892
rect 23992 30880 23998 30932
rect 24673 30923 24731 30929
rect 24673 30889 24685 30923
rect 24719 30889 24731 30923
rect 24673 30883 24731 30889
rect 17037 30855 17095 30861
rect 17037 30821 17049 30855
rect 17083 30821 17095 30855
rect 17037 30815 17095 30821
rect 18141 30855 18199 30861
rect 18141 30821 18153 30855
rect 18187 30852 18199 30855
rect 20346 30852 20352 30864
rect 18187 30824 20352 30852
rect 18187 30821 18199 30824
rect 18141 30815 18199 30821
rect 20346 30812 20352 30824
rect 20404 30812 20410 30864
rect 21266 30852 21272 30864
rect 21227 30824 21272 30852
rect 21266 30812 21272 30824
rect 21324 30812 21330 30864
rect 21637 30855 21695 30861
rect 21637 30821 21649 30855
rect 21683 30852 21695 30855
rect 21726 30852 21732 30864
rect 21683 30824 21732 30852
rect 21683 30821 21695 30824
rect 21637 30815 21695 30821
rect 21726 30812 21732 30824
rect 21784 30812 21790 30864
rect 22373 30855 22431 30861
rect 22373 30821 22385 30855
rect 22419 30852 22431 30855
rect 23106 30852 23112 30864
rect 22419 30824 23112 30852
rect 22419 30821 22431 30824
rect 22373 30815 22431 30821
rect 23106 30812 23112 30824
rect 23164 30852 23170 30864
rect 24688 30852 24716 30883
rect 24854 30880 24860 30932
rect 24912 30920 24918 30932
rect 25961 30923 26019 30929
rect 25961 30920 25973 30923
rect 24912 30892 25973 30920
rect 24912 30880 24918 30892
rect 25961 30889 25973 30892
rect 26007 30889 26019 30923
rect 25961 30883 26019 30889
rect 23164 30824 24716 30852
rect 23164 30812 23170 30824
rect 14458 30784 14464 30796
rect 14016 30756 14464 30784
rect 13909 30747 13967 30753
rect 10045 30719 10103 30725
rect 10045 30685 10057 30719
rect 10091 30716 10103 30719
rect 11609 30719 11667 30725
rect 11609 30716 11621 30719
rect 10091 30688 11621 30716
rect 10091 30685 10103 30688
rect 10045 30679 10103 30685
rect 11609 30685 11621 30688
rect 11655 30685 11667 30719
rect 11609 30679 11667 30685
rect 11698 30676 11704 30728
rect 11756 30716 11762 30728
rect 12069 30719 12127 30725
rect 12069 30716 12081 30719
rect 11756 30688 12081 30716
rect 11756 30676 11762 30688
rect 12069 30685 12081 30688
rect 12115 30685 12127 30719
rect 12069 30679 12127 30685
rect 12713 30719 12771 30725
rect 12713 30685 12725 30719
rect 12759 30716 12771 30719
rect 12894 30716 12900 30728
rect 12759 30688 12900 30716
rect 12759 30685 12771 30688
rect 12713 30679 12771 30685
rect 12894 30676 12900 30688
rect 12952 30676 12958 30728
rect 13173 30719 13231 30725
rect 13173 30685 13185 30719
rect 13219 30716 13231 30719
rect 13633 30719 13691 30725
rect 13633 30716 13645 30719
rect 13219 30688 13645 30716
rect 13219 30685 13231 30688
rect 13173 30679 13231 30685
rect 13633 30685 13645 30688
rect 13679 30716 13691 30719
rect 13722 30716 13728 30728
rect 13679 30688 13728 30716
rect 13679 30685 13691 30688
rect 13633 30679 13691 30685
rect 13722 30676 13728 30688
rect 13780 30676 13786 30728
rect 9180 30620 9996 30648
rect 9180 30608 9186 30620
rect 10226 30608 10232 30660
rect 10284 30648 10290 30660
rect 10284 30620 11100 30648
rect 10284 30608 10290 30620
rect 8113 30583 8171 30589
rect 8113 30549 8125 30583
rect 8159 30580 8171 30583
rect 8294 30580 8300 30592
rect 8159 30552 8300 30580
rect 8159 30549 8171 30552
rect 8113 30543 8171 30549
rect 8294 30540 8300 30552
rect 8352 30540 8358 30592
rect 8478 30580 8484 30592
rect 8439 30552 8484 30580
rect 8478 30540 8484 30552
rect 8536 30540 8542 30592
rect 9306 30540 9312 30592
rect 9364 30580 9370 30592
rect 9401 30583 9459 30589
rect 9401 30580 9413 30583
rect 9364 30552 9413 30580
rect 9364 30540 9370 30552
rect 9401 30549 9413 30552
rect 9447 30549 9459 30583
rect 9401 30543 9459 30549
rect 10873 30583 10931 30589
rect 10873 30549 10885 30583
rect 10919 30580 10931 30583
rect 10962 30580 10968 30592
rect 10919 30552 10968 30580
rect 10919 30549 10931 30552
rect 10873 30543 10931 30549
rect 10962 30540 10968 30552
rect 11020 30540 11026 30592
rect 11072 30580 11100 30620
rect 12802 30608 12808 30660
rect 12860 30648 12866 30660
rect 13078 30648 13084 30660
rect 12860 30620 13084 30648
rect 12860 30608 12866 30620
rect 13078 30608 13084 30620
rect 13136 30608 13142 30660
rect 13924 30648 13952 30747
rect 14458 30744 14464 30756
rect 14516 30744 14522 30796
rect 14826 30744 14832 30796
rect 14884 30784 14890 30796
rect 15013 30787 15071 30793
rect 15013 30784 15025 30787
rect 14884 30756 15025 30784
rect 14884 30744 14890 30756
rect 15013 30753 15025 30756
rect 15059 30753 15071 30787
rect 15013 30747 15071 30753
rect 15289 30787 15347 30793
rect 15289 30753 15301 30787
rect 15335 30784 15347 30787
rect 16206 30784 16212 30796
rect 15335 30756 16212 30784
rect 15335 30753 15347 30756
rect 15289 30747 15347 30753
rect 16206 30744 16212 30756
rect 16264 30784 16270 30796
rect 16485 30787 16543 30793
rect 16485 30784 16497 30787
rect 16264 30756 16497 30784
rect 16264 30744 16270 30756
rect 16485 30753 16497 30756
rect 16531 30753 16543 30787
rect 16485 30747 16543 30753
rect 16577 30787 16635 30793
rect 16577 30753 16589 30787
rect 16623 30784 16635 30787
rect 16758 30784 16764 30796
rect 16623 30756 16764 30784
rect 16623 30753 16635 30756
rect 16577 30747 16635 30753
rect 16758 30744 16764 30756
rect 16816 30784 16822 30796
rect 17126 30784 17132 30796
rect 16816 30756 17132 30784
rect 16816 30744 16822 30756
rect 17126 30744 17132 30756
rect 17184 30784 17190 30796
rect 17313 30787 17371 30793
rect 17313 30784 17325 30787
rect 17184 30756 17325 30784
rect 17184 30744 17190 30756
rect 17313 30753 17325 30756
rect 17359 30753 17371 30787
rect 17313 30747 17371 30753
rect 17954 30744 17960 30796
rect 18012 30784 18018 30796
rect 18012 30756 18552 30784
rect 18012 30744 18018 30756
rect 14737 30719 14795 30725
rect 14737 30685 14749 30719
rect 14783 30716 14795 30719
rect 15102 30716 15108 30728
rect 14783 30688 15108 30716
rect 14783 30685 14795 30688
rect 14737 30679 14795 30685
rect 15102 30676 15108 30688
rect 15160 30676 15166 30728
rect 18230 30676 18236 30728
rect 18288 30676 18294 30728
rect 18524 30725 18552 30756
rect 18598 30744 18604 30796
rect 18656 30784 18662 30796
rect 19613 30787 19671 30793
rect 19613 30784 19625 30787
rect 18656 30756 19625 30784
rect 18656 30744 18662 30756
rect 19613 30753 19625 30756
rect 19659 30753 19671 30787
rect 19613 30747 19671 30753
rect 19797 30787 19855 30793
rect 19797 30753 19809 30787
rect 19843 30784 19855 30787
rect 21085 30787 21143 30793
rect 19843 30756 20392 30784
rect 19843 30753 19855 30756
rect 19797 30747 19855 30753
rect 18509 30719 18567 30725
rect 18509 30685 18521 30719
rect 18555 30716 18567 30719
rect 19978 30716 19984 30728
rect 18555 30688 19984 30716
rect 18555 30685 18567 30688
rect 18509 30679 18567 30685
rect 19978 30676 19984 30688
rect 20036 30676 20042 30728
rect 16942 30648 16948 30660
rect 13924 30620 16948 30648
rect 16942 30608 16948 30620
rect 17000 30608 17006 30660
rect 18248 30648 18276 30676
rect 20364 30660 20392 30756
rect 21085 30753 21097 30787
rect 21131 30784 21143 30787
rect 21358 30784 21364 30796
rect 21131 30756 21364 30784
rect 21131 30753 21143 30756
rect 21085 30747 21143 30753
rect 21358 30744 21364 30756
rect 21416 30744 21422 30796
rect 22278 30744 22284 30796
rect 22336 30784 22342 30796
rect 22465 30787 22523 30793
rect 22465 30784 22477 30787
rect 22336 30756 22477 30784
rect 22336 30744 22342 30756
rect 22465 30753 22477 30756
rect 22511 30753 22523 30787
rect 22465 30747 22523 30753
rect 22741 30787 22799 30793
rect 22741 30753 22753 30787
rect 22787 30784 22799 30787
rect 22830 30784 22836 30796
rect 22787 30756 22836 30784
rect 22787 30753 22799 30756
rect 22741 30747 22799 30753
rect 22830 30744 22836 30756
rect 22888 30744 22894 30796
rect 24029 30787 24087 30793
rect 24029 30753 24041 30787
rect 24075 30784 24087 30787
rect 24486 30784 24492 30796
rect 24075 30756 24492 30784
rect 24075 30753 24087 30756
rect 24029 30747 24087 30753
rect 24486 30744 24492 30756
rect 24544 30784 24550 30796
rect 24854 30784 24860 30796
rect 24544 30756 24860 30784
rect 24544 30744 24550 30756
rect 24854 30744 24860 30756
rect 24912 30744 24918 30796
rect 20714 30676 20720 30728
rect 20772 30716 20778 30728
rect 20901 30719 20959 30725
rect 20901 30716 20913 30719
rect 20772 30688 20913 30716
rect 20772 30676 20778 30688
rect 20901 30685 20913 30688
rect 20947 30716 20959 30719
rect 22002 30716 22008 30728
rect 20947 30688 22008 30716
rect 20947 30685 20959 30688
rect 20901 30679 20959 30685
rect 22002 30676 22008 30688
rect 22060 30676 22066 30728
rect 24397 30719 24455 30725
rect 24397 30685 24409 30719
rect 24443 30716 24455 30719
rect 24670 30716 24676 30728
rect 24443 30688 24676 30716
rect 24443 30685 24455 30688
rect 24397 30679 24455 30685
rect 24670 30676 24676 30688
rect 24728 30676 24734 30728
rect 27157 30719 27215 30725
rect 27157 30685 27169 30719
rect 27203 30716 27215 30719
rect 27338 30716 27344 30728
rect 27203 30688 27344 30716
rect 27203 30685 27215 30688
rect 27157 30679 27215 30685
rect 27338 30676 27344 30688
rect 27396 30676 27402 30728
rect 27433 30719 27491 30725
rect 27433 30685 27445 30719
rect 27479 30716 27491 30719
rect 27522 30716 27528 30728
rect 27479 30688 27528 30716
rect 27479 30685 27491 30688
rect 27433 30679 27491 30685
rect 27522 30676 27528 30688
rect 27580 30676 27586 30728
rect 18417 30651 18475 30657
rect 18417 30648 18429 30651
rect 18248 30620 18429 30648
rect 18417 30617 18429 30620
rect 18463 30617 18475 30651
rect 20346 30648 20352 30660
rect 20307 30620 20352 30648
rect 18417 30611 18475 30617
rect 20346 30608 20352 30620
rect 20404 30608 20410 30660
rect 22554 30648 22560 30660
rect 22515 30620 22560 30648
rect 22554 30608 22560 30620
rect 22612 30608 22618 30660
rect 24302 30648 24308 30660
rect 24263 30620 24308 30648
rect 24302 30608 24308 30620
rect 24360 30608 24366 30660
rect 24486 30608 24492 30660
rect 24544 30648 24550 30660
rect 25593 30651 25651 30657
rect 25593 30648 25605 30651
rect 24544 30620 25605 30648
rect 24544 30608 24550 30620
rect 25593 30617 25605 30620
rect 25639 30617 25651 30651
rect 25593 30611 25651 30617
rect 13446 30580 13452 30592
rect 11072 30552 13452 30580
rect 13446 30540 13452 30552
rect 13504 30540 13510 30592
rect 15746 30580 15752 30592
rect 15707 30552 15752 30580
rect 15746 30540 15752 30552
rect 15804 30540 15810 30592
rect 16206 30580 16212 30592
rect 16167 30552 16212 30580
rect 16206 30540 16212 30552
rect 16264 30580 16270 30592
rect 16574 30580 16580 30592
rect 16264 30552 16580 30580
rect 16264 30540 16270 30552
rect 16574 30540 16580 30552
rect 16632 30540 16638 30592
rect 18306 30583 18364 30589
rect 18306 30549 18318 30583
rect 18352 30580 18364 30583
rect 18782 30580 18788 30592
rect 18352 30552 18788 30580
rect 18352 30549 18364 30552
rect 18306 30543 18364 30549
rect 18782 30540 18788 30552
rect 18840 30540 18846 30592
rect 19334 30540 19340 30592
rect 19392 30580 19398 30592
rect 19981 30583 20039 30589
rect 19981 30580 19993 30583
rect 19392 30552 19993 30580
rect 19392 30540 19398 30552
rect 19981 30549 19993 30552
rect 20027 30580 20039 30583
rect 22462 30580 22468 30592
rect 20027 30552 22468 30580
rect 20027 30549 20039 30552
rect 19981 30543 20039 30549
rect 22462 30540 22468 30552
rect 22520 30540 22526 30592
rect 23750 30540 23756 30592
rect 23808 30580 23814 30592
rect 24210 30589 24216 30592
rect 24167 30583 24216 30589
rect 24167 30580 24179 30583
rect 23808 30552 24179 30580
rect 23808 30540 23814 30552
rect 24167 30549 24179 30552
rect 24213 30549 24216 30583
rect 24167 30543 24216 30549
rect 24210 30540 24216 30543
rect 24268 30580 24274 30592
rect 24268 30552 24315 30580
rect 24268 30540 24274 30552
rect 24946 30540 24952 30592
rect 25004 30580 25010 30592
rect 25317 30583 25375 30589
rect 25317 30580 25329 30583
rect 25004 30552 25329 30580
rect 25004 30540 25010 30552
rect 25317 30549 25329 30552
rect 25363 30580 25375 30583
rect 25406 30580 25412 30592
rect 25363 30552 25412 30580
rect 25363 30549 25375 30552
rect 25317 30543 25375 30549
rect 25406 30540 25412 30552
rect 25464 30540 25470 30592
rect 26418 30540 26424 30592
rect 26476 30580 26482 30592
rect 26697 30583 26755 30589
rect 26697 30580 26709 30583
rect 26476 30552 26709 30580
rect 26476 30540 26482 30552
rect 26697 30549 26709 30552
rect 26743 30549 26755 30583
rect 26697 30543 26755 30549
rect 28166 30540 28172 30592
rect 28224 30580 28230 30592
rect 28534 30580 28540 30592
rect 28224 30552 28540 30580
rect 28224 30540 28230 30552
rect 28534 30540 28540 30552
rect 28592 30540 28598 30592
rect 1104 30490 38824 30512
rect 1104 30438 4246 30490
rect 4298 30438 4310 30490
rect 4362 30438 4374 30490
rect 4426 30438 4438 30490
rect 4490 30438 34966 30490
rect 35018 30438 35030 30490
rect 35082 30438 35094 30490
rect 35146 30438 35158 30490
rect 35210 30438 38824 30490
rect 1104 30416 38824 30438
rect 7558 30376 7564 30388
rect 7519 30348 7564 30376
rect 7558 30336 7564 30348
rect 7616 30336 7622 30388
rect 9122 30376 9128 30388
rect 9083 30348 9128 30376
rect 9122 30336 9128 30348
rect 9180 30336 9186 30388
rect 9674 30336 9680 30388
rect 9732 30376 9738 30388
rect 9950 30376 9956 30388
rect 9732 30348 9956 30376
rect 9732 30336 9738 30348
rect 9950 30336 9956 30348
rect 10008 30336 10014 30388
rect 11238 30336 11244 30388
rect 11296 30376 11302 30388
rect 11793 30379 11851 30385
rect 11793 30376 11805 30379
rect 11296 30348 11805 30376
rect 11296 30336 11302 30348
rect 11793 30345 11805 30348
rect 11839 30376 11851 30379
rect 12066 30376 12072 30388
rect 11839 30348 12072 30376
rect 11839 30345 11851 30348
rect 11793 30339 11851 30345
rect 12066 30336 12072 30348
rect 12124 30376 12130 30388
rect 12618 30376 12624 30388
rect 12124 30348 12624 30376
rect 12124 30336 12130 30348
rect 12618 30336 12624 30348
rect 12676 30336 12682 30388
rect 14182 30376 14188 30388
rect 14143 30348 14188 30376
rect 14182 30336 14188 30348
rect 14240 30336 14246 30388
rect 16298 30376 16304 30388
rect 16259 30348 16304 30376
rect 16298 30336 16304 30348
rect 16356 30336 16362 30388
rect 18230 30376 18236 30388
rect 17880 30348 18236 30376
rect 6273 30311 6331 30317
rect 6273 30277 6285 30311
rect 6319 30308 6331 30311
rect 9582 30308 9588 30320
rect 6319 30280 9588 30308
rect 6319 30277 6331 30280
rect 6273 30271 6331 30277
rect 9582 30268 9588 30280
rect 9640 30268 9646 30320
rect 11330 30268 11336 30320
rect 11388 30308 11394 30320
rect 12161 30311 12219 30317
rect 12161 30308 12173 30311
rect 11388 30280 12173 30308
rect 11388 30268 11394 30280
rect 12161 30277 12173 30280
rect 12207 30277 12219 30311
rect 12710 30308 12716 30320
rect 12623 30280 12716 30308
rect 12161 30271 12219 30277
rect 12710 30268 12716 30280
rect 12768 30308 12774 30320
rect 13722 30308 13728 30320
rect 12768 30280 13728 30308
rect 12768 30268 12774 30280
rect 7650 30240 7656 30252
rect 7611 30212 7656 30240
rect 7650 30200 7656 30212
rect 7708 30200 7714 30252
rect 8110 30240 8116 30252
rect 8071 30212 8116 30240
rect 8110 30200 8116 30212
rect 8168 30200 8174 30252
rect 8202 30200 8208 30252
rect 8260 30240 8266 30252
rect 10594 30240 10600 30252
rect 8260 30212 10600 30240
rect 8260 30200 8266 30212
rect 10594 30200 10600 30212
rect 10652 30200 10658 30252
rect 13188 30249 13216 30280
rect 13722 30268 13728 30280
rect 13780 30308 13786 30320
rect 14826 30308 14832 30320
rect 13780 30280 14832 30308
rect 13780 30268 13786 30280
rect 13173 30243 13231 30249
rect 11164 30212 12940 30240
rect 8294 30172 8300 30184
rect 8255 30144 8300 30172
rect 8294 30132 8300 30144
rect 8352 30132 8358 30184
rect 8478 30132 8484 30184
rect 8536 30172 8542 30184
rect 8665 30175 8723 30181
rect 8665 30172 8677 30175
rect 8536 30144 8677 30172
rect 8536 30132 8542 30144
rect 8665 30141 8677 30144
rect 8711 30141 8723 30175
rect 8665 30135 8723 30141
rect 8757 30175 8815 30181
rect 8757 30141 8769 30175
rect 8803 30141 8815 30175
rect 9769 30175 9827 30181
rect 9769 30172 9781 30175
rect 8757 30135 8815 30141
rect 9692 30144 9781 30172
rect 7193 30107 7251 30113
rect 7193 30073 7205 30107
rect 7239 30104 7251 30107
rect 8772 30104 8800 30135
rect 9214 30104 9220 30116
rect 7239 30076 9220 30104
rect 7239 30073 7251 30076
rect 7193 30067 7251 30073
rect 9214 30064 9220 30076
rect 9272 30064 9278 30116
rect 9692 30048 9720 30144
rect 9769 30141 9781 30144
rect 9815 30141 9827 30175
rect 11057 30175 11115 30181
rect 11057 30172 11069 30175
rect 9769 30135 9827 30141
rect 10336 30144 11069 30172
rect 10336 30048 10364 30144
rect 11057 30141 11069 30144
rect 11103 30141 11115 30175
rect 11057 30135 11115 30141
rect 10778 30104 10784 30116
rect 10691 30076 10784 30104
rect 10778 30064 10784 30076
rect 10836 30104 10842 30116
rect 11164 30113 11192 30212
rect 12912 30184 12940 30212
rect 13173 30209 13185 30243
rect 13219 30209 13231 30243
rect 13173 30203 13231 30209
rect 13262 30200 13268 30252
rect 13320 30240 13326 30252
rect 13814 30240 13820 30252
rect 13320 30212 13820 30240
rect 13320 30200 13326 30212
rect 13814 30200 13820 30212
rect 13872 30200 13878 30252
rect 13909 30243 13967 30249
rect 13909 30209 13921 30243
rect 13955 30240 13967 30243
rect 14642 30240 14648 30252
rect 13955 30212 14648 30240
rect 13955 30209 13967 30212
rect 13909 30203 13967 30209
rect 14642 30200 14648 30212
rect 14700 30200 14706 30252
rect 14752 30249 14780 30280
rect 14826 30268 14832 30280
rect 14884 30308 14890 30320
rect 15562 30308 15568 30320
rect 14884 30280 15568 30308
rect 14884 30268 14890 30280
rect 15562 30268 15568 30280
rect 15620 30268 15626 30320
rect 17402 30268 17408 30320
rect 17460 30308 17466 30320
rect 17586 30308 17592 30320
rect 17460 30280 17592 30308
rect 17460 30268 17466 30280
rect 17586 30268 17592 30280
rect 17644 30268 17650 30320
rect 17880 30317 17908 30348
rect 18230 30336 18236 30348
rect 18288 30336 18294 30388
rect 20438 30336 20444 30388
rect 20496 30376 20502 30388
rect 20496 30348 20760 30376
rect 20496 30336 20502 30348
rect 20732 30320 20760 30348
rect 21174 30336 21180 30388
rect 21232 30376 21238 30388
rect 21232 30348 21312 30376
rect 21232 30336 21238 30348
rect 21284 30320 21312 30348
rect 21358 30336 21364 30388
rect 21416 30376 21422 30388
rect 21416 30348 22140 30376
rect 21416 30336 21422 30348
rect 17865 30311 17923 30317
rect 17865 30277 17877 30311
rect 17911 30277 17923 30311
rect 19058 30308 19064 30320
rect 17865 30271 17923 30277
rect 18248 30280 19064 30308
rect 14737 30243 14795 30249
rect 14737 30209 14749 30243
rect 14783 30209 14795 30243
rect 15473 30243 15531 30249
rect 14737 30203 14795 30209
rect 14844 30212 15148 30240
rect 12894 30132 12900 30184
rect 12952 30132 12958 30184
rect 13078 30172 13084 30184
rect 12991 30144 13084 30172
rect 13078 30132 13084 30144
rect 13136 30172 13142 30184
rect 13357 30175 13415 30181
rect 13357 30172 13369 30175
rect 13136 30144 13369 30172
rect 13136 30132 13142 30144
rect 13357 30141 13369 30144
rect 13403 30172 13415 30175
rect 14182 30172 14188 30184
rect 13403 30144 14188 30172
rect 13403 30141 13415 30144
rect 13357 30135 13415 30141
rect 14182 30132 14188 30144
rect 14240 30132 14246 30184
rect 14461 30175 14519 30181
rect 14461 30141 14473 30175
rect 14507 30172 14519 30175
rect 14844 30172 14872 30212
rect 14507 30144 14872 30172
rect 14921 30175 14979 30181
rect 14507 30141 14519 30144
rect 14461 30135 14519 30141
rect 14921 30141 14933 30175
rect 14967 30172 14979 30175
rect 15010 30172 15016 30184
rect 14967 30144 15016 30172
rect 14967 30141 14979 30144
rect 14921 30135 14979 30141
rect 15010 30132 15016 30144
rect 15068 30132 15074 30184
rect 11149 30107 11207 30113
rect 10836 30076 11100 30104
rect 10836 30064 10842 30076
rect 6641 30039 6699 30045
rect 6641 30005 6653 30039
rect 6687 30036 6699 30039
rect 7466 30036 7472 30048
rect 6687 30008 7472 30036
rect 6687 30005 6699 30008
rect 6641 29999 6699 30005
rect 7466 29996 7472 30008
rect 7524 29996 7530 30048
rect 9674 30036 9680 30048
rect 9635 30008 9680 30036
rect 9674 29996 9680 30008
rect 9732 29996 9738 30048
rect 10318 30036 10324 30048
rect 10279 30008 10324 30036
rect 10318 29996 10324 30008
rect 10376 29996 10382 30048
rect 10689 30039 10747 30045
rect 10689 30005 10701 30039
rect 10735 30036 10747 30039
rect 10962 30036 10968 30048
rect 10735 30008 10968 30036
rect 10735 30005 10747 30008
rect 10689 29999 10747 30005
rect 10962 29996 10968 30008
rect 11020 29996 11026 30048
rect 11072 30036 11100 30076
rect 11149 30073 11161 30107
rect 11195 30104 11207 30107
rect 11330 30104 11336 30116
rect 11195 30076 11336 30104
rect 11195 30073 11207 30076
rect 11149 30067 11207 30073
rect 11330 30064 11336 30076
rect 11388 30064 11394 30116
rect 11517 30107 11575 30113
rect 11517 30073 11529 30107
rect 11563 30104 11575 30107
rect 11974 30104 11980 30116
rect 11563 30076 11980 30104
rect 11563 30073 11575 30076
rect 11517 30067 11575 30073
rect 11974 30064 11980 30076
rect 12032 30064 12038 30116
rect 13541 30107 13599 30113
rect 13541 30073 13553 30107
rect 13587 30104 13599 30107
rect 13722 30104 13728 30116
rect 13587 30076 13728 30104
rect 13587 30073 13599 30076
rect 13541 30067 13599 30073
rect 13722 30064 13728 30076
rect 13780 30064 13786 30116
rect 13906 30064 13912 30116
rect 13964 30104 13970 30116
rect 15120 30113 15148 30212
rect 15473 30209 15485 30243
rect 15519 30240 15531 30243
rect 16390 30240 16396 30252
rect 15519 30212 16396 30240
rect 15519 30209 15531 30212
rect 15473 30203 15531 30209
rect 16390 30200 16396 30212
rect 16448 30200 16454 30252
rect 17129 30243 17187 30249
rect 17129 30209 17141 30243
rect 17175 30240 17187 30243
rect 17770 30240 17776 30252
rect 17175 30212 17776 30240
rect 17175 30209 17187 30212
rect 17129 30203 17187 30209
rect 17770 30200 17776 30212
rect 17828 30200 17834 30252
rect 18046 30240 18052 30252
rect 17880 30212 18052 30240
rect 17497 30175 17555 30181
rect 17497 30141 17509 30175
rect 17543 30172 17555 30175
rect 17880 30172 17908 30212
rect 18046 30200 18052 30212
rect 18104 30200 18110 30252
rect 18248 30181 18276 30280
rect 19058 30268 19064 30280
rect 19116 30268 19122 30320
rect 20070 30268 20076 30320
rect 20128 30308 20134 30320
rect 20128 30280 20484 30308
rect 20128 30268 20134 30280
rect 19978 30240 19984 30252
rect 19939 30212 19984 30240
rect 19978 30200 19984 30212
rect 20036 30200 20042 30252
rect 20456 30184 20484 30280
rect 20714 30268 20720 30320
rect 20772 30268 20778 30320
rect 21266 30268 21272 30320
rect 21324 30268 21330 30320
rect 22002 30308 22008 30320
rect 21963 30280 22008 30308
rect 22002 30268 22008 30280
rect 22060 30268 22066 30320
rect 22112 30308 22140 30348
rect 22554 30336 22560 30388
rect 22612 30376 22618 30388
rect 23293 30379 23351 30385
rect 23293 30376 23305 30379
rect 22612 30348 23305 30376
rect 22612 30336 22618 30348
rect 23293 30345 23305 30348
rect 23339 30345 23351 30379
rect 23293 30339 23351 30345
rect 24121 30379 24179 30385
rect 24121 30345 24133 30379
rect 24167 30345 24179 30379
rect 24121 30339 24179 30345
rect 22281 30311 22339 30317
rect 22281 30308 22293 30311
rect 22112 30280 22293 30308
rect 22281 30277 22293 30280
rect 22327 30277 22339 30311
rect 22281 30271 22339 30277
rect 23842 30268 23848 30320
rect 23900 30308 23906 30320
rect 24136 30308 24164 30339
rect 25866 30336 25872 30388
rect 25924 30376 25930 30388
rect 27522 30376 27528 30388
rect 25924 30348 27528 30376
rect 25924 30336 25930 30348
rect 27522 30336 27528 30348
rect 27580 30336 27586 30388
rect 26602 30308 26608 30320
rect 23900 30280 24164 30308
rect 26563 30280 26608 30308
rect 23900 30268 23906 30280
rect 26602 30268 26608 30280
rect 26660 30268 26666 30320
rect 27614 30268 27620 30320
rect 27672 30308 27678 30320
rect 28721 30311 28779 30317
rect 28721 30308 28733 30311
rect 27672 30280 28733 30308
rect 27672 30268 27678 30280
rect 28721 30277 28733 30280
rect 28767 30277 28779 30311
rect 28721 30271 28779 30277
rect 22186 30200 22192 30252
rect 22244 30200 22250 30252
rect 23661 30243 23719 30249
rect 23661 30209 23673 30243
rect 23707 30240 23719 30243
rect 24762 30240 24768 30252
rect 23707 30212 24768 30240
rect 23707 30209 23719 30212
rect 23661 30203 23719 30209
rect 24762 30200 24768 30212
rect 24820 30200 24826 30252
rect 26620 30240 26648 30268
rect 26620 30212 26924 30240
rect 18233 30175 18291 30181
rect 18233 30172 18245 30175
rect 17543 30144 17908 30172
rect 17972 30144 18245 30172
rect 17543 30141 17555 30144
rect 17497 30135 17555 30141
rect 14553 30107 14611 30113
rect 14553 30104 14565 30107
rect 13964 30076 14565 30104
rect 13964 30064 13970 30076
rect 14553 30073 14565 30076
rect 14599 30104 14611 30107
rect 15105 30107 15163 30113
rect 14599 30076 15056 30104
rect 14599 30073 14611 30076
rect 14553 30067 14611 30073
rect 15028 30048 15056 30076
rect 15105 30073 15117 30107
rect 15151 30073 15163 30107
rect 15105 30067 15163 30073
rect 15286 30064 15292 30116
rect 15344 30104 15350 30116
rect 15654 30104 15660 30116
rect 15344 30076 15660 30104
rect 15344 30064 15350 30076
rect 15654 30064 15660 30076
rect 15712 30104 15718 30116
rect 16393 30107 16451 30113
rect 16393 30104 16405 30107
rect 15712 30076 16405 30104
rect 15712 30064 15718 30076
rect 16393 30073 16405 30076
rect 16439 30073 16451 30107
rect 16393 30067 16451 30073
rect 16761 30107 16819 30113
rect 16761 30073 16773 30107
rect 16807 30104 16819 30107
rect 17034 30104 17040 30116
rect 16807 30076 17040 30104
rect 16807 30073 16819 30076
rect 16761 30067 16819 30073
rect 17034 30064 17040 30076
rect 17092 30064 17098 30116
rect 17126 30064 17132 30116
rect 17184 30104 17190 30116
rect 17862 30104 17868 30116
rect 17184 30076 17868 30104
rect 17184 30064 17190 30076
rect 17862 30064 17868 30076
rect 17920 30104 17926 30116
rect 17972 30104 18000 30144
rect 18233 30141 18245 30144
rect 18279 30141 18291 30175
rect 18966 30172 18972 30184
rect 18233 30135 18291 30141
rect 18432 30144 18972 30172
rect 18432 30116 18460 30144
rect 18966 30132 18972 30144
rect 19024 30132 19030 30184
rect 19889 30175 19947 30181
rect 19889 30141 19901 30175
rect 19935 30172 19947 30175
rect 20070 30172 20076 30184
rect 19935 30144 20076 30172
rect 19935 30141 19947 30144
rect 19889 30135 19947 30141
rect 20070 30132 20076 30144
rect 20128 30132 20134 30184
rect 20165 30175 20223 30181
rect 20165 30141 20177 30175
rect 20211 30141 20223 30175
rect 20438 30172 20444 30184
rect 20351 30144 20444 30172
rect 20165 30135 20223 30141
rect 18414 30104 18420 30116
rect 17920 30076 18000 30104
rect 18327 30076 18420 30104
rect 17920 30064 17926 30076
rect 18414 30064 18420 30076
rect 18472 30064 18478 30116
rect 18782 30104 18788 30116
rect 18743 30076 18788 30104
rect 18782 30064 18788 30076
rect 18840 30064 18846 30116
rect 20180 30104 20208 30135
rect 20438 30132 20444 30144
rect 20496 30172 20502 30184
rect 20533 30175 20591 30181
rect 20533 30172 20545 30175
rect 20496 30144 20545 30172
rect 20496 30132 20502 30144
rect 20533 30141 20545 30144
rect 20579 30141 20591 30175
rect 21174 30172 21180 30184
rect 21135 30144 21180 30172
rect 20533 30135 20591 30141
rect 21174 30132 21180 30144
rect 21232 30132 21238 30184
rect 21637 30175 21695 30181
rect 21637 30141 21649 30175
rect 21683 30172 21695 30175
rect 21726 30172 21732 30184
rect 21683 30144 21732 30172
rect 21683 30141 21695 30144
rect 21637 30135 21695 30141
rect 19536 30076 20208 30104
rect 11238 30036 11244 30048
rect 11072 30008 11244 30036
rect 11238 29996 11244 30008
rect 11296 29996 11302 30048
rect 13078 29996 13084 30048
rect 13136 30036 13142 30048
rect 13354 30036 13360 30048
rect 13136 30008 13360 30036
rect 13136 29996 13142 30008
rect 13354 29996 13360 30008
rect 13412 29996 13418 30048
rect 13449 30039 13507 30045
rect 13449 30005 13461 30039
rect 13495 30036 13507 30039
rect 13814 30036 13820 30048
rect 13495 30008 13820 30036
rect 13495 30005 13507 30008
rect 13449 29999 13507 30005
rect 13814 29996 13820 30008
rect 13872 29996 13878 30048
rect 14461 30039 14519 30045
rect 14461 30005 14473 30039
rect 14507 30036 14519 30039
rect 14642 30036 14648 30048
rect 14507 30008 14648 30036
rect 14507 30005 14519 30008
rect 14461 29999 14519 30005
rect 14642 29996 14648 30008
rect 14700 29996 14706 30048
rect 15010 30036 15016 30048
rect 14923 30008 15016 30036
rect 15010 29996 15016 30008
rect 15068 29996 15074 30048
rect 15470 29996 15476 30048
rect 15528 30036 15534 30048
rect 15841 30039 15899 30045
rect 15841 30036 15853 30039
rect 15528 30008 15853 30036
rect 15528 29996 15534 30008
rect 15841 30005 15853 30008
rect 15887 30036 15899 30039
rect 16206 30036 16212 30048
rect 15887 30008 16212 30036
rect 15887 30005 15899 30008
rect 15841 29999 15899 30005
rect 16206 29996 16212 30008
rect 16264 30036 16270 30048
rect 16577 30039 16635 30045
rect 16577 30036 16589 30039
rect 16264 30008 16589 30036
rect 16264 29996 16270 30008
rect 16577 30005 16589 30008
rect 16623 30005 16635 30039
rect 16577 29999 16635 30005
rect 16666 29996 16672 30048
rect 16724 30036 16730 30048
rect 18322 30036 18328 30048
rect 16724 30008 16769 30036
rect 18235 30008 18328 30036
rect 16724 29996 16730 30008
rect 18322 29996 18328 30008
rect 18380 30036 18386 30048
rect 18874 30036 18880 30048
rect 18380 30008 18880 30036
rect 18380 29996 18386 30008
rect 18874 29996 18880 30008
rect 18932 29996 18938 30048
rect 19242 29996 19248 30048
rect 19300 30036 19306 30048
rect 19536 30045 19564 30076
rect 20714 30064 20720 30116
rect 20772 30104 20778 30116
rect 21652 30104 21680 30135
rect 21726 30132 21732 30144
rect 21784 30132 21790 30184
rect 22204 30172 22232 30200
rect 22465 30175 22523 30181
rect 22465 30172 22477 30175
rect 22204 30144 22477 30172
rect 22465 30141 22477 30144
rect 22511 30172 22523 30175
rect 23382 30172 23388 30184
rect 22511 30144 23388 30172
rect 22511 30141 22523 30144
rect 22465 30135 22523 30141
rect 23382 30132 23388 30144
rect 23440 30132 23446 30184
rect 23934 30172 23940 30184
rect 23895 30144 23940 30172
rect 23934 30132 23940 30144
rect 23992 30172 23998 30184
rect 23992 30144 24164 30172
rect 23992 30132 23998 30144
rect 20772 30076 21680 30104
rect 20772 30064 20778 30076
rect 22186 30064 22192 30116
rect 22244 30104 22250 30116
rect 22830 30104 22836 30116
rect 22244 30076 22836 30104
rect 22244 30064 22250 30076
rect 22830 30064 22836 30076
rect 22888 30104 22894 30116
rect 22925 30107 22983 30113
rect 22925 30104 22937 30107
rect 22888 30076 22937 30104
rect 22888 30064 22894 30076
rect 22925 30073 22937 30076
rect 22971 30073 22983 30107
rect 22925 30067 22983 30073
rect 23845 30107 23903 30113
rect 23845 30073 23857 30107
rect 23891 30104 23903 30107
rect 24026 30104 24032 30116
rect 23891 30076 24032 30104
rect 23891 30073 23903 30076
rect 23845 30067 23903 30073
rect 24026 30064 24032 30076
rect 24084 30064 24090 30116
rect 24136 30104 24164 30144
rect 24210 30132 24216 30184
rect 24268 30172 24274 30184
rect 25961 30175 26019 30181
rect 25961 30172 25973 30175
rect 24268 30144 25973 30172
rect 24268 30132 24274 30144
rect 25961 30141 25973 30144
rect 26007 30141 26019 30175
rect 25961 30135 26019 30141
rect 26602 30132 26608 30184
rect 26660 30172 26666 30184
rect 26896 30181 26924 30212
rect 26789 30175 26847 30181
rect 26789 30172 26801 30175
rect 26660 30144 26801 30172
rect 26660 30132 26666 30144
rect 26789 30141 26801 30144
rect 26835 30141 26847 30175
rect 26789 30135 26847 30141
rect 26881 30175 26939 30181
rect 26881 30141 26893 30175
rect 26927 30141 26939 30175
rect 26881 30135 26939 30141
rect 24486 30104 24492 30116
rect 24136 30076 24492 30104
rect 24486 30064 24492 30076
rect 24544 30064 24550 30116
rect 25225 30107 25283 30113
rect 25225 30073 25237 30107
rect 25271 30073 25283 30107
rect 25225 30067 25283 30073
rect 19521 30039 19579 30045
rect 19521 30036 19533 30039
rect 19300 30008 19533 30036
rect 19300 29996 19306 30008
rect 19521 30005 19533 30008
rect 19567 30005 19579 30039
rect 19521 29999 19579 30005
rect 20806 29996 20812 30048
rect 20864 30036 20870 30048
rect 22554 30036 22560 30048
rect 20864 30008 22560 30036
rect 20864 29996 20870 30008
rect 22554 29996 22560 30008
rect 22612 30036 22618 30048
rect 22649 30039 22707 30045
rect 22649 30036 22661 30039
rect 22612 30008 22661 30036
rect 22612 29996 22618 30008
rect 22649 30005 22661 30008
rect 22695 30005 22707 30039
rect 22649 29999 22707 30005
rect 23658 29996 23664 30048
rect 23716 30036 23722 30048
rect 24118 30036 24124 30048
rect 23716 30008 24124 30036
rect 23716 29996 23722 30008
rect 24118 29996 24124 30008
rect 24176 29996 24182 30048
rect 24670 30036 24676 30048
rect 24631 30008 24676 30036
rect 24670 29996 24676 30008
rect 24728 29996 24734 30048
rect 24946 29996 24952 30048
rect 25004 30036 25010 30048
rect 25041 30039 25099 30045
rect 25041 30036 25053 30039
rect 25004 30008 25053 30036
rect 25004 29996 25010 30008
rect 25041 30005 25053 30008
rect 25087 30036 25099 30039
rect 25240 30036 25268 30067
rect 25314 30064 25320 30116
rect 25372 30104 25378 30116
rect 25409 30107 25467 30113
rect 25409 30104 25421 30107
rect 25372 30076 25421 30104
rect 25372 30064 25378 30076
rect 25409 30073 25421 30076
rect 25455 30073 25467 30107
rect 25409 30067 25467 30073
rect 25593 30107 25651 30113
rect 25593 30073 25605 30107
rect 25639 30104 25651 30107
rect 25866 30104 25872 30116
rect 25639 30076 25872 30104
rect 25639 30073 25651 30076
rect 25593 30067 25651 30073
rect 25866 30064 25872 30076
rect 25924 30064 25930 30116
rect 25498 30036 25504 30048
rect 25087 30008 25268 30036
rect 25459 30008 25504 30036
rect 25087 30005 25099 30008
rect 25041 29999 25099 30005
rect 25498 29996 25504 30008
rect 25556 29996 25562 30048
rect 26234 30036 26240 30048
rect 26195 30008 26240 30036
rect 26234 29996 26240 30008
rect 26292 29996 26298 30048
rect 26804 30036 26832 30135
rect 27338 30104 27344 30116
rect 27299 30076 27344 30104
rect 27338 30064 27344 30076
rect 27396 30064 27402 30116
rect 28074 30104 28080 30116
rect 28035 30076 28080 30104
rect 28074 30064 28080 30076
rect 28132 30064 28138 30116
rect 27617 30039 27675 30045
rect 27617 30036 27629 30039
rect 26804 30008 27629 30036
rect 27617 30005 27629 30008
rect 27663 30005 27675 30039
rect 27617 29999 27675 30005
rect 28445 30039 28503 30045
rect 28445 30005 28457 30039
rect 28491 30036 28503 30039
rect 28718 30036 28724 30048
rect 28491 30008 28724 30036
rect 28491 30005 28503 30008
rect 28445 29999 28503 30005
rect 28718 29996 28724 30008
rect 28776 29996 28782 30048
rect 29454 30036 29460 30048
rect 29415 30008 29460 30036
rect 29454 29996 29460 30008
rect 29512 29996 29518 30048
rect 1104 29946 38824 29968
rect 1104 29894 19606 29946
rect 19658 29894 19670 29946
rect 19722 29894 19734 29946
rect 19786 29894 19798 29946
rect 19850 29894 38824 29946
rect 1104 29872 38824 29894
rect 1670 29832 1676 29844
rect 1412 29804 1676 29832
rect 1412 29705 1440 29804
rect 1670 29792 1676 29804
rect 1728 29792 1734 29844
rect 2866 29792 2872 29844
rect 2924 29832 2930 29844
rect 2961 29835 3019 29841
rect 2961 29832 2973 29835
rect 2924 29804 2973 29832
rect 2924 29792 2930 29804
rect 2961 29801 2973 29804
rect 3007 29801 3019 29835
rect 6730 29832 6736 29844
rect 6691 29804 6736 29832
rect 2961 29795 3019 29801
rect 6730 29792 6736 29804
rect 6788 29792 6794 29844
rect 9490 29832 9496 29844
rect 9451 29804 9496 29832
rect 9490 29792 9496 29804
rect 9548 29792 9554 29844
rect 10321 29835 10379 29841
rect 10321 29801 10333 29835
rect 10367 29832 10379 29835
rect 10870 29832 10876 29844
rect 10367 29804 10876 29832
rect 10367 29801 10379 29804
rect 10321 29795 10379 29801
rect 10870 29792 10876 29804
rect 10928 29792 10934 29844
rect 11054 29792 11060 29844
rect 11112 29792 11118 29844
rect 11238 29792 11244 29844
rect 11296 29832 11302 29844
rect 11425 29835 11483 29841
rect 11425 29832 11437 29835
rect 11296 29804 11437 29832
rect 11296 29792 11302 29804
rect 11425 29801 11437 29804
rect 11471 29801 11483 29835
rect 11425 29795 11483 29801
rect 11882 29792 11888 29844
rect 11940 29792 11946 29844
rect 12066 29792 12072 29844
rect 12124 29832 12130 29844
rect 13262 29832 13268 29844
rect 12124 29804 12204 29832
rect 13223 29804 13268 29832
rect 12124 29792 12130 29804
rect 8478 29764 8484 29776
rect 8439 29736 8484 29764
rect 8478 29724 8484 29736
rect 8536 29724 8542 29776
rect 11072 29764 11100 29792
rect 11900 29764 11928 29792
rect 12176 29773 12204 29804
rect 13262 29792 13268 29804
rect 13320 29792 13326 29844
rect 14826 29832 14832 29844
rect 14787 29804 14832 29832
rect 14826 29792 14832 29804
rect 14884 29792 14890 29844
rect 15470 29832 15476 29844
rect 15431 29804 15476 29832
rect 15470 29792 15476 29804
rect 15528 29792 15534 29844
rect 15654 29792 15660 29844
rect 15712 29832 15718 29844
rect 16025 29835 16083 29841
rect 16025 29832 16037 29835
rect 15712 29804 16037 29832
rect 15712 29792 15718 29804
rect 16025 29801 16037 29804
rect 16071 29801 16083 29835
rect 16025 29795 16083 29801
rect 16390 29792 16396 29844
rect 16448 29792 16454 29844
rect 16666 29792 16672 29844
rect 16724 29832 16730 29844
rect 17221 29835 17279 29841
rect 17221 29832 17233 29835
rect 16724 29804 17233 29832
rect 16724 29792 16730 29804
rect 17221 29801 17233 29804
rect 17267 29801 17279 29835
rect 17221 29795 17279 29801
rect 17681 29835 17739 29841
rect 17681 29801 17693 29835
rect 17727 29832 17739 29835
rect 17862 29832 17868 29844
rect 17727 29804 17868 29832
rect 17727 29801 17739 29804
rect 17681 29795 17739 29801
rect 17862 29792 17868 29804
rect 17920 29792 17926 29844
rect 17957 29835 18015 29841
rect 17957 29801 17969 29835
rect 18003 29832 18015 29835
rect 18690 29832 18696 29844
rect 18003 29804 18696 29832
rect 18003 29801 18015 29804
rect 17957 29795 18015 29801
rect 18690 29792 18696 29804
rect 18748 29792 18754 29844
rect 18969 29835 19027 29841
rect 18969 29801 18981 29835
rect 19015 29832 19027 29835
rect 20070 29832 20076 29844
rect 19015 29804 20076 29832
rect 19015 29801 19027 29804
rect 18969 29795 19027 29801
rect 20070 29792 20076 29804
rect 20128 29792 20134 29844
rect 20165 29835 20223 29841
rect 20165 29801 20177 29835
rect 20211 29832 20223 29835
rect 20349 29835 20407 29841
rect 20349 29832 20361 29835
rect 20211 29804 20361 29832
rect 20211 29801 20223 29804
rect 20165 29795 20223 29801
rect 20349 29801 20361 29804
rect 20395 29832 20407 29835
rect 20714 29832 20720 29844
rect 20395 29804 20720 29832
rect 20395 29801 20407 29804
rect 20349 29795 20407 29801
rect 20714 29792 20720 29804
rect 20772 29792 20778 29844
rect 20990 29792 20996 29844
rect 21048 29832 21054 29844
rect 21177 29835 21235 29841
rect 21177 29832 21189 29835
rect 21048 29804 21189 29832
rect 21048 29792 21054 29804
rect 21177 29801 21189 29804
rect 21223 29801 21235 29835
rect 21177 29795 21235 29801
rect 21634 29792 21640 29844
rect 21692 29832 21698 29844
rect 21821 29835 21879 29841
rect 21821 29832 21833 29835
rect 21692 29804 21833 29832
rect 21692 29792 21698 29804
rect 21821 29801 21833 29804
rect 21867 29832 21879 29835
rect 21913 29835 21971 29841
rect 21913 29832 21925 29835
rect 21867 29804 21925 29832
rect 21867 29801 21879 29804
rect 21821 29795 21879 29801
rect 21913 29801 21925 29804
rect 21959 29801 21971 29835
rect 22278 29832 22284 29844
rect 22239 29804 22284 29832
rect 21913 29795 21971 29801
rect 22278 29792 22284 29804
rect 22336 29792 22342 29844
rect 23569 29835 23627 29841
rect 23569 29801 23581 29835
rect 23615 29832 23627 29835
rect 23750 29832 23756 29844
rect 23615 29804 23756 29832
rect 23615 29801 23627 29804
rect 23569 29795 23627 29801
rect 23750 29792 23756 29804
rect 23808 29792 23814 29844
rect 23937 29835 23995 29841
rect 23937 29801 23949 29835
rect 23983 29832 23995 29835
rect 24302 29832 24308 29844
rect 23983 29804 24308 29832
rect 23983 29801 23995 29804
rect 23937 29795 23995 29801
rect 24302 29792 24308 29804
rect 24360 29792 24366 29844
rect 24854 29792 24860 29844
rect 24912 29832 24918 29844
rect 25593 29835 25651 29841
rect 25593 29832 25605 29835
rect 24912 29804 25605 29832
rect 24912 29792 24918 29804
rect 25593 29801 25605 29804
rect 25639 29801 25651 29835
rect 25593 29795 25651 29801
rect 25682 29792 25688 29844
rect 25740 29832 25746 29844
rect 25961 29835 26019 29841
rect 25961 29832 25973 29835
rect 25740 29804 25973 29832
rect 25740 29792 25746 29804
rect 25961 29801 25973 29804
rect 26007 29801 26019 29835
rect 26697 29835 26755 29841
rect 26697 29832 26709 29835
rect 25961 29795 26019 29801
rect 26160 29804 26709 29832
rect 12161 29767 12219 29773
rect 11072 29736 11192 29764
rect 11900 29736 12112 29764
rect 1397 29699 1455 29705
rect 1397 29665 1409 29699
rect 1443 29665 1455 29699
rect 1397 29659 1455 29665
rect 7101 29699 7159 29705
rect 7101 29665 7113 29699
rect 7147 29696 7159 29699
rect 7190 29696 7196 29708
rect 7147 29668 7196 29696
rect 7147 29665 7159 29668
rect 7101 29659 7159 29665
rect 7190 29656 7196 29668
rect 7248 29696 7254 29708
rect 8110 29696 8116 29708
rect 7248 29668 8116 29696
rect 7248 29656 7254 29668
rect 8110 29656 8116 29668
rect 8168 29656 8174 29708
rect 9122 29696 9128 29708
rect 9083 29668 9128 29696
rect 9122 29656 9128 29668
rect 9180 29656 9186 29708
rect 9766 29696 9772 29708
rect 9727 29668 9772 29696
rect 9766 29656 9772 29668
rect 9824 29656 9830 29708
rect 10781 29699 10839 29705
rect 10781 29665 10793 29699
rect 10827 29696 10839 29699
rect 11054 29696 11060 29708
rect 10827 29668 11060 29696
rect 10827 29665 10839 29668
rect 10781 29659 10839 29665
rect 11054 29656 11060 29668
rect 11112 29656 11118 29708
rect 11164 29696 11192 29736
rect 11238 29696 11244 29708
rect 11164 29668 11244 29696
rect 11238 29656 11244 29668
rect 11296 29656 11302 29708
rect 12084 29705 12112 29736
rect 12161 29733 12173 29767
rect 12207 29733 12219 29767
rect 12161 29727 12219 29733
rect 12529 29767 12587 29773
rect 12529 29733 12541 29767
rect 12575 29764 12587 29767
rect 12618 29764 12624 29776
rect 12575 29736 12624 29764
rect 12575 29733 12587 29736
rect 12529 29727 12587 29733
rect 12618 29724 12624 29736
rect 12676 29724 12682 29776
rect 15010 29724 15016 29776
rect 15068 29764 15074 29776
rect 16209 29767 16267 29773
rect 16209 29764 16221 29767
rect 15068 29736 16221 29764
rect 15068 29724 15074 29736
rect 16209 29733 16221 29736
rect 16255 29764 16267 29767
rect 16298 29764 16304 29776
rect 16255 29736 16304 29764
rect 16255 29733 16267 29736
rect 16209 29727 16267 29733
rect 16298 29724 16304 29736
rect 16356 29724 16362 29776
rect 16408 29764 16436 29792
rect 16574 29764 16580 29776
rect 16408 29736 16580 29764
rect 16574 29724 16580 29736
rect 16632 29724 16638 29776
rect 18141 29767 18199 29773
rect 18141 29733 18153 29767
rect 18187 29764 18199 29767
rect 18414 29764 18420 29776
rect 18187 29736 18420 29764
rect 18187 29733 18199 29736
rect 18141 29727 18199 29733
rect 18414 29724 18420 29736
rect 18472 29724 18478 29776
rect 19337 29767 19395 29773
rect 19337 29733 19349 29767
rect 19383 29764 19395 29767
rect 20438 29764 20444 29776
rect 19383 29736 20444 29764
rect 19383 29733 19395 29736
rect 19337 29727 19395 29733
rect 20438 29724 20444 29736
rect 20496 29724 20502 29776
rect 21269 29767 21327 29773
rect 21269 29733 21281 29767
rect 21315 29764 21327 29767
rect 21542 29764 21548 29776
rect 21315 29736 21548 29764
rect 21315 29733 21327 29736
rect 21269 29727 21327 29733
rect 21542 29724 21548 29736
rect 21600 29724 21606 29776
rect 23382 29764 23388 29776
rect 23032 29736 23388 29764
rect 11977 29699 12035 29705
rect 11977 29696 11989 29699
rect 11900 29668 11989 29696
rect 1670 29628 1676 29640
rect 1631 29600 1676 29628
rect 1670 29588 1676 29600
rect 1728 29588 1734 29640
rect 6638 29588 6644 29640
rect 6696 29628 6702 29640
rect 6825 29631 6883 29637
rect 6825 29628 6837 29631
rect 6696 29600 6837 29628
rect 6696 29588 6702 29600
rect 6825 29597 6837 29600
rect 6871 29597 6883 29631
rect 11698 29628 11704 29640
rect 6825 29591 6883 29597
rect 9968 29600 11704 29628
rect 9968 29569 9996 29600
rect 11698 29588 11704 29600
rect 11756 29588 11762 29640
rect 11793 29631 11851 29637
rect 11793 29597 11805 29631
rect 11839 29597 11851 29631
rect 11793 29591 11851 29597
rect 9953 29563 10011 29569
rect 9953 29529 9965 29563
rect 9999 29529 10011 29563
rect 10962 29560 10968 29572
rect 10923 29532 10968 29560
rect 9953 29523 10011 29529
rect 10962 29520 10968 29532
rect 11020 29520 11026 29572
rect 11333 29563 11391 29569
rect 11333 29529 11345 29563
rect 11379 29560 11391 29563
rect 11425 29563 11483 29569
rect 11425 29560 11437 29563
rect 11379 29532 11437 29560
rect 11379 29529 11391 29532
rect 11333 29523 11391 29529
rect 11425 29529 11437 29532
rect 11471 29560 11483 29563
rect 11808 29560 11836 29591
rect 11900 29572 11928 29668
rect 11977 29665 11989 29668
rect 12023 29665 12035 29699
rect 11977 29659 12035 29665
rect 12069 29699 12127 29705
rect 12069 29665 12081 29699
rect 12115 29665 12127 29699
rect 12069 29659 12127 29665
rect 13722 29656 13728 29708
rect 13780 29696 13786 29708
rect 14090 29696 14096 29708
rect 13780 29668 14096 29696
rect 13780 29656 13786 29668
rect 14090 29656 14096 29668
rect 14148 29696 14154 29708
rect 14185 29699 14243 29705
rect 14185 29696 14197 29699
rect 14148 29668 14197 29696
rect 14148 29656 14154 29668
rect 14185 29665 14197 29668
rect 14231 29665 14243 29699
rect 14185 29659 14243 29665
rect 15194 29656 15200 29708
rect 15252 29696 15258 29708
rect 16393 29699 16451 29705
rect 16393 29696 16405 29699
rect 15252 29668 16405 29696
rect 15252 29656 15258 29668
rect 16393 29665 16405 29668
rect 16439 29665 16451 29699
rect 16393 29659 16451 29665
rect 16485 29699 16543 29705
rect 16485 29665 16497 29699
rect 16531 29665 16543 29699
rect 18046 29696 18052 29708
rect 18007 29668 18052 29696
rect 16485 29659 16543 29665
rect 13354 29628 13360 29640
rect 13315 29600 13360 29628
rect 13354 29588 13360 29600
rect 13412 29588 13418 29640
rect 13909 29631 13967 29637
rect 13909 29597 13921 29631
rect 13955 29628 13967 29631
rect 13998 29628 14004 29640
rect 13955 29600 14004 29628
rect 13955 29597 13967 29600
rect 13909 29591 13967 29597
rect 13998 29588 14004 29600
rect 14056 29588 14062 29640
rect 14369 29631 14427 29637
rect 14369 29597 14381 29631
rect 14415 29597 14427 29631
rect 14369 29591 14427 29597
rect 11471 29532 11836 29560
rect 11471 29529 11483 29532
rect 11425 29523 11483 29529
rect 10689 29495 10747 29501
rect 10689 29461 10701 29495
rect 10735 29492 10747 29495
rect 10870 29492 10876 29504
rect 10735 29464 10876 29492
rect 10735 29461 10747 29464
rect 10689 29455 10747 29461
rect 10870 29452 10876 29464
rect 10928 29452 10934 29504
rect 11698 29492 11704 29504
rect 11659 29464 11704 29492
rect 11698 29452 11704 29464
rect 11756 29452 11762 29504
rect 11808 29492 11836 29532
rect 11882 29520 11888 29572
rect 11940 29520 11946 29572
rect 12894 29520 12900 29572
rect 12952 29560 12958 29572
rect 14090 29560 14096 29572
rect 12952 29532 14096 29560
rect 12952 29520 12958 29532
rect 14090 29520 14096 29532
rect 14148 29560 14154 29572
rect 14384 29560 14412 29591
rect 15654 29588 15660 29640
rect 15712 29628 15718 29640
rect 16500 29628 16528 29659
rect 18046 29656 18052 29668
rect 18104 29656 18110 29708
rect 19518 29696 19524 29708
rect 19479 29668 19524 29696
rect 19518 29656 19524 29668
rect 19576 29656 19582 29708
rect 21085 29699 21143 29705
rect 21085 29665 21097 29699
rect 21131 29696 21143 29699
rect 22002 29696 22008 29708
rect 21131 29668 22008 29696
rect 21131 29665 21143 29668
rect 21085 29659 21143 29665
rect 22002 29656 22008 29668
rect 22060 29656 22066 29708
rect 22094 29656 22100 29708
rect 22152 29696 22158 29708
rect 23032 29705 23060 29736
rect 23382 29724 23388 29736
rect 23440 29724 23446 29776
rect 23474 29724 23480 29776
rect 23532 29764 23538 29776
rect 24762 29764 24768 29776
rect 23532 29736 24348 29764
rect 24723 29736 24768 29764
rect 23532 29724 23538 29736
rect 23017 29699 23075 29705
rect 23017 29696 23029 29699
rect 22152 29668 23029 29696
rect 22152 29656 22158 29668
rect 23017 29665 23029 29668
rect 23063 29665 23075 29699
rect 23017 29659 23075 29665
rect 23106 29656 23112 29708
rect 23164 29696 23170 29708
rect 24320 29705 24348 29736
rect 24762 29724 24768 29736
rect 24820 29724 24826 29776
rect 25314 29764 25320 29776
rect 25275 29736 25320 29764
rect 25314 29724 25320 29736
rect 25372 29764 25378 29776
rect 26160 29764 26188 29804
rect 26697 29801 26709 29804
rect 26743 29801 26755 29835
rect 26697 29795 26755 29801
rect 27617 29835 27675 29841
rect 27617 29801 27629 29835
rect 27663 29832 27675 29835
rect 27706 29832 27712 29844
rect 27663 29804 27712 29832
rect 27663 29801 27675 29804
rect 27617 29795 27675 29801
rect 27706 29792 27712 29804
rect 27764 29792 27770 29844
rect 27890 29792 27896 29844
rect 27948 29832 27954 29844
rect 28261 29835 28319 29841
rect 28261 29832 28273 29835
rect 27948 29804 28273 29832
rect 27948 29792 27954 29804
rect 28261 29801 28273 29804
rect 28307 29801 28319 29835
rect 28261 29795 28319 29801
rect 25372 29736 26188 29764
rect 25372 29724 25378 29736
rect 26326 29724 26332 29776
rect 26384 29764 26390 29776
rect 26881 29767 26939 29773
rect 26384 29736 26832 29764
rect 26384 29724 26390 29736
rect 24029 29699 24087 29705
rect 24029 29696 24041 29699
rect 23164 29668 24041 29696
rect 23164 29656 23170 29668
rect 24029 29665 24041 29668
rect 24075 29665 24087 29699
rect 24029 29659 24087 29665
rect 24305 29699 24363 29705
rect 24305 29665 24317 29699
rect 24351 29665 24363 29699
rect 24305 29659 24363 29665
rect 25682 29656 25688 29708
rect 25740 29696 25746 29708
rect 25866 29696 25872 29708
rect 25740 29668 25872 29696
rect 25740 29656 25746 29668
rect 25866 29656 25872 29668
rect 25924 29656 25930 29708
rect 26510 29696 26516 29708
rect 26471 29668 26516 29696
rect 26510 29656 26516 29668
rect 26568 29656 26574 29708
rect 26804 29705 26832 29736
rect 26881 29733 26893 29767
rect 26927 29764 26939 29767
rect 26970 29764 26976 29776
rect 26927 29736 26976 29764
rect 26927 29733 26939 29736
rect 26881 29727 26939 29733
rect 26970 29724 26976 29736
rect 27028 29724 27034 29776
rect 27246 29764 27252 29776
rect 27207 29736 27252 29764
rect 27246 29724 27252 29736
rect 27304 29724 27310 29776
rect 26789 29699 26847 29705
rect 26789 29665 26801 29699
rect 26835 29696 26847 29699
rect 27890 29696 27896 29708
rect 26835 29668 27896 29696
rect 26835 29665 26847 29668
rect 26789 29659 26847 29665
rect 27890 29656 27896 29668
rect 27948 29656 27954 29708
rect 16942 29628 16948 29640
rect 15712 29600 16528 29628
rect 16903 29600 16948 29628
rect 15712 29588 15718 29600
rect 16942 29588 16948 29600
rect 17000 29588 17006 29640
rect 17770 29628 17776 29640
rect 17731 29600 17776 29628
rect 17770 29588 17776 29600
rect 17828 29588 17834 29640
rect 18509 29631 18567 29637
rect 18509 29597 18521 29631
rect 18555 29628 18567 29631
rect 19058 29628 19064 29640
rect 18555 29600 19064 29628
rect 18555 29597 18567 29600
rect 18509 29591 18567 29597
rect 19058 29588 19064 29600
rect 19116 29588 19122 29640
rect 19429 29631 19487 29637
rect 19429 29597 19441 29631
rect 19475 29628 19487 29631
rect 19702 29628 19708 29640
rect 19475 29600 19708 29628
rect 19475 29597 19487 29600
rect 19429 29591 19487 29597
rect 19702 29588 19708 29600
rect 19760 29588 19766 29640
rect 19981 29631 20039 29637
rect 19981 29597 19993 29631
rect 20027 29597 20039 29631
rect 19981 29591 20039 29597
rect 20901 29631 20959 29637
rect 20901 29597 20913 29631
rect 20947 29628 20959 29631
rect 21174 29628 21180 29640
rect 20947 29600 21180 29628
rect 20947 29597 20959 29600
rect 20901 29591 20959 29597
rect 14148 29532 14412 29560
rect 19996 29560 20024 29591
rect 21174 29588 21180 29600
rect 21232 29588 21238 29640
rect 21358 29588 21364 29640
rect 21416 29628 21422 29640
rect 21637 29631 21695 29637
rect 21637 29628 21649 29631
rect 21416 29600 21649 29628
rect 21416 29588 21422 29600
rect 21637 29597 21649 29600
rect 21683 29597 21695 29631
rect 21637 29591 21695 29597
rect 21726 29588 21732 29640
rect 21784 29628 21790 29640
rect 27614 29628 27620 29640
rect 21784 29600 27620 29628
rect 21784 29588 21790 29600
rect 27614 29588 27620 29600
rect 27672 29588 27678 29640
rect 20438 29560 20444 29572
rect 19996 29532 20444 29560
rect 14148 29520 14154 29532
rect 20438 29520 20444 29532
rect 20496 29560 20502 29572
rect 20496 29532 23060 29560
rect 20496 29520 20502 29532
rect 12434 29492 12440 29504
rect 11808 29464 12440 29492
rect 12434 29452 12440 29464
rect 12492 29452 12498 29504
rect 12802 29492 12808 29504
rect 12763 29464 12808 29492
rect 12802 29452 12808 29464
rect 12860 29452 12866 29504
rect 13262 29452 13268 29504
rect 13320 29492 13326 29504
rect 15746 29492 15752 29504
rect 13320 29464 15752 29492
rect 13320 29452 13326 29464
rect 15746 29452 15752 29464
rect 15804 29452 15810 29504
rect 18782 29452 18788 29504
rect 18840 29492 18846 29504
rect 20165 29495 20223 29501
rect 20165 29492 20177 29495
rect 18840 29464 20177 29492
rect 18840 29452 18846 29464
rect 20165 29461 20177 29464
rect 20211 29461 20223 29495
rect 20622 29492 20628 29504
rect 20583 29464 20628 29492
rect 20165 29455 20223 29461
rect 20622 29452 20628 29464
rect 20680 29452 20686 29504
rect 21174 29452 21180 29504
rect 21232 29492 21238 29504
rect 21542 29492 21548 29504
rect 21232 29464 21548 29492
rect 21232 29452 21238 29464
rect 21542 29452 21548 29464
rect 21600 29452 21606 29504
rect 21821 29495 21879 29501
rect 21821 29461 21833 29495
rect 21867 29492 21879 29495
rect 22462 29492 22468 29504
rect 21867 29464 22468 29492
rect 21867 29461 21879 29464
rect 21821 29455 21879 29461
rect 22462 29452 22468 29464
rect 22520 29452 22526 29504
rect 22922 29492 22928 29504
rect 22883 29464 22928 29492
rect 22922 29452 22928 29464
rect 22980 29452 22986 29504
rect 23032 29492 23060 29532
rect 23934 29520 23940 29572
rect 23992 29560 23998 29572
rect 24121 29563 24179 29569
rect 24121 29560 24133 29563
rect 23992 29532 24133 29560
rect 23992 29520 23998 29532
rect 24121 29529 24133 29532
rect 24167 29560 24179 29563
rect 26602 29560 26608 29572
rect 24167 29532 26608 29560
rect 24167 29529 24179 29532
rect 24121 29523 24179 29529
rect 26602 29520 26608 29532
rect 26660 29560 26666 29572
rect 27246 29560 27252 29572
rect 26660 29532 27252 29560
rect 26660 29520 26666 29532
rect 27246 29520 27252 29532
rect 27304 29520 27310 29572
rect 26326 29492 26332 29504
rect 23032 29464 26332 29492
rect 26326 29452 26332 29464
rect 26384 29452 26390 29504
rect 26970 29452 26976 29504
rect 27028 29492 27034 29504
rect 27893 29495 27951 29501
rect 27893 29492 27905 29495
rect 27028 29464 27905 29492
rect 27028 29452 27034 29464
rect 27893 29461 27905 29464
rect 27939 29492 27951 29495
rect 28258 29492 28264 29504
rect 27939 29464 28264 29492
rect 27939 29461 27951 29464
rect 27893 29455 27951 29461
rect 28258 29452 28264 29464
rect 28316 29452 28322 29504
rect 28718 29492 28724 29504
rect 28679 29464 28724 29492
rect 28718 29452 28724 29464
rect 28776 29452 28782 29504
rect 1104 29402 38824 29424
rect 1104 29350 4246 29402
rect 4298 29350 4310 29402
rect 4362 29350 4374 29402
rect 4426 29350 4438 29402
rect 4490 29350 34966 29402
rect 35018 29350 35030 29402
rect 35082 29350 35094 29402
rect 35146 29350 35158 29402
rect 35210 29350 38824 29402
rect 1104 29328 38824 29350
rect 1762 29248 1768 29300
rect 1820 29288 1826 29300
rect 1949 29291 2007 29297
rect 1949 29288 1961 29291
rect 1820 29260 1961 29288
rect 1820 29248 1826 29260
rect 1949 29257 1961 29260
rect 1995 29288 2007 29291
rect 2774 29288 2780 29300
rect 1995 29260 2780 29288
rect 1995 29257 2007 29260
rect 1949 29251 2007 29257
rect 2774 29248 2780 29260
rect 2832 29248 2838 29300
rect 6638 29288 6644 29300
rect 6599 29260 6644 29288
rect 6638 29248 6644 29260
rect 6696 29248 6702 29300
rect 7006 29248 7012 29300
rect 7064 29288 7070 29300
rect 7101 29291 7159 29297
rect 7101 29288 7113 29291
rect 7064 29260 7113 29288
rect 7064 29248 7070 29260
rect 7101 29257 7113 29260
rect 7147 29288 7159 29291
rect 7190 29288 7196 29300
rect 7147 29260 7196 29288
rect 7147 29257 7159 29260
rect 7101 29251 7159 29257
rect 7190 29248 7196 29260
rect 7248 29288 7254 29300
rect 8478 29288 8484 29300
rect 7248 29260 8248 29288
rect 7248 29248 7254 29260
rect 7282 29180 7288 29232
rect 7340 29180 7346 29232
rect 7300 29152 7328 29180
rect 7300 29124 7420 29152
rect 6638 29044 6644 29096
rect 6696 29084 6702 29096
rect 6914 29084 6920 29096
rect 6696 29056 6920 29084
rect 6696 29044 6702 29056
rect 6914 29044 6920 29056
rect 6972 29084 6978 29096
rect 7285 29087 7343 29093
rect 7285 29084 7297 29087
rect 6972 29056 7297 29084
rect 6972 29044 6978 29056
rect 7285 29053 7297 29056
rect 7331 29053 7343 29087
rect 7285 29047 7343 29053
rect 7392 29028 7420 29124
rect 7466 29112 7472 29164
rect 7524 29152 7530 29164
rect 7561 29155 7619 29161
rect 7561 29152 7573 29155
rect 7524 29124 7573 29152
rect 7524 29112 7530 29124
rect 7561 29121 7573 29124
rect 7607 29152 7619 29155
rect 7607 29124 7880 29152
rect 7607 29121 7619 29124
rect 7561 29115 7619 29121
rect 7852 29096 7880 29124
rect 7834 29044 7840 29096
rect 7892 29044 7898 29096
rect 8018 29044 8024 29096
rect 8076 29084 8082 29096
rect 8220 29084 8248 29260
rect 8404 29260 8484 29288
rect 8404 29084 8432 29260
rect 8478 29248 8484 29260
rect 8536 29248 8542 29300
rect 9214 29288 9220 29300
rect 8588 29260 9220 29288
rect 8588 29084 8616 29260
rect 9214 29248 9220 29260
rect 9272 29248 9278 29300
rect 9306 29248 9312 29300
rect 9364 29288 9370 29300
rect 9401 29291 9459 29297
rect 9401 29288 9413 29291
rect 9364 29260 9413 29288
rect 9364 29248 9370 29260
rect 9401 29257 9413 29260
rect 9447 29257 9459 29291
rect 9766 29288 9772 29300
rect 9727 29260 9772 29288
rect 9401 29251 9459 29257
rect 9766 29248 9772 29260
rect 9824 29248 9830 29300
rect 10226 29288 10232 29300
rect 10187 29260 10232 29288
rect 10226 29248 10232 29260
rect 10284 29248 10290 29300
rect 10502 29288 10508 29300
rect 10463 29260 10508 29288
rect 10502 29248 10508 29260
rect 10560 29248 10566 29300
rect 11882 29288 11888 29300
rect 11843 29260 11888 29288
rect 11882 29248 11888 29260
rect 11940 29248 11946 29300
rect 12250 29288 12256 29300
rect 12211 29260 12256 29288
rect 12250 29248 12256 29260
rect 12308 29248 12314 29300
rect 12434 29248 12440 29300
rect 12492 29288 12498 29300
rect 12713 29291 12771 29297
rect 12713 29288 12725 29291
rect 12492 29260 12725 29288
rect 12492 29248 12498 29260
rect 12713 29257 12725 29260
rect 12759 29288 12771 29291
rect 15286 29288 15292 29300
rect 12759 29260 15292 29288
rect 12759 29257 12771 29260
rect 12713 29251 12771 29257
rect 15286 29248 15292 29260
rect 15344 29248 15350 29300
rect 15470 29248 15476 29300
rect 15528 29288 15534 29300
rect 15565 29291 15623 29297
rect 15565 29288 15577 29291
rect 15528 29260 15577 29288
rect 15528 29248 15534 29260
rect 15565 29257 15577 29260
rect 15611 29257 15623 29291
rect 15565 29251 15623 29257
rect 15746 29248 15752 29300
rect 15804 29288 15810 29300
rect 16209 29291 16267 29297
rect 16209 29288 16221 29291
rect 15804 29260 16221 29288
rect 15804 29248 15810 29260
rect 16209 29257 16221 29260
rect 16255 29288 16267 29291
rect 16393 29291 16451 29297
rect 16393 29288 16405 29291
rect 16255 29260 16405 29288
rect 16255 29257 16267 29260
rect 16209 29251 16267 29257
rect 16393 29257 16405 29260
rect 16439 29288 16451 29291
rect 16666 29288 16672 29300
rect 16439 29260 16672 29288
rect 16439 29257 16451 29260
rect 16393 29251 16451 29257
rect 16666 29248 16672 29260
rect 16724 29248 16730 29300
rect 17034 29248 17040 29300
rect 17092 29288 17098 29300
rect 17092 29260 17264 29288
rect 17092 29248 17098 29260
rect 9582 29220 9588 29232
rect 8076 29056 8248 29084
rect 8312 29056 8432 29084
rect 8496 29056 8616 29084
rect 8680 29192 9588 29220
rect 8076 29044 8082 29056
rect 8312 29028 8340 29056
rect 8496 29028 8524 29056
rect 7374 28976 7380 29028
rect 7432 28976 7438 29028
rect 8294 28976 8300 29028
rect 8352 28976 8358 29028
rect 8478 28976 8484 29028
rect 8536 28976 8542 29028
rect 8570 28976 8576 29028
rect 8628 29016 8634 29028
rect 8680 29016 8708 29192
rect 9582 29180 9588 29192
rect 9640 29180 9646 29232
rect 11517 29223 11575 29229
rect 11517 29189 11529 29223
rect 11563 29220 11575 29223
rect 12158 29220 12164 29232
rect 11563 29192 12164 29220
rect 11563 29189 11575 29192
rect 11517 29183 11575 29189
rect 12158 29180 12164 29192
rect 12216 29180 12222 29232
rect 13265 29223 13323 29229
rect 13265 29189 13277 29223
rect 13311 29220 13323 29223
rect 13722 29220 13728 29232
rect 13311 29192 13728 29220
rect 13311 29189 13323 29192
rect 13265 29183 13323 29189
rect 13722 29180 13728 29192
rect 13780 29180 13786 29232
rect 14366 29220 14372 29232
rect 14108 29192 14372 29220
rect 8754 29112 8760 29164
rect 8812 29152 8818 29164
rect 8812 29124 9260 29152
rect 8812 29112 8818 29124
rect 9232 29096 9260 29124
rect 10594 29112 10600 29164
rect 10652 29152 10658 29164
rect 10652 29124 12848 29152
rect 10652 29112 10658 29124
rect 9214 29044 9220 29096
rect 9272 29044 9278 29096
rect 10318 29084 10324 29096
rect 10231 29056 10324 29084
rect 10318 29044 10324 29056
rect 10376 29084 10382 29096
rect 10870 29084 10876 29096
rect 10376 29056 10876 29084
rect 10376 29044 10382 29056
rect 10870 29044 10876 29056
rect 10928 29044 10934 29096
rect 11333 29087 11391 29093
rect 11333 29053 11345 29087
rect 11379 29084 11391 29087
rect 12250 29084 12256 29096
rect 11379 29056 12256 29084
rect 11379 29053 11391 29056
rect 11333 29047 11391 29053
rect 12250 29044 12256 29056
rect 12308 29044 12314 29096
rect 12820 29084 12848 29124
rect 13354 29112 13360 29164
rect 13412 29152 13418 29164
rect 13412 29124 14044 29152
rect 13412 29112 13418 29124
rect 13814 29084 13820 29096
rect 12820 29056 13676 29084
rect 13775 29056 13820 29084
rect 8628 28988 8708 29016
rect 8628 28976 8634 28988
rect 11054 28976 11060 29028
rect 11112 29016 11118 29028
rect 11241 29019 11299 29025
rect 11241 29016 11253 29019
rect 11112 28988 11253 29016
rect 11112 28976 11118 28988
rect 11241 28985 11253 28988
rect 11287 29016 11299 29019
rect 11287 28988 12480 29016
rect 11287 28985 11299 28988
rect 11241 28979 11299 28985
rect 12452 28960 12480 28988
rect 12986 28976 12992 29028
rect 13044 29016 13050 29028
rect 13357 29019 13415 29025
rect 13357 29016 13369 29019
rect 13044 28988 13369 29016
rect 13044 28976 13050 28988
rect 13357 28985 13369 28988
rect 13403 28985 13415 29019
rect 13648 29016 13676 29056
rect 13814 29044 13820 29056
rect 13872 29044 13878 29096
rect 14016 29093 14044 29124
rect 14108 29096 14136 29192
rect 14366 29180 14372 29192
rect 14424 29180 14430 29232
rect 14921 29223 14979 29229
rect 14921 29189 14933 29223
rect 14967 29220 14979 29223
rect 15654 29220 15660 29232
rect 14967 29192 15660 29220
rect 14967 29189 14979 29192
rect 14921 29183 14979 29189
rect 15654 29180 15660 29192
rect 15712 29180 15718 29232
rect 17126 29220 17132 29232
rect 16500 29192 17132 29220
rect 14182 29112 14188 29164
rect 14240 29152 14246 29164
rect 14277 29155 14335 29161
rect 14277 29152 14289 29155
rect 14240 29124 14289 29152
rect 14240 29112 14246 29124
rect 14277 29121 14289 29124
rect 14323 29152 14335 29155
rect 15010 29152 15016 29164
rect 14323 29124 15016 29152
rect 14323 29121 14335 29124
rect 14277 29115 14335 29121
rect 15010 29112 15016 29124
rect 15068 29112 15074 29164
rect 15746 29112 15752 29164
rect 15804 29152 15810 29164
rect 15930 29152 15936 29164
rect 15804 29124 15936 29152
rect 15804 29112 15810 29124
rect 15930 29112 15936 29124
rect 15988 29112 15994 29164
rect 14001 29087 14059 29093
rect 14001 29053 14013 29087
rect 14047 29053 14059 29087
rect 14001 29047 14059 29053
rect 14090 29044 14096 29096
rect 14148 29044 14154 29096
rect 14366 29084 14372 29096
rect 14327 29056 14372 29084
rect 14366 29044 14372 29056
rect 14424 29044 14430 29096
rect 15102 29044 15108 29096
rect 15160 29084 15166 29096
rect 15381 29087 15439 29093
rect 15381 29084 15393 29087
rect 15160 29056 15393 29084
rect 15160 29044 15166 29056
rect 15381 29053 15393 29056
rect 15427 29084 15439 29087
rect 15841 29087 15899 29093
rect 15841 29084 15853 29087
rect 15427 29056 15853 29084
rect 15427 29053 15439 29056
rect 15381 29047 15439 29053
rect 15841 29053 15853 29056
rect 15887 29084 15899 29087
rect 16500 29084 16528 29192
rect 17126 29180 17132 29192
rect 17184 29180 17190 29232
rect 17236 29220 17264 29260
rect 17402 29248 17408 29300
rect 17460 29288 17466 29300
rect 17497 29291 17555 29297
rect 17497 29288 17509 29291
rect 17460 29260 17509 29288
rect 17460 29248 17466 29260
rect 17497 29257 17509 29260
rect 17543 29288 17555 29291
rect 17770 29288 17776 29300
rect 17543 29260 17776 29288
rect 17543 29257 17555 29260
rect 17497 29251 17555 29257
rect 17770 29248 17776 29260
rect 17828 29248 17834 29300
rect 19150 29288 19156 29300
rect 18984 29260 19156 29288
rect 18984 29220 19012 29260
rect 19150 29248 19156 29260
rect 19208 29248 19214 29300
rect 19702 29288 19708 29300
rect 19663 29260 19708 29288
rect 19702 29248 19708 29260
rect 19760 29248 19766 29300
rect 19794 29248 19800 29300
rect 19852 29288 19858 29300
rect 20165 29291 20223 29297
rect 20165 29288 20177 29291
rect 19852 29260 20177 29288
rect 19852 29248 19858 29260
rect 20165 29257 20177 29260
rect 20211 29288 20223 29291
rect 20211 29260 20392 29288
rect 20211 29257 20223 29260
rect 20165 29251 20223 29257
rect 17236 29192 19012 29220
rect 16574 29112 16580 29164
rect 16632 29152 16638 29164
rect 17773 29155 17831 29161
rect 17773 29152 17785 29155
rect 16632 29124 17785 29152
rect 16632 29112 16638 29124
rect 17773 29121 17785 29124
rect 17819 29152 17831 29155
rect 18046 29152 18052 29164
rect 17819 29124 18052 29152
rect 17819 29121 17831 29124
rect 17773 29115 17831 29121
rect 18046 29112 18052 29124
rect 18104 29112 18110 29164
rect 16666 29084 16672 29096
rect 15887 29056 16528 29084
rect 16627 29056 16672 29084
rect 15887 29053 15899 29056
rect 15841 29047 15899 29053
rect 16666 29044 16672 29056
rect 16724 29044 16730 29096
rect 18782 29084 18788 29096
rect 18432 29056 18788 29084
rect 18432 29028 18460 29056
rect 18782 29044 18788 29056
rect 18840 29044 18846 29096
rect 13906 29016 13912 29028
rect 13648 28988 13912 29016
rect 13357 28979 13415 28985
rect 13906 28976 13912 28988
rect 13964 28976 13970 29028
rect 14182 28976 14188 29028
rect 14240 29016 14246 29028
rect 14642 29016 14648 29028
rect 14240 28988 14648 29016
rect 14240 28976 14246 28988
rect 14642 28976 14648 28988
rect 14700 28976 14706 29028
rect 15289 29019 15347 29025
rect 15289 28985 15301 29019
rect 15335 29016 15347 29019
rect 16206 29016 16212 29028
rect 15335 28988 16212 29016
rect 15335 28985 15347 28988
rect 15289 28979 15347 28985
rect 16206 28976 16212 28988
rect 16264 29016 16270 29028
rect 16577 29019 16635 29025
rect 16577 29016 16589 29019
rect 16264 28988 16589 29016
rect 16264 28976 16270 28988
rect 16577 28985 16589 28988
rect 16623 28985 16635 29019
rect 17126 29016 17132 29028
rect 17087 28988 17132 29016
rect 16577 28979 16635 28985
rect 1670 28948 1676 28960
rect 1631 28920 1676 28948
rect 1670 28908 1676 28920
rect 1728 28908 1734 28960
rect 7650 28908 7656 28960
rect 7708 28948 7714 28960
rect 8386 28948 8392 28960
rect 7708 28920 8392 28948
rect 7708 28908 7714 28920
rect 8386 28908 8392 28920
rect 8444 28908 8450 28960
rect 8662 28948 8668 28960
rect 8623 28920 8668 28948
rect 8662 28908 8668 28920
rect 8720 28908 8726 28960
rect 12434 28908 12440 28960
rect 12492 28948 12498 28960
rect 13538 28948 13544 28960
rect 12492 28920 13544 28948
rect 12492 28908 12498 28920
rect 13538 28908 13544 28920
rect 13596 28908 13602 28960
rect 13924 28948 13952 28976
rect 15930 28948 15936 28960
rect 13924 28920 15936 28948
rect 15930 28908 15936 28920
rect 15988 28908 15994 28960
rect 16592 28948 16620 28979
rect 17126 28976 17132 28988
rect 17184 28976 17190 29028
rect 18414 29016 18420 29028
rect 18375 28988 18420 29016
rect 18414 28976 18420 28988
rect 18472 28976 18478 29028
rect 18598 29016 18604 29028
rect 18559 28988 18604 29016
rect 18598 28976 18604 28988
rect 18656 28976 18662 29028
rect 18800 29016 18828 29044
rect 18984 29025 19012 29192
rect 19150 29112 19156 29164
rect 19208 29112 19214 29164
rect 20364 29161 20392 29260
rect 20898 29248 20904 29300
rect 20956 29288 20962 29300
rect 23106 29288 23112 29300
rect 20956 29260 21864 29288
rect 23067 29260 23112 29288
rect 20956 29248 20962 29260
rect 20990 29180 20996 29232
rect 21048 29220 21054 29232
rect 21361 29223 21419 29229
rect 21361 29220 21373 29223
rect 21048 29192 21373 29220
rect 21048 29180 21054 29192
rect 21361 29189 21373 29192
rect 21407 29220 21419 29223
rect 21542 29220 21548 29232
rect 21407 29192 21548 29220
rect 21407 29189 21419 29192
rect 21361 29183 21419 29189
rect 21542 29180 21548 29192
rect 21600 29180 21606 29232
rect 21836 29229 21864 29260
rect 23106 29248 23112 29260
rect 23164 29248 23170 29300
rect 23474 29288 23480 29300
rect 23435 29260 23480 29288
rect 23474 29248 23480 29260
rect 23532 29248 23538 29300
rect 23584 29260 24624 29288
rect 21821 29223 21879 29229
rect 21821 29189 21833 29223
rect 21867 29220 21879 29223
rect 23584 29220 23612 29260
rect 21867 29192 23612 29220
rect 21867 29189 21879 29192
rect 21821 29183 21879 29189
rect 20349 29155 20407 29161
rect 20349 29121 20361 29155
rect 20395 29121 20407 29155
rect 21910 29152 21916 29164
rect 21871 29124 21916 29152
rect 20349 29115 20407 29121
rect 21910 29112 21916 29124
rect 21968 29112 21974 29164
rect 19168 29084 19196 29112
rect 20533 29087 20591 29093
rect 19168 29056 20024 29084
rect 18969 29019 19027 29025
rect 18800 28988 18920 29016
rect 18046 28948 18052 28960
rect 16592 28920 18052 28948
rect 18046 28908 18052 28920
rect 18104 28908 18110 28960
rect 18690 28908 18696 28960
rect 18748 28948 18754 28960
rect 18892 28957 18920 28988
rect 18969 28985 18981 29019
rect 19015 28985 19027 29019
rect 18969 28979 19027 28985
rect 19150 28976 19156 29028
rect 19208 29016 19214 29028
rect 19337 29019 19395 29025
rect 19337 29016 19349 29019
rect 19208 28988 19349 29016
rect 19208 28976 19214 28988
rect 19337 28985 19349 28988
rect 19383 28985 19395 29019
rect 19996 29016 20024 29056
rect 20533 29053 20545 29087
rect 20579 29084 20591 29087
rect 20622 29084 20628 29096
rect 20579 29056 20628 29084
rect 20579 29053 20591 29056
rect 20533 29047 20591 29053
rect 20622 29044 20628 29056
rect 20680 29044 20686 29096
rect 20717 29019 20775 29025
rect 20717 29016 20729 29019
rect 19996 28988 20729 29016
rect 19337 28979 19395 28985
rect 20717 28985 20729 28988
rect 20763 28985 20775 29019
rect 21082 29016 21088 29028
rect 21043 28988 21088 29016
rect 20717 28979 20775 28985
rect 21082 28976 21088 28988
rect 21140 28976 21146 29028
rect 22112 29016 22140 29192
rect 22646 29112 22652 29164
rect 22704 29152 22710 29164
rect 23474 29152 23480 29164
rect 22704 29124 23480 29152
rect 22704 29112 22710 29124
rect 23474 29112 23480 29124
rect 23532 29112 23538 29164
rect 23842 29112 23848 29164
rect 23900 29152 23906 29164
rect 23937 29155 23995 29161
rect 23937 29152 23949 29155
rect 23900 29124 23949 29152
rect 23900 29112 23906 29124
rect 23937 29121 23949 29124
rect 23983 29121 23995 29155
rect 23937 29115 23995 29121
rect 22189 29087 22247 29093
rect 22189 29053 22201 29087
rect 22235 29084 22247 29087
rect 22462 29084 22468 29096
rect 22235 29056 22468 29084
rect 22235 29053 22247 29056
rect 22189 29047 22247 29053
rect 22462 29044 22468 29056
rect 22520 29044 22526 29096
rect 23661 29087 23719 29093
rect 23661 29053 23673 29087
rect 23707 29084 23719 29087
rect 23750 29084 23756 29096
rect 23707 29056 23756 29084
rect 23707 29053 23719 29056
rect 23661 29047 23719 29053
rect 23750 29044 23756 29056
rect 23808 29044 23814 29096
rect 24596 29084 24624 29260
rect 25314 29248 25320 29300
rect 25372 29288 25378 29300
rect 25593 29291 25651 29297
rect 25593 29288 25605 29291
rect 25372 29260 25605 29288
rect 25372 29248 25378 29260
rect 25593 29257 25605 29260
rect 25639 29288 25651 29291
rect 25866 29288 25872 29300
rect 25639 29260 25872 29288
rect 25639 29257 25651 29260
rect 25593 29251 25651 29257
rect 25866 29248 25872 29260
rect 25924 29248 25930 29300
rect 26053 29291 26111 29297
rect 26053 29257 26065 29291
rect 26099 29288 26111 29291
rect 26510 29288 26516 29300
rect 26099 29260 26516 29288
rect 26099 29257 26111 29260
rect 26053 29251 26111 29257
rect 26510 29248 26516 29260
rect 26568 29248 26574 29300
rect 27985 29291 28043 29297
rect 27985 29288 27997 29291
rect 27172 29260 27997 29288
rect 27062 29220 27068 29232
rect 26252 29192 27068 29220
rect 26252 29164 26280 29192
rect 27062 29180 27068 29192
rect 27120 29180 27126 29232
rect 26234 29152 26240 29164
rect 26147 29124 26240 29152
rect 26234 29112 26240 29124
rect 26292 29112 26298 29164
rect 27172 29161 27200 29260
rect 27985 29257 27997 29260
rect 28031 29288 28043 29291
rect 28350 29288 28356 29300
rect 28031 29260 28356 29288
rect 28031 29257 28043 29260
rect 27985 29251 28043 29257
rect 28350 29248 28356 29260
rect 28408 29248 28414 29300
rect 28718 29248 28724 29300
rect 28776 29288 28782 29300
rect 29457 29291 29515 29297
rect 29457 29288 29469 29291
rect 28776 29260 29469 29288
rect 28776 29248 28782 29260
rect 29457 29257 29469 29260
rect 29503 29257 29515 29291
rect 29457 29251 29515 29257
rect 27617 29223 27675 29229
rect 27617 29189 27629 29223
rect 27663 29220 27675 29223
rect 27890 29220 27896 29232
rect 27663 29192 27896 29220
rect 27663 29189 27675 29192
rect 27617 29183 27675 29189
rect 27890 29180 27896 29192
rect 27948 29180 27954 29232
rect 28166 29180 28172 29232
rect 28224 29220 28230 29232
rect 28261 29223 28319 29229
rect 28261 29220 28273 29223
rect 28224 29192 28273 29220
rect 28224 29180 28230 29192
rect 28261 29189 28273 29192
rect 28307 29189 28319 29223
rect 28261 29183 28319 29189
rect 27157 29155 27215 29161
rect 27157 29121 27169 29155
rect 27203 29121 27215 29155
rect 27157 29115 27215 29121
rect 26786 29084 26792 29096
rect 24596 29056 26792 29084
rect 26786 29044 26792 29056
rect 26844 29044 26850 29096
rect 27065 29087 27123 29093
rect 27065 29053 27077 29087
rect 27111 29053 27123 29087
rect 28074 29084 28080 29096
rect 27987 29056 28080 29084
rect 27065 29047 27123 29053
rect 22281 29019 22339 29025
rect 22281 29016 22293 29019
rect 22112 28988 22293 29016
rect 22281 28985 22293 28988
rect 22327 28985 22339 29019
rect 22646 29016 22652 29028
rect 22607 28988 22652 29016
rect 22281 28979 22339 28985
rect 22646 28976 22652 28988
rect 22704 28976 22710 29028
rect 25314 29016 25320 29028
rect 25275 28988 25320 29016
rect 25314 28976 25320 28988
rect 25372 28976 25378 29028
rect 26326 29016 26332 29028
rect 26287 28988 26332 29016
rect 26326 28976 26332 28988
rect 26384 28976 26390 29028
rect 27080 29016 27108 29047
rect 28074 29044 28080 29056
rect 28132 29084 28138 29096
rect 28537 29087 28595 29093
rect 28537 29084 28549 29087
rect 28132 29056 28549 29084
rect 28132 29044 28138 29056
rect 28537 29053 28549 29056
rect 28583 29053 28595 29087
rect 28537 29047 28595 29053
rect 27430 29016 27436 29028
rect 26436 28988 27436 29016
rect 18785 28951 18843 28957
rect 18785 28948 18797 28951
rect 18748 28920 18797 28948
rect 18748 28908 18754 28920
rect 18785 28917 18797 28920
rect 18831 28917 18843 28951
rect 18785 28911 18843 28917
rect 18877 28951 18935 28957
rect 18877 28917 18889 28951
rect 18923 28917 18935 28951
rect 18877 28911 18935 28917
rect 20438 28908 20444 28960
rect 20496 28948 20502 28960
rect 20625 28951 20683 28957
rect 20625 28948 20637 28951
rect 20496 28920 20637 28948
rect 20496 28908 20502 28920
rect 20625 28917 20637 28920
rect 20671 28917 20683 28951
rect 20625 28911 20683 28917
rect 22094 28908 22100 28960
rect 22152 28948 22158 28960
rect 22152 28920 22197 28948
rect 22152 28908 22158 28920
rect 26050 28908 26056 28960
rect 26108 28948 26114 28960
rect 26436 28948 26464 28988
rect 27430 28976 27436 28988
rect 27488 28976 27494 29028
rect 28718 28976 28724 29028
rect 28776 29016 28782 29028
rect 28994 29016 29000 29028
rect 28776 28988 29000 29016
rect 28776 28976 28782 28988
rect 28994 28976 29000 28988
rect 29052 28976 29058 29028
rect 26108 28920 26464 28948
rect 26108 28908 26114 28920
rect 1104 28858 38824 28880
rect 1104 28806 19606 28858
rect 19658 28806 19670 28858
rect 19722 28806 19734 28858
rect 19786 28806 19798 28858
rect 19850 28806 38824 28858
rect 1104 28784 38824 28806
rect 8018 28704 8024 28756
rect 8076 28744 8082 28756
rect 8478 28744 8484 28756
rect 8076 28716 8484 28744
rect 8076 28704 8082 28716
rect 8478 28704 8484 28716
rect 8536 28704 8542 28756
rect 8938 28704 8944 28756
rect 8996 28744 9002 28756
rect 9401 28747 9459 28753
rect 9401 28744 9413 28747
rect 8996 28716 9413 28744
rect 8996 28704 9002 28716
rect 9401 28713 9413 28716
rect 9447 28713 9459 28747
rect 10594 28744 10600 28756
rect 10555 28716 10600 28744
rect 9401 28707 9459 28713
rect 10594 28704 10600 28716
rect 10652 28704 10658 28756
rect 11790 28744 11796 28756
rect 11751 28716 11796 28744
rect 11790 28704 11796 28716
rect 11848 28704 11854 28756
rect 12342 28744 12348 28756
rect 12303 28716 12348 28744
rect 12342 28704 12348 28716
rect 12400 28704 12406 28756
rect 12894 28704 12900 28756
rect 12952 28744 12958 28756
rect 13446 28744 13452 28756
rect 12952 28716 13452 28744
rect 12952 28704 12958 28716
rect 7558 28676 7564 28688
rect 7519 28648 7564 28676
rect 7558 28636 7564 28648
rect 7616 28636 7622 28688
rect 9122 28676 9128 28688
rect 9083 28648 9128 28676
rect 9122 28636 9128 28648
rect 9180 28636 9186 28688
rect 12250 28636 12256 28688
rect 12308 28676 12314 28688
rect 12802 28676 12808 28688
rect 12308 28648 12808 28676
rect 12308 28636 12314 28648
rect 12802 28636 12808 28648
rect 12860 28636 12866 28688
rect 13280 28676 13308 28716
rect 13446 28704 13452 28716
rect 13504 28704 13510 28756
rect 13817 28747 13875 28753
rect 13817 28713 13829 28747
rect 13863 28744 13875 28747
rect 13998 28744 14004 28756
rect 13863 28716 14004 28744
rect 13863 28713 13875 28716
rect 13817 28707 13875 28713
rect 13998 28704 14004 28716
rect 14056 28704 14062 28756
rect 14737 28747 14795 28753
rect 14737 28713 14749 28747
rect 14783 28744 14795 28747
rect 15102 28744 15108 28756
rect 14783 28716 15108 28744
rect 14783 28713 14795 28716
rect 14737 28707 14795 28713
rect 15102 28704 15108 28716
rect 15160 28704 15166 28756
rect 16298 28704 16304 28756
rect 16356 28744 16362 28756
rect 16945 28747 17003 28753
rect 16945 28744 16957 28747
rect 16356 28716 16957 28744
rect 16356 28704 16362 28716
rect 16945 28713 16957 28716
rect 16991 28713 17003 28747
rect 16945 28707 17003 28713
rect 18601 28747 18659 28753
rect 18601 28713 18613 28747
rect 18647 28744 18659 28747
rect 18690 28744 18696 28756
rect 18647 28716 18696 28744
rect 18647 28713 18659 28716
rect 18601 28707 18659 28713
rect 18690 28704 18696 28716
rect 18748 28704 18754 28756
rect 18874 28704 18880 28756
rect 18932 28744 18938 28756
rect 20349 28747 20407 28753
rect 18932 28716 20024 28744
rect 18932 28704 18938 28716
rect 19996 28688 20024 28716
rect 20349 28713 20361 28747
rect 20395 28744 20407 28747
rect 20438 28744 20444 28756
rect 20395 28716 20444 28744
rect 20395 28713 20407 28716
rect 20349 28707 20407 28713
rect 20438 28704 20444 28716
rect 20496 28704 20502 28756
rect 21174 28744 21180 28756
rect 20548 28716 21180 28744
rect 14366 28676 14372 28688
rect 13280 28648 14372 28676
rect 8018 28568 8024 28620
rect 8076 28608 8082 28620
rect 8205 28611 8263 28617
rect 8205 28608 8217 28611
rect 8076 28580 8217 28608
rect 8076 28568 8082 28580
rect 8205 28577 8217 28580
rect 8251 28577 8263 28611
rect 8205 28571 8263 28577
rect 8573 28611 8631 28617
rect 8573 28577 8585 28611
rect 8619 28608 8631 28611
rect 8662 28608 8668 28620
rect 8619 28580 8668 28608
rect 8619 28577 8631 28580
rect 8573 28571 8631 28577
rect 8662 28568 8668 28580
rect 8720 28568 8726 28620
rect 8757 28611 8815 28617
rect 8757 28577 8769 28611
rect 8803 28608 8815 28611
rect 8938 28608 8944 28620
rect 8803 28580 8944 28608
rect 8803 28577 8815 28580
rect 8757 28571 8815 28577
rect 8938 28568 8944 28580
rect 8996 28568 9002 28620
rect 9766 28568 9772 28620
rect 9824 28608 9830 28620
rect 10778 28608 10784 28620
rect 9824 28580 10784 28608
rect 9824 28568 9830 28580
rect 10778 28568 10784 28580
rect 10836 28568 10842 28620
rect 12897 28611 12955 28617
rect 12897 28577 12909 28611
rect 12943 28608 12955 28611
rect 12986 28608 12992 28620
rect 12943 28580 12992 28608
rect 12943 28577 12955 28580
rect 12897 28571 12955 28577
rect 12986 28568 12992 28580
rect 13044 28568 13050 28620
rect 13280 28617 13308 28648
rect 14366 28636 14372 28648
rect 14424 28636 14430 28688
rect 18785 28679 18843 28685
rect 18785 28645 18797 28679
rect 18831 28676 18843 28679
rect 18966 28676 18972 28688
rect 18831 28648 18972 28676
rect 18831 28645 18843 28648
rect 18785 28639 18843 28645
rect 18966 28636 18972 28648
rect 19024 28636 19030 28688
rect 19978 28676 19984 28688
rect 19891 28648 19984 28676
rect 19978 28636 19984 28648
rect 20036 28676 20042 28688
rect 20548 28676 20576 28716
rect 21174 28704 21180 28716
rect 21232 28704 21238 28756
rect 21910 28744 21916 28756
rect 21871 28716 21916 28744
rect 21910 28704 21916 28716
rect 21968 28704 21974 28756
rect 22462 28704 22468 28756
rect 22520 28744 22526 28756
rect 22649 28747 22707 28753
rect 22649 28744 22661 28747
rect 22520 28716 22661 28744
rect 22520 28704 22526 28716
rect 22649 28713 22661 28716
rect 22695 28713 22707 28747
rect 22649 28707 22707 28713
rect 23106 28704 23112 28756
rect 23164 28704 23170 28756
rect 23569 28747 23627 28753
rect 23569 28713 23581 28747
rect 23615 28744 23627 28747
rect 23658 28744 23664 28756
rect 23615 28716 23664 28744
rect 23615 28713 23627 28716
rect 23569 28707 23627 28713
rect 23658 28704 23664 28716
rect 23716 28704 23722 28756
rect 23934 28744 23940 28756
rect 23895 28716 23940 28744
rect 23934 28704 23940 28716
rect 23992 28704 23998 28756
rect 24854 28704 24860 28756
rect 24912 28744 24918 28756
rect 25133 28747 25191 28753
rect 25133 28744 25145 28747
rect 24912 28716 25145 28744
rect 24912 28704 24918 28716
rect 25133 28713 25145 28716
rect 25179 28744 25191 28747
rect 25590 28744 25596 28756
rect 25179 28716 25596 28744
rect 25179 28713 25191 28716
rect 25133 28707 25191 28713
rect 25590 28704 25596 28716
rect 25648 28704 25654 28756
rect 25869 28747 25927 28753
rect 25869 28713 25881 28747
rect 25915 28744 25927 28747
rect 26050 28744 26056 28756
rect 25915 28716 26056 28744
rect 25915 28713 25927 28716
rect 25869 28707 25927 28713
rect 26050 28704 26056 28716
rect 26108 28704 26114 28756
rect 26234 28744 26240 28756
rect 26195 28716 26240 28744
rect 26234 28704 26240 28716
rect 26292 28704 26298 28756
rect 27338 28744 27344 28756
rect 26344 28716 27344 28744
rect 20714 28676 20720 28688
rect 20036 28648 20576 28676
rect 20627 28648 20720 28676
rect 20036 28636 20042 28648
rect 20714 28636 20720 28648
rect 20772 28676 20778 28688
rect 20898 28676 20904 28688
rect 20772 28648 20904 28676
rect 20772 28636 20778 28648
rect 20898 28636 20904 28648
rect 20956 28676 20962 28688
rect 21085 28679 21143 28685
rect 21085 28676 21097 28679
rect 20956 28648 21097 28676
rect 20956 28636 20962 28648
rect 21085 28645 21097 28648
rect 21131 28645 21143 28679
rect 21085 28639 21143 28645
rect 21269 28679 21327 28685
rect 21269 28645 21281 28679
rect 21315 28676 21327 28679
rect 21450 28676 21456 28688
rect 21315 28648 21456 28676
rect 21315 28645 21327 28648
rect 21269 28639 21327 28645
rect 21450 28636 21456 28648
rect 21508 28636 21514 28688
rect 21729 28679 21787 28685
rect 21729 28645 21741 28679
rect 21775 28676 21787 28679
rect 22094 28676 22100 28688
rect 21775 28648 22100 28676
rect 21775 28645 21787 28648
rect 21729 28639 21787 28645
rect 22094 28636 22100 28648
rect 22152 28636 22158 28688
rect 22833 28679 22891 28685
rect 22572 28648 22784 28676
rect 13265 28611 13323 28617
rect 13265 28577 13277 28611
rect 13311 28577 13323 28611
rect 13265 28571 13323 28577
rect 14458 28568 14464 28620
rect 14516 28608 14522 28620
rect 15194 28608 15200 28620
rect 14516 28580 15200 28608
rect 14516 28568 14522 28580
rect 15194 28568 15200 28580
rect 15252 28568 15258 28620
rect 16117 28611 16175 28617
rect 16117 28577 16129 28611
rect 16163 28608 16175 28611
rect 16758 28608 16764 28620
rect 16163 28580 16764 28608
rect 16163 28577 16175 28580
rect 16117 28571 16175 28577
rect 16758 28568 16764 28580
rect 16816 28568 16822 28620
rect 17405 28611 17463 28617
rect 17405 28577 17417 28611
rect 17451 28608 17463 28611
rect 17770 28608 17776 28620
rect 17451 28580 17776 28608
rect 17451 28577 17463 28580
rect 17405 28571 17463 28577
rect 17770 28568 17776 28580
rect 17828 28568 17834 28620
rect 18322 28568 18328 28620
rect 18380 28608 18386 28620
rect 18693 28611 18751 28617
rect 18693 28608 18705 28611
rect 18380 28580 18705 28608
rect 18380 28568 18386 28580
rect 18693 28577 18705 28580
rect 18739 28608 18751 28611
rect 18874 28608 18880 28620
rect 18739 28580 18880 28608
rect 18739 28577 18751 28580
rect 18693 28571 18751 28577
rect 18874 28568 18880 28580
rect 18932 28568 18938 28620
rect 21174 28568 21180 28620
rect 21232 28608 21238 28620
rect 22572 28608 22600 28648
rect 22756 28617 22784 28648
rect 22833 28645 22845 28679
rect 22879 28676 22891 28679
rect 23124 28676 23152 28704
rect 22879 28648 23152 28676
rect 22879 28645 22891 28648
rect 22833 28639 22891 28645
rect 23382 28636 23388 28688
rect 23440 28676 23446 28688
rect 26344 28676 26372 28716
rect 27338 28704 27344 28716
rect 27396 28704 27402 28756
rect 27617 28747 27675 28753
rect 27617 28713 27629 28747
rect 27663 28744 27675 28747
rect 27706 28744 27712 28756
rect 27663 28716 27712 28744
rect 27663 28713 27675 28716
rect 27617 28707 27675 28713
rect 27706 28704 27712 28716
rect 27764 28704 27770 28756
rect 27985 28747 28043 28753
rect 27985 28713 27997 28747
rect 28031 28744 28043 28747
rect 28902 28744 28908 28756
rect 28031 28716 28908 28744
rect 28031 28713 28043 28716
rect 27985 28707 28043 28713
rect 28902 28704 28908 28716
rect 28960 28704 28966 28756
rect 28994 28704 29000 28756
rect 29052 28744 29058 28756
rect 29052 28716 29097 28744
rect 29052 28704 29058 28716
rect 23440 28648 26372 28676
rect 26513 28679 26571 28685
rect 23440 28636 23446 28648
rect 26513 28645 26525 28679
rect 26559 28676 26571 28679
rect 26602 28676 26608 28688
rect 26559 28648 26608 28676
rect 26559 28645 26571 28648
rect 26513 28639 26571 28645
rect 26602 28636 26608 28648
rect 26660 28676 26666 28688
rect 26786 28676 26792 28688
rect 26660 28648 26792 28676
rect 26660 28636 26666 28648
rect 26786 28636 26792 28648
rect 26844 28636 26850 28688
rect 21232 28580 22600 28608
rect 22741 28611 22799 28617
rect 21232 28568 21238 28580
rect 22741 28577 22753 28611
rect 22787 28608 22799 28611
rect 23106 28608 23112 28620
rect 22787 28580 23112 28608
rect 22787 28577 22799 28580
rect 22741 28571 22799 28577
rect 23106 28568 23112 28580
rect 23164 28568 23170 28620
rect 24210 28608 24216 28620
rect 24171 28580 24216 28608
rect 24210 28568 24216 28580
rect 24268 28568 24274 28620
rect 28077 28611 28135 28617
rect 28077 28577 28089 28611
rect 28123 28608 28135 28611
rect 28166 28608 28172 28620
rect 28123 28580 28172 28608
rect 28123 28577 28135 28580
rect 28077 28571 28135 28577
rect 28166 28568 28172 28580
rect 28224 28568 28230 28620
rect 32030 28568 32036 28620
rect 32088 28608 32094 28620
rect 32490 28608 32496 28620
rect 32088 28580 32496 28608
rect 32088 28568 32094 28580
rect 32490 28568 32496 28580
rect 32548 28608 32554 28620
rect 32677 28611 32735 28617
rect 32677 28608 32689 28611
rect 32548 28580 32689 28608
rect 32548 28568 32554 28580
rect 32677 28577 32689 28580
rect 32723 28577 32735 28611
rect 32677 28571 32735 28577
rect 7834 28500 7840 28552
rect 7892 28540 7898 28552
rect 8297 28543 8355 28549
rect 8297 28540 8309 28543
rect 7892 28512 8309 28540
rect 7892 28500 7898 28512
rect 8297 28509 8309 28512
rect 8343 28540 8355 28543
rect 8386 28540 8392 28552
rect 8343 28512 8392 28540
rect 8343 28509 8355 28512
rect 8297 28503 8355 28509
rect 8386 28500 8392 28512
rect 8444 28500 8450 28552
rect 12802 28540 12808 28552
rect 12763 28512 12808 28540
rect 12802 28500 12808 28512
rect 12860 28500 12866 28552
rect 13173 28543 13231 28549
rect 13173 28509 13185 28543
rect 13219 28540 13231 28543
rect 13446 28540 13452 28552
rect 13219 28512 13452 28540
rect 13219 28509 13231 28512
rect 13173 28503 13231 28509
rect 13446 28500 13452 28512
rect 13504 28500 13510 28552
rect 14642 28500 14648 28552
rect 14700 28540 14706 28552
rect 15289 28543 15347 28549
rect 15289 28540 15301 28543
rect 14700 28512 15301 28540
rect 14700 28500 14706 28512
rect 15289 28509 15301 28512
rect 15335 28509 15347 28543
rect 15289 28503 15347 28509
rect 15841 28543 15899 28549
rect 15841 28509 15853 28543
rect 15887 28509 15899 28543
rect 15841 28503 15899 28509
rect 10229 28475 10287 28481
rect 10229 28441 10241 28475
rect 10275 28472 10287 28475
rect 13722 28472 13728 28484
rect 10275 28444 13728 28472
rect 10275 28441 10287 28444
rect 10229 28435 10287 28441
rect 13722 28432 13728 28444
rect 13780 28432 13786 28484
rect 13998 28432 14004 28484
rect 14056 28472 14062 28484
rect 15856 28472 15884 28503
rect 15930 28500 15936 28552
rect 15988 28540 15994 28552
rect 16301 28543 16359 28549
rect 16301 28540 16313 28543
rect 15988 28512 16313 28540
rect 15988 28500 15994 28512
rect 16301 28509 16313 28512
rect 16347 28509 16359 28543
rect 16301 28503 16359 28509
rect 18417 28543 18475 28549
rect 18417 28509 18429 28543
rect 18463 28540 18475 28543
rect 18598 28540 18604 28552
rect 18463 28512 18604 28540
rect 18463 28509 18475 28512
rect 18417 28503 18475 28509
rect 18598 28500 18604 28512
rect 18656 28500 18662 28552
rect 18966 28500 18972 28552
rect 19024 28540 19030 28552
rect 19153 28543 19211 28549
rect 19153 28540 19165 28543
rect 19024 28512 19165 28540
rect 19024 28500 19030 28512
rect 19153 28509 19165 28512
rect 19199 28509 19211 28543
rect 19153 28503 19211 28509
rect 19334 28500 19340 28552
rect 19392 28540 19398 28552
rect 19392 28512 20208 28540
rect 19392 28500 19398 28512
rect 14056 28444 15884 28472
rect 18325 28475 18383 28481
rect 14056 28432 14062 28444
rect 18325 28441 18337 28475
rect 18371 28472 18383 28475
rect 19794 28472 19800 28484
rect 18371 28444 19800 28472
rect 18371 28441 18383 28444
rect 18325 28435 18383 28441
rect 19794 28432 19800 28444
rect 19852 28432 19858 28484
rect 20180 28472 20208 28512
rect 20438 28500 20444 28552
rect 20496 28540 20502 28552
rect 20901 28543 20959 28549
rect 20901 28540 20913 28543
rect 20496 28512 20913 28540
rect 20496 28500 20502 28512
rect 20901 28509 20913 28512
rect 20947 28540 20959 28543
rect 21266 28540 21272 28552
rect 20947 28512 21272 28540
rect 20947 28509 20959 28512
rect 20901 28503 20959 28509
rect 21266 28500 21272 28512
rect 21324 28500 21330 28552
rect 21634 28540 21640 28552
rect 21595 28512 21640 28540
rect 21634 28500 21640 28512
rect 21692 28500 21698 28552
rect 21910 28500 21916 28552
rect 21968 28540 21974 28552
rect 22465 28543 22523 28549
rect 22465 28540 22477 28543
rect 21968 28512 22477 28540
rect 21968 28500 21974 28512
rect 22465 28509 22477 28512
rect 22511 28509 22523 28543
rect 22465 28503 22523 28509
rect 22554 28500 22560 28552
rect 22612 28540 22618 28552
rect 23201 28543 23259 28549
rect 23201 28540 23213 28543
rect 22612 28512 23213 28540
rect 22612 28500 22618 28512
rect 23201 28509 23213 28512
rect 23247 28509 23259 28543
rect 23201 28503 23259 28509
rect 26786 28500 26792 28552
rect 26844 28540 26850 28552
rect 26881 28543 26939 28549
rect 26881 28540 26893 28543
rect 26844 28512 26893 28540
rect 26844 28500 26850 28512
rect 26881 28509 26893 28512
rect 26927 28509 26939 28543
rect 26881 28503 26939 28509
rect 32401 28543 32459 28549
rect 32401 28509 32413 28543
rect 32447 28540 32459 28543
rect 32766 28540 32772 28552
rect 32447 28512 32772 28540
rect 32447 28509 32459 28512
rect 32401 28503 32459 28509
rect 32766 28500 32772 28512
rect 32824 28500 32830 28552
rect 21729 28475 21787 28481
rect 21729 28472 21741 28475
rect 20180 28444 21741 28472
rect 21729 28441 21741 28444
rect 21775 28441 21787 28475
rect 21729 28435 21787 28441
rect 22002 28432 22008 28484
rect 22060 28472 22066 28484
rect 22281 28475 22339 28481
rect 22281 28472 22293 28475
rect 22060 28444 22293 28472
rect 22060 28432 22066 28444
rect 22281 28441 22293 28444
rect 22327 28441 22339 28475
rect 22281 28435 22339 28441
rect 26510 28432 26516 28484
rect 26568 28472 26574 28484
rect 26678 28475 26736 28481
rect 26678 28472 26690 28475
rect 26568 28444 26690 28472
rect 26568 28432 26574 28444
rect 26678 28441 26690 28444
rect 26724 28472 26736 28475
rect 27338 28472 27344 28484
rect 26724 28444 27344 28472
rect 26724 28441 26736 28444
rect 26678 28435 26736 28441
rect 27338 28432 27344 28444
rect 27396 28432 27402 28484
rect 27614 28432 27620 28484
rect 27672 28472 27678 28484
rect 28261 28475 28319 28481
rect 28261 28472 28273 28475
rect 27672 28444 28273 28472
rect 27672 28432 27678 28444
rect 28261 28441 28273 28444
rect 28307 28441 28319 28475
rect 28261 28435 28319 28441
rect 6914 28404 6920 28416
rect 6875 28376 6920 28404
rect 6914 28364 6920 28376
rect 6972 28364 6978 28416
rect 7282 28404 7288 28416
rect 7243 28376 7288 28404
rect 7282 28364 7288 28376
rect 7340 28364 7346 28416
rect 11054 28364 11060 28416
rect 11112 28404 11118 28416
rect 11149 28407 11207 28413
rect 11149 28404 11161 28407
rect 11112 28376 11161 28404
rect 11112 28364 11118 28376
rect 11149 28373 11161 28376
rect 11195 28373 11207 28407
rect 11149 28367 11207 28373
rect 13906 28364 13912 28416
rect 13964 28404 13970 28416
rect 14277 28407 14335 28413
rect 14277 28404 14289 28407
rect 13964 28376 14289 28404
rect 13964 28364 13970 28376
rect 14277 28373 14289 28376
rect 14323 28373 14335 28407
rect 14277 28367 14335 28373
rect 15105 28407 15163 28413
rect 15105 28373 15117 28407
rect 15151 28404 15163 28407
rect 15470 28404 15476 28416
rect 15151 28376 15476 28404
rect 15151 28373 15163 28376
rect 15105 28367 15163 28373
rect 15470 28364 15476 28376
rect 15528 28364 15534 28416
rect 16666 28404 16672 28416
rect 16627 28376 16672 28404
rect 16666 28364 16672 28376
rect 16724 28364 16730 28416
rect 17586 28404 17592 28416
rect 17547 28376 17592 28404
rect 17586 28364 17592 28376
rect 17644 28364 17650 28416
rect 17954 28404 17960 28416
rect 17915 28376 17960 28404
rect 17954 28364 17960 28376
rect 18012 28364 18018 28416
rect 18598 28364 18604 28416
rect 18656 28404 18662 28416
rect 19429 28407 19487 28413
rect 19429 28404 19441 28407
rect 18656 28376 19441 28404
rect 18656 28364 18662 28376
rect 19429 28373 19441 28376
rect 19475 28373 19487 28407
rect 19429 28367 19487 28373
rect 21266 28364 21272 28416
rect 21324 28404 21330 28416
rect 23934 28404 23940 28416
rect 21324 28376 23940 28404
rect 21324 28364 21330 28376
rect 23934 28364 23940 28376
rect 23992 28364 23998 28416
rect 24302 28404 24308 28416
rect 24263 28376 24308 28404
rect 24302 28364 24308 28376
rect 24360 28404 24366 28416
rect 24762 28404 24768 28416
rect 24360 28376 24768 28404
rect 24360 28364 24366 28376
rect 24762 28364 24768 28376
rect 24820 28364 24826 28416
rect 25038 28364 25044 28416
rect 25096 28404 25102 28416
rect 25501 28407 25559 28413
rect 25501 28404 25513 28407
rect 25096 28376 25513 28404
rect 25096 28364 25102 28376
rect 25501 28373 25513 28376
rect 25547 28404 25559 28407
rect 25590 28404 25596 28416
rect 25547 28376 25596 28404
rect 25547 28373 25559 28376
rect 25501 28367 25559 28373
rect 25590 28364 25596 28376
rect 25648 28364 25654 28416
rect 25866 28364 25872 28416
rect 25924 28404 25930 28416
rect 26789 28407 26847 28413
rect 26789 28404 26801 28407
rect 25924 28376 26801 28404
rect 25924 28364 25930 28376
rect 26789 28373 26801 28376
rect 26835 28373 26847 28407
rect 27154 28404 27160 28416
rect 27115 28376 27160 28404
rect 26789 28367 26847 28373
rect 27154 28364 27160 28376
rect 27212 28364 27218 28416
rect 28534 28404 28540 28416
rect 28495 28376 28540 28404
rect 28534 28364 28540 28376
rect 28592 28364 28598 28416
rect 33778 28404 33784 28416
rect 33739 28376 33784 28404
rect 33778 28364 33784 28376
rect 33836 28364 33842 28416
rect 1104 28314 38824 28336
rect 1104 28262 4246 28314
rect 4298 28262 4310 28314
rect 4362 28262 4374 28314
rect 4426 28262 4438 28314
rect 4490 28262 34966 28314
rect 35018 28262 35030 28314
rect 35082 28262 35094 28314
rect 35146 28262 35158 28314
rect 35210 28262 38824 28314
rect 1104 28240 38824 28262
rect 1670 28200 1676 28212
rect 1631 28172 1676 28200
rect 1670 28160 1676 28172
rect 1728 28160 1734 28212
rect 2222 28200 2228 28212
rect 2183 28172 2228 28200
rect 2222 28160 2228 28172
rect 2280 28160 2286 28212
rect 8389 28203 8447 28209
rect 8389 28169 8401 28203
rect 8435 28200 8447 28203
rect 8662 28200 8668 28212
rect 8435 28172 8668 28200
rect 8435 28169 8447 28172
rect 8389 28163 8447 28169
rect 8662 28160 8668 28172
rect 8720 28160 8726 28212
rect 9490 28200 9496 28212
rect 9451 28172 9496 28200
rect 9490 28160 9496 28172
rect 9548 28160 9554 28212
rect 10229 28203 10287 28209
rect 10229 28169 10241 28203
rect 10275 28200 10287 28203
rect 10318 28200 10324 28212
rect 10275 28172 10324 28200
rect 10275 28169 10287 28172
rect 10229 28163 10287 28169
rect 10318 28160 10324 28172
rect 10376 28160 10382 28212
rect 10502 28200 10508 28212
rect 10463 28172 10508 28200
rect 10502 28160 10508 28172
rect 10560 28160 10566 28212
rect 10778 28200 10784 28212
rect 10739 28172 10784 28200
rect 10778 28160 10784 28172
rect 10836 28160 10842 28212
rect 12434 28160 12440 28212
rect 12492 28200 12498 28212
rect 12897 28203 12955 28209
rect 12897 28200 12909 28203
rect 12492 28172 12909 28200
rect 12492 28160 12498 28172
rect 12897 28169 12909 28172
rect 12943 28169 12955 28203
rect 12897 28163 12955 28169
rect 14001 28203 14059 28209
rect 14001 28169 14013 28203
rect 14047 28200 14059 28203
rect 14734 28200 14740 28212
rect 14047 28172 14740 28200
rect 14047 28169 14059 28172
rect 14001 28163 14059 28169
rect 14734 28160 14740 28172
rect 14792 28160 14798 28212
rect 15102 28160 15108 28212
rect 15160 28160 15166 28212
rect 17770 28200 17776 28212
rect 17731 28172 17776 28200
rect 17770 28160 17776 28172
rect 17828 28160 17834 28212
rect 18230 28160 18236 28212
rect 18288 28200 18294 28212
rect 18509 28203 18567 28209
rect 18509 28200 18521 28203
rect 18288 28172 18521 28200
rect 18288 28160 18294 28172
rect 18509 28169 18521 28172
rect 18555 28169 18567 28203
rect 18874 28200 18880 28212
rect 18835 28172 18880 28200
rect 18509 28163 18567 28169
rect 18874 28160 18880 28172
rect 18932 28160 18938 28212
rect 19794 28160 19800 28212
rect 19852 28200 19858 28212
rect 20622 28200 20628 28212
rect 19852 28172 20628 28200
rect 19852 28160 19858 28172
rect 20622 28160 20628 28172
rect 20680 28160 20686 28212
rect 20990 28160 20996 28212
rect 21048 28200 21054 28212
rect 21269 28203 21327 28209
rect 21269 28200 21281 28203
rect 21048 28172 21281 28200
rect 21048 28160 21054 28172
rect 21269 28169 21281 28172
rect 21315 28169 21327 28203
rect 21269 28163 21327 28169
rect 21910 28160 21916 28212
rect 21968 28200 21974 28212
rect 22649 28203 22707 28209
rect 22649 28200 22661 28203
rect 21968 28172 22661 28200
rect 21968 28160 21974 28172
rect 22649 28169 22661 28172
rect 22695 28169 22707 28203
rect 23934 28200 23940 28212
rect 23895 28172 23940 28200
rect 22649 28163 22707 28169
rect 23934 28160 23940 28172
rect 23992 28160 23998 28212
rect 25866 28200 25872 28212
rect 25827 28172 25872 28200
rect 25866 28160 25872 28172
rect 25924 28160 25930 28212
rect 26237 28203 26295 28209
rect 26237 28169 26249 28203
rect 26283 28200 26295 28203
rect 26602 28200 26608 28212
rect 26283 28172 26608 28200
rect 26283 28169 26295 28172
rect 26237 28163 26295 28169
rect 26602 28160 26608 28172
rect 26660 28160 26666 28212
rect 27430 28160 27436 28212
rect 27488 28200 27494 28212
rect 28077 28203 28135 28209
rect 28077 28200 28089 28203
rect 27488 28172 28089 28200
rect 27488 28160 27494 28172
rect 28077 28169 28089 28172
rect 28123 28169 28135 28203
rect 28077 28163 28135 28169
rect 28166 28160 28172 28212
rect 28224 28200 28230 28212
rect 28629 28203 28687 28209
rect 28629 28200 28641 28203
rect 28224 28172 28641 28200
rect 28224 28160 28230 28172
rect 28629 28169 28641 28172
rect 28675 28169 28687 28203
rect 28629 28163 28687 28169
rect 29089 28203 29147 28209
rect 29089 28169 29101 28203
rect 29135 28200 29147 28203
rect 29178 28200 29184 28212
rect 29135 28172 29184 28200
rect 29135 28169 29147 28172
rect 29089 28163 29147 28169
rect 29178 28160 29184 28172
rect 29236 28200 29242 28212
rect 30006 28200 30012 28212
rect 29236 28172 30012 28200
rect 29236 28160 29242 28172
rect 30006 28160 30012 28172
rect 30064 28160 30070 28212
rect 32490 28200 32496 28212
rect 32451 28172 32496 28200
rect 32490 28160 32496 28172
rect 32548 28160 32554 28212
rect 32766 28200 32772 28212
rect 32727 28172 32772 28200
rect 32766 28160 32772 28172
rect 32824 28160 32830 28212
rect 2240 28064 2268 28160
rect 8570 28092 8576 28144
rect 8628 28132 8634 28144
rect 8757 28135 8815 28141
rect 8757 28132 8769 28135
rect 8628 28104 8769 28132
rect 8628 28092 8634 28104
rect 8757 28101 8769 28104
rect 8803 28101 8815 28135
rect 11606 28132 11612 28144
rect 11519 28104 11612 28132
rect 8757 28095 8815 28101
rect 11606 28092 11612 28104
rect 11664 28132 11670 28144
rect 11885 28135 11943 28141
rect 11885 28132 11897 28135
rect 11664 28104 11897 28132
rect 11664 28092 11670 28104
rect 11885 28101 11897 28104
rect 11931 28132 11943 28135
rect 14182 28132 14188 28144
rect 11931 28104 14188 28132
rect 11931 28101 11943 28104
rect 11885 28095 11943 28101
rect 14182 28092 14188 28104
rect 14240 28092 14246 28144
rect 15120 28132 15148 28160
rect 16758 28132 16764 28144
rect 15120 28104 15240 28132
rect 1412 28036 2268 28064
rect 1412 28005 1440 28036
rect 8478 28024 8484 28076
rect 8536 28064 8542 28076
rect 9122 28064 9128 28076
rect 8536 28036 9128 28064
rect 8536 28024 8542 28036
rect 9122 28024 9128 28036
rect 9180 28024 9186 28076
rect 9582 28024 9588 28076
rect 9640 28064 9646 28076
rect 9640 28036 10364 28064
rect 9640 28024 9646 28036
rect 1397 27999 1455 28005
rect 1397 27965 1409 27999
rect 1443 27965 1455 27999
rect 1578 27996 1584 28008
rect 1539 27968 1584 27996
rect 1397 27959 1455 27965
rect 1578 27956 1584 27968
rect 1636 27956 1642 28008
rect 7653 27999 7711 28005
rect 7653 27965 7665 27999
rect 7699 27996 7711 27999
rect 8938 27996 8944 28008
rect 7699 27968 8944 27996
rect 7699 27965 7711 27968
rect 7653 27959 7711 27965
rect 8938 27956 8944 27968
rect 8996 27956 9002 28008
rect 10336 28005 10364 28036
rect 10962 28024 10968 28076
rect 11020 28064 11026 28076
rect 13170 28064 13176 28076
rect 11020 28036 13176 28064
rect 11020 28024 11026 28036
rect 13170 28024 13176 28036
rect 13228 28024 13234 28076
rect 13538 28024 13544 28076
rect 13596 28064 13602 28076
rect 13633 28067 13691 28073
rect 13633 28064 13645 28067
rect 13596 28036 13645 28064
rect 13596 28024 13602 28036
rect 13633 28033 13645 28036
rect 13679 28064 13691 28067
rect 13998 28064 14004 28076
rect 13679 28036 14004 28064
rect 13679 28033 13691 28036
rect 13633 28027 13691 28033
rect 13998 28024 14004 28036
rect 14056 28024 14062 28076
rect 15102 28064 15108 28076
rect 14200 28036 15108 28064
rect 9309 27999 9367 28005
rect 9309 27965 9321 27999
rect 9355 27996 9367 27999
rect 10321 27999 10379 28005
rect 9355 27968 9904 27996
rect 9355 27965 9367 27968
rect 9309 27959 9367 27965
rect 7282 27928 7288 27940
rect 7195 27900 7288 27928
rect 7282 27888 7288 27900
rect 7340 27928 7346 27940
rect 8386 27928 8392 27940
rect 7340 27900 8392 27928
rect 7340 27888 7346 27900
rect 8386 27888 8392 27900
rect 8444 27888 8450 27940
rect 9876 27872 9904 27968
rect 10321 27965 10333 27999
rect 10367 27996 10379 27999
rect 11333 27999 11391 28005
rect 10367 27968 11284 27996
rect 10367 27965 10379 27968
rect 10321 27959 10379 27965
rect 8018 27860 8024 27872
rect 7979 27832 8024 27860
rect 8018 27820 8024 27832
rect 8076 27820 8082 27872
rect 9858 27860 9864 27872
rect 9819 27832 9864 27860
rect 9858 27820 9864 27832
rect 9916 27820 9922 27872
rect 11256 27869 11284 27968
rect 11333 27965 11345 27999
rect 11379 27996 11391 27999
rect 11609 27999 11667 28005
rect 11609 27996 11621 27999
rect 11379 27968 11621 27996
rect 11379 27965 11391 27968
rect 11333 27959 11391 27965
rect 11609 27965 11621 27968
rect 11655 27965 11667 27999
rect 11609 27959 11667 27965
rect 12158 27956 12164 28008
rect 12216 27996 12222 28008
rect 12713 27999 12771 28005
rect 12713 27996 12725 27999
rect 12216 27968 12725 27996
rect 12216 27956 12222 27968
rect 12713 27965 12725 27968
rect 12759 27996 12771 27999
rect 12759 27968 13492 27996
rect 12759 27965 12771 27968
rect 12713 27959 12771 27965
rect 13464 27872 13492 27968
rect 13722 27956 13728 28008
rect 13780 27996 13786 28008
rect 14200 28005 14228 28036
rect 15102 28024 15108 28036
rect 15160 28024 15166 28076
rect 14185 27999 14243 28005
rect 14185 27996 14197 27999
rect 13780 27968 14197 27996
rect 13780 27956 13786 27968
rect 14185 27965 14197 27968
rect 14231 27965 14243 27999
rect 14185 27959 14243 27965
rect 14369 27999 14427 28005
rect 14369 27965 14381 27999
rect 14415 27996 14427 27999
rect 14642 27996 14648 28008
rect 14415 27968 14648 27996
rect 14415 27965 14427 27968
rect 14369 27959 14427 27965
rect 13998 27888 14004 27940
rect 14056 27928 14062 27940
rect 14384 27928 14412 27959
rect 14642 27956 14648 27968
rect 14700 27956 14706 28008
rect 14737 27999 14795 28005
rect 14737 27965 14749 27999
rect 14783 27965 14795 27999
rect 14737 27959 14795 27965
rect 14056 27900 14412 27928
rect 14056 27888 14062 27900
rect 14458 27888 14464 27940
rect 14516 27928 14522 27940
rect 14752 27928 14780 27959
rect 14826 27956 14832 28008
rect 14884 27996 14890 28008
rect 14921 27999 14979 28005
rect 14921 27996 14933 27999
rect 14884 27968 14933 27996
rect 14884 27956 14890 27968
rect 14921 27965 14933 27968
rect 14967 27996 14979 27999
rect 15212 27996 15240 28104
rect 14967 27968 15240 27996
rect 15304 28104 16764 28132
rect 14967 27965 14979 27968
rect 14921 27959 14979 27965
rect 14516 27900 14780 27928
rect 14516 27888 14522 27900
rect 11241 27863 11299 27869
rect 11241 27829 11253 27863
rect 11287 27860 11299 27863
rect 11330 27860 11336 27872
rect 11287 27832 11336 27860
rect 11287 27829 11299 27832
rect 11241 27823 11299 27829
rect 11330 27820 11336 27832
rect 11388 27820 11394 27872
rect 11422 27820 11428 27872
rect 11480 27860 11486 27872
rect 11517 27863 11575 27869
rect 11517 27860 11529 27863
rect 11480 27832 11529 27860
rect 11480 27820 11486 27832
rect 11517 27829 11529 27832
rect 11563 27829 11575 27863
rect 11517 27823 11575 27829
rect 12253 27863 12311 27869
rect 12253 27829 12265 27863
rect 12299 27860 12311 27863
rect 12434 27860 12440 27872
rect 12299 27832 12440 27860
rect 12299 27829 12311 27832
rect 12253 27823 12311 27829
rect 12434 27820 12440 27832
rect 12492 27860 12498 27872
rect 12894 27860 12900 27872
rect 12492 27832 12900 27860
rect 12492 27820 12498 27832
rect 12894 27820 12900 27832
rect 12952 27820 12958 27872
rect 13265 27863 13323 27869
rect 13265 27829 13277 27863
rect 13311 27860 13323 27863
rect 13446 27860 13452 27872
rect 13311 27832 13452 27860
rect 13311 27829 13323 27832
rect 13265 27823 13323 27829
rect 13446 27820 13452 27832
rect 13504 27820 13510 27872
rect 14182 27820 14188 27872
rect 14240 27860 14246 27872
rect 15304 27869 15332 28104
rect 16758 28092 16764 28104
rect 16816 28092 16822 28144
rect 17954 28092 17960 28144
rect 18012 28132 18018 28144
rect 20717 28135 20775 28141
rect 18012 28104 20392 28132
rect 18012 28092 18018 28104
rect 15749 28067 15807 28073
rect 15749 28033 15761 28067
rect 15795 28064 15807 28067
rect 16114 28064 16120 28076
rect 15795 28036 16120 28064
rect 15795 28033 15807 28036
rect 15749 28027 15807 28033
rect 16114 28024 16120 28036
rect 16172 28024 16178 28076
rect 16298 28064 16304 28076
rect 16259 28036 16304 28064
rect 16298 28024 16304 28036
rect 16356 28064 16362 28076
rect 17218 28064 17224 28076
rect 16356 28036 17224 28064
rect 16356 28024 16362 28036
rect 17218 28024 17224 28036
rect 17276 28064 17282 28076
rect 17405 28067 17463 28073
rect 17405 28064 17417 28067
rect 17276 28036 17417 28064
rect 17276 28024 17282 28036
rect 17405 28033 17417 28036
rect 17451 28033 17463 28067
rect 17405 28027 17463 28033
rect 19245 28067 19303 28073
rect 19245 28033 19257 28067
rect 19291 28064 19303 28067
rect 20254 28064 20260 28076
rect 19291 28036 20260 28064
rect 19291 28033 19303 28036
rect 19245 28027 19303 28033
rect 16577 27999 16635 28005
rect 16577 27965 16589 27999
rect 16623 27996 16635 27999
rect 16666 27996 16672 28008
rect 16623 27968 16672 27996
rect 16623 27965 16635 27968
rect 16577 27959 16635 27965
rect 16666 27956 16672 27968
rect 16724 27956 16730 28008
rect 16761 27999 16819 28005
rect 16761 27965 16773 27999
rect 16807 27965 16819 27999
rect 16761 27959 16819 27965
rect 18325 27999 18383 28005
rect 18325 27965 18337 27999
rect 18371 27996 18383 27999
rect 18874 27996 18880 28008
rect 18371 27968 18880 27996
rect 18371 27965 18383 27968
rect 18325 27959 18383 27965
rect 15289 27863 15347 27869
rect 15289 27860 15301 27863
rect 14240 27832 15301 27860
rect 14240 27820 14246 27832
rect 15289 27829 15301 27832
rect 15335 27829 15347 27863
rect 15289 27823 15347 27829
rect 15930 27820 15936 27872
rect 15988 27860 15994 27872
rect 16776 27860 16804 27959
rect 18874 27956 18880 27968
rect 18932 27956 18938 28008
rect 19628 28005 19656 28036
rect 20254 28024 20260 28036
rect 20312 28024 20318 28076
rect 20364 28064 20392 28104
rect 20717 28101 20729 28135
rect 20763 28132 20775 28135
rect 20806 28132 20812 28144
rect 20763 28104 20812 28132
rect 20763 28101 20775 28104
rect 20717 28095 20775 28101
rect 20806 28092 20812 28104
rect 20864 28092 20870 28144
rect 23106 28132 23112 28144
rect 23067 28104 23112 28132
rect 23106 28092 23112 28104
rect 23164 28092 23170 28144
rect 24026 28092 24032 28144
rect 24084 28132 24090 28144
rect 25501 28135 25559 28141
rect 25501 28132 25513 28135
rect 24084 28104 25513 28132
rect 24084 28092 24090 28104
rect 25501 28101 25513 28104
rect 25547 28132 25559 28135
rect 25547 28104 25728 28132
rect 25547 28101 25559 28104
rect 25501 28095 25559 28101
rect 20990 28064 20996 28076
rect 20364 28036 20996 28064
rect 19613 27999 19671 28005
rect 19613 27965 19625 27999
rect 19659 27965 19671 27999
rect 19794 27996 19800 28008
rect 19755 27968 19800 27996
rect 19613 27959 19671 27965
rect 19794 27956 19800 27968
rect 19852 27956 19858 28008
rect 20364 28005 20392 28036
rect 20990 28024 20996 28036
rect 21048 28024 21054 28076
rect 21545 28067 21603 28073
rect 21545 28033 21557 28067
rect 21591 28064 21603 28067
rect 21637 28067 21695 28073
rect 21637 28064 21649 28067
rect 21591 28036 21649 28064
rect 21591 28033 21603 28036
rect 21545 28027 21603 28033
rect 21637 28033 21649 28036
rect 21683 28064 21695 28067
rect 21726 28064 21732 28076
rect 21683 28036 21732 28064
rect 21683 28033 21695 28036
rect 21637 28027 21695 28033
rect 21726 28024 21732 28036
rect 21784 28024 21790 28076
rect 23290 28064 23296 28076
rect 23124 28036 23296 28064
rect 23124 28008 23152 28036
rect 23290 28024 23296 28036
rect 23348 28064 23354 28076
rect 24121 28067 24179 28073
rect 24121 28064 24133 28067
rect 23348 28036 24133 28064
rect 23348 28024 23354 28036
rect 24121 28033 24133 28036
rect 24167 28064 24179 28067
rect 25133 28067 25191 28073
rect 25133 28064 25145 28067
rect 24167 28036 25145 28064
rect 24167 28033 24179 28036
rect 24121 28027 24179 28033
rect 25133 28033 25145 28036
rect 25179 28033 25191 28067
rect 25590 28064 25596 28076
rect 25133 28027 25191 28033
rect 25240 28036 25596 28064
rect 20349 27999 20407 28005
rect 20349 27965 20361 27999
rect 20395 27965 20407 27999
rect 20625 27999 20683 28005
rect 20625 27996 20637 27999
rect 20349 27959 20407 27965
rect 20456 27968 20637 27996
rect 20456 27872 20484 27968
rect 20625 27965 20637 27968
rect 20671 27996 20683 27999
rect 20806 27996 20812 28008
rect 20671 27968 20812 27996
rect 20671 27965 20683 27968
rect 20625 27959 20683 27965
rect 20806 27956 20812 27968
rect 20864 27956 20870 28008
rect 21269 27999 21327 28005
rect 21269 27965 21281 27999
rect 21315 27996 21327 27999
rect 21989 27999 22047 28005
rect 21989 27996 22001 27999
rect 21315 27968 22001 27996
rect 21315 27965 21327 27968
rect 21269 27959 21327 27965
rect 21989 27965 22001 27968
rect 22035 27965 22047 27999
rect 21989 27959 22047 27965
rect 23106 27956 23112 28008
rect 23164 27956 23170 28008
rect 24305 27999 24363 28005
rect 24305 27965 24317 27999
rect 24351 27965 24363 27999
rect 24670 27996 24676 28008
rect 24631 27968 24676 27996
rect 24305 27959 24363 27965
rect 20898 27888 20904 27940
rect 20956 27928 20962 27940
rect 21726 27928 21732 27940
rect 20956 27900 21732 27928
rect 20956 27888 20962 27900
rect 21726 27888 21732 27900
rect 21784 27928 21790 27940
rect 21821 27931 21879 27937
rect 21821 27928 21833 27931
rect 21784 27900 21833 27928
rect 21784 27888 21790 27900
rect 21821 27897 21833 27900
rect 21867 27928 21879 27931
rect 21867 27900 22032 27928
rect 21867 27897 21879 27900
rect 21821 27891 21879 27897
rect 17034 27860 17040 27872
rect 15988 27832 17040 27860
rect 15988 27820 15994 27832
rect 17034 27820 17040 27832
rect 17092 27820 17098 27872
rect 20070 27820 20076 27872
rect 20128 27860 20134 27872
rect 20254 27860 20260 27872
rect 20128 27832 20260 27860
rect 20128 27820 20134 27832
rect 20254 27820 20260 27832
rect 20312 27820 20318 27872
rect 20438 27820 20444 27872
rect 20496 27820 20502 27872
rect 20806 27820 20812 27872
rect 20864 27860 20870 27872
rect 21085 27863 21143 27869
rect 21085 27860 21097 27863
rect 20864 27832 21097 27860
rect 20864 27820 20870 27832
rect 21085 27829 21097 27832
rect 21131 27860 21143 27863
rect 21174 27860 21180 27872
rect 21131 27832 21180 27860
rect 21131 27829 21143 27832
rect 21085 27823 21143 27829
rect 21174 27820 21180 27832
rect 21232 27820 21238 27872
rect 21910 27860 21916 27872
rect 21871 27832 21916 27860
rect 21910 27820 21916 27832
rect 21968 27820 21974 27872
rect 22004 27860 22032 27900
rect 22186 27888 22192 27940
rect 22244 27928 22250 27940
rect 22373 27931 22431 27937
rect 22373 27928 22385 27931
rect 22244 27900 22385 27928
rect 22244 27888 22250 27900
rect 22373 27897 22385 27900
rect 22419 27897 22431 27931
rect 22373 27891 22431 27897
rect 22922 27888 22928 27940
rect 22980 27928 22986 27940
rect 23934 27928 23940 27940
rect 22980 27900 23940 27928
rect 22980 27888 22986 27900
rect 23934 27888 23940 27900
rect 23992 27888 23998 27940
rect 24320 27928 24348 27959
rect 24670 27956 24676 27968
rect 24728 27956 24734 28008
rect 24854 27996 24860 28008
rect 24815 27968 24860 27996
rect 24854 27956 24860 27968
rect 24912 27956 24918 28008
rect 25240 27928 25268 28036
rect 25590 28024 25596 28036
rect 25648 28024 25654 28076
rect 25700 28005 25728 28104
rect 26697 28067 26755 28073
rect 26697 28033 26709 28067
rect 26743 28064 26755 28067
rect 27062 28064 27068 28076
rect 26743 28036 27068 28064
rect 26743 28033 26755 28036
rect 26697 28027 26755 28033
rect 27062 28024 27068 28036
rect 27120 28024 27126 28076
rect 25685 27999 25743 28005
rect 25685 27965 25697 27999
rect 25731 27965 25743 27999
rect 26973 27999 27031 28005
rect 26973 27996 26985 27999
rect 25685 27959 25743 27965
rect 26528 27968 26985 27996
rect 24320 27900 25268 27928
rect 26528 27872 26556 27968
rect 26973 27965 26985 27968
rect 27019 27965 27031 27999
rect 29270 27996 29276 28008
rect 29231 27968 29276 27996
rect 26973 27959 27031 27965
rect 29270 27956 29276 27968
rect 29328 27996 29334 28008
rect 29733 27999 29791 28005
rect 29733 27996 29745 27999
rect 29328 27968 29745 27996
rect 29328 27956 29334 27968
rect 29733 27965 29745 27968
rect 29779 27965 29791 27999
rect 29733 27959 29791 27965
rect 22462 27860 22468 27872
rect 22004 27832 22468 27860
rect 22462 27820 22468 27832
rect 22520 27860 22526 27872
rect 23477 27863 23535 27869
rect 23477 27860 23489 27863
rect 22520 27832 23489 27860
rect 22520 27820 22526 27832
rect 23477 27829 23489 27832
rect 23523 27860 23535 27863
rect 25038 27860 25044 27872
rect 23523 27832 25044 27860
rect 23523 27829 23535 27832
rect 23477 27823 23535 27829
rect 25038 27820 25044 27832
rect 25096 27820 25102 27872
rect 26510 27860 26516 27872
rect 26471 27832 26516 27860
rect 26510 27820 26516 27832
rect 26568 27820 26574 27872
rect 29454 27860 29460 27872
rect 29415 27832 29460 27860
rect 29454 27820 29460 27832
rect 29512 27820 29518 27872
rect 1104 27770 38824 27792
rect 1104 27718 19606 27770
rect 19658 27718 19670 27770
rect 19722 27718 19734 27770
rect 19786 27718 19798 27770
rect 19850 27718 38824 27770
rect 1104 27696 38824 27718
rect 8294 27616 8300 27668
rect 8352 27656 8358 27668
rect 8665 27659 8723 27665
rect 8665 27656 8677 27659
rect 8352 27628 8677 27656
rect 8352 27616 8358 27628
rect 8665 27625 8677 27628
rect 8711 27625 8723 27659
rect 10778 27656 10784 27668
rect 10739 27628 10784 27656
rect 8665 27619 8723 27625
rect 10778 27616 10784 27628
rect 10836 27616 10842 27668
rect 12434 27656 12440 27668
rect 12395 27628 12440 27656
rect 12434 27616 12440 27628
rect 12492 27616 12498 27668
rect 12897 27659 12955 27665
rect 12897 27625 12909 27659
rect 12943 27656 12955 27659
rect 13354 27656 13360 27668
rect 12943 27628 13360 27656
rect 12943 27625 12955 27628
rect 12897 27619 12955 27625
rect 13354 27616 13360 27628
rect 13412 27656 13418 27668
rect 14090 27656 14096 27668
rect 13412 27628 14096 27656
rect 13412 27616 13418 27628
rect 14090 27616 14096 27628
rect 14148 27616 14154 27668
rect 17310 27616 17316 27668
rect 17368 27656 17374 27668
rect 17368 27628 17540 27656
rect 17368 27616 17374 27628
rect 10502 27588 10508 27600
rect 10463 27560 10508 27588
rect 10502 27548 10508 27560
rect 10560 27548 10566 27600
rect 11149 27591 11207 27597
rect 11149 27557 11161 27591
rect 11195 27588 11207 27591
rect 12986 27588 12992 27600
rect 11195 27560 12848 27588
rect 12947 27560 12992 27588
rect 11195 27557 11207 27560
rect 11149 27551 11207 27557
rect 5994 27480 6000 27532
rect 6052 27520 6058 27532
rect 6733 27523 6791 27529
rect 6733 27520 6745 27523
rect 6052 27492 6745 27520
rect 6052 27480 6058 27492
rect 6733 27489 6745 27492
rect 6779 27520 6791 27523
rect 6822 27520 6828 27532
rect 6779 27492 6828 27520
rect 6779 27489 6791 27492
rect 6733 27483 6791 27489
rect 6822 27480 6828 27492
rect 6880 27480 6886 27532
rect 10594 27520 10600 27532
rect 10555 27492 10600 27520
rect 10594 27480 10600 27492
rect 10652 27480 10658 27532
rect 11698 27520 11704 27532
rect 11611 27492 11704 27520
rect 11698 27480 11704 27492
rect 11756 27520 11762 27532
rect 12618 27520 12624 27532
rect 11756 27492 12624 27520
rect 11756 27480 11762 27492
rect 12618 27480 12624 27492
rect 12676 27480 12682 27532
rect 12820 27520 12848 27560
rect 12986 27548 12992 27560
rect 13044 27548 13050 27600
rect 14829 27591 14887 27597
rect 14829 27557 14841 27591
rect 14875 27588 14887 27591
rect 14918 27588 14924 27600
rect 14875 27560 14924 27588
rect 14875 27557 14887 27560
rect 14829 27551 14887 27557
rect 14918 27548 14924 27560
rect 14976 27548 14982 27600
rect 15102 27548 15108 27600
rect 15160 27588 15166 27600
rect 16209 27591 16267 27597
rect 16209 27588 16221 27591
rect 15160 27560 16221 27588
rect 15160 27548 15166 27560
rect 16209 27557 16221 27560
rect 16255 27588 16267 27591
rect 16850 27588 16856 27600
rect 16255 27560 16856 27588
rect 16255 27557 16267 27560
rect 16209 27551 16267 27557
rect 16850 27548 16856 27560
rect 16908 27548 16914 27600
rect 17402 27588 17408 27600
rect 17363 27560 17408 27588
rect 17402 27548 17408 27560
rect 17460 27548 17466 27600
rect 17512 27588 17540 27628
rect 18322 27616 18328 27668
rect 18380 27656 18386 27668
rect 18417 27659 18475 27665
rect 18417 27656 18429 27659
rect 18380 27628 18429 27656
rect 18380 27616 18386 27628
rect 18417 27625 18429 27628
rect 18463 27625 18475 27659
rect 18417 27619 18475 27625
rect 18598 27616 18604 27668
rect 18656 27656 18662 27668
rect 18877 27659 18935 27665
rect 18877 27656 18889 27659
rect 18656 27628 18889 27656
rect 18656 27616 18662 27628
rect 18877 27625 18889 27628
rect 18923 27656 18935 27659
rect 20254 27656 20260 27668
rect 18923 27628 20260 27656
rect 18923 27625 18935 27628
rect 18877 27619 18935 27625
rect 20254 27616 20260 27628
rect 20312 27616 20318 27668
rect 20346 27616 20352 27668
rect 20404 27656 20410 27668
rect 20717 27659 20775 27665
rect 20717 27656 20729 27659
rect 20404 27628 20729 27656
rect 20404 27616 20410 27628
rect 20717 27625 20729 27628
rect 20763 27625 20775 27659
rect 21266 27656 21272 27668
rect 20717 27619 20775 27625
rect 20805 27628 21272 27656
rect 17770 27588 17776 27600
rect 17512 27560 17776 27588
rect 17770 27548 17776 27560
rect 17828 27548 17834 27600
rect 18046 27548 18052 27600
rect 18104 27588 18110 27600
rect 18104 27560 19104 27588
rect 18104 27548 18110 27560
rect 13722 27520 13728 27532
rect 12820 27492 13728 27520
rect 13722 27480 13728 27492
rect 13780 27480 13786 27532
rect 13814 27480 13820 27532
rect 13872 27520 13878 27532
rect 14001 27523 14059 27529
rect 13872 27492 13917 27520
rect 13872 27480 13878 27492
rect 14001 27489 14013 27523
rect 14047 27520 14059 27523
rect 14734 27520 14740 27532
rect 14047 27492 14740 27520
rect 14047 27489 14059 27492
rect 14001 27483 14059 27489
rect 7009 27455 7067 27461
rect 7009 27421 7021 27455
rect 7055 27452 7067 27455
rect 7098 27452 7104 27464
rect 7055 27424 7104 27452
rect 7055 27421 7067 27424
rect 7009 27415 7067 27421
rect 7098 27412 7104 27424
rect 7156 27412 7162 27464
rect 7466 27412 7472 27464
rect 7524 27452 7530 27464
rect 9033 27455 9091 27461
rect 9033 27452 9045 27455
rect 7524 27424 9045 27452
rect 7524 27412 7530 27424
rect 9033 27421 9045 27424
rect 9079 27452 9091 27455
rect 9122 27452 9128 27464
rect 9079 27424 9128 27452
rect 9079 27421 9091 27424
rect 9033 27415 9091 27421
rect 9122 27412 9128 27424
rect 9180 27412 9186 27464
rect 10134 27452 10140 27464
rect 10095 27424 10140 27452
rect 10134 27412 10140 27424
rect 10192 27412 10198 27464
rect 11609 27455 11667 27461
rect 11609 27421 11621 27455
rect 11655 27452 11667 27455
rect 12250 27452 12256 27464
rect 11655 27424 12256 27452
rect 11655 27421 11667 27424
rect 11609 27415 11667 27421
rect 12250 27412 12256 27424
rect 12308 27412 12314 27464
rect 13538 27452 13544 27464
rect 13499 27424 13544 27452
rect 13538 27412 13544 27424
rect 13596 27412 13602 27464
rect 1578 27316 1584 27328
rect 1539 27288 1584 27316
rect 1578 27276 1584 27288
rect 1636 27276 1642 27328
rect 8294 27316 8300 27328
rect 8255 27288 8300 27316
rect 8294 27276 8300 27288
rect 8352 27276 8358 27328
rect 8386 27276 8392 27328
rect 8444 27316 8450 27328
rect 8938 27316 8944 27328
rect 8444 27288 8944 27316
rect 8444 27276 8450 27288
rect 8938 27276 8944 27288
rect 8996 27316 9002 27328
rect 9401 27319 9459 27325
rect 9401 27316 9413 27319
rect 8996 27288 9413 27316
rect 8996 27276 9002 27288
rect 9401 27285 9413 27288
rect 9447 27285 9459 27319
rect 9401 27279 9459 27285
rect 11517 27319 11575 27325
rect 11517 27285 11529 27319
rect 11563 27316 11575 27319
rect 11882 27316 11888 27328
rect 11563 27288 11888 27316
rect 11563 27285 11575 27288
rect 11517 27279 11575 27285
rect 11882 27276 11888 27288
rect 11940 27276 11946 27328
rect 13538 27276 13544 27328
rect 13596 27316 13602 27328
rect 14200 27316 14228 27492
rect 14734 27480 14740 27492
rect 14792 27480 14798 27532
rect 15838 27520 15844 27532
rect 15799 27492 15844 27520
rect 15838 27480 15844 27492
rect 15896 27480 15902 27532
rect 16025 27523 16083 27529
rect 16025 27489 16037 27523
rect 16071 27489 16083 27523
rect 16025 27483 16083 27489
rect 14458 27452 14464 27464
rect 14419 27424 14464 27452
rect 14458 27412 14464 27424
rect 14516 27412 14522 27464
rect 16040 27452 16068 27483
rect 16114 27480 16120 27532
rect 16172 27520 16178 27532
rect 17313 27523 17371 27529
rect 16172 27492 16217 27520
rect 16172 27480 16178 27492
rect 17313 27489 17325 27523
rect 17359 27520 17371 27523
rect 17586 27520 17592 27532
rect 17359 27492 17592 27520
rect 17359 27489 17371 27492
rect 17313 27483 17371 27489
rect 16206 27452 16212 27464
rect 16040 27424 16212 27452
rect 16206 27412 16212 27424
rect 16264 27412 16270 27464
rect 16298 27412 16304 27464
rect 16356 27452 16362 27464
rect 16577 27455 16635 27461
rect 16577 27452 16589 27455
rect 16356 27424 16589 27452
rect 16356 27412 16362 27424
rect 16577 27421 16589 27424
rect 16623 27421 16635 27455
rect 16577 27415 16635 27421
rect 14642 27344 14648 27396
rect 14700 27384 14706 27396
rect 15470 27384 15476 27396
rect 14700 27356 15476 27384
rect 14700 27344 14706 27356
rect 15470 27344 15476 27356
rect 15528 27384 15534 27396
rect 15749 27387 15807 27393
rect 15749 27384 15761 27387
rect 15528 27356 15761 27384
rect 15528 27344 15534 27356
rect 15749 27353 15761 27356
rect 15795 27384 15807 27387
rect 17328 27384 17356 27483
rect 17586 27480 17592 27492
rect 17644 27480 17650 27532
rect 17681 27523 17739 27529
rect 17681 27489 17693 27523
rect 17727 27520 17739 27523
rect 17862 27520 17868 27532
rect 17727 27492 17868 27520
rect 17727 27489 17739 27492
rect 17681 27483 17739 27489
rect 17862 27480 17868 27492
rect 17920 27480 17926 27532
rect 18966 27520 18972 27532
rect 18927 27492 18972 27520
rect 18966 27480 18972 27492
rect 19024 27480 19030 27532
rect 19076 27520 19104 27560
rect 19426 27548 19432 27600
rect 19484 27588 19490 27600
rect 19978 27588 19984 27600
rect 19484 27560 19984 27588
rect 19484 27548 19490 27560
rect 19978 27548 19984 27560
rect 20036 27548 20042 27600
rect 20622 27548 20628 27600
rect 20680 27588 20686 27600
rect 20732 27588 20760 27619
rect 20680 27560 20760 27588
rect 20680 27548 20686 27560
rect 19518 27520 19524 27532
rect 19076 27492 19524 27520
rect 19518 27480 19524 27492
rect 19576 27520 19582 27532
rect 20805 27520 20833 27628
rect 21266 27616 21272 27628
rect 21324 27616 21330 27668
rect 21910 27616 21916 27668
rect 21968 27656 21974 27668
rect 22097 27659 22155 27665
rect 22097 27656 22109 27659
rect 21968 27628 22109 27656
rect 21968 27616 21974 27628
rect 22097 27625 22109 27628
rect 22143 27625 22155 27659
rect 22097 27619 22155 27625
rect 22189 27659 22247 27665
rect 22189 27625 22201 27659
rect 22235 27656 22247 27659
rect 22554 27656 22560 27668
rect 22235 27628 22560 27656
rect 22235 27625 22247 27628
rect 22189 27619 22247 27625
rect 22554 27616 22560 27628
rect 22612 27616 22618 27668
rect 24118 27656 24124 27668
rect 23584 27628 24124 27656
rect 20901 27591 20959 27597
rect 20901 27557 20913 27591
rect 20947 27588 20959 27591
rect 21634 27588 21640 27600
rect 20947 27560 21640 27588
rect 20947 27557 20959 27560
rect 20901 27551 20959 27557
rect 21634 27548 21640 27560
rect 21692 27588 21698 27600
rect 23477 27591 23535 27597
rect 23477 27588 23489 27591
rect 21692 27560 23489 27588
rect 21692 27548 21698 27560
rect 23477 27557 23489 27560
rect 23523 27557 23535 27591
rect 23477 27551 23535 27557
rect 21082 27529 21088 27532
rect 19576 27492 20833 27520
rect 21048 27523 21088 27529
rect 19576 27480 19582 27492
rect 21048 27489 21060 27523
rect 21048 27483 21088 27489
rect 21082 27480 21088 27483
rect 21140 27480 21146 27532
rect 21726 27480 21732 27532
rect 21784 27520 21790 27532
rect 21913 27523 21971 27529
rect 21913 27520 21925 27523
rect 21784 27492 21925 27520
rect 21784 27480 21790 27492
rect 21913 27489 21925 27492
rect 21959 27489 21971 27523
rect 22465 27523 22523 27529
rect 22465 27520 22477 27523
rect 21913 27483 21971 27489
rect 22020 27492 22477 27520
rect 22020 27464 22048 27492
rect 22465 27489 22477 27492
rect 22511 27520 22523 27523
rect 22511 27492 22692 27520
rect 22511 27489 22523 27492
rect 22465 27483 22523 27489
rect 18046 27412 18052 27464
rect 18104 27452 18110 27464
rect 18141 27455 18199 27461
rect 18141 27452 18153 27455
rect 18104 27424 18153 27452
rect 18104 27412 18110 27424
rect 18141 27421 18153 27424
rect 18187 27452 18199 27455
rect 19337 27455 19395 27461
rect 19337 27452 19349 27455
rect 18187 27424 19349 27452
rect 18187 27421 18199 27424
rect 18141 27415 18199 27421
rect 19337 27421 19349 27424
rect 19383 27421 19395 27455
rect 21266 27452 21272 27464
rect 21227 27424 21272 27452
rect 19337 27415 19395 27421
rect 21266 27412 21272 27424
rect 21324 27412 21330 27464
rect 22002 27412 22008 27464
rect 22060 27412 22066 27464
rect 22278 27412 22284 27464
rect 22336 27452 22342 27464
rect 22336 27424 22508 27452
rect 22336 27412 22342 27424
rect 19150 27393 19156 27396
rect 15795 27356 17356 27384
rect 19134 27387 19156 27393
rect 15795 27353 15807 27356
rect 15749 27347 15807 27353
rect 19134 27353 19146 27387
rect 19134 27347 19156 27353
rect 19150 27344 19156 27347
rect 19208 27344 19214 27396
rect 21177 27387 21235 27393
rect 21177 27353 21189 27387
rect 21223 27384 21235 27387
rect 22189 27387 22247 27393
rect 22189 27384 22201 27387
rect 21223 27356 22201 27384
rect 21223 27353 21235 27356
rect 21177 27347 21235 27353
rect 22189 27353 22201 27356
rect 22235 27353 22247 27387
rect 22189 27347 22247 27353
rect 22480 27328 22508 27424
rect 22664 27384 22692 27492
rect 22738 27480 22744 27532
rect 22796 27520 22802 27532
rect 23201 27523 23259 27529
rect 23201 27520 23213 27523
rect 22796 27492 23213 27520
rect 22796 27480 22802 27492
rect 23201 27489 23213 27492
rect 23247 27489 23259 27523
rect 23201 27483 23259 27489
rect 22833 27455 22891 27461
rect 22833 27421 22845 27455
rect 22879 27452 22891 27455
rect 23382 27452 23388 27464
rect 22879 27424 23388 27452
rect 22879 27421 22891 27424
rect 22833 27415 22891 27421
rect 23382 27412 23388 27424
rect 23440 27412 23446 27464
rect 23584 27452 23612 27628
rect 24118 27616 24124 27628
rect 24176 27616 24182 27668
rect 24670 27616 24676 27668
rect 24728 27656 24734 27668
rect 24728 27628 24808 27656
rect 24728 27616 24734 27628
rect 23658 27548 23664 27600
rect 23716 27588 23722 27600
rect 24026 27588 24032 27600
rect 23716 27560 24032 27588
rect 23716 27548 23722 27560
rect 24026 27548 24032 27560
rect 24084 27548 24090 27600
rect 24397 27591 24455 27597
rect 24397 27557 24409 27591
rect 24443 27588 24455 27591
rect 24486 27588 24492 27600
rect 24443 27560 24492 27588
rect 24443 27557 24455 27560
rect 24397 27551 24455 27557
rect 24486 27548 24492 27560
rect 24544 27548 24550 27600
rect 24780 27588 24808 27628
rect 25866 27616 25872 27668
rect 25924 27656 25930 27668
rect 26237 27659 26295 27665
rect 26237 27656 26249 27659
rect 25924 27628 26249 27656
rect 25924 27616 25930 27628
rect 26237 27625 26249 27628
rect 26283 27625 26295 27659
rect 26237 27619 26295 27625
rect 26697 27659 26755 27665
rect 26697 27625 26709 27659
rect 26743 27656 26755 27659
rect 26786 27656 26792 27668
rect 26743 27628 26792 27656
rect 26743 27625 26755 27628
rect 26697 27619 26755 27625
rect 26786 27616 26792 27628
rect 26844 27656 26850 27668
rect 26973 27659 27031 27665
rect 26973 27656 26985 27659
rect 26844 27628 26985 27656
rect 26844 27616 26850 27628
rect 26973 27625 26985 27628
rect 27019 27625 27031 27659
rect 26973 27619 27031 27625
rect 27062 27616 27068 27668
rect 27120 27656 27126 27668
rect 27120 27628 27660 27656
rect 27120 27616 27126 27628
rect 25314 27588 25320 27600
rect 24780 27560 25320 27588
rect 25314 27548 25320 27560
rect 25372 27588 25378 27600
rect 25777 27591 25835 27597
rect 25777 27588 25789 27591
rect 25372 27560 25789 27588
rect 25372 27548 25378 27560
rect 25777 27557 25789 27560
rect 25823 27557 25835 27591
rect 27338 27588 27344 27600
rect 27299 27560 27344 27588
rect 25777 27551 25835 27557
rect 27338 27548 27344 27560
rect 27396 27548 27402 27600
rect 27632 27588 27660 27628
rect 28813 27591 28871 27597
rect 28813 27588 28825 27591
rect 27632 27560 28825 27588
rect 28813 27557 28825 27560
rect 28859 27588 28871 27591
rect 28902 27588 28908 27600
rect 28859 27560 28908 27588
rect 28859 27557 28871 27560
rect 28813 27551 28871 27557
rect 28902 27548 28908 27560
rect 28960 27548 28966 27600
rect 23842 27480 23848 27532
rect 23900 27520 23906 27532
rect 24213 27523 24271 27529
rect 24213 27520 24225 27523
rect 23900 27492 24225 27520
rect 23900 27480 23906 27492
rect 24213 27489 24225 27492
rect 24259 27489 24271 27523
rect 24213 27483 24271 27489
rect 24305 27523 24363 27529
rect 24305 27489 24317 27523
rect 24351 27520 24363 27523
rect 24670 27520 24676 27532
rect 24351 27492 24676 27520
rect 24351 27489 24363 27492
rect 24305 27483 24363 27489
rect 24670 27480 24676 27492
rect 24728 27480 24734 27532
rect 26513 27523 26571 27529
rect 26513 27489 26525 27523
rect 26559 27520 26571 27523
rect 27062 27520 27068 27532
rect 26559 27492 27068 27520
rect 26559 27489 26571 27492
rect 26513 27483 26571 27489
rect 27062 27480 27068 27492
rect 27120 27480 27126 27532
rect 27525 27523 27583 27529
rect 27525 27489 27537 27523
rect 27571 27520 27583 27523
rect 28074 27520 28080 27532
rect 27571 27492 28080 27520
rect 27571 27489 27583 27492
rect 27525 27483 27583 27489
rect 28074 27480 28080 27492
rect 28132 27480 28138 27532
rect 28258 27480 28264 27532
rect 28316 27520 28322 27532
rect 28353 27523 28411 27529
rect 28353 27520 28365 27523
rect 28316 27492 28365 27520
rect 28316 27480 28322 27492
rect 28353 27489 28365 27492
rect 28399 27489 28411 27523
rect 28353 27483 28411 27489
rect 23658 27452 23664 27464
rect 23584 27424 23664 27452
rect 23658 27412 23664 27424
rect 23716 27412 23722 27464
rect 24118 27412 24124 27464
rect 24176 27452 24182 27464
rect 24765 27455 24823 27461
rect 24765 27452 24777 27455
rect 24176 27424 24777 27452
rect 24176 27412 24182 27424
rect 24765 27421 24777 27424
rect 24811 27421 24823 27455
rect 24765 27415 24823 27421
rect 25409 27387 25467 27393
rect 25409 27384 25421 27387
rect 22664 27356 25421 27384
rect 25409 27353 25421 27356
rect 25455 27353 25467 27387
rect 25409 27347 25467 27353
rect 16850 27316 16856 27328
rect 13596 27288 14228 27316
rect 16811 27288 16856 27316
rect 13596 27276 13602 27288
rect 16850 27276 16856 27288
rect 16908 27276 16914 27328
rect 19242 27316 19248 27328
rect 19203 27288 19248 27316
rect 19242 27276 19248 27288
rect 19300 27276 19306 27328
rect 19613 27319 19671 27325
rect 19613 27285 19625 27319
rect 19659 27316 19671 27319
rect 20898 27316 20904 27328
rect 19659 27288 20904 27316
rect 19659 27285 19671 27288
rect 19613 27279 19671 27285
rect 20898 27276 20904 27288
rect 20956 27276 20962 27328
rect 21542 27316 21548 27328
rect 21503 27288 21548 27316
rect 21542 27276 21548 27288
rect 21600 27276 21606 27328
rect 22097 27319 22155 27325
rect 22097 27285 22109 27319
rect 22143 27316 22155 27319
rect 22278 27316 22284 27328
rect 22143 27288 22284 27316
rect 22143 27285 22155 27288
rect 22097 27279 22155 27285
rect 22278 27276 22284 27288
rect 22336 27276 22342 27328
rect 22462 27316 22468 27328
rect 22375 27288 22468 27316
rect 22462 27276 22468 27288
rect 22520 27316 22526 27328
rect 22603 27319 22661 27325
rect 22603 27316 22615 27319
rect 22520 27288 22615 27316
rect 22520 27276 22526 27288
rect 22603 27285 22615 27288
rect 22649 27285 22661 27319
rect 22738 27316 22744 27328
rect 22699 27288 22744 27316
rect 22603 27279 22661 27285
rect 22738 27276 22744 27288
rect 22796 27276 22802 27328
rect 23842 27316 23848 27328
rect 23803 27288 23848 27316
rect 23842 27276 23848 27288
rect 23900 27276 23906 27328
rect 24854 27276 24860 27328
rect 24912 27316 24918 27328
rect 25041 27319 25099 27325
rect 25041 27316 25053 27319
rect 24912 27288 25053 27316
rect 24912 27276 24918 27288
rect 25041 27285 25053 27288
rect 25087 27285 25099 27319
rect 25041 27279 25099 27285
rect 25314 27276 25320 27328
rect 25372 27316 25378 27328
rect 27709 27319 27767 27325
rect 27709 27316 27721 27319
rect 25372 27288 27721 27316
rect 25372 27276 25378 27288
rect 27709 27285 27721 27288
rect 27755 27285 27767 27319
rect 27709 27279 27767 27285
rect 27798 27276 27804 27328
rect 27856 27316 27862 27328
rect 27985 27319 28043 27325
rect 27985 27316 27997 27319
rect 27856 27288 27997 27316
rect 27856 27276 27862 27288
rect 27985 27285 27997 27288
rect 28031 27285 28043 27319
rect 27985 27279 28043 27285
rect 1104 27226 38824 27248
rect 1104 27174 4246 27226
rect 4298 27174 4310 27226
rect 4362 27174 4374 27226
rect 4426 27174 4438 27226
rect 4490 27174 34966 27226
rect 35018 27174 35030 27226
rect 35082 27174 35094 27226
rect 35146 27174 35158 27226
rect 35210 27174 38824 27226
rect 1104 27152 38824 27174
rect 6914 27072 6920 27124
rect 6972 27112 6978 27124
rect 7377 27115 7435 27121
rect 7377 27112 7389 27115
rect 6972 27084 7389 27112
rect 6972 27072 6978 27084
rect 7377 27081 7389 27084
rect 7423 27081 7435 27115
rect 7377 27075 7435 27081
rect 9493 27115 9551 27121
rect 9493 27081 9505 27115
rect 9539 27112 9551 27115
rect 9582 27112 9588 27124
rect 9539 27084 9588 27112
rect 9539 27081 9551 27084
rect 9493 27075 9551 27081
rect 9582 27072 9588 27084
rect 9640 27072 9646 27124
rect 14642 27112 14648 27124
rect 14603 27084 14648 27112
rect 14642 27072 14648 27084
rect 14700 27072 14706 27124
rect 15654 27072 15660 27124
rect 15712 27112 15718 27124
rect 15712 27084 15792 27112
rect 15712 27072 15718 27084
rect 9217 27047 9275 27053
rect 9217 27013 9229 27047
rect 9263 27044 9275 27047
rect 9263 27016 11100 27044
rect 9263 27013 9275 27016
rect 9217 27007 9275 27013
rect 1854 26976 1860 26988
rect 1815 26948 1860 26976
rect 1854 26936 1860 26948
rect 1912 26936 1918 26988
rect 10410 26976 10416 26988
rect 10371 26948 10416 26976
rect 10410 26936 10416 26948
rect 10468 26936 10474 26988
rect 10870 26976 10876 26988
rect 10831 26948 10876 26976
rect 10870 26936 10876 26948
rect 10928 26936 10934 26988
rect 1581 26911 1639 26917
rect 1581 26877 1593 26911
rect 1627 26908 1639 26911
rect 1670 26908 1676 26920
rect 1627 26880 1676 26908
rect 1627 26877 1639 26880
rect 1581 26871 1639 26877
rect 1670 26868 1676 26880
rect 1728 26868 1734 26920
rect 8297 26911 8355 26917
rect 8297 26877 8309 26911
rect 8343 26908 8355 26911
rect 9309 26911 9367 26917
rect 8343 26880 8708 26908
rect 8343 26877 8355 26880
rect 8297 26871 8355 26877
rect 8680 26852 8708 26880
rect 9309 26877 9321 26911
rect 9355 26908 9367 26911
rect 9355 26880 9904 26908
rect 9355 26877 9367 26880
rect 9309 26871 9367 26877
rect 3237 26843 3295 26849
rect 3237 26809 3249 26843
rect 3283 26840 3295 26843
rect 4062 26840 4068 26852
rect 3283 26812 4068 26840
rect 3283 26809 3295 26812
rect 3237 26803 3295 26809
rect 4062 26800 4068 26812
rect 4120 26800 4126 26852
rect 8662 26800 8668 26852
rect 8720 26840 8726 26852
rect 8849 26843 8907 26849
rect 8849 26840 8861 26843
rect 8720 26812 8861 26840
rect 8720 26800 8726 26812
rect 8849 26809 8861 26812
rect 8895 26840 8907 26843
rect 9766 26840 9772 26852
rect 8895 26812 9772 26840
rect 8895 26809 8907 26812
rect 8849 26803 8907 26809
rect 9766 26800 9772 26812
rect 9824 26800 9830 26852
rect 9876 26784 9904 26880
rect 10134 26868 10140 26920
rect 10192 26908 10198 26920
rect 10962 26908 10968 26920
rect 10192 26880 10968 26908
rect 10192 26868 10198 26880
rect 10962 26868 10968 26880
rect 11020 26868 11026 26920
rect 11072 26908 11100 27016
rect 11698 27004 11704 27056
rect 11756 27044 11762 27056
rect 11793 27047 11851 27053
rect 11793 27044 11805 27047
rect 11756 27016 11805 27044
rect 11756 27004 11762 27016
rect 11793 27013 11805 27016
rect 11839 27013 11851 27047
rect 12250 27044 12256 27056
rect 12163 27016 12256 27044
rect 11793 27007 11851 27013
rect 12250 27004 12256 27016
rect 12308 27044 12314 27056
rect 15102 27044 15108 27056
rect 12308 27016 15108 27044
rect 12308 27004 12314 27016
rect 15102 27004 15108 27016
rect 15160 27004 15166 27056
rect 15764 27044 15792 27084
rect 15838 27072 15844 27124
rect 15896 27112 15902 27124
rect 16025 27115 16083 27121
rect 16025 27112 16037 27115
rect 15896 27084 16037 27112
rect 15896 27072 15902 27084
rect 16025 27081 16037 27084
rect 16071 27081 16083 27115
rect 16025 27075 16083 27081
rect 16206 27072 16212 27124
rect 16264 27112 16270 27124
rect 16393 27115 16451 27121
rect 16393 27112 16405 27115
rect 16264 27084 16405 27112
rect 16264 27072 16270 27084
rect 16393 27081 16405 27084
rect 16439 27081 16451 27115
rect 16393 27075 16451 27081
rect 16758 27072 16764 27124
rect 16816 27112 16822 27124
rect 16853 27115 16911 27121
rect 16853 27112 16865 27115
rect 16816 27084 16865 27112
rect 16816 27072 16822 27084
rect 16853 27081 16865 27084
rect 16899 27081 16911 27115
rect 16853 27075 16911 27081
rect 17402 27072 17408 27124
rect 17460 27112 17466 27124
rect 17773 27115 17831 27121
rect 17773 27112 17785 27115
rect 17460 27084 17785 27112
rect 17460 27072 17466 27084
rect 17773 27081 17785 27084
rect 17819 27081 17831 27115
rect 18782 27112 18788 27124
rect 18743 27084 18788 27112
rect 17773 27075 17831 27081
rect 18782 27072 18788 27084
rect 18840 27072 18846 27124
rect 21082 27072 21088 27124
rect 21140 27112 21146 27124
rect 22925 27115 22983 27121
rect 22925 27112 22937 27115
rect 21140 27084 22937 27112
rect 21140 27072 21146 27084
rect 22925 27081 22937 27084
rect 22971 27081 22983 27115
rect 22925 27075 22983 27081
rect 23032 27084 24072 27112
rect 17586 27044 17592 27056
rect 15764 27016 17592 27044
rect 17586 27004 17592 27016
rect 17644 27004 17650 27056
rect 18417 27047 18475 27053
rect 18417 27013 18429 27047
rect 18463 27044 18475 27047
rect 22373 27047 22431 27053
rect 18463 27016 20392 27044
rect 18463 27013 18475 27016
rect 18417 27007 18475 27013
rect 11882 26936 11888 26988
rect 11940 26976 11946 26988
rect 13587 26979 13645 26985
rect 13587 26976 13599 26979
rect 11940 26948 13599 26976
rect 11940 26936 11946 26948
rect 13587 26945 13599 26948
rect 13633 26945 13645 26979
rect 13587 26939 13645 26945
rect 14458 26936 14464 26988
rect 14516 26976 14522 26988
rect 14918 26976 14924 26988
rect 14516 26948 14924 26976
rect 14516 26936 14522 26948
rect 14918 26936 14924 26948
rect 14976 26976 14982 26988
rect 16574 26976 16580 26988
rect 14976 26948 15608 26976
rect 16535 26948 16580 26976
rect 14976 26936 14982 26948
rect 11238 26908 11244 26920
rect 11072 26880 11244 26908
rect 11238 26868 11244 26880
rect 11296 26908 11302 26920
rect 11333 26911 11391 26917
rect 11333 26908 11345 26911
rect 11296 26880 11345 26908
rect 11296 26868 11302 26880
rect 11333 26877 11345 26880
rect 11379 26877 11391 26911
rect 11333 26871 11391 26877
rect 11425 26911 11483 26917
rect 11425 26877 11437 26911
rect 11471 26877 11483 26911
rect 11425 26871 11483 26877
rect 10318 26800 10324 26852
rect 10376 26840 10382 26852
rect 11440 26840 11468 26871
rect 12802 26868 12808 26920
rect 12860 26908 12866 26920
rect 12897 26911 12955 26917
rect 12897 26908 12909 26911
rect 12860 26880 12909 26908
rect 12860 26868 12866 26880
rect 12897 26877 12909 26880
rect 12943 26877 12955 26911
rect 12897 26871 12955 26877
rect 13354 26868 13360 26920
rect 13412 26908 13418 26920
rect 13449 26911 13507 26917
rect 13449 26908 13461 26911
rect 13412 26880 13461 26908
rect 13412 26868 13418 26880
rect 13449 26877 13461 26880
rect 13495 26877 13507 26911
rect 13722 26908 13728 26920
rect 13683 26880 13728 26908
rect 13449 26871 13507 26877
rect 13722 26868 13728 26880
rect 13780 26908 13786 26920
rect 15580 26917 15608 26948
rect 16574 26936 16580 26948
rect 16632 26936 16638 26988
rect 20254 26976 20260 26988
rect 20215 26948 20260 26976
rect 20254 26936 20260 26948
rect 20312 26936 20318 26988
rect 20364 26920 20392 27016
rect 22373 27013 22385 27047
rect 22419 27044 22431 27047
rect 23032 27044 23060 27084
rect 22419 27016 23060 27044
rect 23477 27047 23535 27053
rect 22419 27013 22431 27016
rect 22373 27007 22431 27013
rect 23477 27013 23489 27047
rect 23523 27044 23535 27047
rect 23934 27044 23940 27056
rect 23523 27016 23796 27044
rect 23895 27016 23940 27044
rect 23523 27013 23535 27016
rect 23477 27007 23535 27013
rect 20622 26936 20628 26988
rect 20680 26936 20686 26988
rect 20898 26936 20904 26988
rect 20956 26976 20962 26988
rect 21082 26976 21088 26988
rect 20956 26948 21088 26976
rect 20956 26936 20962 26948
rect 21082 26936 21088 26948
rect 21140 26936 21146 26988
rect 23382 26976 23388 26988
rect 23216 26948 23388 26976
rect 14737 26911 14795 26917
rect 14737 26908 14749 26911
rect 13780 26880 14749 26908
rect 13780 26868 13786 26880
rect 14737 26877 14749 26880
rect 14783 26877 14795 26911
rect 14737 26871 14795 26877
rect 15197 26911 15255 26917
rect 15197 26877 15209 26911
rect 15243 26877 15255 26911
rect 15197 26871 15255 26877
rect 15565 26911 15623 26917
rect 15565 26877 15577 26911
rect 15611 26877 15623 26911
rect 15565 26871 15623 26877
rect 11606 26840 11612 26852
rect 10376 26812 11612 26840
rect 10376 26800 10382 26812
rect 11606 26800 11612 26812
rect 11664 26800 11670 26852
rect 15212 26840 15240 26871
rect 15654 26868 15660 26920
rect 15712 26908 15718 26920
rect 16390 26908 16396 26920
rect 15712 26880 16396 26908
rect 15712 26868 15718 26880
rect 16390 26868 16396 26880
rect 16448 26868 16454 26920
rect 16666 26908 16672 26920
rect 16627 26880 16672 26908
rect 16666 26868 16672 26880
rect 16724 26908 16730 26920
rect 17405 26911 17463 26917
rect 17405 26908 17417 26911
rect 16724 26880 17417 26908
rect 16724 26868 16730 26880
rect 17405 26877 17417 26880
rect 17451 26877 17463 26911
rect 17405 26871 17463 26877
rect 18233 26911 18291 26917
rect 18233 26877 18245 26911
rect 18279 26908 18291 26911
rect 18782 26908 18788 26920
rect 18279 26880 18788 26908
rect 18279 26877 18291 26880
rect 18233 26871 18291 26877
rect 18782 26868 18788 26880
rect 18840 26868 18846 26920
rect 19426 26908 19432 26920
rect 19387 26880 19432 26908
rect 19426 26868 19432 26880
rect 19484 26868 19490 26920
rect 19613 26911 19671 26917
rect 19613 26877 19625 26911
rect 19659 26877 19671 26911
rect 19978 26908 19984 26920
rect 19939 26880 19984 26908
rect 19613 26871 19671 26877
rect 14752 26812 15240 26840
rect 14752 26784 14780 26812
rect 7098 26772 7104 26784
rect 7059 26744 7104 26772
rect 7098 26732 7104 26744
rect 7156 26732 7162 26784
rect 8478 26772 8484 26784
rect 8439 26744 8484 26772
rect 8478 26732 8484 26744
rect 8536 26732 8542 26784
rect 9858 26772 9864 26784
rect 9819 26744 9864 26772
rect 9858 26732 9864 26744
rect 9916 26732 9922 26784
rect 9950 26732 9956 26784
rect 10008 26772 10014 26784
rect 10229 26775 10287 26781
rect 10229 26772 10241 26775
rect 10008 26744 10241 26772
rect 10008 26732 10014 26744
rect 10229 26741 10241 26744
rect 10275 26772 10287 26775
rect 10594 26772 10600 26784
rect 10275 26744 10600 26772
rect 10275 26741 10287 26744
rect 10229 26735 10287 26741
rect 10594 26732 10600 26744
rect 10652 26772 10658 26784
rect 10962 26772 10968 26784
rect 10652 26744 10968 26772
rect 10652 26732 10658 26744
rect 10962 26732 10968 26744
rect 11020 26732 11026 26784
rect 12805 26775 12863 26781
rect 12805 26741 12817 26775
rect 12851 26772 12863 26775
rect 13170 26772 13176 26784
rect 12851 26744 13176 26772
rect 12851 26741 12863 26744
rect 12805 26735 12863 26741
rect 13170 26732 13176 26744
rect 13228 26772 13234 26784
rect 13814 26772 13820 26784
rect 13228 26744 13820 26772
rect 13228 26732 13234 26744
rect 13814 26732 13820 26744
rect 13872 26732 13878 26784
rect 14277 26775 14335 26781
rect 14277 26741 14289 26775
rect 14323 26772 14335 26775
rect 14734 26772 14740 26784
rect 14323 26744 14740 26772
rect 14323 26741 14335 26744
rect 14277 26735 14335 26741
rect 14734 26732 14740 26744
rect 14792 26732 14798 26784
rect 18874 26732 18880 26784
rect 18932 26772 18938 26784
rect 19061 26775 19119 26781
rect 19061 26772 19073 26775
rect 18932 26744 19073 26772
rect 18932 26732 18938 26744
rect 19061 26741 19073 26744
rect 19107 26772 19119 26775
rect 19628 26772 19656 26871
rect 19978 26868 19984 26880
rect 20036 26868 20042 26920
rect 20346 26868 20352 26920
rect 20404 26908 20410 26920
rect 20533 26911 20591 26917
rect 20533 26908 20545 26911
rect 20404 26880 20545 26908
rect 20404 26868 20410 26880
rect 20533 26877 20545 26880
rect 20579 26908 20591 26911
rect 20640 26908 20668 26936
rect 20579 26880 20668 26908
rect 20993 26911 21051 26917
rect 20579 26877 20591 26880
rect 20533 26871 20591 26877
rect 20993 26877 21005 26911
rect 21039 26908 21051 26911
rect 21450 26908 21456 26920
rect 21039 26880 21456 26908
rect 21039 26877 21051 26880
rect 20993 26871 21051 26877
rect 19996 26840 20024 26868
rect 20622 26840 20628 26852
rect 19996 26812 20628 26840
rect 20622 26800 20628 26812
rect 20680 26800 20686 26852
rect 20898 26800 20904 26852
rect 20956 26840 20962 26852
rect 21008 26840 21036 26871
rect 21450 26868 21456 26880
rect 21508 26908 21514 26920
rect 21508 26880 21772 26908
rect 21508 26868 21514 26880
rect 20956 26812 21036 26840
rect 21545 26843 21603 26849
rect 20956 26800 20962 26812
rect 21545 26809 21557 26843
rect 21591 26809 21603 26843
rect 21744 26840 21772 26880
rect 21928 26880 22600 26908
rect 21928 26849 21956 26880
rect 21821 26843 21879 26849
rect 21821 26840 21833 26843
rect 21744 26812 21833 26840
rect 21545 26803 21603 26809
rect 21821 26809 21833 26812
rect 21867 26809 21879 26843
rect 21821 26803 21879 26809
rect 21913 26843 21971 26849
rect 21913 26809 21925 26843
rect 21959 26809 21971 26843
rect 22278 26840 22284 26852
rect 22239 26812 22284 26840
rect 21913 26803 21971 26809
rect 20806 26772 20812 26784
rect 19107 26744 20812 26772
rect 19107 26741 19119 26744
rect 19061 26735 19119 26741
rect 20806 26732 20812 26744
rect 20864 26732 20870 26784
rect 21174 26732 21180 26784
rect 21232 26772 21238 26784
rect 21361 26775 21419 26781
rect 21361 26772 21373 26775
rect 21232 26744 21373 26772
rect 21232 26732 21238 26744
rect 21361 26741 21373 26744
rect 21407 26772 21419 26775
rect 21560 26772 21588 26803
rect 22278 26800 22284 26812
rect 22336 26800 22342 26852
rect 21726 26772 21732 26784
rect 21407 26744 21588 26772
rect 21639 26744 21732 26772
rect 21407 26741 21419 26744
rect 21361 26735 21419 26741
rect 21726 26732 21732 26744
rect 21784 26772 21790 26784
rect 22094 26772 22100 26784
rect 21784 26744 22100 26772
rect 21784 26732 21790 26744
rect 22094 26732 22100 26744
rect 22152 26772 22158 26784
rect 22373 26775 22431 26781
rect 22373 26772 22385 26775
rect 22152 26744 22385 26772
rect 22152 26732 22158 26744
rect 22373 26741 22385 26744
rect 22419 26741 22431 26775
rect 22572 26772 22600 26880
rect 22649 26843 22707 26849
rect 22649 26809 22661 26843
rect 22695 26840 22707 26843
rect 23216 26840 23244 26948
rect 23382 26936 23388 26948
rect 23440 26936 23446 26988
rect 23768 26976 23796 27016
rect 23934 27004 23940 27016
rect 23992 27004 23998 27056
rect 24044 27044 24072 27084
rect 25038 27072 25044 27124
rect 25096 27112 25102 27124
rect 25409 27115 25467 27121
rect 25409 27112 25421 27115
rect 25096 27084 25421 27112
rect 25096 27072 25102 27084
rect 25409 27081 25421 27084
rect 25455 27081 25467 27115
rect 25409 27075 25467 27081
rect 25777 27115 25835 27121
rect 25777 27081 25789 27115
rect 25823 27112 25835 27115
rect 25866 27112 25872 27124
rect 25823 27084 25872 27112
rect 25823 27081 25835 27084
rect 25777 27075 25835 27081
rect 25866 27072 25872 27084
rect 25924 27072 25930 27124
rect 26050 27112 26056 27124
rect 26011 27084 26056 27112
rect 26050 27072 26056 27084
rect 26108 27072 26114 27124
rect 27062 27112 27068 27124
rect 27023 27084 27068 27112
rect 27062 27072 27068 27084
rect 27120 27072 27126 27124
rect 28350 27072 28356 27124
rect 28408 27112 28414 27124
rect 28445 27115 28503 27121
rect 28445 27112 28457 27115
rect 28408 27084 28457 27112
rect 28408 27072 28414 27084
rect 28445 27081 28457 27084
rect 28491 27112 28503 27115
rect 28718 27112 28724 27124
rect 28491 27084 28724 27112
rect 28491 27081 28503 27084
rect 28445 27075 28503 27081
rect 28718 27072 28724 27084
rect 28776 27072 28782 27124
rect 25314 27044 25320 27056
rect 24044 27016 25320 27044
rect 25314 27004 25320 27016
rect 25372 27004 25378 27056
rect 24029 26979 24087 26985
rect 24029 26976 24041 26979
rect 23768 26948 24041 26976
rect 24029 26945 24041 26948
rect 24075 26976 24087 26979
rect 24302 26976 24308 26988
rect 24075 26948 24308 26976
rect 24075 26945 24087 26948
rect 24029 26939 24087 26945
rect 24302 26936 24308 26948
rect 24360 26976 24366 26988
rect 27080 26976 27108 27072
rect 24360 26948 27108 26976
rect 24360 26936 24366 26948
rect 23290 26868 23296 26920
rect 23348 26908 23354 26920
rect 23661 26911 23719 26917
rect 23661 26908 23673 26911
rect 23348 26880 23673 26908
rect 23348 26868 23354 26880
rect 23661 26877 23673 26880
rect 23707 26877 23719 26911
rect 23661 26871 23719 26877
rect 23808 26911 23866 26917
rect 23808 26877 23820 26911
rect 23854 26908 23866 26911
rect 24670 26908 24676 26920
rect 23854 26880 24676 26908
rect 23854 26877 23866 26880
rect 23808 26871 23866 26877
rect 24670 26868 24676 26880
rect 24728 26868 24734 26920
rect 25225 26911 25283 26917
rect 25225 26877 25237 26911
rect 25271 26908 25283 26911
rect 25866 26908 25872 26920
rect 25271 26880 25872 26908
rect 25271 26877 25283 26880
rect 25225 26871 25283 26877
rect 25866 26868 25872 26880
rect 25924 26868 25930 26920
rect 26237 26911 26295 26917
rect 26237 26877 26249 26911
rect 26283 26877 26295 26911
rect 26237 26871 26295 26877
rect 22695 26812 23244 26840
rect 22695 26809 22707 26812
rect 22649 26803 22707 26809
rect 24026 26800 24032 26852
rect 24084 26840 24090 26852
rect 25041 26843 25099 26849
rect 25041 26840 25053 26843
rect 24084 26812 25053 26840
rect 24084 26800 24090 26812
rect 25041 26809 25053 26812
rect 25087 26809 25099 26843
rect 26252 26840 26280 26871
rect 26694 26868 26700 26920
rect 26752 26908 26758 26920
rect 27062 26908 27068 26920
rect 26752 26880 27068 26908
rect 26752 26868 26758 26880
rect 27062 26868 27068 26880
rect 27120 26868 27126 26920
rect 27249 26911 27307 26917
rect 27249 26877 27261 26911
rect 27295 26908 27307 26911
rect 27709 26911 27767 26917
rect 27709 26908 27721 26911
rect 27295 26880 27721 26908
rect 27295 26877 27307 26880
rect 27249 26871 27307 26877
rect 27709 26877 27721 26880
rect 27755 26877 27767 26911
rect 28074 26908 28080 26920
rect 28035 26880 28080 26908
rect 27709 26871 27767 26877
rect 26252 26812 26740 26840
rect 25041 26803 25099 26809
rect 26712 26784 26740 26812
rect 26786 26800 26792 26852
rect 26844 26840 26850 26852
rect 27264 26840 27292 26871
rect 28074 26868 28080 26880
rect 28132 26868 28138 26920
rect 26844 26812 27292 26840
rect 26844 26800 26850 26812
rect 23474 26772 23480 26784
rect 22572 26744 23480 26772
rect 22373 26735 22431 26741
rect 23474 26732 23480 26744
rect 23532 26732 23538 26784
rect 24302 26772 24308 26784
rect 24263 26744 24308 26772
rect 24302 26732 24308 26744
rect 24360 26732 24366 26784
rect 24762 26772 24768 26784
rect 24675 26744 24768 26772
rect 24762 26732 24768 26744
rect 24820 26772 24826 26784
rect 25866 26772 25872 26784
rect 24820 26744 25872 26772
rect 24820 26732 24826 26744
rect 25866 26732 25872 26744
rect 25924 26732 25930 26784
rect 26234 26732 26240 26784
rect 26292 26772 26298 26784
rect 26421 26775 26479 26781
rect 26421 26772 26433 26775
rect 26292 26744 26433 26772
rect 26292 26732 26298 26744
rect 26421 26741 26433 26744
rect 26467 26741 26479 26775
rect 26694 26772 26700 26784
rect 26655 26744 26700 26772
rect 26421 26735 26479 26741
rect 26694 26732 26700 26744
rect 26752 26732 26758 26784
rect 27246 26732 27252 26784
rect 27304 26772 27310 26784
rect 27433 26775 27491 26781
rect 27433 26772 27445 26775
rect 27304 26744 27445 26772
rect 27304 26732 27310 26744
rect 27433 26741 27445 26744
rect 27479 26741 27491 26775
rect 27433 26735 27491 26741
rect 1104 26682 38824 26704
rect 1104 26630 19606 26682
rect 19658 26630 19670 26682
rect 19722 26630 19734 26682
rect 19786 26630 19798 26682
rect 19850 26630 38824 26682
rect 1104 26608 38824 26630
rect 1673 26571 1731 26577
rect 1673 26537 1685 26571
rect 1719 26568 1731 26571
rect 1854 26568 1860 26580
rect 1719 26540 1860 26568
rect 1719 26537 1731 26540
rect 1673 26531 1731 26537
rect 1854 26528 1860 26540
rect 1912 26528 1918 26580
rect 7374 26528 7380 26580
rect 7432 26568 7438 26580
rect 7469 26571 7527 26577
rect 7469 26568 7481 26571
rect 7432 26540 7481 26568
rect 7432 26528 7438 26540
rect 7469 26537 7481 26540
rect 7515 26537 7527 26571
rect 7469 26531 7527 26537
rect 10045 26571 10103 26577
rect 10045 26537 10057 26571
rect 10091 26568 10103 26571
rect 10134 26568 10140 26580
rect 10091 26540 10140 26568
rect 10091 26537 10103 26540
rect 10045 26531 10103 26537
rect 10134 26528 10140 26540
rect 10192 26528 10198 26580
rect 11238 26528 11244 26580
rect 11296 26568 11302 26580
rect 11885 26571 11943 26577
rect 11885 26568 11897 26571
rect 11296 26540 11897 26568
rect 11296 26528 11302 26540
rect 11885 26537 11897 26540
rect 11931 26537 11943 26571
rect 11885 26531 11943 26537
rect 13081 26571 13139 26577
rect 13081 26537 13093 26571
rect 13127 26568 13139 26571
rect 13446 26568 13452 26580
rect 13127 26540 13452 26568
rect 13127 26537 13139 26540
rect 13081 26531 13139 26537
rect 13446 26528 13452 26540
rect 13504 26528 13510 26580
rect 14642 26568 14648 26580
rect 14603 26540 14648 26568
rect 14642 26528 14648 26540
rect 14700 26568 14706 26580
rect 16114 26568 16120 26580
rect 14700 26540 16120 26568
rect 14700 26528 14706 26540
rect 16114 26528 16120 26540
rect 16172 26568 16178 26580
rect 16393 26571 16451 26577
rect 16393 26568 16405 26571
rect 16172 26540 16405 26568
rect 16172 26528 16178 26540
rect 16393 26537 16405 26540
rect 16439 26537 16451 26571
rect 16393 26531 16451 26537
rect 16666 26528 16672 26580
rect 16724 26568 16730 26580
rect 17218 26568 17224 26580
rect 16724 26540 17224 26568
rect 16724 26528 16730 26540
rect 17218 26528 17224 26540
rect 17276 26528 17282 26580
rect 18506 26528 18512 26580
rect 18564 26568 18570 26580
rect 20349 26571 20407 26577
rect 18564 26540 19288 26568
rect 18564 26528 18570 26540
rect 13262 26460 13268 26512
rect 13320 26500 13326 26512
rect 13357 26503 13415 26509
rect 13357 26500 13369 26503
rect 13320 26472 13369 26500
rect 13320 26460 13326 26472
rect 13357 26469 13369 26472
rect 13403 26469 13415 26503
rect 14734 26500 14740 26512
rect 13357 26463 13415 26469
rect 13740 26472 14740 26500
rect 1670 26392 1676 26444
rect 1728 26432 1734 26444
rect 1949 26435 2007 26441
rect 1949 26432 1961 26435
rect 1728 26404 1961 26432
rect 1728 26392 1734 26404
rect 1949 26401 1961 26404
rect 1995 26432 2007 26435
rect 2038 26432 2044 26444
rect 1995 26404 2044 26432
rect 1995 26401 2007 26404
rect 1949 26395 2007 26401
rect 2038 26392 2044 26404
rect 2096 26432 2102 26444
rect 2774 26432 2780 26444
rect 2096 26404 2780 26432
rect 2096 26392 2102 26404
rect 2774 26392 2780 26404
rect 2832 26432 2838 26444
rect 5994 26432 6000 26444
rect 2832 26404 6000 26432
rect 2832 26392 2838 26404
rect 5994 26392 6000 26404
rect 6052 26432 6058 26444
rect 6089 26435 6147 26441
rect 6089 26432 6101 26435
rect 6052 26404 6101 26432
rect 6052 26392 6058 26404
rect 6089 26401 6101 26404
rect 6135 26401 6147 26435
rect 6089 26395 6147 26401
rect 6178 26392 6184 26444
rect 6236 26432 6242 26444
rect 6365 26435 6423 26441
rect 6365 26432 6377 26435
rect 6236 26404 6377 26432
rect 6236 26392 6242 26404
rect 6365 26401 6377 26404
rect 6411 26401 6423 26435
rect 6365 26395 6423 26401
rect 8573 26435 8631 26441
rect 8573 26401 8585 26435
rect 8619 26432 8631 26435
rect 8662 26432 8668 26444
rect 8619 26404 8668 26432
rect 8619 26401 8631 26404
rect 8573 26395 8631 26401
rect 8662 26392 8668 26404
rect 8720 26392 8726 26444
rect 9125 26435 9183 26441
rect 9125 26401 9137 26435
rect 9171 26432 9183 26435
rect 9490 26432 9496 26444
rect 9171 26404 9496 26432
rect 9171 26401 9183 26404
rect 9125 26395 9183 26401
rect 9490 26392 9496 26404
rect 9548 26432 9554 26444
rect 10781 26435 10839 26441
rect 10781 26432 10793 26435
rect 9548 26404 10793 26432
rect 9548 26392 9554 26404
rect 10781 26401 10793 26404
rect 10827 26432 10839 26435
rect 10870 26432 10876 26444
rect 10827 26404 10876 26432
rect 10827 26401 10839 26404
rect 10781 26395 10839 26401
rect 10870 26392 10876 26404
rect 10928 26392 10934 26444
rect 12529 26435 12587 26441
rect 12529 26401 12541 26435
rect 12575 26432 12587 26435
rect 12618 26432 12624 26444
rect 12575 26404 12624 26432
rect 12575 26401 12587 26404
rect 12529 26395 12587 26401
rect 12618 26392 12624 26404
rect 12676 26432 12682 26444
rect 13740 26432 13768 26472
rect 14734 26460 14740 26472
rect 14792 26460 14798 26512
rect 15102 26500 15108 26512
rect 15063 26472 15108 26500
rect 15102 26460 15108 26472
rect 15160 26460 15166 26512
rect 17310 26500 17316 26512
rect 15580 26472 17316 26500
rect 12676 26404 13768 26432
rect 12676 26392 12682 26404
rect 13814 26392 13820 26444
rect 13872 26432 13878 26444
rect 14185 26435 14243 26441
rect 14185 26432 14197 26435
rect 13872 26404 14197 26432
rect 13872 26392 13878 26404
rect 14185 26401 14197 26404
rect 14231 26401 14243 26435
rect 14185 26395 14243 26401
rect 14550 26392 14556 26444
rect 14608 26432 14614 26444
rect 15010 26432 15016 26444
rect 14608 26404 15016 26432
rect 14608 26392 14614 26404
rect 15010 26392 15016 26404
rect 15068 26392 15074 26444
rect 15286 26392 15292 26444
rect 15344 26432 15350 26444
rect 15580 26441 15608 26472
rect 17310 26460 17316 26472
rect 17368 26460 17374 26512
rect 18966 26500 18972 26512
rect 18879 26472 18972 26500
rect 18966 26460 18972 26472
rect 19024 26500 19030 26512
rect 19260 26509 19288 26540
rect 20349 26537 20361 26571
rect 20395 26568 20407 26571
rect 20438 26568 20444 26580
rect 20395 26540 20444 26568
rect 20395 26537 20407 26540
rect 20349 26531 20407 26537
rect 20438 26528 20444 26540
rect 20496 26528 20502 26580
rect 20717 26571 20775 26577
rect 20717 26537 20729 26571
rect 20763 26568 20775 26571
rect 21266 26568 21272 26580
rect 20763 26540 21272 26568
rect 20763 26537 20775 26540
rect 20717 26531 20775 26537
rect 21266 26528 21272 26540
rect 21324 26528 21330 26580
rect 21726 26528 21732 26580
rect 21784 26568 21790 26580
rect 21910 26568 21916 26580
rect 21784 26540 21916 26568
rect 21784 26528 21790 26540
rect 21910 26528 21916 26540
rect 21968 26528 21974 26580
rect 22373 26571 22431 26577
rect 22373 26537 22385 26571
rect 22419 26568 22431 26571
rect 22554 26568 22560 26580
rect 22419 26540 22560 26568
rect 22419 26537 22431 26540
rect 22373 26531 22431 26537
rect 22554 26528 22560 26540
rect 22612 26528 22618 26580
rect 23474 26528 23480 26580
rect 23532 26568 23538 26580
rect 23532 26540 24808 26568
rect 23532 26528 23538 26540
rect 19153 26503 19211 26509
rect 19153 26500 19165 26503
rect 19024 26472 19165 26500
rect 19024 26460 19030 26472
rect 19153 26469 19165 26472
rect 19199 26469 19211 26503
rect 19153 26463 19211 26469
rect 19245 26503 19303 26509
rect 19245 26469 19257 26503
rect 19291 26469 19303 26503
rect 19245 26463 19303 26469
rect 20806 26460 20812 26512
rect 20864 26500 20870 26512
rect 21174 26500 21180 26512
rect 20864 26472 21180 26500
rect 20864 26460 20870 26472
rect 21174 26460 21180 26472
rect 21232 26460 21238 26512
rect 21637 26503 21695 26509
rect 21637 26469 21649 26503
rect 21683 26500 21695 26503
rect 22002 26500 22008 26512
rect 21683 26472 22008 26500
rect 21683 26469 21695 26472
rect 21637 26463 21695 26469
rect 22002 26460 22008 26472
rect 22060 26460 22066 26512
rect 22465 26503 22523 26509
rect 22465 26469 22477 26503
rect 22511 26500 22523 26503
rect 22922 26500 22928 26512
rect 22511 26472 22928 26500
rect 22511 26469 22523 26472
rect 22465 26463 22523 26469
rect 22922 26460 22928 26472
rect 22980 26500 22986 26512
rect 23753 26503 23811 26509
rect 23753 26500 23765 26503
rect 22980 26472 23765 26500
rect 22980 26460 22986 26472
rect 23753 26469 23765 26472
rect 23799 26500 23811 26503
rect 23934 26500 23940 26512
rect 23799 26472 23940 26500
rect 23799 26469 23811 26472
rect 23753 26463 23811 26469
rect 23934 26460 23940 26472
rect 23992 26460 23998 26512
rect 24670 26500 24676 26512
rect 24412 26472 24676 26500
rect 15565 26435 15623 26441
rect 15565 26432 15577 26435
rect 15344 26404 15577 26432
rect 15344 26392 15350 26404
rect 15565 26401 15577 26404
rect 15611 26401 15623 26435
rect 16666 26432 16672 26444
rect 16627 26404 16672 26432
rect 15565 26395 15623 26401
rect 16666 26392 16672 26404
rect 16724 26392 16730 26444
rect 16850 26432 16856 26444
rect 16763 26404 16856 26432
rect 9674 26324 9680 26376
rect 9732 26364 9738 26376
rect 10502 26364 10508 26376
rect 9732 26336 10508 26364
rect 9732 26324 9738 26336
rect 10502 26324 10508 26336
rect 10560 26324 10566 26376
rect 13354 26324 13360 26376
rect 13412 26364 13418 26376
rect 13909 26367 13967 26373
rect 13909 26364 13921 26367
rect 13412 26336 13921 26364
rect 13412 26324 13418 26336
rect 13909 26333 13921 26336
rect 13955 26333 13967 26367
rect 13909 26327 13967 26333
rect 8757 26299 8815 26305
rect 8757 26265 8769 26299
rect 8803 26296 8815 26299
rect 10318 26296 10324 26308
rect 8803 26268 10324 26296
rect 8803 26265 8815 26268
rect 8757 26259 8815 26265
rect 10318 26256 10324 26268
rect 10376 26256 10382 26308
rect 13924 26296 13952 26327
rect 13998 26324 14004 26376
rect 14056 26364 14062 26376
rect 14369 26367 14427 26373
rect 14369 26364 14381 26367
rect 14056 26336 14381 26364
rect 14056 26324 14062 26336
rect 14369 26333 14381 26336
rect 14415 26333 14427 26367
rect 14369 26327 14427 26333
rect 16390 26324 16396 26376
rect 16448 26364 16454 26376
rect 16776 26364 16804 26404
rect 16850 26392 16856 26404
rect 16908 26432 16914 26444
rect 17405 26435 17463 26441
rect 17405 26432 17417 26435
rect 16908 26404 17417 26432
rect 16908 26392 16914 26404
rect 17405 26401 17417 26404
rect 17451 26401 17463 26435
rect 17586 26432 17592 26444
rect 17547 26404 17592 26432
rect 17405 26395 17463 26401
rect 17586 26392 17592 26404
rect 17644 26392 17650 26444
rect 18506 26392 18512 26444
rect 18564 26432 18570 26444
rect 18877 26435 18935 26441
rect 18877 26432 18889 26435
rect 18564 26404 18889 26432
rect 18564 26392 18570 26404
rect 18877 26401 18889 26404
rect 18923 26401 18935 26435
rect 18877 26395 18935 26401
rect 16448 26336 16804 26364
rect 16448 26324 16454 26336
rect 17310 26324 17316 26376
rect 17368 26364 17374 26376
rect 17770 26364 17776 26376
rect 17368 26336 17776 26364
rect 17368 26324 17374 26336
rect 17770 26324 17776 26336
rect 17828 26324 17834 26376
rect 18598 26324 18604 26376
rect 18656 26364 18662 26376
rect 18693 26367 18751 26373
rect 18693 26364 18705 26367
rect 18656 26336 18705 26364
rect 18656 26324 18662 26336
rect 18693 26333 18705 26336
rect 18739 26364 18751 26367
rect 18984 26364 19012 26460
rect 19061 26435 19119 26441
rect 19061 26401 19073 26435
rect 19107 26432 19119 26435
rect 19981 26435 20039 26441
rect 19107 26404 19932 26432
rect 19107 26401 19119 26404
rect 19061 26395 19119 26401
rect 18739 26336 19012 26364
rect 18739 26333 18751 26336
rect 18693 26327 18751 26333
rect 19242 26324 19248 26376
rect 19300 26364 19306 26376
rect 19610 26364 19616 26376
rect 19300 26336 19616 26364
rect 19300 26324 19306 26336
rect 19610 26324 19616 26336
rect 19668 26324 19674 26376
rect 19904 26364 19932 26404
rect 19981 26401 19993 26435
rect 20027 26432 20039 26435
rect 20346 26432 20352 26444
rect 20027 26404 20352 26432
rect 20027 26401 20039 26404
rect 19981 26395 20039 26401
rect 20346 26392 20352 26404
rect 20404 26392 20410 26444
rect 20901 26435 20959 26441
rect 20901 26401 20913 26435
rect 20947 26432 20959 26435
rect 21450 26432 21456 26444
rect 20947 26404 21456 26432
rect 20947 26401 20959 26404
rect 20901 26395 20959 26401
rect 21450 26392 21456 26404
rect 21508 26392 21514 26444
rect 22094 26432 22100 26444
rect 22020 26404 22100 26432
rect 20622 26364 20628 26376
rect 19904 26336 20628 26364
rect 20622 26324 20628 26336
rect 20680 26324 20686 26376
rect 21082 26373 21088 26376
rect 21048 26367 21088 26373
rect 21048 26333 21060 26367
rect 21048 26327 21088 26333
rect 21082 26324 21088 26327
rect 21140 26324 21146 26376
rect 21269 26367 21327 26373
rect 21269 26333 21281 26367
rect 21315 26364 21327 26367
rect 21910 26364 21916 26376
rect 21315 26336 21916 26364
rect 21315 26333 21327 26336
rect 21269 26327 21327 26333
rect 14550 26296 14556 26308
rect 13924 26268 14556 26296
rect 14550 26256 14556 26268
rect 14608 26256 14614 26308
rect 14734 26256 14740 26308
rect 14792 26296 14798 26308
rect 15102 26296 15108 26308
rect 14792 26268 15108 26296
rect 14792 26256 14798 26268
rect 15102 26256 15108 26268
rect 15160 26256 15166 26308
rect 15749 26299 15807 26305
rect 15749 26265 15761 26299
rect 15795 26296 15807 26299
rect 15838 26296 15844 26308
rect 15795 26268 15844 26296
rect 15795 26265 15807 26268
rect 15749 26259 15807 26265
rect 15838 26256 15844 26268
rect 15896 26256 15902 26308
rect 17218 26256 17224 26308
rect 17276 26296 17282 26308
rect 17405 26299 17463 26305
rect 17405 26296 17417 26299
rect 17276 26268 17417 26296
rect 17276 26256 17282 26268
rect 17405 26265 17417 26268
rect 17451 26265 17463 26299
rect 17405 26259 17463 26265
rect 17862 26256 17868 26308
rect 17920 26296 17926 26308
rect 18049 26299 18107 26305
rect 18049 26296 18061 26299
rect 17920 26268 18061 26296
rect 17920 26256 17926 26268
rect 18049 26265 18061 26268
rect 18095 26296 18107 26299
rect 18095 26268 19288 26296
rect 18095 26265 18107 26268
rect 18049 26259 18107 26265
rect 8202 26188 8208 26240
rect 8260 26228 8266 26240
rect 15562 26228 15568 26240
rect 8260 26200 15568 26228
rect 8260 26188 8266 26200
rect 15562 26188 15568 26200
rect 15620 26188 15626 26240
rect 16114 26228 16120 26240
rect 16075 26200 16120 26228
rect 16114 26188 16120 26200
rect 16172 26188 16178 26240
rect 18230 26188 18236 26240
rect 18288 26228 18294 26240
rect 18325 26231 18383 26237
rect 18325 26228 18337 26231
rect 18288 26200 18337 26228
rect 18288 26188 18294 26200
rect 18325 26197 18337 26200
rect 18371 26197 18383 26231
rect 19260 26228 19288 26268
rect 20898 26256 20904 26308
rect 20956 26296 20962 26308
rect 21174 26296 21180 26308
rect 20956 26268 21036 26296
rect 21135 26268 21180 26296
rect 20956 26256 20962 26268
rect 19334 26228 19340 26240
rect 19260 26200 19340 26228
rect 18325 26191 18383 26197
rect 19334 26188 19340 26200
rect 19392 26188 19398 26240
rect 21008 26228 21036 26268
rect 21174 26256 21180 26268
rect 21232 26256 21238 26308
rect 21284 26228 21312 26327
rect 21910 26324 21916 26336
rect 21968 26324 21974 26376
rect 22020 26373 22048 26404
rect 22094 26392 22100 26404
rect 22152 26392 22158 26444
rect 22612 26435 22670 26441
rect 22612 26401 22624 26435
rect 22658 26432 22670 26435
rect 24210 26432 24216 26444
rect 22658 26404 24216 26432
rect 22658 26401 22670 26404
rect 22612 26395 22670 26401
rect 24210 26392 24216 26404
rect 24268 26392 24274 26444
rect 24412 26441 24440 26472
rect 24670 26460 24676 26472
rect 24728 26460 24734 26512
rect 24780 26500 24808 26540
rect 25130 26528 25136 26580
rect 25188 26568 25194 26580
rect 25777 26571 25835 26577
rect 25777 26568 25789 26571
rect 25188 26540 25789 26568
rect 25188 26528 25194 26540
rect 25777 26537 25789 26540
rect 25823 26537 25835 26571
rect 25777 26531 25835 26537
rect 26418 26528 26424 26580
rect 26476 26568 26482 26580
rect 28077 26571 28135 26577
rect 26476 26540 27200 26568
rect 26476 26528 26482 26540
rect 25682 26500 25688 26512
rect 24780 26472 25688 26500
rect 25682 26460 25688 26472
rect 25740 26500 25746 26512
rect 26145 26503 26203 26509
rect 26145 26500 26157 26503
rect 25740 26472 26157 26500
rect 25740 26460 25746 26472
rect 26145 26469 26157 26472
rect 26191 26469 26203 26503
rect 26145 26463 26203 26469
rect 26252 26472 27108 26500
rect 24397 26435 24455 26441
rect 24397 26401 24409 26435
rect 24443 26401 24455 26435
rect 24397 26395 24455 26401
rect 24486 26392 24492 26444
rect 24544 26432 24550 26444
rect 26252 26432 26280 26472
rect 24544 26404 26280 26432
rect 26513 26435 26571 26441
rect 24544 26392 24550 26404
rect 26513 26401 26525 26435
rect 26559 26401 26571 26435
rect 26513 26395 26571 26401
rect 22005 26367 22063 26373
rect 22005 26333 22017 26367
rect 22051 26333 22063 26367
rect 22830 26364 22836 26376
rect 22791 26336 22836 26364
rect 22005 26327 22063 26333
rect 22830 26324 22836 26336
rect 22888 26324 22894 26376
rect 23474 26324 23480 26376
rect 23532 26364 23538 26376
rect 24029 26367 24087 26373
rect 24029 26364 24041 26367
rect 23532 26336 24041 26364
rect 23532 26324 23538 26336
rect 24029 26333 24041 26336
rect 24075 26364 24087 26367
rect 26528 26364 26556 26395
rect 26970 26364 26976 26376
rect 24075 26336 26976 26364
rect 24075 26333 24087 26336
rect 24029 26327 24087 26333
rect 26970 26324 26976 26336
rect 27028 26324 27034 26376
rect 27080 26373 27108 26472
rect 27172 26432 27200 26540
rect 28077 26537 28089 26571
rect 28123 26568 28135 26571
rect 28442 26568 28448 26580
rect 28123 26540 28448 26568
rect 28123 26537 28135 26540
rect 28077 26531 28135 26537
rect 28442 26528 28448 26540
rect 28500 26528 28506 26580
rect 27522 26432 27528 26444
rect 27172 26404 27528 26432
rect 27522 26392 27528 26404
rect 27580 26392 27586 26444
rect 27065 26367 27123 26373
rect 27065 26333 27077 26367
rect 27111 26364 27123 26367
rect 27433 26367 27491 26373
rect 27433 26364 27445 26367
rect 27111 26336 27445 26364
rect 27111 26333 27123 26336
rect 27065 26327 27123 26333
rect 27433 26333 27445 26336
rect 27479 26364 27491 26367
rect 27614 26364 27620 26376
rect 27479 26336 27620 26364
rect 27479 26333 27491 26336
rect 27433 26327 27491 26333
rect 27614 26324 27620 26336
rect 27672 26324 27678 26376
rect 22094 26256 22100 26308
rect 22152 26296 22158 26308
rect 22925 26299 22983 26305
rect 22925 26296 22937 26299
rect 22152 26268 22937 26296
rect 22152 26256 22158 26268
rect 22925 26265 22937 26268
rect 22971 26265 22983 26299
rect 24118 26296 24124 26308
rect 22925 26259 22983 26265
rect 23400 26268 24124 26296
rect 21008 26200 21312 26228
rect 22741 26231 22799 26237
rect 22741 26197 22753 26231
rect 22787 26228 22799 26231
rect 22830 26228 22836 26240
rect 22787 26200 22836 26228
rect 22787 26197 22799 26200
rect 22741 26191 22799 26197
rect 22830 26188 22836 26200
rect 22888 26188 22894 26240
rect 23290 26188 23296 26240
rect 23348 26228 23354 26240
rect 23400 26228 23428 26268
rect 24118 26256 24124 26268
rect 24176 26256 24182 26308
rect 25038 26296 25044 26308
rect 24999 26268 25044 26296
rect 25038 26256 25044 26268
rect 25096 26256 25102 26308
rect 25498 26296 25504 26308
rect 25459 26268 25504 26296
rect 25498 26256 25504 26268
rect 25556 26256 25562 26308
rect 25866 26256 25872 26308
rect 25924 26296 25930 26308
rect 27709 26299 27767 26305
rect 27709 26296 27721 26299
rect 25924 26268 27721 26296
rect 25924 26256 25930 26268
rect 27709 26265 27721 26268
rect 27755 26265 27767 26299
rect 27709 26259 27767 26265
rect 23348 26200 23428 26228
rect 23348 26188 23354 26200
rect 26050 26188 26056 26240
rect 26108 26228 26114 26240
rect 26697 26231 26755 26237
rect 26697 26228 26709 26231
rect 26108 26200 26709 26228
rect 26108 26188 26114 26200
rect 26697 26197 26709 26200
rect 26743 26197 26755 26231
rect 26697 26191 26755 26197
rect 1104 26138 38824 26160
rect 1104 26086 4246 26138
rect 4298 26086 4310 26138
rect 4362 26086 4374 26138
rect 4426 26086 4438 26138
rect 4490 26086 34966 26138
rect 35018 26086 35030 26138
rect 35082 26086 35094 26138
rect 35146 26086 35158 26138
rect 35210 26086 38824 26138
rect 1104 26064 38824 26086
rect 5994 25984 6000 26036
rect 6052 26024 6058 26036
rect 6457 26027 6515 26033
rect 6457 26024 6469 26027
rect 6052 25996 6469 26024
rect 6052 25984 6058 25996
rect 6457 25993 6469 25996
rect 6503 25993 6515 26027
rect 8662 26024 8668 26036
rect 8623 25996 8668 26024
rect 6457 25987 6515 25993
rect 8662 25984 8668 25996
rect 8720 25984 8726 26036
rect 13449 26027 13507 26033
rect 13449 25993 13461 26027
rect 13495 26024 13507 26027
rect 13998 26024 14004 26036
rect 13495 25996 14004 26024
rect 13495 25993 13507 25996
rect 13449 25987 13507 25993
rect 13998 25984 14004 25996
rect 14056 25984 14062 26036
rect 14921 26027 14979 26033
rect 14921 25993 14933 26027
rect 14967 26024 14979 26027
rect 15286 26024 15292 26036
rect 14967 25996 15292 26024
rect 14967 25993 14979 25996
rect 14921 25987 14979 25993
rect 11514 25956 11520 25968
rect 11475 25928 11520 25956
rect 11514 25916 11520 25928
rect 11572 25916 11578 25968
rect 12618 25916 12624 25968
rect 12676 25916 12682 25968
rect 14366 25956 14372 25968
rect 13832 25928 14372 25956
rect 9214 25848 9220 25900
rect 9272 25888 9278 25900
rect 9309 25891 9367 25897
rect 9309 25888 9321 25891
rect 9272 25860 9321 25888
rect 9272 25848 9278 25860
rect 9309 25857 9321 25860
rect 9355 25857 9367 25891
rect 12636 25888 12664 25916
rect 9309 25851 9367 25857
rect 12452 25860 12664 25888
rect 8297 25823 8355 25829
rect 8297 25789 8309 25823
rect 8343 25820 8355 25823
rect 9033 25823 9091 25829
rect 9033 25820 9045 25823
rect 8343 25792 9045 25820
rect 8343 25789 8355 25792
rect 8297 25783 8355 25789
rect 9033 25789 9045 25792
rect 9079 25820 9091 25823
rect 9674 25820 9680 25832
rect 9079 25792 9680 25820
rect 9079 25789 9091 25792
rect 9033 25783 9091 25789
rect 9674 25780 9680 25792
rect 9732 25780 9738 25832
rect 12452 25829 12480 25860
rect 12253 25823 12311 25829
rect 12253 25789 12265 25823
rect 12299 25820 12311 25823
rect 12437 25823 12495 25829
rect 12299 25792 12388 25820
rect 12299 25789 12311 25792
rect 12253 25783 12311 25789
rect 11885 25755 11943 25761
rect 11885 25721 11897 25755
rect 11931 25752 11943 25755
rect 12360 25752 12388 25792
rect 12437 25789 12449 25823
rect 12483 25789 12495 25823
rect 12618 25820 12624 25832
rect 12437 25783 12495 25789
rect 12544 25792 12624 25820
rect 12544 25752 12572 25792
rect 12618 25780 12624 25792
rect 12676 25780 12682 25832
rect 13832 25829 13860 25928
rect 14366 25916 14372 25928
rect 14424 25956 14430 25968
rect 14936 25956 14964 25987
rect 15286 25984 15292 25996
rect 15344 25984 15350 26036
rect 16666 26024 16672 26036
rect 16627 25996 16672 26024
rect 16666 25984 16672 25996
rect 16724 25984 16730 26036
rect 17862 26024 17868 26036
rect 17823 25996 17868 26024
rect 17862 25984 17868 25996
rect 17920 25984 17926 26036
rect 19058 25984 19064 26036
rect 19116 26024 19122 26036
rect 21085 26027 21143 26033
rect 21085 26024 21097 26027
rect 19116 25996 21097 26024
rect 19116 25984 19122 25996
rect 21085 25993 21097 25996
rect 21131 26024 21143 26027
rect 21266 26024 21272 26036
rect 21131 25996 21272 26024
rect 21131 25993 21143 25996
rect 21085 25987 21143 25993
rect 21266 25984 21272 25996
rect 21324 25984 21330 26036
rect 21450 26024 21456 26036
rect 21411 25996 21456 26024
rect 21450 25984 21456 25996
rect 21508 25984 21514 26036
rect 22554 25984 22560 26036
rect 22612 26024 22618 26036
rect 23201 26027 23259 26033
rect 23201 26024 23213 26027
rect 22612 25996 23213 26024
rect 22612 25984 22618 25996
rect 23201 25993 23213 25996
rect 23247 26024 23259 26027
rect 23474 26024 23480 26036
rect 23247 25996 23480 26024
rect 23247 25993 23259 25996
rect 23201 25987 23259 25993
rect 23474 25984 23480 25996
rect 23532 25984 23538 26036
rect 25314 26024 25320 26036
rect 25275 25996 25320 26024
rect 25314 25984 25320 25996
rect 25372 25984 25378 26036
rect 26970 25984 26976 26036
rect 27028 26024 27034 26036
rect 27065 26027 27123 26033
rect 27065 26024 27077 26027
rect 27028 25996 27077 26024
rect 27028 25984 27034 25996
rect 27065 25993 27077 25996
rect 27111 25993 27123 26027
rect 27614 26024 27620 26036
rect 27575 25996 27620 26024
rect 27065 25987 27123 25993
rect 27614 25984 27620 25996
rect 27672 25984 27678 26036
rect 14424 25928 14964 25956
rect 14424 25916 14430 25928
rect 18506 25916 18512 25968
rect 18564 25956 18570 25968
rect 19886 25956 19892 25968
rect 18564 25928 19892 25956
rect 18564 25916 18570 25928
rect 19886 25916 19892 25928
rect 19944 25956 19950 25968
rect 20165 25959 20223 25965
rect 20165 25956 20177 25959
rect 19944 25928 20177 25956
rect 19944 25916 19950 25928
rect 20165 25925 20177 25928
rect 20211 25925 20223 25959
rect 20165 25919 20223 25925
rect 20622 25916 20628 25968
rect 20680 25956 20686 25968
rect 20717 25959 20775 25965
rect 20717 25956 20729 25959
rect 20680 25928 20729 25956
rect 20680 25916 20686 25928
rect 20717 25925 20729 25928
rect 20763 25956 20775 25959
rect 21726 25956 21732 25968
rect 20763 25928 21732 25956
rect 20763 25925 20775 25928
rect 20717 25919 20775 25925
rect 21726 25916 21732 25928
rect 21784 25916 21790 25968
rect 22281 25959 22339 25965
rect 22281 25925 22293 25959
rect 22327 25956 22339 25959
rect 22922 25956 22928 25968
rect 22327 25928 22928 25956
rect 22327 25925 22339 25928
rect 22281 25919 22339 25925
rect 22922 25916 22928 25928
rect 22980 25916 22986 25968
rect 23492 25956 23520 25984
rect 25685 25959 25743 25965
rect 25685 25956 25697 25959
rect 23492 25928 25697 25956
rect 25685 25925 25697 25928
rect 25731 25925 25743 25959
rect 25685 25919 25743 25925
rect 14550 25848 14556 25900
rect 14608 25888 14614 25900
rect 14608 25860 15148 25888
rect 14608 25848 14614 25860
rect 13817 25823 13875 25829
rect 13817 25789 13829 25823
rect 13863 25789 13875 25823
rect 13817 25783 13875 25789
rect 14001 25823 14059 25829
rect 14001 25789 14013 25823
rect 14047 25820 14059 25823
rect 14642 25820 14648 25832
rect 14047 25792 14648 25820
rect 14047 25789 14059 25792
rect 14001 25783 14059 25789
rect 14642 25780 14648 25792
rect 14700 25780 14706 25832
rect 13722 25752 13728 25764
rect 11931 25724 12296 25752
rect 12360 25724 12572 25752
rect 12636 25724 13728 25752
rect 11931 25721 11943 25724
rect 11885 25715 11943 25721
rect 6086 25684 6092 25696
rect 6047 25656 6092 25684
rect 6086 25644 6092 25656
rect 6144 25644 6150 25696
rect 10594 25684 10600 25696
rect 10555 25656 10600 25684
rect 10594 25644 10600 25656
rect 10652 25644 10658 25696
rect 11146 25684 11152 25696
rect 11107 25656 11152 25684
rect 11146 25644 11152 25656
rect 11204 25644 11210 25696
rect 12268 25684 12296 25724
rect 12636 25684 12664 25724
rect 13722 25712 13728 25724
rect 13780 25712 13786 25764
rect 14185 25755 14243 25761
rect 14185 25721 14197 25755
rect 14231 25752 14243 25755
rect 14366 25752 14372 25764
rect 14231 25724 14372 25752
rect 14231 25721 14243 25724
rect 14185 25715 14243 25721
rect 14366 25712 14372 25724
rect 14424 25712 14430 25764
rect 14550 25752 14556 25764
rect 14511 25724 14556 25752
rect 14550 25712 14556 25724
rect 14608 25712 14614 25764
rect 15120 25752 15148 25860
rect 15286 25848 15292 25900
rect 15344 25888 15350 25900
rect 16114 25888 16120 25900
rect 15344 25860 16120 25888
rect 15344 25848 15350 25860
rect 16114 25848 16120 25860
rect 16172 25888 16178 25900
rect 16393 25891 16451 25897
rect 16393 25888 16405 25891
rect 16172 25860 16405 25888
rect 16172 25848 16178 25860
rect 16393 25857 16405 25860
rect 16439 25888 16451 25891
rect 18230 25888 18236 25900
rect 16439 25860 18236 25888
rect 16439 25857 16451 25860
rect 16393 25851 16451 25857
rect 15194 25780 15200 25832
rect 15252 25820 15258 25832
rect 15381 25823 15439 25829
rect 15381 25820 15393 25823
rect 15252 25792 15393 25820
rect 15252 25780 15258 25792
rect 15381 25789 15393 25792
rect 15427 25789 15439 25823
rect 15381 25783 15439 25789
rect 15933 25823 15991 25829
rect 15933 25789 15945 25823
rect 15979 25789 15991 25823
rect 16206 25820 16212 25832
rect 16167 25792 16212 25820
rect 15933 25783 15991 25789
rect 15948 25752 15976 25783
rect 16206 25780 16212 25792
rect 16264 25820 16270 25832
rect 16574 25820 16580 25832
rect 16264 25792 16580 25820
rect 16264 25780 16270 25792
rect 16574 25780 16580 25792
rect 16632 25780 16638 25832
rect 18156 25829 18184 25860
rect 18230 25848 18236 25860
rect 18288 25848 18294 25900
rect 18325 25891 18383 25897
rect 18325 25857 18337 25891
rect 18371 25888 18383 25891
rect 19334 25888 19340 25900
rect 18371 25860 19340 25888
rect 18371 25857 18383 25860
rect 18325 25851 18383 25857
rect 19334 25848 19340 25860
rect 19392 25848 19398 25900
rect 20070 25848 20076 25900
rect 20128 25888 20134 25900
rect 21177 25891 21235 25897
rect 21177 25888 21189 25891
rect 20128 25860 21189 25888
rect 20128 25848 20134 25860
rect 21177 25857 21189 25860
rect 21223 25857 21235 25891
rect 21177 25851 21235 25857
rect 21450 25848 21456 25900
rect 21508 25888 21514 25900
rect 21634 25888 21640 25900
rect 21508 25860 21640 25888
rect 21508 25848 21514 25860
rect 21634 25848 21640 25860
rect 21692 25848 21698 25900
rect 23934 25848 23940 25900
rect 23992 25888 23998 25900
rect 24305 25891 24363 25897
rect 24305 25888 24317 25891
rect 23992 25860 24317 25888
rect 23992 25848 23998 25860
rect 24305 25857 24317 25860
rect 24351 25857 24363 25891
rect 24305 25851 24363 25857
rect 24765 25891 24823 25897
rect 24765 25857 24777 25891
rect 24811 25888 24823 25891
rect 24946 25888 24952 25900
rect 24811 25860 24952 25888
rect 24811 25857 24823 25860
rect 24765 25851 24823 25857
rect 24946 25848 24952 25860
rect 25004 25848 25010 25900
rect 18141 25823 18199 25829
rect 18141 25789 18153 25823
rect 18187 25789 18199 25823
rect 18690 25820 18696 25832
rect 18651 25792 18696 25820
rect 18141 25783 18199 25789
rect 18690 25780 18696 25792
rect 18748 25780 18754 25832
rect 18782 25780 18788 25832
rect 18840 25820 18846 25832
rect 18877 25823 18935 25829
rect 18877 25820 18889 25823
rect 18840 25792 18889 25820
rect 18840 25780 18846 25792
rect 18877 25789 18889 25792
rect 18923 25789 18935 25823
rect 18877 25783 18935 25789
rect 19245 25823 19303 25829
rect 19245 25789 19257 25823
rect 19291 25820 19303 25823
rect 19291 25792 19380 25820
rect 19291 25789 19303 25792
rect 19245 25783 19303 25789
rect 15120 25724 15976 25752
rect 17497 25755 17555 25761
rect 17497 25721 17509 25755
rect 17543 25752 17555 25755
rect 18708 25752 18736 25780
rect 17543 25724 18736 25752
rect 19352 25752 19380 25792
rect 19426 25780 19432 25832
rect 19484 25820 19490 25832
rect 19613 25823 19671 25829
rect 19613 25820 19625 25823
rect 19484 25792 19625 25820
rect 19484 25780 19490 25792
rect 19613 25789 19625 25792
rect 19659 25789 19671 25823
rect 19613 25783 19671 25789
rect 20956 25823 21014 25829
rect 20956 25789 20968 25823
rect 21002 25820 21014 25823
rect 21358 25820 21364 25832
rect 21002 25792 21364 25820
rect 21002 25789 21014 25792
rect 20956 25783 21014 25789
rect 21358 25780 21364 25792
rect 21416 25820 21422 25832
rect 21726 25820 21732 25832
rect 21416 25792 21732 25820
rect 21416 25780 21422 25792
rect 21726 25780 21732 25792
rect 21784 25780 21790 25832
rect 21913 25823 21971 25829
rect 21913 25789 21925 25823
rect 21959 25820 21971 25823
rect 22373 25823 22431 25829
rect 22373 25820 22385 25823
rect 21959 25792 22385 25820
rect 21959 25789 21971 25792
rect 21913 25783 21971 25789
rect 22373 25789 22385 25792
rect 22419 25820 22431 25823
rect 22462 25820 22468 25832
rect 22419 25792 22468 25820
rect 22419 25789 22431 25792
rect 22373 25783 22431 25789
rect 22462 25780 22468 25792
rect 22520 25780 22526 25832
rect 24026 25780 24032 25832
rect 24084 25820 24090 25832
rect 24489 25823 24547 25829
rect 24489 25820 24501 25823
rect 24084 25792 24501 25820
rect 24084 25780 24090 25792
rect 24489 25789 24501 25792
rect 24535 25789 24547 25823
rect 24854 25820 24860 25832
rect 24815 25792 24860 25820
rect 24489 25783 24547 25789
rect 24854 25780 24860 25792
rect 24912 25780 24918 25832
rect 20346 25752 20352 25764
rect 19352 25724 20352 25752
rect 17543 25721 17555 25724
rect 17497 25715 17555 25721
rect 20346 25712 20352 25724
rect 20404 25712 20410 25764
rect 20806 25752 20812 25764
rect 20767 25724 20812 25752
rect 20806 25712 20812 25724
rect 20864 25712 20870 25764
rect 25700 25752 25728 25919
rect 26694 25888 26700 25900
rect 25884 25860 26700 25888
rect 25884 25832 25912 25860
rect 26694 25848 26700 25860
rect 26752 25848 26758 25900
rect 25866 25820 25872 25832
rect 25827 25792 25872 25820
rect 25866 25780 25872 25792
rect 25924 25780 25930 25832
rect 26050 25820 26056 25832
rect 25963 25792 26056 25820
rect 26050 25780 26056 25792
rect 26108 25780 26114 25832
rect 26068 25752 26096 25780
rect 26418 25752 26424 25764
rect 20971 25724 24256 25752
rect 25700 25724 26096 25752
rect 26379 25724 26424 25752
rect 12268 25656 12664 25684
rect 12713 25687 12771 25693
rect 12713 25653 12725 25687
rect 12759 25684 12771 25687
rect 13906 25684 13912 25696
rect 12759 25656 13912 25684
rect 12759 25653 12771 25656
rect 12713 25647 12771 25653
rect 13906 25644 13912 25656
rect 13964 25644 13970 25696
rect 14093 25687 14151 25693
rect 14093 25653 14105 25687
rect 14139 25684 14151 25687
rect 14734 25684 14740 25696
rect 14139 25656 14740 25684
rect 14139 25653 14151 25656
rect 14093 25647 14151 25653
rect 14734 25644 14740 25656
rect 14792 25684 14798 25696
rect 17129 25687 17187 25693
rect 17129 25684 17141 25687
rect 14792 25656 17141 25684
rect 14792 25644 14798 25656
rect 17129 25653 17141 25656
rect 17175 25684 17187 25687
rect 17586 25684 17592 25696
rect 17175 25656 17592 25684
rect 17175 25653 17187 25656
rect 17129 25647 17187 25653
rect 17586 25644 17592 25656
rect 17644 25644 17650 25696
rect 20165 25687 20223 25693
rect 20165 25653 20177 25687
rect 20211 25684 20223 25687
rect 20257 25687 20315 25693
rect 20257 25684 20269 25687
rect 20211 25656 20269 25684
rect 20211 25653 20223 25656
rect 20165 25647 20223 25653
rect 20257 25653 20269 25656
rect 20303 25684 20315 25687
rect 20971 25684 20999 25724
rect 20303 25656 20999 25684
rect 20303 25653 20315 25656
rect 20257 25647 20315 25653
rect 21634 25644 21640 25696
rect 21692 25684 21698 25696
rect 22557 25687 22615 25693
rect 22557 25684 22569 25687
rect 21692 25656 22569 25684
rect 21692 25644 21698 25656
rect 22557 25653 22569 25656
rect 22603 25653 22615 25687
rect 22830 25684 22836 25696
rect 22791 25656 22836 25684
rect 22557 25647 22615 25653
rect 22830 25644 22836 25656
rect 22888 25644 22894 25696
rect 24118 25684 24124 25696
rect 24079 25656 24124 25684
rect 24118 25644 24124 25656
rect 24176 25644 24182 25696
rect 24228 25684 24256 25724
rect 26418 25712 26424 25724
rect 26476 25712 26482 25764
rect 27246 25684 27252 25696
rect 24228 25656 27252 25684
rect 27246 25644 27252 25656
rect 27304 25644 27310 25696
rect 1104 25594 38824 25616
rect 1104 25542 19606 25594
rect 19658 25542 19670 25594
rect 19722 25542 19734 25594
rect 19786 25542 19798 25594
rect 19850 25542 38824 25594
rect 1104 25520 38824 25542
rect 9125 25483 9183 25489
rect 9125 25449 9137 25483
rect 9171 25480 9183 25483
rect 9214 25480 9220 25492
rect 9171 25452 9220 25480
rect 9171 25449 9183 25452
rect 9125 25443 9183 25449
rect 9214 25440 9220 25452
rect 9272 25440 9278 25492
rect 9490 25480 9496 25492
rect 9451 25452 9496 25480
rect 9490 25440 9496 25452
rect 9548 25440 9554 25492
rect 11330 25480 11336 25492
rect 11291 25452 11336 25480
rect 11330 25440 11336 25452
rect 11388 25440 11394 25492
rect 12158 25480 12164 25492
rect 12119 25452 12164 25480
rect 12158 25440 12164 25452
rect 12216 25440 12222 25492
rect 12342 25440 12348 25492
rect 12400 25480 12406 25492
rect 12437 25483 12495 25489
rect 12437 25480 12449 25483
rect 12400 25452 12449 25480
rect 12400 25440 12406 25452
rect 12437 25449 12449 25452
rect 12483 25449 12495 25483
rect 12437 25443 12495 25449
rect 12897 25483 12955 25489
rect 12897 25449 12909 25483
rect 12943 25480 12955 25483
rect 13265 25483 13323 25489
rect 13265 25480 13277 25483
rect 12943 25452 13277 25480
rect 12943 25449 12955 25452
rect 12897 25443 12955 25449
rect 13265 25449 13277 25452
rect 13311 25480 13323 25483
rect 13354 25480 13360 25492
rect 13311 25452 13360 25480
rect 13311 25449 13323 25452
rect 13265 25443 13323 25449
rect 13354 25440 13360 25452
rect 13412 25440 13418 25492
rect 14734 25480 14740 25492
rect 14695 25452 14740 25480
rect 14734 25440 14740 25452
rect 14792 25440 14798 25492
rect 15562 25480 15568 25492
rect 15523 25452 15568 25480
rect 15562 25440 15568 25452
rect 15620 25440 15626 25492
rect 16482 25480 16488 25492
rect 16443 25452 16488 25480
rect 16482 25440 16488 25452
rect 16540 25440 16546 25492
rect 16942 25440 16948 25492
rect 17000 25480 17006 25492
rect 17678 25480 17684 25492
rect 17000 25452 17684 25480
rect 17000 25440 17006 25452
rect 17678 25440 17684 25452
rect 17736 25440 17742 25492
rect 20070 25480 20076 25492
rect 20031 25452 20076 25480
rect 20070 25440 20076 25452
rect 20128 25480 20134 25492
rect 21085 25483 21143 25489
rect 21085 25480 21097 25483
rect 20128 25452 21097 25480
rect 20128 25440 20134 25452
rect 21085 25449 21097 25452
rect 21131 25449 21143 25483
rect 22738 25480 22744 25492
rect 22699 25452 22744 25480
rect 21085 25443 21143 25449
rect 22738 25440 22744 25452
rect 22796 25440 22802 25492
rect 25314 25480 25320 25492
rect 25275 25452 25320 25480
rect 25314 25440 25320 25452
rect 25372 25440 25378 25492
rect 26697 25483 26755 25489
rect 26697 25449 26709 25483
rect 26743 25480 26755 25483
rect 27338 25480 27344 25492
rect 26743 25452 27344 25480
rect 26743 25449 26755 25452
rect 26697 25443 26755 25449
rect 27338 25440 27344 25452
rect 27396 25440 27402 25492
rect 9232 25344 9260 25440
rect 10594 25372 10600 25424
rect 10652 25372 10658 25424
rect 18506 25412 18512 25424
rect 15396 25384 18512 25412
rect 10137 25347 10195 25353
rect 10137 25344 10149 25347
rect 9232 25316 10149 25344
rect 10137 25313 10149 25316
rect 10183 25313 10195 25347
rect 10137 25307 10195 25313
rect 10226 25304 10232 25356
rect 10284 25344 10290 25356
rect 10321 25347 10379 25353
rect 10321 25344 10333 25347
rect 10284 25316 10333 25344
rect 10284 25304 10290 25316
rect 10321 25313 10333 25316
rect 10367 25313 10379 25347
rect 10612 25344 10640 25372
rect 15396 25356 15424 25384
rect 18506 25372 18512 25384
rect 18564 25372 18570 25424
rect 19426 25372 19432 25424
rect 19484 25412 19490 25424
rect 19610 25412 19616 25424
rect 19484 25384 19616 25412
rect 19484 25372 19490 25384
rect 19610 25372 19616 25384
rect 19668 25412 19674 25424
rect 22465 25415 22523 25421
rect 19668 25384 19748 25412
rect 19668 25372 19674 25384
rect 10689 25347 10747 25353
rect 10689 25344 10701 25347
rect 10612 25316 10701 25344
rect 10321 25307 10379 25313
rect 10689 25313 10701 25316
rect 10735 25313 10747 25347
rect 10689 25307 10747 25313
rect 10778 25304 10784 25356
rect 10836 25344 10842 25356
rect 10836 25316 10881 25344
rect 10836 25304 10842 25316
rect 11054 25304 11060 25356
rect 11112 25344 11118 25356
rect 11882 25344 11888 25356
rect 11112 25316 11888 25344
rect 11112 25304 11118 25316
rect 11882 25304 11888 25316
rect 11940 25344 11946 25356
rect 12253 25347 12311 25353
rect 12253 25344 12265 25347
rect 11940 25316 12265 25344
rect 11940 25304 11946 25316
rect 12253 25313 12265 25316
rect 12299 25313 12311 25347
rect 12253 25307 12311 25313
rect 13817 25347 13875 25353
rect 13817 25313 13829 25347
rect 13863 25344 13875 25347
rect 14090 25344 14096 25356
rect 13863 25316 14096 25344
rect 13863 25313 13875 25316
rect 13817 25307 13875 25313
rect 14090 25304 14096 25316
rect 14148 25304 14154 25356
rect 14185 25347 14243 25353
rect 14185 25313 14197 25347
rect 14231 25344 14243 25347
rect 14458 25344 14464 25356
rect 14231 25316 14464 25344
rect 14231 25313 14243 25316
rect 14185 25307 14243 25313
rect 9674 25276 9680 25288
rect 9635 25248 9680 25276
rect 9674 25236 9680 25248
rect 9732 25236 9738 25288
rect 13906 25236 13912 25288
rect 13964 25276 13970 25288
rect 14200 25276 14228 25307
rect 14458 25304 14464 25316
rect 14516 25304 14522 25356
rect 15378 25344 15384 25356
rect 15339 25316 15384 25344
rect 15378 25304 15384 25316
rect 15436 25304 15442 25356
rect 16666 25304 16672 25356
rect 16724 25344 16730 25356
rect 16942 25344 16948 25356
rect 16724 25316 16948 25344
rect 16724 25304 16730 25316
rect 16942 25304 16948 25316
rect 17000 25304 17006 25356
rect 17034 25304 17040 25356
rect 17092 25344 17098 25356
rect 17218 25344 17224 25356
rect 17092 25316 17137 25344
rect 17179 25316 17224 25344
rect 17092 25304 17098 25316
rect 17218 25304 17224 25316
rect 17276 25304 17282 25356
rect 17494 25344 17500 25356
rect 17455 25316 17500 25344
rect 17494 25304 17500 25316
rect 17552 25304 17558 25356
rect 17862 25344 17868 25356
rect 17823 25316 17868 25344
rect 17862 25304 17868 25316
rect 17920 25304 17926 25356
rect 18969 25347 19027 25353
rect 18969 25313 18981 25347
rect 19015 25344 19027 25347
rect 19242 25344 19248 25356
rect 19015 25316 19248 25344
rect 19015 25313 19027 25316
rect 18969 25307 19027 25313
rect 19242 25304 19248 25316
rect 19300 25304 19306 25356
rect 19334 25304 19340 25356
rect 19392 25344 19398 25356
rect 19720 25353 19748 25384
rect 22465 25381 22477 25415
rect 22511 25412 22523 25415
rect 22830 25412 22836 25424
rect 22511 25384 22836 25412
rect 22511 25381 22523 25384
rect 22465 25375 22523 25381
rect 22830 25372 22836 25384
rect 22888 25372 22894 25424
rect 26786 25372 26792 25424
rect 26844 25412 26850 25424
rect 26973 25415 27031 25421
rect 26973 25412 26985 25415
rect 26844 25384 26985 25412
rect 26844 25372 26850 25384
rect 26973 25381 26985 25384
rect 27019 25381 27031 25415
rect 26973 25375 27031 25381
rect 19521 25347 19579 25353
rect 19521 25344 19533 25347
rect 19392 25316 19533 25344
rect 19392 25304 19398 25316
rect 19521 25313 19533 25316
rect 19567 25313 19579 25347
rect 19521 25307 19579 25313
rect 19705 25347 19763 25353
rect 19705 25313 19717 25347
rect 19751 25313 19763 25347
rect 19705 25307 19763 25313
rect 21082 25304 21088 25356
rect 21140 25344 21146 25356
rect 21266 25344 21272 25356
rect 21140 25316 21272 25344
rect 21140 25304 21146 25316
rect 21266 25304 21272 25316
rect 21324 25304 21330 25356
rect 22281 25347 22339 25353
rect 22281 25344 22293 25347
rect 22204 25316 22293 25344
rect 13964 25248 14228 25276
rect 14277 25279 14335 25285
rect 13964 25236 13970 25248
rect 14277 25245 14289 25279
rect 14323 25276 14335 25279
rect 14366 25276 14372 25288
rect 14323 25248 14372 25276
rect 14323 25245 14335 25248
rect 14277 25239 14335 25245
rect 14366 25236 14372 25248
rect 14424 25236 14430 25288
rect 16301 25279 16359 25285
rect 16301 25245 16313 25279
rect 16347 25276 16359 25279
rect 17880 25276 17908 25304
rect 22204 25288 22232 25316
rect 22281 25313 22293 25316
rect 22327 25313 22339 25347
rect 22281 25307 22339 25313
rect 22554 25304 22560 25356
rect 22612 25344 22618 25356
rect 23109 25347 23167 25353
rect 23109 25344 23121 25347
rect 22612 25316 23121 25344
rect 22612 25304 22618 25316
rect 23109 25313 23121 25316
rect 23155 25313 23167 25347
rect 23109 25307 23167 25313
rect 23385 25347 23443 25353
rect 23385 25313 23397 25347
rect 23431 25344 23443 25347
rect 23750 25344 23756 25356
rect 23431 25316 23756 25344
rect 23431 25313 23443 25316
rect 23385 25307 23443 25313
rect 23750 25304 23756 25316
rect 23808 25304 23814 25356
rect 23934 25304 23940 25356
rect 23992 25304 23998 25356
rect 24026 25304 24032 25356
rect 24084 25344 24090 25356
rect 25590 25344 25596 25356
rect 24084 25316 25596 25344
rect 24084 25304 24090 25316
rect 25590 25304 25596 25316
rect 25648 25344 25654 25356
rect 25685 25347 25743 25353
rect 25685 25344 25697 25347
rect 25648 25316 25697 25344
rect 25648 25304 25654 25316
rect 25685 25313 25697 25316
rect 25731 25313 25743 25347
rect 25685 25307 25743 25313
rect 26513 25347 26571 25353
rect 26513 25313 26525 25347
rect 26559 25344 26571 25347
rect 26602 25344 26608 25356
rect 26559 25316 26608 25344
rect 26559 25313 26571 25316
rect 26513 25307 26571 25313
rect 26602 25304 26608 25316
rect 26660 25304 26666 25356
rect 16347 25248 17908 25276
rect 16347 25245 16359 25248
rect 16301 25239 16359 25245
rect 22186 25236 22192 25288
rect 22244 25236 22250 25288
rect 23661 25279 23719 25285
rect 23661 25245 23673 25279
rect 23707 25276 23719 25279
rect 23952 25276 23980 25304
rect 24762 25276 24768 25288
rect 23707 25248 24768 25276
rect 23707 25245 23719 25248
rect 23661 25239 23719 25245
rect 24762 25236 24768 25248
rect 24820 25276 24826 25288
rect 26050 25276 26056 25288
rect 24820 25248 26056 25276
rect 24820 25236 24826 25248
rect 26050 25236 26056 25248
rect 26108 25236 26114 25288
rect 11793 25211 11851 25217
rect 11793 25177 11805 25211
rect 11839 25208 11851 25211
rect 12342 25208 12348 25220
rect 11839 25180 12348 25208
rect 11839 25177 11851 25180
rect 11793 25171 11851 25177
rect 12342 25168 12348 25180
rect 12400 25168 12406 25220
rect 13633 25211 13691 25217
rect 13633 25177 13645 25211
rect 13679 25208 13691 25211
rect 13722 25208 13728 25220
rect 13679 25180 13728 25208
rect 13679 25177 13691 25180
rect 13633 25171 13691 25177
rect 13722 25168 13728 25180
rect 13780 25168 13786 25220
rect 15562 25168 15568 25220
rect 15620 25208 15626 25220
rect 17862 25208 17868 25220
rect 15620 25180 17868 25208
rect 15620 25168 15626 25180
rect 17862 25168 17868 25180
rect 17920 25168 17926 25220
rect 18046 25168 18052 25220
rect 18104 25208 18110 25220
rect 18509 25211 18567 25217
rect 18509 25208 18521 25211
rect 18104 25180 18521 25208
rect 18104 25168 18110 25180
rect 18509 25177 18521 25180
rect 18555 25177 18567 25211
rect 19518 25208 19524 25220
rect 19479 25180 19524 25208
rect 18509 25171 18567 25177
rect 19518 25168 19524 25180
rect 19576 25168 19582 25220
rect 15102 25140 15108 25152
rect 15063 25112 15108 25140
rect 15102 25100 15108 25112
rect 15160 25100 15166 25152
rect 15930 25140 15936 25152
rect 15843 25112 15936 25140
rect 15930 25100 15936 25112
rect 15988 25140 15994 25152
rect 16482 25140 16488 25152
rect 15988 25112 16488 25140
rect 15988 25100 15994 25112
rect 16482 25100 16488 25112
rect 16540 25100 16546 25152
rect 18233 25143 18291 25149
rect 18233 25109 18245 25143
rect 18279 25140 18291 25143
rect 18782 25140 18788 25152
rect 18279 25112 18788 25140
rect 18279 25109 18291 25112
rect 18233 25103 18291 25109
rect 18782 25100 18788 25112
rect 18840 25100 18846 25152
rect 20438 25140 20444 25152
rect 20399 25112 20444 25140
rect 20438 25100 20444 25112
rect 20496 25100 20502 25152
rect 21450 25140 21456 25152
rect 21411 25112 21456 25140
rect 21450 25100 21456 25112
rect 21508 25100 21514 25152
rect 24854 25100 24860 25152
rect 24912 25140 24918 25152
rect 24949 25143 25007 25149
rect 24949 25140 24961 25143
rect 24912 25112 24961 25140
rect 24912 25100 24918 25112
rect 24949 25109 24961 25112
rect 24995 25109 25007 25143
rect 24949 25103 25007 25109
rect 1104 25050 38824 25072
rect 1104 24998 4246 25050
rect 4298 24998 4310 25050
rect 4362 24998 4374 25050
rect 4426 24998 4438 25050
rect 4490 24998 34966 25050
rect 35018 24998 35030 25050
rect 35082 24998 35094 25050
rect 35146 24998 35158 25050
rect 35210 24998 38824 25050
rect 1104 24976 38824 24998
rect 11882 24936 11888 24948
rect 11843 24908 11888 24936
rect 11882 24896 11888 24908
rect 11940 24896 11946 24948
rect 14182 24896 14188 24948
rect 14240 24936 14246 24948
rect 14737 24939 14795 24945
rect 14737 24936 14749 24939
rect 14240 24908 14749 24936
rect 14240 24896 14246 24908
rect 14737 24905 14749 24908
rect 14783 24905 14795 24939
rect 15378 24936 15384 24948
rect 15339 24908 15384 24936
rect 14737 24899 14795 24905
rect 15378 24896 15384 24908
rect 15436 24896 15442 24948
rect 19610 24936 19616 24948
rect 19571 24908 19616 24936
rect 19610 24896 19616 24908
rect 19668 24896 19674 24948
rect 20070 24896 20076 24948
rect 20128 24896 20134 24948
rect 21174 24896 21180 24948
rect 21232 24936 21238 24948
rect 23017 24939 23075 24945
rect 23017 24936 23029 24939
rect 21232 24908 23029 24936
rect 21232 24896 21238 24908
rect 23017 24905 23029 24908
rect 23063 24905 23075 24939
rect 23474 24936 23480 24948
rect 23435 24908 23480 24936
rect 23017 24899 23075 24905
rect 23474 24896 23480 24908
rect 23532 24896 23538 24948
rect 26602 24936 26608 24948
rect 26563 24908 26608 24936
rect 26602 24896 26608 24908
rect 26660 24896 26666 24948
rect 10594 24828 10600 24880
rect 10652 24868 10658 24880
rect 14090 24868 14096 24880
rect 10652 24840 11008 24868
rect 14003 24840 14096 24868
rect 10652 24828 10658 24840
rect 2682 24760 2688 24812
rect 2740 24800 2746 24812
rect 8941 24803 8999 24809
rect 8941 24800 8953 24803
rect 2740 24772 8953 24800
rect 2740 24760 2746 24772
rect 8941 24769 8953 24772
rect 8987 24800 8999 24803
rect 9401 24803 9459 24809
rect 9401 24800 9413 24803
rect 8987 24772 9413 24800
rect 8987 24769 8999 24772
rect 8941 24763 8999 24769
rect 9401 24769 9413 24772
rect 9447 24769 9459 24803
rect 9401 24763 9459 24769
rect 10042 24760 10048 24812
rect 10100 24800 10106 24812
rect 10505 24803 10563 24809
rect 10505 24800 10517 24803
rect 10100 24772 10517 24800
rect 10100 24760 10106 24772
rect 10505 24769 10517 24772
rect 10551 24769 10563 24803
rect 10980 24800 11008 24840
rect 14090 24828 14096 24840
rect 14148 24868 14154 24880
rect 15102 24868 15108 24880
rect 14148 24840 15108 24868
rect 14148 24828 14154 24840
rect 15102 24828 15108 24840
rect 15160 24828 15166 24880
rect 16942 24828 16948 24880
rect 17000 24868 17006 24880
rect 17494 24868 17500 24880
rect 17000 24840 17500 24868
rect 17000 24828 17006 24840
rect 17494 24828 17500 24840
rect 17552 24868 17558 24880
rect 20088 24868 20116 24896
rect 20349 24871 20407 24877
rect 20349 24868 20361 24871
rect 17552 24840 17908 24868
rect 17552 24828 17558 24840
rect 11057 24803 11115 24809
rect 11057 24800 11069 24803
rect 10980 24772 11069 24800
rect 10505 24763 10563 24769
rect 11057 24769 11069 24772
rect 11103 24769 11115 24803
rect 11057 24763 11115 24769
rect 12434 24760 12440 24812
rect 12492 24800 12498 24812
rect 14458 24800 14464 24812
rect 12492 24772 13584 24800
rect 14419 24772 14464 24800
rect 12492 24760 12498 24772
rect 9125 24735 9183 24741
rect 9125 24732 9137 24735
rect 8680 24704 9137 24732
rect 8680 24608 8708 24704
rect 9125 24701 9137 24704
rect 9171 24701 9183 24735
rect 9125 24695 9183 24701
rect 12618 24692 12624 24744
rect 12676 24732 12682 24744
rect 12989 24735 13047 24741
rect 12989 24732 13001 24735
rect 12676 24704 13001 24732
rect 12676 24692 12682 24704
rect 12989 24701 13001 24704
rect 13035 24732 13047 24735
rect 13078 24732 13084 24744
rect 13035 24704 13084 24732
rect 13035 24701 13047 24704
rect 12989 24695 13047 24701
rect 13078 24692 13084 24704
rect 13136 24692 13142 24744
rect 13556 24741 13584 24772
rect 14458 24760 14464 24772
rect 14516 24760 14522 24812
rect 14918 24760 14924 24812
rect 14976 24800 14982 24812
rect 16206 24800 16212 24812
rect 14976 24772 16212 24800
rect 14976 24760 14982 24772
rect 16206 24760 16212 24772
rect 16264 24760 16270 24812
rect 17880 24800 17908 24840
rect 19260 24840 20116 24868
rect 20272 24840 20361 24868
rect 18049 24803 18107 24809
rect 18049 24800 18061 24803
rect 17880 24772 18061 24800
rect 18049 24769 18061 24772
rect 18095 24769 18107 24803
rect 18049 24763 18107 24769
rect 18785 24803 18843 24809
rect 18785 24769 18797 24803
rect 18831 24800 18843 24803
rect 19260 24800 19288 24840
rect 18831 24772 19288 24800
rect 18831 24769 18843 24772
rect 18785 24763 18843 24769
rect 20070 24760 20076 24812
rect 20128 24800 20134 24812
rect 20272 24800 20300 24840
rect 20349 24837 20361 24840
rect 20395 24868 20407 24871
rect 21450 24868 21456 24880
rect 20395 24840 21456 24868
rect 20395 24837 20407 24840
rect 20349 24831 20407 24837
rect 21450 24828 21456 24840
rect 21508 24828 21514 24880
rect 20438 24800 20444 24812
rect 20128 24772 20300 24800
rect 20399 24772 20444 24800
rect 20128 24760 20134 24772
rect 20438 24760 20444 24772
rect 20496 24760 20502 24812
rect 22278 24800 22284 24812
rect 20548 24772 22284 24800
rect 13173 24735 13231 24741
rect 13173 24701 13185 24735
rect 13219 24701 13231 24735
rect 13173 24695 13231 24701
rect 13541 24735 13599 24741
rect 13541 24701 13553 24735
rect 13587 24701 13599 24735
rect 13722 24732 13728 24744
rect 13683 24704 13728 24732
rect 13541 24695 13599 24701
rect 13188 24664 13216 24695
rect 11440 24636 13216 24664
rect 13556 24664 13584 24695
rect 13722 24692 13728 24704
rect 13780 24692 13786 24744
rect 14553 24735 14611 24741
rect 14553 24701 14565 24735
rect 14599 24732 14611 24735
rect 14599 24704 14964 24732
rect 14599 24701 14611 24704
rect 14553 24695 14611 24701
rect 13814 24664 13820 24676
rect 13556 24636 13820 24664
rect 8662 24596 8668 24608
rect 8623 24568 8668 24596
rect 8662 24556 8668 24568
rect 8720 24556 8726 24608
rect 10962 24556 10968 24608
rect 11020 24596 11026 24608
rect 11440 24605 11468 24636
rect 13814 24624 13820 24636
rect 13872 24624 13878 24676
rect 14936 24608 14964 24704
rect 15194 24692 15200 24744
rect 15252 24732 15258 24744
rect 15470 24732 15476 24744
rect 15252 24704 15476 24732
rect 15252 24692 15258 24704
rect 15470 24692 15476 24704
rect 15528 24692 15534 24744
rect 16117 24735 16175 24741
rect 16117 24701 16129 24735
rect 16163 24732 16175 24735
rect 16482 24732 16488 24744
rect 16163 24704 16488 24732
rect 16163 24701 16175 24704
rect 16117 24695 16175 24701
rect 16482 24692 16488 24704
rect 16540 24692 16546 24744
rect 16669 24735 16727 24741
rect 16669 24701 16681 24735
rect 16715 24732 16727 24735
rect 16758 24732 16764 24744
rect 16715 24704 16764 24732
rect 16715 24701 16727 24704
rect 16669 24695 16727 24701
rect 16758 24692 16764 24704
rect 16816 24692 16822 24744
rect 16853 24735 16911 24741
rect 16853 24701 16865 24735
rect 16899 24732 16911 24735
rect 17310 24732 17316 24744
rect 16899 24704 17316 24732
rect 16899 24701 16911 24704
rect 16853 24695 16911 24701
rect 17310 24692 17316 24704
rect 17368 24692 17374 24744
rect 18690 24732 18696 24744
rect 18651 24704 18696 24732
rect 18690 24692 18696 24704
rect 18748 24692 18754 24744
rect 19058 24732 19064 24744
rect 19019 24704 19064 24732
rect 19058 24692 19064 24704
rect 19116 24692 19122 24744
rect 19153 24735 19211 24741
rect 19153 24701 19165 24735
rect 19199 24701 19211 24735
rect 19153 24695 19211 24701
rect 18046 24624 18052 24676
rect 18104 24664 18110 24676
rect 19168 24664 19196 24695
rect 19242 24692 19248 24744
rect 19300 24732 19306 24744
rect 19889 24735 19947 24741
rect 19889 24732 19901 24735
rect 19300 24704 19901 24732
rect 19300 24692 19306 24704
rect 19889 24701 19901 24704
rect 19935 24732 19947 24735
rect 19978 24732 19984 24744
rect 19935 24704 19984 24732
rect 19935 24701 19947 24704
rect 19889 24695 19947 24701
rect 19978 24692 19984 24704
rect 20036 24692 20042 24744
rect 20220 24735 20278 24741
rect 20220 24701 20232 24735
rect 20266 24732 20278 24735
rect 20548 24732 20576 24772
rect 22278 24760 22284 24772
rect 22336 24800 22342 24812
rect 22649 24803 22707 24809
rect 22649 24800 22661 24803
rect 22336 24772 22661 24800
rect 22336 24760 22342 24772
rect 22649 24769 22661 24772
rect 22695 24769 22707 24803
rect 23492 24800 23520 24896
rect 23661 24803 23719 24809
rect 23661 24800 23673 24803
rect 23492 24772 23673 24800
rect 22649 24763 22707 24769
rect 23661 24769 23673 24772
rect 23707 24769 23719 24803
rect 24581 24803 24639 24809
rect 24581 24800 24593 24803
rect 23661 24763 23719 24769
rect 23768 24772 24593 24800
rect 23768 24744 23796 24772
rect 24581 24769 24593 24772
rect 24627 24800 24639 24803
rect 24670 24800 24676 24812
rect 24627 24772 24676 24800
rect 24627 24769 24639 24772
rect 24581 24763 24639 24769
rect 24670 24760 24676 24772
rect 24728 24760 24734 24812
rect 24946 24800 24952 24812
rect 24907 24772 24952 24800
rect 24946 24760 24952 24772
rect 25004 24760 25010 24812
rect 25774 24760 25780 24812
rect 25832 24800 25838 24812
rect 25869 24803 25927 24809
rect 25869 24800 25881 24803
rect 25832 24772 25881 24800
rect 25832 24760 25838 24772
rect 25869 24769 25881 24772
rect 25915 24769 25927 24803
rect 25869 24763 25927 24769
rect 20806 24732 20812 24744
rect 20266 24704 20576 24732
rect 20767 24704 20812 24732
rect 20266 24701 20278 24704
rect 20220 24695 20278 24701
rect 20806 24692 20812 24704
rect 20864 24692 20870 24744
rect 21082 24732 21088 24744
rect 21043 24704 21088 24732
rect 21082 24692 21088 24704
rect 21140 24692 21146 24744
rect 21450 24692 21456 24744
rect 21508 24732 21514 24744
rect 21637 24735 21695 24741
rect 21637 24732 21649 24735
rect 21508 24704 21649 24732
rect 21508 24692 21514 24704
rect 21637 24701 21649 24704
rect 21683 24701 21695 24735
rect 21637 24695 21695 24701
rect 21729 24735 21787 24741
rect 21729 24701 21741 24735
rect 21775 24701 21787 24735
rect 21729 24695 21787 24701
rect 18104 24636 19196 24664
rect 18104 24624 18110 24636
rect 19794 24624 19800 24676
rect 19852 24624 19858 24676
rect 20073 24667 20131 24673
rect 20073 24633 20085 24667
rect 20119 24664 20131 24667
rect 21542 24664 21548 24676
rect 20119 24636 21548 24664
rect 20119 24633 20131 24636
rect 20073 24627 20131 24633
rect 21542 24624 21548 24636
rect 21600 24624 21606 24676
rect 21744 24664 21772 24695
rect 23750 24692 23756 24744
rect 23808 24732 23814 24744
rect 25038 24732 25044 24744
rect 23808 24704 23901 24732
rect 24951 24704 25044 24732
rect 23808 24692 23814 24704
rect 25038 24692 25044 24704
rect 25096 24732 25102 24744
rect 25501 24735 25559 24741
rect 25501 24732 25513 24735
rect 25096 24704 25513 24732
rect 25096 24692 25102 24704
rect 25501 24701 25513 24704
rect 25547 24701 25559 24735
rect 25501 24695 25559 24701
rect 22002 24664 22008 24676
rect 21744 24636 22008 24664
rect 11425 24599 11483 24605
rect 11425 24596 11437 24599
rect 11020 24568 11437 24596
rect 11020 24556 11026 24568
rect 11425 24565 11437 24568
rect 11471 24565 11483 24599
rect 11425 24559 11483 24565
rect 11974 24556 11980 24608
rect 12032 24596 12038 24608
rect 12253 24599 12311 24605
rect 12253 24596 12265 24599
rect 12032 24568 12265 24596
rect 12032 24556 12038 24568
rect 12253 24565 12265 24568
rect 12299 24596 12311 24599
rect 12618 24596 12624 24608
rect 12299 24568 12624 24596
rect 12299 24565 12311 24568
rect 12253 24559 12311 24565
rect 12618 24556 12624 24568
rect 12676 24556 12682 24608
rect 12802 24596 12808 24608
rect 12763 24568 12808 24596
rect 12802 24556 12808 24568
rect 12860 24556 12866 24608
rect 14918 24556 14924 24608
rect 14976 24596 14982 24608
rect 15013 24599 15071 24605
rect 15013 24596 15025 24599
rect 14976 24568 15025 24596
rect 14976 24556 14982 24568
rect 15013 24565 15025 24568
rect 15059 24565 15071 24599
rect 15013 24559 15071 24565
rect 16117 24599 16175 24605
rect 16117 24565 16129 24599
rect 16163 24596 16175 24599
rect 16390 24596 16396 24608
rect 16163 24568 16396 24596
rect 16163 24565 16175 24568
rect 16117 24559 16175 24565
rect 16390 24556 16396 24568
rect 16448 24556 16454 24608
rect 17494 24596 17500 24608
rect 17455 24568 17500 24596
rect 17494 24556 17500 24568
rect 17552 24556 17558 24608
rect 17770 24596 17776 24608
rect 17731 24568 17776 24596
rect 17770 24556 17776 24568
rect 17828 24596 17834 24608
rect 19058 24596 19064 24608
rect 17828 24568 19064 24596
rect 17828 24556 17834 24568
rect 19058 24556 19064 24568
rect 19116 24556 19122 24608
rect 19812 24596 19840 24624
rect 19978 24596 19984 24608
rect 19812 24568 19984 24596
rect 19978 24556 19984 24568
rect 20036 24556 20042 24608
rect 20806 24556 20812 24608
rect 20864 24596 20870 24608
rect 21453 24599 21511 24605
rect 21453 24596 21465 24599
rect 20864 24568 21465 24596
rect 20864 24556 20870 24568
rect 21453 24565 21465 24568
rect 21499 24596 21511 24599
rect 21744 24596 21772 24636
rect 22002 24624 22008 24636
rect 22060 24624 22066 24676
rect 24210 24664 24216 24676
rect 24171 24636 24216 24664
rect 24210 24624 24216 24636
rect 24268 24624 24274 24676
rect 25222 24596 25228 24608
rect 21499 24568 21772 24596
rect 25183 24568 25228 24596
rect 21499 24565 21511 24568
rect 21453 24559 21511 24565
rect 25222 24556 25228 24568
rect 25280 24556 25286 24608
rect 1104 24506 38824 24528
rect 1104 24454 19606 24506
rect 19658 24454 19670 24506
rect 19722 24454 19734 24506
rect 19786 24454 19798 24506
rect 19850 24454 38824 24506
rect 1104 24432 38824 24454
rect 7926 24392 7932 24404
rect 7887 24364 7932 24392
rect 7926 24352 7932 24364
rect 7984 24352 7990 24404
rect 9214 24352 9220 24404
rect 9272 24392 9278 24404
rect 9401 24395 9459 24401
rect 9401 24392 9413 24395
rect 9272 24364 9413 24392
rect 9272 24352 9278 24364
rect 9401 24361 9413 24364
rect 9447 24392 9459 24395
rect 10042 24392 10048 24404
rect 9447 24364 10048 24392
rect 9447 24361 9459 24364
rect 9401 24355 9459 24361
rect 10042 24352 10048 24364
rect 10100 24352 10106 24404
rect 10226 24392 10232 24404
rect 10187 24364 10232 24392
rect 10226 24352 10232 24364
rect 10284 24352 10290 24404
rect 10502 24352 10508 24404
rect 10560 24392 10566 24404
rect 10597 24395 10655 24401
rect 10597 24392 10609 24395
rect 10560 24364 10609 24392
rect 10560 24352 10566 24364
rect 10597 24361 10609 24364
rect 10643 24361 10655 24395
rect 10962 24392 10968 24404
rect 10875 24364 10968 24392
rect 10597 24355 10655 24361
rect 10962 24352 10968 24364
rect 11020 24352 11026 24404
rect 11974 24392 11980 24404
rect 11935 24364 11980 24392
rect 11974 24352 11980 24364
rect 12032 24352 12038 24404
rect 13357 24395 13415 24401
rect 13357 24361 13369 24395
rect 13403 24392 13415 24395
rect 13906 24392 13912 24404
rect 13403 24364 13912 24392
rect 13403 24361 13415 24364
rect 13357 24355 13415 24361
rect 13906 24352 13912 24364
rect 13964 24352 13970 24404
rect 14734 24392 14740 24404
rect 14695 24364 14740 24392
rect 14734 24352 14740 24364
rect 14792 24352 14798 24404
rect 15749 24395 15807 24401
rect 15749 24361 15761 24395
rect 15795 24392 15807 24395
rect 16942 24392 16948 24404
rect 15795 24364 16948 24392
rect 15795 24361 15807 24364
rect 15749 24355 15807 24361
rect 16942 24352 16948 24364
rect 17000 24352 17006 24404
rect 17954 24352 17960 24404
rect 18012 24392 18018 24404
rect 18141 24395 18199 24401
rect 18141 24392 18153 24395
rect 18012 24364 18153 24392
rect 18012 24352 18018 24364
rect 18141 24361 18153 24364
rect 18187 24361 18199 24395
rect 18141 24355 18199 24361
rect 19334 24352 19340 24404
rect 19392 24392 19398 24404
rect 19429 24395 19487 24401
rect 19429 24392 19441 24395
rect 19392 24364 19441 24392
rect 19392 24352 19398 24364
rect 19429 24361 19441 24364
rect 19475 24361 19487 24395
rect 19429 24355 19487 24361
rect 19889 24395 19947 24401
rect 19889 24361 19901 24395
rect 19935 24392 19947 24395
rect 19978 24392 19984 24404
rect 19935 24364 19984 24392
rect 19935 24361 19947 24364
rect 19889 24355 19947 24361
rect 19978 24352 19984 24364
rect 20036 24352 20042 24404
rect 20622 24392 20628 24404
rect 20583 24364 20628 24392
rect 20622 24352 20628 24364
rect 20680 24392 20686 24404
rect 21085 24395 21143 24401
rect 21085 24392 21097 24395
rect 20680 24364 21097 24392
rect 20680 24352 20686 24364
rect 21085 24361 21097 24364
rect 21131 24361 21143 24395
rect 21450 24392 21456 24404
rect 21085 24355 21143 24361
rect 21192 24364 21456 24392
rect 10244 24324 10272 24352
rect 10980 24324 11008 24352
rect 13630 24324 13636 24336
rect 10244 24296 11008 24324
rect 13591 24296 13636 24324
rect 13630 24284 13636 24296
rect 13688 24284 13694 24336
rect 14369 24327 14427 24333
rect 14369 24293 14381 24327
rect 14415 24324 14427 24327
rect 15286 24324 15292 24336
rect 14415 24296 15292 24324
rect 14415 24293 14427 24296
rect 14369 24287 14427 24293
rect 15286 24284 15292 24296
rect 15344 24284 15350 24336
rect 17494 24284 17500 24336
rect 17552 24324 17558 24336
rect 18782 24324 18788 24336
rect 17552 24296 18788 24324
rect 17552 24284 17558 24296
rect 18782 24284 18788 24296
rect 18840 24324 18846 24336
rect 18840 24296 18920 24324
rect 18840 24284 18846 24296
rect 8110 24256 8116 24268
rect 8071 24228 8116 24256
rect 8110 24216 8116 24228
rect 8168 24216 8174 24268
rect 10781 24259 10839 24265
rect 10781 24225 10793 24259
rect 10827 24256 10839 24259
rect 10870 24256 10876 24268
rect 10827 24228 10876 24256
rect 10827 24225 10839 24228
rect 10781 24219 10839 24225
rect 10870 24216 10876 24228
rect 10928 24216 10934 24268
rect 11793 24259 11851 24265
rect 11793 24225 11805 24259
rect 11839 24256 11851 24259
rect 12526 24256 12532 24268
rect 11839 24228 12532 24256
rect 11839 24225 11851 24228
rect 11793 24219 11851 24225
rect 12526 24216 12532 24228
rect 12584 24216 12590 24268
rect 12802 24256 12808 24268
rect 12763 24228 12808 24256
rect 12802 24216 12808 24228
rect 12860 24216 12866 24268
rect 12894 24216 12900 24268
rect 12952 24256 12958 24268
rect 13906 24256 13912 24268
rect 12952 24228 13912 24256
rect 12952 24216 12958 24228
rect 13906 24216 13912 24228
rect 13964 24216 13970 24268
rect 15194 24216 15200 24268
rect 15252 24256 15258 24268
rect 16025 24259 16083 24265
rect 16025 24256 16037 24259
rect 15252 24228 16037 24256
rect 15252 24216 15258 24228
rect 16025 24225 16037 24228
rect 16071 24225 16083 24259
rect 16025 24219 16083 24225
rect 16390 24216 16396 24268
rect 16448 24256 16454 24268
rect 16485 24259 16543 24265
rect 16485 24256 16497 24259
rect 16448 24228 16497 24256
rect 16448 24216 16454 24228
rect 16485 24225 16497 24228
rect 16531 24225 16543 24259
rect 16485 24219 16543 24225
rect 16577 24259 16635 24265
rect 16577 24225 16589 24259
rect 16623 24256 16635 24259
rect 16666 24256 16672 24268
rect 16623 24228 16672 24256
rect 16623 24225 16635 24228
rect 16577 24219 16635 24225
rect 16666 24216 16672 24228
rect 16724 24216 16730 24268
rect 17586 24256 17592 24268
rect 17547 24228 17592 24256
rect 17586 24216 17592 24228
rect 17644 24216 17650 24268
rect 17862 24216 17868 24268
rect 17920 24256 17926 24268
rect 18892 24265 18920 24296
rect 18966 24284 18972 24336
rect 19024 24324 19030 24336
rect 21192 24324 21220 24364
rect 21450 24352 21456 24364
rect 21508 24352 21514 24404
rect 21542 24352 21548 24404
rect 21600 24392 21606 24404
rect 21913 24395 21971 24401
rect 21913 24392 21925 24395
rect 21600 24364 21925 24392
rect 21600 24352 21606 24364
rect 21913 24361 21925 24364
rect 21959 24361 21971 24395
rect 21913 24355 21971 24361
rect 22462 24352 22468 24404
rect 22520 24392 22526 24404
rect 22741 24395 22799 24401
rect 22741 24392 22753 24395
rect 22520 24364 22753 24392
rect 22520 24352 22526 24364
rect 22741 24361 22753 24364
rect 22787 24361 22799 24395
rect 22741 24355 22799 24361
rect 23106 24352 23112 24404
rect 23164 24392 23170 24404
rect 23293 24395 23351 24401
rect 23293 24392 23305 24395
rect 23164 24364 23305 24392
rect 23164 24352 23170 24364
rect 23293 24361 23305 24364
rect 23339 24361 23351 24395
rect 23750 24392 23756 24404
rect 23663 24364 23756 24392
rect 23293 24355 23351 24361
rect 23750 24352 23756 24364
rect 23808 24392 23814 24404
rect 24670 24392 24676 24404
rect 23808 24364 24676 24392
rect 23808 24352 23814 24364
rect 24670 24352 24676 24364
rect 24728 24352 24734 24404
rect 24765 24395 24823 24401
rect 24765 24361 24777 24395
rect 24811 24392 24823 24395
rect 24854 24392 24860 24404
rect 24811 24364 24860 24392
rect 24811 24361 24823 24364
rect 24765 24355 24823 24361
rect 24854 24352 24860 24364
rect 24912 24352 24918 24404
rect 19024 24296 21220 24324
rect 21269 24327 21327 24333
rect 19024 24284 19030 24296
rect 21269 24293 21281 24327
rect 21315 24324 21327 24327
rect 22002 24324 22008 24336
rect 21315 24296 22008 24324
rect 21315 24293 21327 24296
rect 21269 24287 21327 24293
rect 22002 24284 22008 24296
rect 22060 24284 22066 24336
rect 24397 24327 24455 24333
rect 24397 24293 24409 24327
rect 24443 24324 24455 24327
rect 25038 24324 25044 24336
rect 24443 24296 25044 24324
rect 24443 24293 24455 24296
rect 24397 24287 24455 24293
rect 25038 24284 25044 24296
rect 25096 24284 25102 24336
rect 18049 24259 18107 24265
rect 18049 24256 18061 24259
rect 17920 24228 18061 24256
rect 17920 24216 17926 24228
rect 18049 24225 18061 24228
rect 18095 24225 18107 24259
rect 18049 24219 18107 24225
rect 18877 24259 18935 24265
rect 18877 24225 18889 24259
rect 18923 24225 18935 24259
rect 18877 24219 18935 24225
rect 19061 24259 19119 24265
rect 19061 24225 19073 24259
rect 19107 24256 19119 24259
rect 19978 24256 19984 24268
rect 19107 24228 19984 24256
rect 19107 24225 19119 24228
rect 19061 24219 19119 24225
rect 19978 24216 19984 24228
rect 20036 24216 20042 24268
rect 20714 24216 20720 24268
rect 20772 24256 20778 24268
rect 21177 24259 21235 24265
rect 20772 24228 21036 24256
rect 20772 24216 20778 24228
rect 7650 24148 7656 24200
rect 7708 24188 7714 24200
rect 8478 24188 8484 24200
rect 7708 24160 8484 24188
rect 7708 24148 7714 24160
rect 8478 24148 8484 24160
rect 8536 24148 8542 24200
rect 8754 24148 8760 24200
rect 8812 24188 8818 24200
rect 9582 24188 9588 24200
rect 8812 24160 9588 24188
rect 8812 24148 8818 24160
rect 9582 24148 9588 24160
rect 9640 24148 9646 24200
rect 11146 24148 11152 24200
rect 11204 24188 11210 24200
rect 11609 24191 11667 24197
rect 11609 24188 11621 24191
rect 11204 24160 11621 24188
rect 11204 24148 11210 24160
rect 11609 24157 11621 24160
rect 11655 24188 11667 24191
rect 13081 24191 13139 24197
rect 13081 24188 13093 24191
rect 11655 24160 13093 24188
rect 11655 24157 11667 24160
rect 11609 24151 11667 24157
rect 13081 24157 13093 24160
rect 13127 24157 13139 24191
rect 13081 24151 13139 24157
rect 13817 24191 13875 24197
rect 13817 24157 13829 24191
rect 13863 24188 13875 24191
rect 14550 24188 14556 24200
rect 13863 24160 14556 24188
rect 13863 24157 13875 24160
rect 13817 24151 13875 24157
rect 14550 24148 14556 24160
rect 14608 24188 14614 24200
rect 14826 24188 14832 24200
rect 14608 24160 14832 24188
rect 14608 24148 14614 24160
rect 14826 24148 14832 24160
rect 14884 24148 14890 24200
rect 15838 24188 15844 24200
rect 15799 24160 15844 24188
rect 15838 24148 15844 24160
rect 15896 24148 15902 24200
rect 20898 24188 20904 24200
rect 20272 24160 20904 24188
rect 9953 24123 10011 24129
rect 9953 24089 9965 24123
rect 9999 24120 10011 24123
rect 10778 24120 10784 24132
rect 9999 24092 10784 24120
rect 9999 24089 10011 24092
rect 9953 24083 10011 24089
rect 10778 24080 10784 24092
rect 10836 24120 10842 24132
rect 12529 24123 12587 24129
rect 12529 24120 12541 24123
rect 10836 24092 12541 24120
rect 10836 24080 10842 24092
rect 12529 24089 12541 24092
rect 12575 24120 12587 24123
rect 13722 24120 13728 24132
rect 12575 24092 13728 24120
rect 12575 24089 12587 24092
rect 12529 24083 12587 24089
rect 13722 24080 13728 24092
rect 13780 24080 13786 24132
rect 16574 24080 16580 24132
rect 16632 24120 16638 24132
rect 16945 24123 17003 24129
rect 16945 24120 16957 24123
rect 16632 24092 16957 24120
rect 16632 24080 16638 24092
rect 16945 24089 16957 24092
rect 16991 24089 17003 24123
rect 16945 24083 17003 24089
rect 19334 24080 19340 24132
rect 19392 24120 19398 24132
rect 20272 24129 20300 24160
rect 20898 24148 20904 24160
rect 20956 24148 20962 24200
rect 21008 24188 21036 24228
rect 21177 24225 21189 24259
rect 21223 24256 21235 24259
rect 21542 24256 21548 24268
rect 21223 24228 21548 24256
rect 21223 24225 21235 24228
rect 21177 24219 21235 24225
rect 21542 24216 21548 24228
rect 21600 24216 21606 24268
rect 22186 24216 22192 24268
rect 22244 24256 22250 24268
rect 22462 24256 22468 24268
rect 22244 24228 22468 24256
rect 22244 24216 22250 24228
rect 22462 24216 22468 24228
rect 22520 24216 22526 24268
rect 22554 24216 22560 24268
rect 22612 24256 22618 24268
rect 22649 24259 22707 24265
rect 22649 24256 22661 24259
rect 22612 24228 22661 24256
rect 22612 24216 22618 24228
rect 22649 24225 22661 24228
rect 22695 24256 22707 24259
rect 23382 24256 23388 24268
rect 22695 24228 23388 24256
rect 22695 24225 22707 24228
rect 22649 24219 22707 24225
rect 23382 24216 23388 24228
rect 23440 24216 23446 24268
rect 23474 24216 23480 24268
rect 23532 24256 23538 24268
rect 23937 24259 23995 24265
rect 23937 24256 23949 24259
rect 23532 24228 23949 24256
rect 23532 24216 23538 24228
rect 23937 24225 23949 24228
rect 23983 24256 23995 24259
rect 24210 24256 24216 24268
rect 23983 24228 24216 24256
rect 23983 24225 23995 24228
rect 23937 24219 23995 24225
rect 24210 24216 24216 24228
rect 24268 24216 24274 24268
rect 25222 24256 25228 24268
rect 25183 24228 25228 24256
rect 25222 24216 25228 24228
rect 25280 24216 25286 24268
rect 21637 24191 21695 24197
rect 21637 24188 21649 24191
rect 21008 24160 21649 24188
rect 21637 24157 21649 24160
rect 21683 24157 21695 24191
rect 21637 24151 21695 24157
rect 21910 24148 21916 24200
rect 21968 24188 21974 24200
rect 22281 24191 22339 24197
rect 22281 24188 22293 24191
rect 21968 24160 22293 24188
rect 21968 24148 21974 24160
rect 22281 24157 22293 24160
rect 22327 24157 22339 24191
rect 22281 24151 22339 24157
rect 23566 24148 23572 24200
rect 23624 24188 23630 24200
rect 23845 24191 23903 24197
rect 23845 24188 23857 24191
rect 23624 24160 23857 24188
rect 23624 24148 23630 24160
rect 23845 24157 23857 24160
rect 23891 24157 23903 24191
rect 23845 24151 23903 24157
rect 20257 24123 20315 24129
rect 20257 24120 20269 24123
rect 19392 24092 20269 24120
rect 19392 24080 19398 24092
rect 20257 24089 20269 24092
rect 20303 24089 20315 24123
rect 20257 24083 20315 24089
rect 23934 24080 23940 24132
rect 23992 24120 23998 24132
rect 25590 24120 25596 24132
rect 23992 24092 25596 24120
rect 23992 24080 23998 24092
rect 25590 24080 25596 24092
rect 25648 24120 25654 24132
rect 25685 24123 25743 24129
rect 25685 24120 25697 24123
rect 25648 24092 25697 24120
rect 25648 24080 25654 24092
rect 25685 24089 25697 24092
rect 25731 24089 25743 24123
rect 25685 24083 25743 24089
rect 11330 24052 11336 24064
rect 11291 24024 11336 24052
rect 11330 24012 11336 24024
rect 11388 24012 11394 24064
rect 12986 24052 12992 24064
rect 12947 24024 12992 24052
rect 12986 24012 12992 24024
rect 13044 24012 13050 24064
rect 13081 24055 13139 24061
rect 13081 24021 13093 24055
rect 13127 24052 13139 24055
rect 14366 24052 14372 24064
rect 13127 24024 14372 24052
rect 13127 24021 13139 24024
rect 13081 24015 13139 24021
rect 14366 24012 14372 24024
rect 14424 24012 14430 24064
rect 15102 24052 15108 24064
rect 15063 24024 15108 24052
rect 15102 24012 15108 24024
rect 15160 24012 15166 24064
rect 17954 24052 17960 24064
rect 17915 24024 17960 24052
rect 17954 24012 17960 24024
rect 18012 24012 18018 24064
rect 22462 24012 22468 24064
rect 22520 24052 22526 24064
rect 25041 24055 25099 24061
rect 25041 24052 25053 24055
rect 22520 24024 25053 24052
rect 22520 24012 22526 24024
rect 25041 24021 25053 24024
rect 25087 24021 25099 24055
rect 25406 24052 25412 24064
rect 25367 24024 25412 24052
rect 25041 24015 25099 24021
rect 25406 24012 25412 24024
rect 25464 24012 25470 24064
rect 1104 23962 38824 23984
rect 1104 23910 4246 23962
rect 4298 23910 4310 23962
rect 4362 23910 4374 23962
rect 4426 23910 4438 23962
rect 4490 23910 34966 23962
rect 35018 23910 35030 23962
rect 35082 23910 35094 23962
rect 35146 23910 35158 23962
rect 35210 23910 38824 23962
rect 1104 23888 38824 23910
rect 3605 23851 3663 23857
rect 3605 23817 3617 23851
rect 3651 23848 3663 23851
rect 7006 23848 7012 23860
rect 3651 23820 7012 23848
rect 3651 23817 3663 23820
rect 3605 23811 3663 23817
rect 7006 23808 7012 23820
rect 7064 23808 7070 23860
rect 8021 23851 8079 23857
rect 8021 23817 8033 23851
rect 8067 23848 8079 23851
rect 8110 23848 8116 23860
rect 8067 23820 8116 23848
rect 8067 23817 8079 23820
rect 8021 23811 8079 23817
rect 8110 23808 8116 23820
rect 8168 23808 8174 23860
rect 10870 23808 10876 23860
rect 10928 23848 10934 23860
rect 11793 23851 11851 23857
rect 11793 23848 11805 23851
rect 10928 23820 11805 23848
rect 10928 23808 10934 23820
rect 11793 23817 11805 23820
rect 11839 23848 11851 23851
rect 12434 23848 12440 23860
rect 11839 23820 12440 23848
rect 11839 23817 11851 23820
rect 11793 23811 11851 23817
rect 12434 23808 12440 23820
rect 12492 23848 12498 23860
rect 13814 23848 13820 23860
rect 12492 23820 13676 23848
rect 13775 23820 13820 23848
rect 12492 23808 12498 23820
rect 12253 23783 12311 23789
rect 12253 23749 12265 23783
rect 12299 23780 12311 23783
rect 12342 23780 12348 23792
rect 12299 23752 12348 23780
rect 12299 23749 12311 23752
rect 12253 23743 12311 23749
rect 12342 23740 12348 23752
rect 12400 23740 12406 23792
rect 13648 23780 13676 23820
rect 13814 23808 13820 23820
rect 13872 23808 13878 23860
rect 13906 23808 13912 23860
rect 13964 23848 13970 23860
rect 14461 23851 14519 23857
rect 14461 23848 14473 23851
rect 13964 23820 14473 23848
rect 13964 23808 13970 23820
rect 14461 23817 14473 23820
rect 14507 23848 14519 23851
rect 15102 23848 15108 23860
rect 14507 23820 15108 23848
rect 14507 23817 14519 23820
rect 14461 23811 14519 23817
rect 15102 23808 15108 23820
rect 15160 23808 15166 23860
rect 16758 23848 16764 23860
rect 16719 23820 16764 23848
rect 16758 23808 16764 23820
rect 16816 23808 16822 23860
rect 17862 23848 17868 23860
rect 17823 23820 17868 23848
rect 17862 23808 17868 23820
rect 17920 23808 17926 23860
rect 18322 23808 18328 23860
rect 18380 23848 18386 23860
rect 19981 23851 20039 23857
rect 19981 23848 19993 23851
rect 18380 23820 19993 23848
rect 18380 23808 18386 23820
rect 19981 23817 19993 23820
rect 20027 23848 20039 23851
rect 21542 23848 21548 23860
rect 20027 23820 21548 23848
rect 20027 23817 20039 23820
rect 19981 23811 20039 23817
rect 21542 23808 21548 23820
rect 21600 23808 21606 23860
rect 22554 23848 22560 23860
rect 22515 23820 22560 23848
rect 22554 23808 22560 23820
rect 22612 23808 22618 23860
rect 22925 23851 22983 23857
rect 22925 23817 22937 23851
rect 22971 23848 22983 23851
rect 23290 23848 23296 23860
rect 22971 23820 23296 23848
rect 22971 23817 22983 23820
rect 22925 23811 22983 23817
rect 23290 23808 23296 23820
rect 23348 23808 23354 23860
rect 23842 23848 23848 23860
rect 23803 23820 23848 23848
rect 23842 23808 23848 23820
rect 23900 23808 23906 23860
rect 24210 23848 24216 23860
rect 24171 23820 24216 23848
rect 24210 23808 24216 23820
rect 24268 23808 24274 23860
rect 26234 23808 26240 23860
rect 26292 23848 26298 23860
rect 26329 23851 26387 23857
rect 26329 23848 26341 23851
rect 26292 23820 26341 23848
rect 26292 23808 26298 23820
rect 26329 23817 26341 23820
rect 26375 23817 26387 23851
rect 26329 23811 26387 23817
rect 14182 23780 14188 23792
rect 13648 23752 14188 23780
rect 14182 23740 14188 23752
rect 14240 23740 14246 23792
rect 16025 23783 16083 23789
rect 16025 23749 16037 23783
rect 16071 23780 16083 23783
rect 16666 23780 16672 23792
rect 16071 23752 16672 23780
rect 16071 23749 16083 23752
rect 16025 23743 16083 23749
rect 16666 23740 16672 23752
rect 16724 23780 16730 23792
rect 17586 23780 17592 23792
rect 16724 23752 17592 23780
rect 16724 23740 16730 23752
rect 17586 23740 17592 23752
rect 17644 23740 17650 23792
rect 19518 23740 19524 23792
rect 19576 23780 19582 23792
rect 21634 23780 21640 23792
rect 19576 23752 21640 23780
rect 19576 23740 19582 23752
rect 21634 23740 21640 23752
rect 21692 23740 21698 23792
rect 2038 23712 2044 23724
rect 1999 23684 2044 23712
rect 2038 23672 2044 23684
rect 2096 23672 2102 23724
rect 9674 23672 9680 23724
rect 9732 23712 9738 23724
rect 10045 23715 10103 23721
rect 10045 23712 10057 23715
rect 9732 23684 10057 23712
rect 9732 23672 9738 23684
rect 10045 23681 10057 23684
rect 10091 23681 10103 23715
rect 10045 23675 10103 23681
rect 11330 23672 11336 23724
rect 11388 23712 11394 23724
rect 12437 23715 12495 23721
rect 12437 23712 12449 23715
rect 11388 23684 12449 23712
rect 11388 23672 11394 23684
rect 12437 23681 12449 23684
rect 12483 23712 12495 23715
rect 13630 23712 13636 23724
rect 12483 23684 13636 23712
rect 12483 23681 12495 23684
rect 12437 23675 12495 23681
rect 13630 23672 13636 23684
rect 13688 23672 13694 23724
rect 14829 23715 14887 23721
rect 14829 23681 14841 23715
rect 14875 23712 14887 23715
rect 14875 23684 15608 23712
rect 14875 23681 14887 23684
rect 14829 23675 14887 23681
rect 15580 23656 15608 23684
rect 16206 23672 16212 23724
rect 16264 23712 16270 23724
rect 16485 23715 16543 23721
rect 16485 23712 16497 23715
rect 16264 23684 16497 23712
rect 16264 23672 16270 23684
rect 16485 23681 16497 23684
rect 16531 23681 16543 23715
rect 16485 23675 16543 23681
rect 17954 23672 17960 23724
rect 18012 23712 18018 23724
rect 20714 23712 20720 23724
rect 18012 23684 19196 23712
rect 20675 23684 20720 23712
rect 18012 23672 18018 23684
rect 2317 23647 2375 23653
rect 2317 23644 2329 23647
rect 1872 23616 2329 23644
rect 1762 23468 1768 23520
rect 1820 23508 1826 23520
rect 1872 23517 1900 23616
rect 2317 23613 2329 23616
rect 2363 23613 2375 23647
rect 2317 23607 2375 23613
rect 9769 23647 9827 23653
rect 9769 23613 9781 23647
rect 9815 23644 9827 23647
rect 9815 23616 9849 23644
rect 9815 23613 9827 23616
rect 9769 23607 9827 23613
rect 8662 23536 8668 23588
rect 8720 23576 8726 23588
rect 9309 23579 9367 23585
rect 9309 23576 9321 23579
rect 8720 23548 9321 23576
rect 8720 23536 8726 23548
rect 9309 23545 9321 23548
rect 9355 23576 9367 23579
rect 9784 23576 9812 23607
rect 12526 23604 12532 23656
rect 12584 23644 12590 23656
rect 12713 23647 12771 23653
rect 12713 23644 12725 23647
rect 12584 23616 12725 23644
rect 12584 23604 12590 23616
rect 12713 23613 12725 23616
rect 12759 23613 12771 23647
rect 12713 23607 12771 23613
rect 12802 23604 12808 23656
rect 12860 23644 12866 23656
rect 14918 23644 14924 23656
rect 12860 23616 14924 23644
rect 12860 23604 12866 23616
rect 14918 23604 14924 23616
rect 14976 23604 14982 23656
rect 15562 23644 15568 23656
rect 15523 23616 15568 23644
rect 15562 23604 15568 23616
rect 15620 23604 15626 23656
rect 9858 23576 9864 23588
rect 9355 23548 9864 23576
rect 9355 23545 9367 23548
rect 9309 23539 9367 23545
rect 9858 23536 9864 23548
rect 9916 23536 9922 23588
rect 15102 23536 15108 23588
rect 15160 23576 15166 23588
rect 16224 23576 16252 23672
rect 19168 23656 19196 23684
rect 20714 23672 20720 23684
rect 20772 23672 20778 23724
rect 21450 23712 21456 23724
rect 21284 23684 21456 23712
rect 16574 23604 16580 23656
rect 16632 23644 16638 23656
rect 18506 23644 18512 23656
rect 16632 23616 16677 23644
rect 18467 23616 18512 23644
rect 16632 23604 16638 23616
rect 18506 23604 18512 23616
rect 18564 23604 18570 23656
rect 18693 23647 18751 23653
rect 18693 23613 18705 23647
rect 18739 23613 18751 23647
rect 19150 23644 19156 23656
rect 19111 23616 19156 23644
rect 18693 23607 18751 23613
rect 15160 23548 16252 23576
rect 17497 23579 17555 23585
rect 15160 23536 15166 23548
rect 17497 23545 17509 23579
rect 17543 23576 17555 23579
rect 18708 23576 18736 23607
rect 19150 23604 19156 23616
rect 19208 23604 19214 23656
rect 19426 23644 19432 23656
rect 19387 23616 19432 23644
rect 19426 23604 19432 23616
rect 19484 23604 19490 23656
rect 20809 23647 20867 23653
rect 20809 23613 20821 23647
rect 20855 23644 20867 23647
rect 20898 23644 20904 23656
rect 20855 23616 20904 23644
rect 20855 23613 20867 23616
rect 20809 23607 20867 23613
rect 20898 23604 20904 23616
rect 20956 23604 20962 23656
rect 21284 23653 21312 23684
rect 21450 23672 21456 23684
rect 21508 23672 21514 23724
rect 24673 23715 24731 23721
rect 24673 23681 24685 23715
rect 24719 23712 24731 23715
rect 24719 23684 25084 23712
rect 24719 23681 24731 23684
rect 24673 23675 24731 23681
rect 25056 23656 25084 23684
rect 21269 23647 21327 23653
rect 21269 23613 21281 23647
rect 21315 23613 21327 23647
rect 21542 23644 21548 23656
rect 21503 23616 21548 23644
rect 21269 23607 21327 23613
rect 21542 23604 21548 23616
rect 21600 23604 21606 23656
rect 21729 23647 21787 23653
rect 21729 23613 21741 23647
rect 21775 23613 21787 23647
rect 21729 23607 21787 23613
rect 23477 23647 23535 23653
rect 23477 23613 23489 23647
rect 23523 23644 23535 23647
rect 23658 23644 23664 23656
rect 23523 23616 23664 23644
rect 23523 23613 23535 23616
rect 23477 23607 23535 23613
rect 18874 23576 18880 23588
rect 17543 23548 18880 23576
rect 17543 23545 17555 23548
rect 17497 23539 17555 23545
rect 18874 23536 18880 23548
rect 18932 23536 18938 23588
rect 20441 23579 20499 23585
rect 20441 23545 20453 23579
rect 20487 23576 20499 23579
rect 20990 23576 20996 23588
rect 20487 23548 20996 23576
rect 20487 23545 20499 23548
rect 20441 23539 20499 23545
rect 20990 23536 20996 23548
rect 21048 23576 21054 23588
rect 21744 23576 21772 23607
rect 23658 23604 23664 23616
rect 23716 23604 23722 23656
rect 23934 23604 23940 23656
rect 23992 23644 23998 23656
rect 24765 23647 24823 23653
rect 24765 23644 24777 23647
rect 23992 23616 24777 23644
rect 23992 23604 23998 23616
rect 24765 23613 24777 23616
rect 24811 23613 24823 23647
rect 25038 23644 25044 23656
rect 24999 23616 25044 23644
rect 24765 23607 24823 23613
rect 25038 23604 25044 23616
rect 25096 23604 25102 23656
rect 21910 23576 21916 23588
rect 21048 23548 21916 23576
rect 21048 23536 21054 23548
rect 21910 23536 21916 23548
rect 21968 23536 21974 23588
rect 1857 23511 1915 23517
rect 1857 23508 1869 23511
rect 1820 23480 1869 23508
rect 1820 23468 1826 23480
rect 1857 23477 1869 23480
rect 1903 23477 1915 23511
rect 9674 23508 9680 23520
rect 9635 23480 9680 23508
rect 1857 23471 1915 23477
rect 9674 23468 9680 23480
rect 9732 23468 9738 23520
rect 11146 23508 11152 23520
rect 11107 23480 11152 23508
rect 11146 23468 11152 23480
rect 11204 23468 11210 23520
rect 15654 23468 15660 23520
rect 15712 23508 15718 23520
rect 16206 23508 16212 23520
rect 15712 23480 16212 23508
rect 15712 23468 15718 23480
rect 16206 23468 16212 23480
rect 16264 23468 16270 23520
rect 16390 23508 16396 23520
rect 16351 23480 16396 23508
rect 16390 23468 16396 23480
rect 16448 23468 16454 23520
rect 19242 23468 19248 23520
rect 19300 23508 19306 23520
rect 19429 23511 19487 23517
rect 19429 23508 19441 23511
rect 19300 23480 19441 23508
rect 19300 23468 19306 23480
rect 19429 23477 19441 23480
rect 19475 23477 19487 23511
rect 19429 23471 19487 23477
rect 21542 23468 21548 23520
rect 21600 23508 21606 23520
rect 22186 23508 22192 23520
rect 21600 23480 22192 23508
rect 21600 23468 21606 23480
rect 22186 23468 22192 23480
rect 22244 23468 22250 23520
rect 1104 23418 38824 23440
rect 1104 23366 19606 23418
rect 19658 23366 19670 23418
rect 19722 23366 19734 23418
rect 19786 23366 19798 23418
rect 19850 23366 38824 23418
rect 1104 23344 38824 23366
rect 2038 23304 2044 23316
rect 1999 23276 2044 23304
rect 2038 23264 2044 23276
rect 2096 23264 2102 23316
rect 11146 23264 11152 23316
rect 11204 23264 11210 23316
rect 12802 23304 12808 23316
rect 12763 23276 12808 23304
rect 12802 23264 12808 23276
rect 12860 23264 12866 23316
rect 14090 23264 14096 23316
rect 14148 23304 14154 23316
rect 15013 23307 15071 23313
rect 15013 23304 15025 23307
rect 14148 23276 15025 23304
rect 14148 23264 14154 23276
rect 15013 23273 15025 23276
rect 15059 23273 15071 23307
rect 15013 23267 15071 23273
rect 16298 23264 16304 23316
rect 16356 23304 16362 23316
rect 16574 23304 16580 23316
rect 16356 23276 16580 23304
rect 16356 23264 16362 23276
rect 16574 23264 16580 23276
rect 16632 23264 16638 23316
rect 18325 23307 18383 23313
rect 18325 23273 18337 23307
rect 18371 23304 18383 23307
rect 18506 23304 18512 23316
rect 18371 23276 18512 23304
rect 18371 23273 18383 23276
rect 18325 23267 18383 23273
rect 18506 23264 18512 23276
rect 18564 23304 18570 23316
rect 18564 23276 21680 23304
rect 18564 23264 18570 23276
rect 11164 23236 11192 23264
rect 14826 23236 14832 23248
rect 11164 23208 11284 23236
rect 10962 23128 10968 23180
rect 11020 23168 11026 23180
rect 11149 23171 11207 23177
rect 11149 23168 11161 23171
rect 11020 23140 11161 23168
rect 11020 23128 11026 23140
rect 11149 23137 11161 23140
rect 11195 23137 11207 23171
rect 11256 23168 11284 23208
rect 13832 23208 14832 23236
rect 11471 23171 11529 23177
rect 11471 23168 11483 23171
rect 11256 23140 11483 23168
rect 11149 23131 11207 23137
rect 11471 23137 11483 23140
rect 11517 23137 11529 23171
rect 11606 23168 11612 23180
rect 11567 23140 11612 23168
rect 11471 23131 11529 23137
rect 11606 23128 11612 23140
rect 11664 23128 11670 23180
rect 13354 23128 13360 23180
rect 13412 23168 13418 23180
rect 13832 23177 13860 23208
rect 14826 23196 14832 23208
rect 14884 23196 14890 23248
rect 13817 23171 13875 23177
rect 13817 23168 13829 23171
rect 13412 23140 13829 23168
rect 13412 23128 13418 23140
rect 13817 23137 13829 23140
rect 13863 23137 13875 23171
rect 13817 23131 13875 23137
rect 13998 23128 14004 23180
rect 14056 23168 14062 23180
rect 14185 23171 14243 23177
rect 14185 23168 14197 23171
rect 14056 23140 14197 23168
rect 14056 23128 14062 23140
rect 14185 23137 14197 23140
rect 14231 23137 14243 23171
rect 14185 23131 14243 23137
rect 15473 23171 15531 23177
rect 15473 23137 15485 23171
rect 15519 23168 15531 23171
rect 15562 23168 15568 23180
rect 15519 23140 15568 23168
rect 15519 23137 15531 23140
rect 15473 23131 15531 23137
rect 15562 23128 15568 23140
rect 15620 23168 15626 23180
rect 16316 23168 16344 23264
rect 18782 23236 18788 23248
rect 18743 23208 18788 23236
rect 18782 23196 18788 23208
rect 18840 23196 18846 23248
rect 20806 23236 20812 23248
rect 19812 23208 20812 23236
rect 19812 23180 19840 23208
rect 20806 23196 20812 23208
rect 20864 23196 20870 23248
rect 21269 23239 21327 23245
rect 21269 23205 21281 23239
rect 21315 23236 21327 23239
rect 21542 23236 21548 23248
rect 21315 23208 21548 23236
rect 21315 23205 21327 23208
rect 21269 23199 21327 23205
rect 21542 23196 21548 23208
rect 21600 23196 21606 23248
rect 21652 23245 21680 23276
rect 21726 23264 21732 23316
rect 21784 23304 21790 23316
rect 22281 23307 22339 23313
rect 22281 23304 22293 23307
rect 21784 23276 22293 23304
rect 21784 23264 21790 23276
rect 22281 23273 22293 23276
rect 22327 23273 22339 23307
rect 22281 23267 22339 23273
rect 23661 23307 23719 23313
rect 23661 23273 23673 23307
rect 23707 23273 23719 23307
rect 25590 23304 25596 23316
rect 25551 23276 25596 23304
rect 23661 23267 23719 23273
rect 21637 23239 21695 23245
rect 21637 23205 21649 23239
rect 21683 23205 21695 23239
rect 21637 23199 21695 23205
rect 21821 23239 21879 23245
rect 21821 23205 21833 23239
rect 21867 23236 21879 23239
rect 23676 23236 23704 23267
rect 25590 23264 25596 23276
rect 25648 23264 25654 23316
rect 21867 23208 23704 23236
rect 21867 23205 21879 23208
rect 21821 23199 21879 23205
rect 17218 23168 17224 23180
rect 15620 23140 16344 23168
rect 17179 23140 17224 23168
rect 15620 23128 15626 23140
rect 17218 23128 17224 23140
rect 17276 23128 17282 23180
rect 17494 23128 17500 23180
rect 17552 23168 17558 23180
rect 17589 23171 17647 23177
rect 17589 23168 17601 23171
rect 17552 23140 17601 23168
rect 17552 23128 17558 23140
rect 17589 23137 17601 23140
rect 17635 23137 17647 23171
rect 19426 23168 19432 23180
rect 19387 23140 19432 23168
rect 17589 23131 17647 23137
rect 19426 23128 19432 23140
rect 19484 23128 19490 23180
rect 19794 23168 19800 23180
rect 19755 23140 19800 23168
rect 19794 23128 19800 23140
rect 19852 23128 19858 23180
rect 19886 23128 19892 23180
rect 19944 23168 19950 23180
rect 19944 23140 19989 23168
rect 19944 23128 19950 23140
rect 20622 23128 20628 23180
rect 20680 23168 20686 23180
rect 21085 23171 21143 23177
rect 21085 23168 21097 23171
rect 20680 23140 21097 23168
rect 20680 23128 20686 23140
rect 21085 23137 21097 23140
rect 21131 23137 21143 23171
rect 21085 23131 21143 23137
rect 21177 23171 21235 23177
rect 21177 23137 21189 23171
rect 21223 23168 21235 23171
rect 21358 23168 21364 23180
rect 21223 23140 21364 23168
rect 21223 23137 21235 23140
rect 21177 23131 21235 23137
rect 10594 23100 10600 23112
rect 10555 23072 10600 23100
rect 10594 23060 10600 23072
rect 10652 23060 10658 23112
rect 11241 23103 11299 23109
rect 11241 23069 11253 23103
rect 11287 23069 11299 23103
rect 13262 23100 13268 23112
rect 13223 23072 13268 23100
rect 11241 23063 11299 23069
rect 10778 22992 10784 23044
rect 10836 23032 10842 23044
rect 11256 23032 11284 23063
rect 13262 23060 13268 23072
rect 13320 23060 13326 23112
rect 13906 23100 13912 23112
rect 13867 23072 13912 23100
rect 13906 23060 13912 23072
rect 13964 23060 13970 23112
rect 14093 23103 14151 23109
rect 14093 23069 14105 23103
rect 14139 23069 14151 23103
rect 14093 23063 14151 23069
rect 12618 23032 12624 23044
rect 10836 23004 12624 23032
rect 10836 22992 10842 23004
rect 12618 22992 12624 23004
rect 12676 23032 12682 23044
rect 13170 23032 13176 23044
rect 12676 23004 13176 23032
rect 12676 22992 12682 23004
rect 13170 22992 13176 23004
rect 13228 22992 13234 23044
rect 13722 22992 13728 23044
rect 13780 23032 13786 23044
rect 14108 23032 14136 23063
rect 15286 23060 15292 23112
rect 15344 23100 15350 23112
rect 15381 23103 15439 23109
rect 15381 23100 15393 23103
rect 15344 23072 15393 23100
rect 15344 23060 15350 23072
rect 15381 23069 15393 23072
rect 15427 23069 15439 23103
rect 15381 23063 15439 23069
rect 17681 23103 17739 23109
rect 17681 23069 17693 23103
rect 17727 23100 17739 23103
rect 17862 23100 17868 23112
rect 17727 23072 17868 23100
rect 17727 23069 17739 23072
rect 17681 23063 17739 23069
rect 17862 23060 17868 23072
rect 17920 23060 17926 23112
rect 19334 23100 19340 23112
rect 19295 23072 19340 23100
rect 19334 23060 19340 23072
rect 19392 23060 19398 23112
rect 19978 23060 19984 23112
rect 20036 23100 20042 23112
rect 20901 23103 20959 23109
rect 20901 23100 20913 23103
rect 20036 23072 20913 23100
rect 20036 23060 20042 23072
rect 20901 23069 20913 23072
rect 20947 23069 20959 23103
rect 20901 23063 20959 23069
rect 15194 23032 15200 23044
rect 13780 23004 14136 23032
rect 14660 23004 15200 23032
rect 13780 22992 13786 23004
rect 14660 22976 14688 23004
rect 15194 22992 15200 23004
rect 15252 22992 15258 23044
rect 17034 23032 17040 23044
rect 16995 23004 17040 23032
rect 17034 22992 17040 23004
rect 17092 22992 17098 23044
rect 1394 22924 1400 22976
rect 1452 22964 1458 22976
rect 1581 22967 1639 22973
rect 1581 22964 1593 22967
rect 1452 22936 1593 22964
rect 1452 22924 1458 22936
rect 1581 22933 1593 22936
rect 1627 22933 1639 22967
rect 1581 22927 1639 22933
rect 12069 22967 12127 22973
rect 12069 22933 12081 22967
rect 12115 22964 12127 22967
rect 12526 22964 12532 22976
rect 12115 22936 12532 22964
rect 12115 22933 12127 22936
rect 12069 22927 12127 22933
rect 12526 22924 12532 22936
rect 12584 22924 12590 22976
rect 14642 22964 14648 22976
rect 14603 22936 14648 22964
rect 14642 22924 14648 22936
rect 14700 22924 14706 22976
rect 15470 22924 15476 22976
rect 15528 22964 15534 22976
rect 15657 22967 15715 22973
rect 15657 22964 15669 22967
rect 15528 22936 15669 22964
rect 15528 22924 15534 22936
rect 15657 22933 15669 22936
rect 15703 22933 15715 22967
rect 18598 22964 18604 22976
rect 18559 22936 18604 22964
rect 15657 22927 15715 22933
rect 18598 22924 18604 22936
rect 18656 22924 18662 22976
rect 20625 22967 20683 22973
rect 20625 22933 20637 22967
rect 20671 22964 20683 22967
rect 20898 22964 20904 22976
rect 20671 22936 20904 22964
rect 20671 22933 20683 22936
rect 20625 22927 20683 22933
rect 20898 22924 20904 22936
rect 20956 22924 20962 22976
rect 21100 22964 21128 23131
rect 21358 23128 21364 23140
rect 21416 23128 21422 23180
rect 21910 23128 21916 23180
rect 21968 23168 21974 23180
rect 22465 23171 22523 23177
rect 22465 23168 22477 23171
rect 21968 23140 22477 23168
rect 21968 23128 21974 23140
rect 22465 23137 22477 23140
rect 22511 23168 22523 23171
rect 22738 23168 22744 23180
rect 22511 23140 22744 23168
rect 22511 23137 22523 23140
rect 22465 23131 22523 23137
rect 22738 23128 22744 23140
rect 22796 23168 22802 23180
rect 23382 23168 23388 23180
rect 22796 23140 23388 23168
rect 22796 23128 22802 23140
rect 23382 23128 23388 23140
rect 23440 23128 23446 23180
rect 23477 23171 23535 23177
rect 23477 23137 23489 23171
rect 23523 23137 23535 23171
rect 23477 23131 23535 23137
rect 21376 23100 21404 23128
rect 21376 23072 22692 23100
rect 22664 23041 22692 23072
rect 22922 23060 22928 23112
rect 22980 23100 22986 23112
rect 23492 23100 23520 23131
rect 23566 23128 23572 23180
rect 23624 23168 23630 23180
rect 23937 23171 23995 23177
rect 23937 23168 23949 23171
rect 23624 23140 23949 23168
rect 23624 23128 23630 23140
rect 23937 23137 23949 23140
rect 23983 23137 23995 23171
rect 24670 23168 24676 23180
rect 24631 23140 24676 23168
rect 23937 23131 23995 23137
rect 24670 23128 24676 23140
rect 24728 23128 24734 23180
rect 23842 23100 23848 23112
rect 22980 23072 23848 23100
rect 22980 23060 22986 23072
rect 23842 23060 23848 23072
rect 23900 23060 23906 23112
rect 22649 23035 22707 23041
rect 22649 23001 22661 23035
rect 22695 23001 22707 23035
rect 22649 22995 22707 23001
rect 22830 22992 22836 23044
rect 22888 23032 22894 23044
rect 23017 23035 23075 23041
rect 23017 23032 23029 23035
rect 22888 23004 23029 23032
rect 22888 22992 22894 23004
rect 23017 23001 23029 23004
rect 23063 23001 23075 23035
rect 24486 23032 24492 23044
rect 24447 23004 24492 23032
rect 23017 22995 23075 23001
rect 24486 22992 24492 23004
rect 24544 22992 24550 23044
rect 21174 22964 21180 22976
rect 21087 22936 21180 22964
rect 21174 22924 21180 22936
rect 21232 22964 21238 22976
rect 21821 22967 21879 22973
rect 21821 22964 21833 22967
rect 21232 22936 21833 22964
rect 21232 22924 21238 22936
rect 21821 22933 21833 22936
rect 21867 22964 21879 22967
rect 21913 22967 21971 22973
rect 21913 22964 21925 22967
rect 21867 22936 21925 22964
rect 21867 22933 21879 22936
rect 21821 22927 21879 22933
rect 21913 22933 21925 22936
rect 21959 22933 21971 22967
rect 21913 22927 21971 22933
rect 22186 22924 22192 22976
rect 22244 22964 22250 22976
rect 23293 22967 23351 22973
rect 23293 22964 23305 22967
rect 22244 22936 23305 22964
rect 22244 22924 22250 22936
rect 23293 22933 23305 22936
rect 23339 22933 23351 22967
rect 25222 22964 25228 22976
rect 25183 22936 25228 22964
rect 23293 22927 23351 22933
rect 25222 22924 25228 22936
rect 25280 22924 25286 22976
rect 1104 22874 38824 22896
rect 1104 22822 4246 22874
rect 4298 22822 4310 22874
rect 4362 22822 4374 22874
rect 4426 22822 4438 22874
rect 4490 22822 34966 22874
rect 35018 22822 35030 22874
rect 35082 22822 35094 22874
rect 35146 22822 35158 22874
rect 35210 22822 38824 22874
rect 1104 22800 38824 22822
rect 3142 22760 3148 22772
rect 3103 22732 3148 22760
rect 3142 22720 3148 22732
rect 3200 22720 3206 22772
rect 10229 22763 10287 22769
rect 10229 22729 10241 22763
rect 10275 22760 10287 22763
rect 11146 22760 11152 22772
rect 10275 22732 11152 22760
rect 10275 22729 10287 22732
rect 10229 22723 10287 22729
rect 11146 22720 11152 22732
rect 11204 22720 11210 22772
rect 11790 22760 11796 22772
rect 11751 22732 11796 22760
rect 11790 22720 11796 22732
rect 11848 22720 11854 22772
rect 12618 22760 12624 22772
rect 12579 22732 12624 22760
rect 12618 22720 12624 22732
rect 12676 22720 12682 22772
rect 13265 22763 13323 22769
rect 13265 22729 13277 22763
rect 13311 22760 13323 22763
rect 13354 22760 13360 22772
rect 13311 22732 13360 22760
rect 13311 22729 13323 22732
rect 13265 22723 13323 22729
rect 13354 22720 13360 22732
rect 13412 22720 13418 22772
rect 15562 22760 15568 22772
rect 15523 22732 15568 22760
rect 15562 22720 15568 22732
rect 15620 22720 15626 22772
rect 15746 22720 15752 22772
rect 15804 22760 15810 22772
rect 16025 22763 16083 22769
rect 16025 22760 16037 22763
rect 15804 22732 16037 22760
rect 15804 22720 15810 22732
rect 16025 22729 16037 22732
rect 16071 22729 16083 22763
rect 16025 22723 16083 22729
rect 10597 22695 10655 22701
rect 10597 22661 10609 22695
rect 10643 22692 10655 22695
rect 10778 22692 10784 22704
rect 10643 22664 10784 22692
rect 10643 22661 10655 22664
rect 10597 22655 10655 22661
rect 10778 22652 10784 22664
rect 10836 22652 10842 22704
rect 10962 22692 10968 22704
rect 10923 22664 10968 22692
rect 10962 22652 10968 22664
rect 11020 22652 11026 22704
rect 11238 22652 11244 22704
rect 11296 22692 11302 22704
rect 11333 22695 11391 22701
rect 11333 22692 11345 22695
rect 11296 22664 11345 22692
rect 11296 22652 11302 22664
rect 11333 22661 11345 22664
rect 11379 22692 11391 22695
rect 11606 22692 11612 22704
rect 11379 22664 11612 22692
rect 11379 22661 11391 22664
rect 11333 22655 11391 22661
rect 11606 22652 11612 22664
rect 11664 22652 11670 22704
rect 15470 22652 15476 22704
rect 15528 22692 15534 22704
rect 15764 22692 15792 22720
rect 15528 22664 15792 22692
rect 15528 22652 15534 22664
rect 13998 22584 14004 22636
rect 14056 22624 14062 22636
rect 15013 22627 15071 22633
rect 15013 22624 15025 22627
rect 14056 22596 15025 22624
rect 14056 22584 14062 22596
rect 15013 22593 15025 22596
rect 15059 22593 15071 22627
rect 16040 22624 16068 22723
rect 17586 22720 17592 22772
rect 17644 22760 17650 22772
rect 19153 22763 19211 22769
rect 19153 22760 19165 22763
rect 17644 22732 19165 22760
rect 17644 22720 17650 22732
rect 19153 22729 19165 22732
rect 19199 22760 19211 22763
rect 19794 22760 19800 22772
rect 19199 22732 19800 22760
rect 19199 22729 19211 22732
rect 19153 22723 19211 22729
rect 19794 22720 19800 22732
rect 19852 22720 19858 22772
rect 20806 22720 20812 22772
rect 20864 22760 20870 22772
rect 21358 22760 21364 22772
rect 20864 22732 21364 22760
rect 20864 22720 20870 22732
rect 21358 22720 21364 22732
rect 21416 22760 21422 22772
rect 21453 22763 21511 22769
rect 21453 22760 21465 22763
rect 21416 22732 21465 22760
rect 21416 22720 21422 22732
rect 21453 22729 21465 22732
rect 21499 22729 21511 22763
rect 22738 22760 22744 22772
rect 22699 22732 22744 22760
rect 21453 22723 21511 22729
rect 22738 22720 22744 22732
rect 22796 22720 22802 22772
rect 23842 22760 23848 22772
rect 23803 22732 23848 22760
rect 23842 22720 23848 22732
rect 23900 22720 23906 22772
rect 24581 22763 24639 22769
rect 24581 22729 24593 22763
rect 24627 22760 24639 22763
rect 24670 22760 24676 22772
rect 24627 22732 24676 22760
rect 24627 22729 24639 22732
rect 24581 22723 24639 22729
rect 24670 22720 24676 22732
rect 24728 22720 24734 22772
rect 16114 22652 16120 22704
rect 16172 22692 16178 22704
rect 16390 22692 16396 22704
rect 16172 22664 16396 22692
rect 16172 22652 16178 22664
rect 16390 22652 16396 22664
rect 16448 22692 16454 22704
rect 16485 22695 16543 22701
rect 16485 22692 16497 22695
rect 16448 22664 16497 22692
rect 16448 22652 16454 22664
rect 16485 22661 16497 22664
rect 16531 22692 16543 22695
rect 18414 22692 18420 22704
rect 16531 22664 18420 22692
rect 16531 22661 16543 22664
rect 16485 22655 16543 22661
rect 18414 22652 18420 22664
rect 18472 22652 18478 22704
rect 19613 22695 19671 22701
rect 19613 22661 19625 22695
rect 19659 22692 19671 22695
rect 19978 22692 19984 22704
rect 19659 22664 19984 22692
rect 19659 22661 19671 22664
rect 19613 22655 19671 22661
rect 19978 22652 19984 22664
rect 20036 22652 20042 22704
rect 22002 22652 22008 22704
rect 22060 22692 22066 22704
rect 23106 22692 23112 22704
rect 22060 22664 23112 22692
rect 22060 22652 22066 22664
rect 23106 22652 23112 22664
rect 23164 22652 23170 22704
rect 16577 22627 16635 22633
rect 16577 22624 16589 22627
rect 16040 22596 16589 22624
rect 15013 22587 15071 22593
rect 16577 22593 16589 22596
rect 16623 22593 16635 22627
rect 17497 22627 17555 22633
rect 17497 22624 17509 22627
rect 16577 22587 16635 22593
rect 16684 22596 17509 22624
rect 1394 22516 1400 22568
rect 1452 22556 1458 22568
rect 1581 22559 1639 22565
rect 1581 22556 1593 22559
rect 1452 22528 1593 22556
rect 1452 22516 1458 22528
rect 1581 22525 1593 22528
rect 1627 22525 1639 22559
rect 1854 22556 1860 22568
rect 1815 22528 1860 22556
rect 1581 22519 1639 22525
rect 1854 22516 1860 22528
rect 1912 22516 1918 22568
rect 11790 22516 11796 22568
rect 11848 22556 11854 22568
rect 12434 22556 12440 22568
rect 11848 22528 12440 22556
rect 11848 22516 11854 22528
rect 12434 22516 12440 22528
rect 12492 22556 12498 22568
rect 13630 22556 13636 22568
rect 12492 22528 12537 22556
rect 13591 22528 13636 22556
rect 12492 22516 12498 22528
rect 13630 22516 13636 22528
rect 13688 22516 13694 22568
rect 13906 22556 13912 22568
rect 13740 22528 13912 22556
rect 12253 22491 12311 22497
rect 12253 22457 12265 22491
rect 12299 22488 12311 22491
rect 13740 22488 13768 22528
rect 13906 22516 13912 22528
rect 13964 22516 13970 22568
rect 16298 22516 16304 22568
rect 16356 22556 16362 22568
rect 16684 22565 16712 22596
rect 17497 22593 17509 22596
rect 17543 22624 17555 22627
rect 18874 22624 18880 22636
rect 17543 22596 18736 22624
rect 18835 22596 18880 22624
rect 17543 22593 17555 22596
rect 17497 22587 17555 22593
rect 16669 22559 16727 22565
rect 16669 22556 16681 22559
rect 16356 22528 16681 22556
rect 16356 22516 16362 22528
rect 16669 22525 16681 22528
rect 16715 22525 16727 22559
rect 16669 22519 16727 22525
rect 17862 22516 17868 22568
rect 17920 22556 17926 22568
rect 18417 22559 18475 22565
rect 18417 22556 18429 22559
rect 17920 22528 18429 22556
rect 17920 22516 17926 22528
rect 18417 22525 18429 22528
rect 18463 22556 18475 22559
rect 18598 22556 18604 22568
rect 18463 22528 18604 22556
rect 18463 22525 18475 22528
rect 18417 22519 18475 22525
rect 18598 22516 18604 22528
rect 18656 22516 18662 22568
rect 12299 22460 13768 22488
rect 17129 22491 17187 22497
rect 12299 22457 12311 22460
rect 12253 22451 12311 22457
rect 17129 22457 17141 22491
rect 17175 22488 17187 22491
rect 17678 22488 17684 22500
rect 17175 22460 17684 22488
rect 17175 22457 17187 22460
rect 17129 22451 17187 22457
rect 17678 22448 17684 22460
rect 17736 22448 17742 22500
rect 18046 22448 18052 22500
rect 18104 22488 18110 22500
rect 18141 22491 18199 22497
rect 18141 22488 18153 22491
rect 18104 22460 18153 22488
rect 18104 22448 18110 22460
rect 18141 22457 18153 22460
rect 18187 22457 18199 22491
rect 18322 22488 18328 22500
rect 18283 22460 18328 22488
rect 18141 22451 18199 22457
rect 18322 22448 18328 22460
rect 18380 22448 18386 22500
rect 18506 22488 18512 22500
rect 18467 22460 18512 22488
rect 18506 22448 18512 22460
rect 18564 22448 18570 22500
rect 18708 22488 18736 22596
rect 18874 22584 18880 22596
rect 18932 22584 18938 22636
rect 19058 22516 19064 22568
rect 19116 22556 19122 22568
rect 19996 22565 20024 22652
rect 20438 22624 20444 22636
rect 20399 22596 20444 22624
rect 20438 22584 20444 22596
rect 20496 22584 20502 22636
rect 20898 22584 20904 22636
rect 20956 22624 20962 22636
rect 22373 22627 22431 22633
rect 22373 22624 22385 22627
rect 20956 22596 22385 22624
rect 20956 22584 20962 22596
rect 22373 22593 22385 22596
rect 22419 22624 22431 22627
rect 25222 22624 25228 22636
rect 22419 22596 25228 22624
rect 22419 22593 22431 22596
rect 22373 22587 22431 22593
rect 25222 22584 25228 22596
rect 25280 22584 25286 22636
rect 19981 22559 20039 22565
rect 19981 22556 19993 22559
rect 19116 22528 19993 22556
rect 19116 22516 19122 22528
rect 19981 22525 19993 22528
rect 20027 22525 20039 22559
rect 19981 22519 20039 22525
rect 20533 22559 20591 22565
rect 20533 22525 20545 22559
rect 20579 22556 20591 22559
rect 20622 22556 20628 22568
rect 20579 22528 20628 22556
rect 20579 22525 20591 22528
rect 20533 22519 20591 22525
rect 19150 22488 19156 22500
rect 18708 22460 19156 22488
rect 19150 22448 19156 22460
rect 19208 22448 19214 22500
rect 19996 22488 20024 22519
rect 20622 22516 20628 22528
rect 20680 22516 20686 22568
rect 21726 22556 21732 22568
rect 21687 22528 21732 22556
rect 21726 22516 21732 22528
rect 21784 22516 21790 22568
rect 23106 22556 23112 22568
rect 23067 22528 23112 22556
rect 23106 22516 23112 22528
rect 23164 22516 23170 22568
rect 21085 22491 21143 22497
rect 21085 22488 21097 22491
rect 19996 22460 21097 22488
rect 21085 22457 21097 22460
rect 21131 22457 21143 22491
rect 21085 22451 21143 22457
rect 14366 22380 14372 22432
rect 14424 22420 14430 22432
rect 16666 22420 16672 22432
rect 14424 22392 16672 22420
rect 14424 22380 14430 22392
rect 16666 22380 16672 22392
rect 16724 22380 16730 22432
rect 17865 22423 17923 22429
rect 17865 22389 17877 22423
rect 17911 22420 17923 22423
rect 18340 22420 18368 22448
rect 19978 22420 19984 22432
rect 17911 22392 18368 22420
rect 19939 22392 19984 22420
rect 17911 22389 17923 22392
rect 17865 22383 17923 22389
rect 19978 22380 19984 22392
rect 20036 22380 20042 22432
rect 1104 22330 38824 22352
rect 1104 22278 19606 22330
rect 19658 22278 19670 22330
rect 19722 22278 19734 22330
rect 19786 22278 19798 22330
rect 19850 22278 38824 22330
rect 1104 22256 38824 22278
rect 11330 22176 11336 22228
rect 11388 22216 11394 22228
rect 11882 22216 11888 22228
rect 11388 22188 11888 22216
rect 11388 22176 11394 22188
rect 11882 22176 11888 22188
rect 11940 22176 11946 22228
rect 13265 22219 13323 22225
rect 13265 22185 13277 22219
rect 13311 22216 13323 22219
rect 13722 22216 13728 22228
rect 13311 22188 13728 22216
rect 13311 22185 13323 22188
rect 13265 22179 13323 22185
rect 13722 22176 13728 22188
rect 13780 22176 13786 22228
rect 14369 22219 14427 22225
rect 14369 22185 14381 22219
rect 14415 22216 14427 22219
rect 14826 22216 14832 22228
rect 14415 22188 14832 22216
rect 14415 22185 14427 22188
rect 14369 22179 14427 22185
rect 14826 22176 14832 22188
rect 14884 22176 14890 22228
rect 17034 22176 17040 22228
rect 17092 22216 17098 22228
rect 17678 22216 17684 22228
rect 17092 22188 17684 22216
rect 17092 22176 17098 22188
rect 17678 22176 17684 22188
rect 17736 22176 17742 22228
rect 18046 22176 18052 22228
rect 18104 22216 18110 22228
rect 18233 22219 18291 22225
rect 18233 22216 18245 22219
rect 18104 22188 18245 22216
rect 18104 22176 18110 22188
rect 18233 22185 18245 22188
rect 18279 22216 18291 22219
rect 19242 22216 19248 22228
rect 18279 22188 19248 22216
rect 18279 22185 18291 22188
rect 18233 22179 18291 22185
rect 19242 22176 19248 22188
rect 19300 22176 19306 22228
rect 20165 22219 20223 22225
rect 20165 22185 20177 22219
rect 20211 22216 20223 22219
rect 20622 22216 20628 22228
rect 20211 22188 20628 22216
rect 20211 22185 20223 22188
rect 20165 22179 20223 22185
rect 20622 22176 20628 22188
rect 20680 22176 20686 22228
rect 21726 22216 21732 22228
rect 21687 22188 21732 22216
rect 21726 22176 21732 22188
rect 21784 22176 21790 22228
rect 5442 22108 5448 22160
rect 5500 22148 5506 22160
rect 9858 22148 9864 22160
rect 5500 22120 9864 22148
rect 5500 22108 5506 22120
rect 9858 22108 9864 22120
rect 9916 22108 9922 22160
rect 13998 22148 14004 22160
rect 13832 22120 14004 22148
rect 10134 22040 10140 22092
rect 10192 22080 10198 22092
rect 11330 22080 11336 22092
rect 10192 22052 11336 22080
rect 10192 22040 10198 22052
rect 11330 22040 11336 22052
rect 11388 22080 11394 22092
rect 12253 22083 12311 22089
rect 12253 22080 12265 22083
rect 11388 22052 12265 22080
rect 11388 22040 11394 22052
rect 12253 22049 12265 22052
rect 12299 22049 12311 22083
rect 12253 22043 12311 22049
rect 12621 22083 12679 22089
rect 12621 22049 12633 22083
rect 12667 22080 12679 22083
rect 13078 22080 13084 22092
rect 12667 22052 13084 22080
rect 12667 22049 12679 22052
rect 12621 22043 12679 22049
rect 13078 22040 13084 22052
rect 13136 22040 13142 22092
rect 13633 22083 13691 22089
rect 13633 22049 13645 22083
rect 13679 22080 13691 22083
rect 13832 22080 13860 22120
rect 13998 22108 14004 22120
rect 14056 22108 14062 22160
rect 15105 22151 15163 22157
rect 15105 22117 15117 22151
rect 15151 22148 15163 22151
rect 15194 22148 15200 22160
rect 15151 22120 15200 22148
rect 15151 22117 15163 22120
rect 15105 22111 15163 22117
rect 15194 22108 15200 22120
rect 15252 22108 15258 22160
rect 16577 22151 16635 22157
rect 16577 22117 16589 22151
rect 16623 22148 16635 22151
rect 16850 22148 16856 22160
rect 16623 22120 16856 22148
rect 16623 22117 16635 22120
rect 16577 22111 16635 22117
rect 16850 22108 16856 22120
rect 16908 22148 16914 22160
rect 17218 22148 17224 22160
rect 16908 22120 17224 22148
rect 16908 22108 16914 22120
rect 17218 22108 17224 22120
rect 17276 22108 17282 22160
rect 17310 22108 17316 22160
rect 17368 22148 17374 22160
rect 17957 22151 18015 22157
rect 17957 22148 17969 22151
rect 17368 22120 17969 22148
rect 17368 22108 17374 22120
rect 17957 22117 17969 22120
rect 18003 22117 18015 22151
rect 19426 22148 19432 22160
rect 17957 22111 18015 22117
rect 18800 22120 19432 22148
rect 14182 22080 14188 22092
rect 13679 22052 13860 22080
rect 14143 22052 14188 22080
rect 13679 22049 13691 22052
rect 13633 22043 13691 22049
rect 14182 22040 14188 22052
rect 14240 22040 14246 22092
rect 14734 22080 14740 22092
rect 14695 22052 14740 22080
rect 14734 22040 14740 22052
rect 14792 22040 14798 22092
rect 16022 22080 16028 22092
rect 15983 22052 16028 22080
rect 16022 22040 16028 22052
rect 16080 22040 16086 22092
rect 16117 22083 16175 22089
rect 16117 22049 16129 22083
rect 16163 22080 16175 22083
rect 16298 22080 16304 22092
rect 16163 22052 16304 22080
rect 16163 22049 16175 22052
rect 16117 22043 16175 22049
rect 16298 22040 16304 22052
rect 16356 22040 16362 22092
rect 17494 22080 17500 22092
rect 17407 22052 17500 22080
rect 17494 22040 17500 22052
rect 17552 22080 17558 22092
rect 17862 22080 17868 22092
rect 17552 22052 17868 22080
rect 17552 22040 17558 22052
rect 17862 22040 17868 22052
rect 17920 22040 17926 22092
rect 18693 22083 18751 22089
rect 18693 22049 18705 22083
rect 18739 22080 18751 22083
rect 18800 22080 18828 22120
rect 19426 22108 19432 22120
rect 19484 22108 19490 22160
rect 19797 22151 19855 22157
rect 19797 22117 19809 22151
rect 19843 22148 19855 22151
rect 20438 22148 20444 22160
rect 19843 22120 20444 22148
rect 19843 22117 19855 22120
rect 19797 22111 19855 22117
rect 20438 22108 20444 22120
rect 20496 22108 20502 22160
rect 21542 22108 21548 22160
rect 21600 22148 21606 22160
rect 21600 22120 22048 22148
rect 21600 22108 21606 22120
rect 18739 22052 18828 22080
rect 18739 22049 18751 22052
rect 18693 22043 18751 22049
rect 18874 22040 18880 22092
rect 18932 22080 18938 22092
rect 20990 22080 20996 22092
rect 18932 22052 18977 22080
rect 20951 22052 20996 22080
rect 18932 22040 18938 22052
rect 20990 22040 20996 22052
rect 21048 22040 21054 22092
rect 22020 22080 22048 22120
rect 22097 22083 22155 22089
rect 22097 22080 22109 22083
rect 22020 22052 22109 22080
rect 22097 22049 22109 22052
rect 22143 22049 22155 22083
rect 22097 22043 22155 22049
rect 11606 22012 11612 22024
rect 11567 21984 11612 22012
rect 11606 21972 11612 21984
rect 11664 21972 11670 22024
rect 12342 22012 12348 22024
rect 12303 21984 12348 22012
rect 12342 21972 12348 21984
rect 12400 21972 12406 22024
rect 12526 22012 12532 22024
rect 12487 21984 12532 22012
rect 12526 21972 12532 21984
rect 12584 21972 12590 22024
rect 15930 22012 15936 22024
rect 15891 21984 15936 22012
rect 15930 21972 15936 21984
rect 15988 21972 15994 22024
rect 17405 22015 17463 22021
rect 17405 21981 17417 22015
rect 17451 22012 17463 22015
rect 18046 22012 18052 22024
rect 17451 21984 18052 22012
rect 17451 21981 17463 21984
rect 17405 21975 17463 21981
rect 18046 21972 18052 21984
rect 18104 22012 18110 22024
rect 18230 22012 18236 22024
rect 18104 21984 18236 22012
rect 18104 21972 18110 21984
rect 18230 21972 18236 21984
rect 18288 21972 18294 22024
rect 18782 22012 18788 22024
rect 18743 21984 18788 22012
rect 18782 21972 18788 21984
rect 18840 21972 18846 22024
rect 20901 22015 20959 22021
rect 20901 21981 20913 22015
rect 20947 22012 20959 22015
rect 21910 22012 21916 22024
rect 20947 21984 21916 22012
rect 20947 21981 20959 21984
rect 20901 21975 20959 21981
rect 21910 21972 21916 21984
rect 21968 21972 21974 22024
rect 23106 22012 23112 22024
rect 23067 21984 23112 22012
rect 23106 21972 23112 21984
rect 23164 21972 23170 22024
rect 23382 22012 23388 22024
rect 23343 21984 23388 22012
rect 23382 21972 23388 21984
rect 23440 21972 23446 22024
rect 16945 21947 17003 21953
rect 16945 21913 16957 21947
rect 16991 21944 17003 21947
rect 17954 21944 17960 21956
rect 16991 21916 17960 21944
rect 16991 21913 17003 21916
rect 16945 21907 17003 21913
rect 17954 21904 17960 21916
rect 18012 21904 18018 21956
rect 1673 21879 1731 21885
rect 1673 21845 1685 21879
rect 1719 21876 1731 21879
rect 1854 21876 1860 21888
rect 1719 21848 1860 21876
rect 1719 21845 1731 21848
rect 1673 21839 1731 21845
rect 1854 21836 1860 21848
rect 1912 21836 1918 21888
rect 13906 21836 13912 21888
rect 13964 21876 13970 21888
rect 14001 21879 14059 21885
rect 14001 21876 14013 21879
rect 13964 21848 14013 21876
rect 13964 21836 13970 21848
rect 14001 21845 14013 21848
rect 14047 21876 14059 21879
rect 15102 21876 15108 21888
rect 14047 21848 15108 21876
rect 14047 21845 14059 21848
rect 14001 21839 14059 21845
rect 15102 21836 15108 21848
rect 15160 21876 15166 21888
rect 15562 21876 15568 21888
rect 15160 21848 15568 21876
rect 15160 21836 15166 21848
rect 15562 21836 15568 21848
rect 15620 21836 15626 21888
rect 17313 21879 17371 21885
rect 17313 21845 17325 21879
rect 17359 21876 17371 21879
rect 17586 21876 17592 21888
rect 17359 21848 17592 21876
rect 17359 21845 17371 21848
rect 17313 21839 17371 21845
rect 17586 21836 17592 21848
rect 17644 21836 17650 21888
rect 18690 21836 18696 21888
rect 18748 21876 18754 21888
rect 19061 21879 19119 21885
rect 19061 21876 19073 21879
rect 18748 21848 19073 21876
rect 18748 21836 18754 21848
rect 19061 21845 19073 21848
rect 19107 21845 19119 21879
rect 20438 21876 20444 21888
rect 20399 21848 20444 21876
rect 19061 21839 19119 21845
rect 20438 21836 20444 21848
rect 20496 21836 20502 21888
rect 21082 21836 21088 21888
rect 21140 21876 21146 21888
rect 21177 21879 21235 21885
rect 21177 21876 21189 21879
rect 21140 21848 21189 21876
rect 21140 21836 21146 21848
rect 21177 21845 21189 21848
rect 21223 21845 21235 21879
rect 22462 21876 22468 21888
rect 22423 21848 22468 21876
rect 21177 21839 21235 21845
rect 22462 21836 22468 21848
rect 22520 21836 22526 21888
rect 24486 21876 24492 21888
rect 24447 21848 24492 21876
rect 24486 21836 24492 21848
rect 24544 21836 24550 21888
rect 1104 21786 38824 21808
rect 1104 21734 4246 21786
rect 4298 21734 4310 21786
rect 4362 21734 4374 21786
rect 4426 21734 4438 21786
rect 4490 21734 34966 21786
rect 35018 21734 35030 21786
rect 35082 21734 35094 21786
rect 35146 21734 35158 21786
rect 35210 21734 38824 21786
rect 1104 21712 38824 21734
rect 11330 21672 11336 21684
rect 11291 21644 11336 21672
rect 11330 21632 11336 21644
rect 11388 21632 11394 21684
rect 11701 21675 11759 21681
rect 11701 21641 11713 21675
rect 11747 21672 11759 21675
rect 12250 21672 12256 21684
rect 11747 21644 12256 21672
rect 11747 21641 11759 21644
rect 11701 21635 11759 21641
rect 12250 21632 12256 21644
rect 12308 21632 12314 21684
rect 13630 21672 13636 21684
rect 13591 21644 13636 21672
rect 13630 21632 13636 21644
rect 13688 21632 13694 21684
rect 14182 21672 14188 21684
rect 14143 21644 14188 21672
rect 14182 21632 14188 21644
rect 14240 21672 14246 21684
rect 15378 21672 15384 21684
rect 14240 21644 15384 21672
rect 14240 21632 14246 21644
rect 15378 21632 15384 21644
rect 15436 21632 15442 21684
rect 15746 21672 15752 21684
rect 15659 21644 15752 21672
rect 15746 21632 15752 21644
rect 15804 21672 15810 21684
rect 16022 21672 16028 21684
rect 15804 21644 16028 21672
rect 15804 21632 15810 21644
rect 16022 21632 16028 21644
rect 16080 21632 16086 21684
rect 16117 21675 16175 21681
rect 16117 21641 16129 21675
rect 16163 21672 16175 21675
rect 16298 21672 16304 21684
rect 16163 21644 16304 21672
rect 16163 21641 16175 21644
rect 16117 21635 16175 21641
rect 16298 21632 16304 21644
rect 16356 21632 16362 21684
rect 17494 21672 17500 21684
rect 17455 21644 17500 21672
rect 17494 21632 17500 21644
rect 17552 21632 17558 21684
rect 18874 21632 18880 21684
rect 18932 21672 18938 21684
rect 19153 21675 19211 21681
rect 19153 21672 19165 21675
rect 18932 21644 19165 21672
rect 18932 21632 18938 21644
rect 19153 21641 19165 21644
rect 19199 21641 19211 21675
rect 19153 21635 19211 21641
rect 20990 21632 20996 21684
rect 21048 21672 21054 21684
rect 21361 21675 21419 21681
rect 21361 21672 21373 21675
rect 21048 21644 21373 21672
rect 21048 21632 21054 21644
rect 21361 21641 21373 21644
rect 21407 21641 21419 21675
rect 21361 21635 21419 21641
rect 21821 21675 21879 21681
rect 21821 21641 21833 21675
rect 21867 21672 21879 21675
rect 21910 21672 21916 21684
rect 21867 21644 21916 21672
rect 21867 21641 21879 21644
rect 21821 21635 21879 21641
rect 21910 21632 21916 21644
rect 21968 21632 21974 21684
rect 23201 21675 23259 21681
rect 23201 21641 23213 21675
rect 23247 21672 23259 21675
rect 23382 21672 23388 21684
rect 23247 21644 23388 21672
rect 23247 21641 23259 21644
rect 23201 21635 23259 21641
rect 23382 21632 23388 21644
rect 23440 21632 23446 21684
rect 26418 21672 26424 21684
rect 26379 21644 26424 21672
rect 26418 21632 26424 21644
rect 26476 21632 26482 21684
rect 11238 21564 11244 21616
rect 11296 21604 11302 21616
rect 11977 21607 12035 21613
rect 11977 21604 11989 21607
rect 11296 21576 11989 21604
rect 11296 21564 11302 21576
rect 11977 21573 11989 21576
rect 12023 21604 12035 21607
rect 12526 21604 12532 21616
rect 12023 21576 12532 21604
rect 12023 21573 12035 21576
rect 11977 21567 12035 21573
rect 12526 21564 12532 21576
rect 12584 21604 12590 21616
rect 12802 21604 12808 21616
rect 12584 21576 12808 21604
rect 12584 21564 12590 21576
rect 12802 21564 12808 21576
rect 12860 21564 12866 21616
rect 19886 21564 19892 21616
rect 19944 21604 19950 21616
rect 19944 21576 20116 21604
rect 19944 21564 19950 21576
rect 14550 21496 14556 21548
rect 14608 21536 14614 21548
rect 16390 21536 16396 21548
rect 14608 21508 16396 21536
rect 14608 21496 14614 21508
rect 16390 21496 16396 21508
rect 16448 21536 16454 21548
rect 16577 21539 16635 21545
rect 16577 21536 16589 21539
rect 16448 21508 16589 21536
rect 16448 21496 16454 21508
rect 16577 21505 16589 21508
rect 16623 21505 16635 21539
rect 16577 21499 16635 21505
rect 17129 21539 17187 21545
rect 17129 21505 17141 21539
rect 17175 21536 17187 21539
rect 17770 21536 17776 21548
rect 17175 21508 17776 21536
rect 17175 21505 17187 21508
rect 17129 21499 17187 21505
rect 17770 21496 17776 21508
rect 17828 21496 17834 21548
rect 17954 21496 17960 21548
rect 18012 21536 18018 21548
rect 18141 21539 18199 21545
rect 18141 21536 18153 21539
rect 18012 21508 18153 21536
rect 18012 21496 18018 21508
rect 18141 21505 18153 21508
rect 18187 21505 18199 21539
rect 19610 21536 19616 21548
rect 19523 21508 19616 21536
rect 18141 21499 18199 21505
rect 19610 21496 19616 21508
rect 19668 21536 19674 21548
rect 19668 21508 19932 21536
rect 19668 21496 19674 21508
rect 16485 21471 16543 21477
rect 16485 21437 16497 21471
rect 16531 21468 16543 21471
rect 16666 21468 16672 21480
rect 16531 21440 16672 21468
rect 16531 21437 16543 21440
rect 16485 21431 16543 21437
rect 16666 21428 16672 21440
rect 16724 21428 16730 21480
rect 17865 21471 17923 21477
rect 17865 21437 17877 21471
rect 17911 21468 17923 21471
rect 18782 21468 18788 21480
rect 17911 21440 18788 21468
rect 17911 21437 17923 21440
rect 17865 21431 17923 21437
rect 18782 21428 18788 21440
rect 18840 21428 18846 21480
rect 19904 21477 19932 21508
rect 19705 21471 19763 21477
rect 19705 21437 19717 21471
rect 19751 21437 19763 21471
rect 19705 21431 19763 21437
rect 19889 21471 19947 21477
rect 19889 21437 19901 21471
rect 19935 21437 19947 21471
rect 20088 21468 20116 21576
rect 20993 21539 21051 21545
rect 20993 21505 21005 21539
rect 21039 21536 21051 21539
rect 21266 21536 21272 21548
rect 21039 21508 21272 21536
rect 21039 21505 21051 21508
rect 20993 21499 21051 21505
rect 21266 21496 21272 21508
rect 21324 21496 21330 21548
rect 20346 21468 20352 21480
rect 20088 21440 20352 21468
rect 19889 21431 19947 21437
rect 10962 21400 10968 21412
rect 10923 21372 10968 21400
rect 10962 21360 10968 21372
rect 11020 21360 11026 21412
rect 19426 21292 19432 21344
rect 19484 21332 19490 21344
rect 19720 21332 19748 21431
rect 19904 21400 19932 21431
rect 20346 21428 20352 21440
rect 20404 21428 20410 21480
rect 20438 21428 20444 21480
rect 20496 21468 20502 21480
rect 24857 21471 24915 21477
rect 20496 21440 20541 21468
rect 20496 21428 20502 21440
rect 24857 21437 24869 21471
rect 24903 21437 24915 21471
rect 24857 21431 24915 21437
rect 25133 21471 25191 21477
rect 25133 21437 25145 21471
rect 25179 21468 25191 21471
rect 25222 21468 25228 21480
rect 25179 21440 25228 21468
rect 25179 21437 25191 21440
rect 25133 21431 25191 21437
rect 22646 21400 22652 21412
rect 19904 21372 22652 21400
rect 22646 21360 22652 21372
rect 22704 21360 22710 21412
rect 23106 21360 23112 21412
rect 23164 21400 23170 21412
rect 23937 21403 23995 21409
rect 23937 21400 23949 21403
rect 23164 21372 23949 21400
rect 23164 21360 23170 21372
rect 23937 21369 23949 21372
rect 23983 21400 23995 21403
rect 24872 21400 24900 21431
rect 25222 21428 25228 21440
rect 25280 21428 25286 21480
rect 24946 21400 24952 21412
rect 23983 21372 24952 21400
rect 23983 21369 23995 21372
rect 23937 21363 23995 21369
rect 24946 21360 24952 21372
rect 25004 21360 25010 21412
rect 22186 21332 22192 21344
rect 19484 21304 22192 21332
rect 19484 21292 19490 21304
rect 22186 21292 22192 21304
rect 22244 21292 22250 21344
rect 24670 21332 24676 21344
rect 24631 21304 24676 21332
rect 24670 21292 24676 21304
rect 24728 21332 24734 21344
rect 25222 21332 25228 21344
rect 24728 21304 25228 21332
rect 24728 21292 24734 21304
rect 25222 21292 25228 21304
rect 25280 21292 25286 21344
rect 1104 21242 38824 21264
rect 1104 21190 19606 21242
rect 19658 21190 19670 21242
rect 19722 21190 19734 21242
rect 19786 21190 19798 21242
rect 19850 21190 38824 21242
rect 1104 21168 38824 21190
rect 13078 21128 13084 21140
rect 13039 21100 13084 21128
rect 13078 21088 13084 21100
rect 13136 21088 13142 21140
rect 16390 21128 16396 21140
rect 16351 21100 16396 21128
rect 16390 21088 16396 21100
rect 16448 21088 16454 21140
rect 16850 21128 16856 21140
rect 16811 21100 16856 21128
rect 16850 21088 16856 21100
rect 16908 21088 16914 21140
rect 18046 21128 18052 21140
rect 18007 21100 18052 21128
rect 18046 21088 18052 21100
rect 18104 21088 18110 21140
rect 18509 21131 18567 21137
rect 18509 21097 18521 21131
rect 18555 21128 18567 21131
rect 18598 21128 18604 21140
rect 18555 21100 18604 21128
rect 18555 21097 18567 21100
rect 18509 21091 18567 21097
rect 18598 21088 18604 21100
rect 18656 21088 18662 21140
rect 19978 21088 19984 21140
rect 20036 21128 20042 21140
rect 20257 21131 20315 21137
rect 20257 21128 20269 21131
rect 20036 21100 20269 21128
rect 20036 21088 20042 21100
rect 20257 21097 20269 21100
rect 20303 21128 20315 21131
rect 20622 21128 20628 21140
rect 20303 21100 20628 21128
rect 20303 21097 20315 21100
rect 20257 21091 20315 21097
rect 20622 21088 20628 21100
rect 20680 21088 20686 21140
rect 21082 21128 21088 21140
rect 21043 21100 21088 21128
rect 21082 21088 21088 21100
rect 21140 21088 21146 21140
rect 21358 21128 21364 21140
rect 21319 21100 21364 21128
rect 21358 21088 21364 21100
rect 21416 21088 21422 21140
rect 19058 21060 19064 21072
rect 18892 21032 19064 21060
rect 11701 20995 11759 21001
rect 11701 20961 11713 20995
rect 11747 20992 11759 20995
rect 12066 20992 12072 21004
rect 11747 20964 12072 20992
rect 11747 20961 11759 20964
rect 11701 20955 11759 20961
rect 12066 20952 12072 20964
rect 12124 20992 12130 21004
rect 13630 20992 13636 21004
rect 12124 20964 13636 20992
rect 12124 20952 12130 20964
rect 13630 20952 13636 20964
rect 13688 20952 13694 21004
rect 17678 20992 17684 21004
rect 17639 20964 17684 20992
rect 17678 20952 17684 20964
rect 17736 20952 17742 21004
rect 18892 21001 18920 21032
rect 19058 21020 19064 21032
rect 19116 21020 19122 21072
rect 19150 21020 19156 21072
rect 19208 21060 19214 21072
rect 20438 21060 20444 21072
rect 19208 21032 20444 21060
rect 19208 21020 19214 21032
rect 19352 21001 19380 21032
rect 20438 21020 20444 21032
rect 20496 21020 20502 21072
rect 18785 20995 18843 21001
rect 18785 20961 18797 20995
rect 18831 20961 18843 20995
rect 18785 20955 18843 20961
rect 18877 20995 18935 21001
rect 18877 20961 18889 20995
rect 18923 20961 18935 20995
rect 18877 20955 18935 20961
rect 19337 20995 19395 21001
rect 19337 20961 19349 20995
rect 19383 20961 19395 20995
rect 19337 20955 19395 20961
rect 19521 20995 19579 21001
rect 19521 20961 19533 20995
rect 19567 20992 19579 20995
rect 19702 20992 19708 21004
rect 19567 20964 19708 20992
rect 19567 20961 19579 20964
rect 19521 20955 19579 20961
rect 11974 20924 11980 20936
rect 11935 20896 11980 20924
rect 11974 20884 11980 20896
rect 12032 20884 12038 20936
rect 17773 20927 17831 20933
rect 17773 20893 17785 20927
rect 17819 20924 17831 20927
rect 18322 20924 18328 20936
rect 17819 20896 18328 20924
rect 17819 20893 17831 20896
rect 17773 20887 17831 20893
rect 18322 20884 18328 20896
rect 18380 20884 18386 20936
rect 18800 20856 18828 20955
rect 19702 20952 19708 20964
rect 19760 20952 19766 21004
rect 20346 20952 20352 21004
rect 20404 20992 20410 21004
rect 20625 20995 20683 21001
rect 20625 20992 20637 20995
rect 20404 20964 20637 20992
rect 20404 20952 20410 20964
rect 20625 20961 20637 20964
rect 20671 20961 20683 20995
rect 20625 20955 20683 20961
rect 20901 20995 20959 21001
rect 20901 20961 20913 20995
rect 20947 20992 20959 20995
rect 21174 20992 21180 21004
rect 20947 20964 21180 20992
rect 20947 20961 20959 20964
rect 20901 20955 20959 20961
rect 21174 20952 21180 20964
rect 21232 20992 21238 21004
rect 21358 20992 21364 21004
rect 21232 20964 21364 20992
rect 21232 20952 21238 20964
rect 21358 20952 21364 20964
rect 21416 20952 21422 21004
rect 19889 20927 19947 20933
rect 19889 20893 19901 20927
rect 19935 20924 19947 20927
rect 20530 20924 20536 20936
rect 19935 20896 20536 20924
rect 19935 20893 19947 20896
rect 19889 20887 19947 20893
rect 20530 20884 20536 20896
rect 20588 20884 20594 20936
rect 19334 20856 19340 20868
rect 18800 20828 19340 20856
rect 19334 20816 19340 20828
rect 19392 20856 19398 20868
rect 20806 20856 20812 20868
rect 19392 20828 20812 20856
rect 19392 20816 19398 20828
rect 20806 20816 20812 20828
rect 20864 20816 20870 20868
rect 1854 20748 1860 20800
rect 1912 20788 1918 20800
rect 2682 20788 2688 20800
rect 1912 20760 2688 20788
rect 1912 20748 1918 20760
rect 2682 20748 2688 20760
rect 2740 20748 2746 20800
rect 17954 20748 17960 20800
rect 18012 20788 18018 20800
rect 19702 20788 19708 20800
rect 18012 20760 19708 20788
rect 18012 20748 18018 20760
rect 19702 20748 19708 20760
rect 19760 20748 19766 20800
rect 24946 20788 24952 20800
rect 24907 20760 24952 20788
rect 24946 20748 24952 20760
rect 25004 20748 25010 20800
rect 1104 20698 38824 20720
rect 1104 20646 4246 20698
rect 4298 20646 4310 20698
rect 4362 20646 4374 20698
rect 4426 20646 4438 20698
rect 4490 20646 34966 20698
rect 35018 20646 35030 20698
rect 35082 20646 35094 20698
rect 35146 20646 35158 20698
rect 35210 20646 38824 20698
rect 1104 20624 38824 20646
rect 12066 20584 12072 20596
rect 12027 20556 12072 20584
rect 12066 20544 12072 20556
rect 12124 20544 12130 20596
rect 12250 20544 12256 20596
rect 12308 20584 12314 20596
rect 13541 20587 13599 20593
rect 13541 20584 13553 20587
rect 12308 20556 13553 20584
rect 12308 20544 12314 20556
rect 13541 20553 13553 20556
rect 13587 20584 13599 20587
rect 13722 20584 13728 20596
rect 13587 20556 13728 20584
rect 13587 20553 13599 20556
rect 13541 20547 13599 20553
rect 13722 20544 13728 20556
rect 13780 20544 13786 20596
rect 15562 20584 15568 20596
rect 15523 20556 15568 20584
rect 15562 20544 15568 20556
rect 15620 20544 15626 20596
rect 17497 20587 17555 20593
rect 17497 20553 17509 20587
rect 17543 20584 17555 20587
rect 17678 20584 17684 20596
rect 17543 20556 17684 20584
rect 17543 20553 17555 20556
rect 17497 20547 17555 20553
rect 17678 20544 17684 20556
rect 17736 20544 17742 20596
rect 17862 20584 17868 20596
rect 17823 20556 17868 20584
rect 17862 20544 17868 20556
rect 17920 20544 17926 20596
rect 19058 20584 19064 20596
rect 19019 20556 19064 20584
rect 19058 20544 19064 20556
rect 19116 20544 19122 20596
rect 19334 20544 19340 20596
rect 19392 20584 19398 20596
rect 19429 20587 19487 20593
rect 19429 20584 19441 20587
rect 19392 20556 19441 20584
rect 19392 20544 19398 20556
rect 19429 20553 19441 20556
rect 19475 20553 19487 20587
rect 19429 20547 19487 20553
rect 13906 20516 13912 20528
rect 13867 20488 13912 20516
rect 13906 20476 13912 20488
rect 13964 20476 13970 20528
rect 20714 20476 20720 20528
rect 20772 20516 20778 20528
rect 21545 20519 21603 20525
rect 21545 20516 21557 20519
rect 20772 20488 21557 20516
rect 20772 20476 20778 20488
rect 21545 20485 21557 20488
rect 21591 20485 21603 20519
rect 21545 20479 21603 20485
rect 11793 20383 11851 20389
rect 11793 20349 11805 20383
rect 11839 20380 11851 20383
rect 11974 20380 11980 20392
rect 11839 20352 11980 20380
rect 11839 20349 11851 20352
rect 11793 20343 11851 20349
rect 11974 20340 11980 20352
rect 12032 20380 12038 20392
rect 13357 20383 13415 20389
rect 13357 20380 13369 20383
rect 12032 20352 13369 20380
rect 12032 20340 12038 20352
rect 13357 20349 13369 20352
rect 13403 20380 13415 20383
rect 13924 20380 13952 20476
rect 15654 20448 15660 20460
rect 15396 20420 15660 20448
rect 15396 20389 15424 20420
rect 15654 20408 15660 20420
rect 15712 20448 15718 20460
rect 15841 20451 15899 20457
rect 15841 20448 15853 20451
rect 15712 20420 15853 20448
rect 15712 20408 15718 20420
rect 15841 20417 15853 20420
rect 15887 20448 15899 20451
rect 16022 20448 16028 20460
rect 15887 20420 16028 20448
rect 15887 20417 15899 20420
rect 15841 20411 15899 20417
rect 16022 20408 16028 20420
rect 16080 20408 16086 20460
rect 16114 20408 16120 20460
rect 16172 20448 16178 20460
rect 16393 20451 16451 20457
rect 16393 20448 16405 20451
rect 16172 20420 16405 20448
rect 16172 20408 16178 20420
rect 16393 20417 16405 20420
rect 16439 20417 16451 20451
rect 16393 20411 16451 20417
rect 17586 20408 17592 20460
rect 17644 20448 17650 20460
rect 18049 20451 18107 20457
rect 18049 20448 18061 20451
rect 17644 20420 18061 20448
rect 17644 20408 17650 20420
rect 18049 20417 18061 20420
rect 18095 20448 18107 20451
rect 19426 20448 19432 20460
rect 18095 20420 19432 20448
rect 18095 20417 18107 20420
rect 18049 20411 18107 20417
rect 19426 20408 19432 20420
rect 19484 20408 19490 20460
rect 20530 20408 20536 20460
rect 20588 20448 20594 20460
rect 20588 20420 21404 20448
rect 20588 20408 20594 20420
rect 13403 20352 13952 20380
rect 15381 20383 15439 20389
rect 13403 20349 13415 20352
rect 13357 20343 13415 20349
rect 15381 20349 15393 20383
rect 15427 20349 15439 20383
rect 15381 20343 15439 20349
rect 16301 20383 16359 20389
rect 16301 20349 16313 20383
rect 16347 20380 16359 20383
rect 16942 20380 16948 20392
rect 16347 20352 16948 20380
rect 16347 20349 16359 20352
rect 16301 20343 16359 20349
rect 16942 20340 16948 20352
rect 17000 20340 17006 20392
rect 17310 20340 17316 20392
rect 17368 20380 17374 20392
rect 18141 20383 18199 20389
rect 18141 20380 18153 20383
rect 17368 20352 18153 20380
rect 17368 20340 17374 20352
rect 18141 20349 18153 20352
rect 18187 20349 18199 20383
rect 18141 20343 18199 20349
rect 20165 20383 20223 20389
rect 20165 20349 20177 20383
rect 20211 20349 20223 20383
rect 20165 20343 20223 20349
rect 19978 20244 19984 20256
rect 19939 20216 19984 20244
rect 19978 20204 19984 20216
rect 20036 20244 20042 20256
rect 20180 20244 20208 20343
rect 20254 20340 20260 20392
rect 20312 20380 20318 20392
rect 20625 20383 20683 20389
rect 20625 20380 20637 20383
rect 20312 20352 20637 20380
rect 20312 20340 20318 20352
rect 20625 20349 20637 20352
rect 20671 20349 20683 20383
rect 20625 20343 20683 20349
rect 20714 20340 20720 20392
rect 20772 20380 20778 20392
rect 21376 20389 21404 20420
rect 20993 20383 21051 20389
rect 20993 20380 21005 20383
rect 20772 20352 21005 20380
rect 20772 20340 20778 20352
rect 20993 20349 21005 20352
rect 21039 20349 21051 20383
rect 20993 20343 21051 20349
rect 21361 20383 21419 20389
rect 21361 20349 21373 20383
rect 21407 20349 21419 20383
rect 21361 20343 21419 20349
rect 20036 20216 20208 20244
rect 20036 20204 20042 20216
rect 1104 20154 38824 20176
rect 1104 20102 19606 20154
rect 19658 20102 19670 20154
rect 19722 20102 19734 20154
rect 19786 20102 19798 20154
rect 19850 20102 38824 20154
rect 1104 20080 38824 20102
rect 12066 20000 12072 20052
rect 12124 20040 12130 20052
rect 12434 20040 12440 20052
rect 12124 20012 12440 20040
rect 12124 20000 12130 20012
rect 12434 20000 12440 20012
rect 12492 20040 12498 20052
rect 13909 20043 13967 20049
rect 12492 20012 12585 20040
rect 12492 20000 12498 20012
rect 13909 20009 13921 20043
rect 13955 20040 13967 20043
rect 14734 20040 14740 20052
rect 13955 20012 14740 20040
rect 13955 20009 13967 20012
rect 13909 20003 13967 20009
rect 14734 20000 14740 20012
rect 14792 20040 14798 20052
rect 15470 20040 15476 20052
rect 14792 20012 15476 20040
rect 14792 20000 14798 20012
rect 15470 20000 15476 20012
rect 15528 20000 15534 20052
rect 19150 20040 19156 20052
rect 19111 20012 19156 20040
rect 19150 20000 19156 20012
rect 19208 20000 19214 20052
rect 19426 20040 19432 20052
rect 19387 20012 19432 20040
rect 19426 20000 19432 20012
rect 19484 20000 19490 20052
rect 20254 20040 20260 20052
rect 20215 20012 20260 20040
rect 20254 20000 20260 20012
rect 20312 20000 20318 20052
rect 20530 20040 20536 20052
rect 20491 20012 20536 20040
rect 20530 20000 20536 20012
rect 20588 20000 20594 20052
rect 21358 20040 21364 20052
rect 21319 20012 21364 20040
rect 21358 20000 21364 20012
rect 21416 20000 21422 20052
rect 6089 19975 6147 19981
rect 6089 19941 6101 19975
rect 6135 19972 6147 19975
rect 7834 19972 7840 19984
rect 6135 19944 7840 19972
rect 6135 19941 6147 19944
rect 6089 19935 6147 19941
rect 7834 19932 7840 19944
rect 7892 19932 7898 19984
rect 17678 19932 17684 19984
rect 17736 19972 17742 19984
rect 18693 19975 18751 19981
rect 17736 19944 18368 19972
rect 17736 19932 17742 19944
rect 18340 19916 18368 19944
rect 18693 19941 18705 19975
rect 18739 19972 18751 19975
rect 19978 19972 19984 19984
rect 18739 19944 19984 19972
rect 18739 19941 18751 19944
rect 18693 19935 18751 19941
rect 19978 19932 19984 19944
rect 20036 19932 20042 19984
rect 4433 19907 4491 19913
rect 4433 19873 4445 19907
rect 4479 19904 4491 19907
rect 5442 19904 5448 19916
rect 4479 19876 5448 19904
rect 4479 19873 4491 19876
rect 4433 19867 4491 19873
rect 4908 19848 4936 19876
rect 5442 19864 5448 19876
rect 5500 19864 5506 19916
rect 13630 19864 13636 19916
rect 13688 19904 13694 19916
rect 13725 19907 13783 19913
rect 13725 19904 13737 19907
rect 13688 19876 13737 19904
rect 13688 19864 13694 19876
rect 13725 19873 13737 19876
rect 13771 19873 13783 19907
rect 16022 19904 16028 19916
rect 15983 19876 16028 19904
rect 13725 19867 13783 19873
rect 16022 19864 16028 19876
rect 16080 19864 16086 19916
rect 16298 19864 16304 19916
rect 16356 19904 16362 19916
rect 17589 19907 17647 19913
rect 17589 19904 17601 19907
rect 16356 19876 17601 19904
rect 16356 19864 16362 19876
rect 17589 19873 17601 19876
rect 17635 19904 17647 19907
rect 17954 19904 17960 19916
rect 17635 19876 17960 19904
rect 17635 19873 17647 19876
rect 17589 19867 17647 19873
rect 17954 19864 17960 19876
rect 18012 19864 18018 19916
rect 18138 19904 18144 19916
rect 18099 19876 18144 19904
rect 18138 19864 18144 19876
rect 18196 19864 18202 19916
rect 18322 19904 18328 19916
rect 18283 19876 18328 19904
rect 18322 19864 18328 19876
rect 18380 19864 18386 19916
rect 20901 19907 20959 19913
rect 20901 19873 20913 19907
rect 20947 19904 20959 19907
rect 20990 19904 20996 19916
rect 20947 19876 20996 19904
rect 20947 19873 20959 19876
rect 20901 19867 20959 19873
rect 20990 19864 20996 19876
rect 21048 19904 21054 19916
rect 22002 19904 22008 19916
rect 21048 19876 22008 19904
rect 21048 19864 21054 19876
rect 22002 19864 22008 19876
rect 22060 19864 22066 19916
rect 4706 19836 4712 19848
rect 4667 19808 4712 19836
rect 4706 19796 4712 19808
rect 4764 19796 4770 19848
rect 4890 19796 4896 19848
rect 4948 19796 4954 19848
rect 15933 19839 15991 19845
rect 15933 19805 15945 19839
rect 15979 19836 15991 19839
rect 16206 19836 16212 19848
rect 15979 19808 16212 19836
rect 15979 19805 15991 19808
rect 15933 19799 15991 19805
rect 16206 19796 16212 19808
rect 16264 19836 16270 19848
rect 16761 19839 16819 19845
rect 16761 19836 16773 19839
rect 16264 19808 16773 19836
rect 16264 19796 16270 19808
rect 16761 19805 16773 19808
rect 16807 19836 16819 19839
rect 17405 19839 17463 19845
rect 17405 19836 17417 19839
rect 16807 19808 17417 19836
rect 16807 19805 16819 19808
rect 16761 19799 16819 19805
rect 17405 19805 17417 19808
rect 17451 19836 17463 19839
rect 17770 19836 17776 19848
rect 17451 19808 17776 19836
rect 17451 19805 17463 19808
rect 17405 19799 17463 19805
rect 17770 19796 17776 19808
rect 17828 19796 17834 19848
rect 21082 19768 21088 19780
rect 21043 19740 21088 19768
rect 21082 19728 21088 19740
rect 21140 19728 21146 19780
rect 14918 19700 14924 19712
rect 14879 19672 14924 19700
rect 14918 19660 14924 19672
rect 14976 19660 14982 19712
rect 15930 19660 15936 19712
rect 15988 19700 15994 19712
rect 16209 19703 16267 19709
rect 16209 19700 16221 19703
rect 15988 19672 16221 19700
rect 15988 19660 15994 19672
rect 16209 19669 16221 19672
rect 16255 19669 16267 19703
rect 16209 19663 16267 19669
rect 16758 19660 16764 19712
rect 16816 19700 16822 19712
rect 17221 19703 17279 19709
rect 17221 19700 17233 19703
rect 16816 19672 17233 19700
rect 16816 19660 16822 19672
rect 17221 19669 17233 19672
rect 17267 19700 17279 19703
rect 17310 19700 17316 19712
rect 17267 19672 17316 19700
rect 17267 19669 17279 19672
rect 17221 19663 17279 19669
rect 17310 19660 17316 19672
rect 17368 19660 17374 19712
rect 1104 19610 38824 19632
rect 1104 19558 4246 19610
rect 4298 19558 4310 19610
rect 4362 19558 4374 19610
rect 4426 19558 4438 19610
rect 4490 19558 34966 19610
rect 35018 19558 35030 19610
rect 35082 19558 35094 19610
rect 35146 19558 35158 19610
rect 35210 19558 38824 19610
rect 1104 19536 38824 19558
rect 16022 19496 16028 19508
rect 15983 19468 16028 19496
rect 16022 19456 16028 19468
rect 16080 19456 16086 19508
rect 20070 19496 20076 19508
rect 20031 19468 20076 19496
rect 20070 19456 20076 19468
rect 20128 19456 20134 19508
rect 20990 19496 20996 19508
rect 20951 19468 20996 19496
rect 20990 19456 20996 19468
rect 21048 19456 21054 19508
rect 31478 19496 31484 19508
rect 31439 19468 31484 19496
rect 31478 19456 31484 19468
rect 31536 19456 31542 19508
rect 12434 19320 12440 19372
rect 12492 19360 12498 19372
rect 12713 19363 12771 19369
rect 12492 19332 12537 19360
rect 12492 19320 12498 19332
rect 12713 19329 12725 19363
rect 12759 19360 12771 19363
rect 13630 19360 13636 19372
rect 12759 19332 13636 19360
rect 12759 19329 12771 19332
rect 12713 19323 12771 19329
rect 12253 19295 12311 19301
rect 12253 19261 12265 19295
rect 12299 19292 12311 19295
rect 12728 19292 12756 19323
rect 13630 19320 13636 19332
rect 13688 19320 13694 19372
rect 14182 19320 14188 19372
rect 14240 19360 14246 19372
rect 14918 19360 14924 19372
rect 14240 19332 14924 19360
rect 14240 19320 14246 19332
rect 14918 19320 14924 19332
rect 14976 19320 14982 19372
rect 12299 19264 12756 19292
rect 12299 19261 12311 19264
rect 12253 19255 12311 19261
rect 14274 19252 14280 19304
rect 14332 19292 14338 19304
rect 14737 19295 14795 19301
rect 14737 19292 14749 19295
rect 14332 19264 14749 19292
rect 14332 19252 14338 19264
rect 14737 19261 14749 19264
rect 14783 19261 14795 19295
rect 14737 19255 14795 19261
rect 15013 19295 15071 19301
rect 15013 19261 15025 19295
rect 15059 19261 15071 19295
rect 16574 19292 16580 19304
rect 16535 19264 16580 19292
rect 15013 19255 15071 19261
rect 14458 19224 14464 19236
rect 14419 19196 14464 19224
rect 14458 19184 14464 19196
rect 14516 19184 14522 19236
rect 14752 19224 14780 19255
rect 15028 19224 15056 19255
rect 16574 19252 16580 19264
rect 16632 19252 16638 19304
rect 17865 19295 17923 19301
rect 17865 19261 17877 19295
rect 17911 19292 17923 19295
rect 18138 19292 18144 19304
rect 17911 19264 18144 19292
rect 17911 19261 17923 19264
rect 17865 19255 17923 19261
rect 18138 19252 18144 19264
rect 18196 19252 18202 19304
rect 18782 19292 18788 19304
rect 18743 19264 18788 19292
rect 18782 19252 18788 19264
rect 18840 19252 18846 19304
rect 18966 19252 18972 19304
rect 19024 19301 19030 19304
rect 19024 19295 19073 19301
rect 19024 19261 19027 19295
rect 19061 19261 19073 19295
rect 19150 19292 19156 19304
rect 19111 19264 19156 19292
rect 19024 19255 19073 19261
rect 19024 19252 19030 19255
rect 19150 19252 19156 19264
rect 19208 19252 19214 19304
rect 19426 19252 19432 19304
rect 19484 19292 19490 19304
rect 19521 19295 19579 19301
rect 19521 19292 19533 19295
rect 19484 19264 19533 19292
rect 19484 19252 19490 19264
rect 19521 19261 19533 19264
rect 19567 19261 19579 19295
rect 19521 19255 19579 19261
rect 19613 19295 19671 19301
rect 19613 19261 19625 19295
rect 19659 19261 19671 19295
rect 30098 19292 30104 19304
rect 30059 19264 30104 19292
rect 19613 19255 19671 19261
rect 15470 19224 15476 19236
rect 14752 19196 15056 19224
rect 15431 19196 15476 19224
rect 15470 19184 15476 19196
rect 15528 19184 15534 19236
rect 17129 19227 17187 19233
rect 17129 19193 17141 19227
rect 17175 19224 17187 19227
rect 18414 19224 18420 19236
rect 17175 19196 18420 19224
rect 17175 19193 17187 19196
rect 17129 19187 17187 19193
rect 18414 19184 18420 19196
rect 18472 19184 18478 19236
rect 18800 19224 18828 19252
rect 19628 19224 19656 19255
rect 30098 19252 30104 19264
rect 30156 19252 30162 19304
rect 30377 19295 30435 19301
rect 30377 19292 30389 19295
rect 30208 19264 30389 19292
rect 18800 19196 19656 19224
rect 30009 19227 30067 19233
rect 30009 19193 30021 19227
rect 30055 19224 30067 19227
rect 30208 19224 30236 19264
rect 30377 19261 30389 19264
rect 30423 19292 30435 19295
rect 31662 19292 31668 19304
rect 30423 19264 31668 19292
rect 30423 19261 30435 19264
rect 30377 19255 30435 19261
rect 31662 19252 31668 19264
rect 31720 19252 31726 19304
rect 30055 19196 30236 19224
rect 30055 19193 30067 19196
rect 30009 19187 30067 19193
rect 4430 19156 4436 19168
rect 4391 19128 4436 19156
rect 4430 19116 4436 19128
rect 4488 19156 4494 19168
rect 4706 19156 4712 19168
rect 4488 19128 4712 19156
rect 4488 19116 4494 19128
rect 4706 19116 4712 19128
rect 4764 19116 4770 19168
rect 4890 19156 4896 19168
rect 4851 19128 4896 19156
rect 4890 19116 4896 19128
rect 4948 19116 4954 19168
rect 13814 19156 13820 19168
rect 13775 19128 13820 19156
rect 13814 19116 13820 19128
rect 13872 19116 13878 19168
rect 16666 19116 16672 19168
rect 16724 19156 16730 19168
rect 17405 19159 17463 19165
rect 17405 19156 17417 19159
rect 16724 19128 17417 19156
rect 16724 19116 16730 19128
rect 17405 19125 17417 19128
rect 17451 19156 17463 19159
rect 17678 19156 17684 19168
rect 17451 19128 17684 19156
rect 17451 19125 17463 19128
rect 17405 19119 17463 19125
rect 17678 19116 17684 19128
rect 17736 19116 17742 19168
rect 17954 19116 17960 19168
rect 18012 19156 18018 19168
rect 18233 19159 18291 19165
rect 18233 19156 18245 19159
rect 18012 19128 18245 19156
rect 18012 19116 18018 19128
rect 18233 19125 18245 19128
rect 18279 19125 18291 19159
rect 18233 19119 18291 19125
rect 18966 19116 18972 19168
rect 19024 19156 19030 19168
rect 20533 19159 20591 19165
rect 20533 19156 20545 19159
rect 19024 19128 20545 19156
rect 19024 19116 19030 19128
rect 20533 19125 20545 19128
rect 20579 19125 20591 19159
rect 20533 19119 20591 19125
rect 1104 19066 38824 19088
rect 1104 19014 19606 19066
rect 19658 19014 19670 19066
rect 19722 19014 19734 19066
rect 19786 19014 19798 19066
rect 19850 19014 38824 19066
rect 1104 18992 38824 19014
rect 14185 18955 14243 18961
rect 14185 18921 14197 18955
rect 14231 18921 14243 18955
rect 14185 18915 14243 18921
rect 15013 18955 15071 18961
rect 15013 18921 15025 18955
rect 15059 18952 15071 18955
rect 15470 18952 15476 18964
rect 15059 18924 15476 18952
rect 15059 18921 15071 18924
rect 15013 18915 15071 18921
rect 12342 18844 12348 18896
rect 12400 18884 12406 18896
rect 12400 18856 12940 18884
rect 12400 18844 12406 18856
rect 11330 18776 11336 18828
rect 11388 18816 11394 18828
rect 11793 18819 11851 18825
rect 11793 18816 11805 18819
rect 11388 18788 11805 18816
rect 11388 18776 11394 18788
rect 11793 18785 11805 18788
rect 11839 18816 11851 18819
rect 12526 18816 12532 18828
rect 11839 18788 12532 18816
rect 11839 18785 11851 18788
rect 11793 18779 11851 18785
rect 12526 18776 12532 18788
rect 12584 18776 12590 18828
rect 12912 18825 12940 18856
rect 13906 18844 13912 18896
rect 13964 18884 13970 18896
rect 14200 18884 14228 18915
rect 15470 18912 15476 18924
rect 15528 18912 15534 18964
rect 16574 18912 16580 18964
rect 16632 18952 16638 18964
rect 16761 18955 16819 18961
rect 16761 18952 16773 18955
rect 16632 18924 16773 18952
rect 16632 18912 16638 18924
rect 16761 18921 16773 18924
rect 16807 18921 16819 18955
rect 17770 18952 17776 18964
rect 17731 18924 17776 18952
rect 16761 18915 16819 18921
rect 17770 18912 17776 18924
rect 17828 18912 17834 18964
rect 17954 18912 17960 18964
rect 18012 18952 18018 18964
rect 18417 18955 18475 18961
rect 18417 18952 18429 18955
rect 18012 18924 18429 18952
rect 18012 18912 18018 18924
rect 18417 18921 18429 18924
rect 18463 18952 18475 18955
rect 19150 18952 19156 18964
rect 18463 18924 19156 18952
rect 18463 18921 18475 18924
rect 18417 18915 18475 18921
rect 19150 18912 19156 18924
rect 19208 18912 19214 18964
rect 23842 18952 23848 18964
rect 23803 18924 23848 18952
rect 23842 18912 23848 18924
rect 23900 18912 23906 18964
rect 15746 18884 15752 18896
rect 13964 18856 15752 18884
rect 13964 18844 13970 18856
rect 15746 18844 15752 18856
rect 15804 18844 15810 18896
rect 19613 18887 19671 18893
rect 19613 18853 19625 18887
rect 19659 18884 19671 18887
rect 20254 18884 20260 18896
rect 19659 18856 20260 18884
rect 19659 18853 19671 18856
rect 19613 18847 19671 18853
rect 20254 18844 20260 18856
rect 20312 18844 20318 18896
rect 12897 18819 12955 18825
rect 12897 18785 12909 18819
rect 12943 18816 12955 18819
rect 13814 18816 13820 18828
rect 12943 18788 13820 18816
rect 12943 18785 12955 18788
rect 12897 18779 12955 18785
rect 13814 18776 13820 18788
rect 13872 18776 13878 18828
rect 14001 18819 14059 18825
rect 14001 18785 14013 18819
rect 14047 18816 14059 18819
rect 14458 18816 14464 18828
rect 14047 18788 14464 18816
rect 14047 18785 14059 18788
rect 14001 18779 14059 18785
rect 11882 18748 11888 18760
rect 11843 18720 11888 18748
rect 11882 18708 11888 18720
rect 11940 18708 11946 18760
rect 12621 18751 12679 18757
rect 12621 18717 12633 18751
rect 12667 18717 12679 18751
rect 12802 18748 12808 18760
rect 12763 18720 12808 18748
rect 12621 18711 12679 18717
rect 12066 18640 12072 18692
rect 12124 18680 12130 18692
rect 12636 18680 12664 18711
rect 12802 18708 12808 18720
rect 12860 18708 12866 18760
rect 13446 18748 13452 18760
rect 13359 18720 13452 18748
rect 13446 18708 13452 18720
rect 13504 18748 13510 18760
rect 14016 18748 14044 18779
rect 14458 18776 14464 18788
rect 14516 18776 14522 18828
rect 15930 18816 15936 18828
rect 15891 18788 15936 18816
rect 15930 18776 15936 18788
rect 15988 18776 15994 18828
rect 16298 18816 16304 18828
rect 16259 18788 16304 18816
rect 16298 18776 16304 18788
rect 16356 18776 16362 18828
rect 17310 18816 17316 18828
rect 17271 18788 17316 18816
rect 17310 18776 17316 18788
rect 17368 18776 17374 18828
rect 18414 18776 18420 18828
rect 18472 18816 18478 18828
rect 18509 18819 18567 18825
rect 18509 18816 18521 18819
rect 18472 18788 18521 18816
rect 18472 18776 18478 18788
rect 18509 18785 18521 18788
rect 18555 18785 18567 18819
rect 18509 18779 18567 18785
rect 18782 18776 18788 18828
rect 18840 18816 18846 18828
rect 18877 18819 18935 18825
rect 18877 18816 18889 18819
rect 18840 18788 18889 18816
rect 18840 18776 18846 18788
rect 18877 18785 18889 18788
rect 18923 18785 18935 18819
rect 18877 18779 18935 18785
rect 19334 18776 19340 18828
rect 19392 18816 19398 18828
rect 19429 18819 19487 18825
rect 19429 18816 19441 18819
rect 19392 18788 19441 18816
rect 19392 18776 19398 18788
rect 19429 18785 19441 18788
rect 19475 18816 19487 18819
rect 20438 18816 20444 18828
rect 19475 18788 20444 18816
rect 19475 18785 19487 18788
rect 19429 18779 19487 18785
rect 20438 18776 20444 18788
rect 20496 18776 20502 18828
rect 22738 18816 22744 18828
rect 22699 18788 22744 18816
rect 22738 18776 22744 18788
rect 22796 18776 22802 18828
rect 16390 18748 16396 18760
rect 13504 18720 14044 18748
rect 16351 18720 16396 18748
rect 13504 18708 13510 18720
rect 16390 18708 16396 18720
rect 16448 18708 16454 18760
rect 22462 18748 22468 18760
rect 22423 18720 22468 18748
rect 22462 18708 22468 18720
rect 22520 18708 22526 18760
rect 14734 18680 14740 18692
rect 12124 18652 14740 18680
rect 12124 18640 12130 18652
rect 14734 18640 14740 18652
rect 14792 18640 14798 18692
rect 15746 18680 15752 18692
rect 15707 18652 15752 18680
rect 15746 18640 15752 18652
rect 15804 18640 15810 18692
rect 12434 18572 12440 18624
rect 12492 18612 12498 18624
rect 13354 18612 13360 18624
rect 12492 18584 13360 18612
rect 12492 18572 12498 18584
rect 13354 18572 13360 18584
rect 13412 18612 13418 18624
rect 13725 18615 13783 18621
rect 13725 18612 13737 18615
rect 13412 18584 13737 18612
rect 13412 18572 13418 18584
rect 13725 18581 13737 18584
rect 13771 18581 13783 18615
rect 17494 18612 17500 18624
rect 17455 18584 17500 18612
rect 13725 18575 13783 18581
rect 17494 18572 17500 18584
rect 17552 18572 17558 18624
rect 30098 18612 30104 18624
rect 30059 18584 30104 18612
rect 30098 18572 30104 18584
rect 30156 18572 30162 18624
rect 1104 18522 38824 18544
rect 1104 18470 4246 18522
rect 4298 18470 4310 18522
rect 4362 18470 4374 18522
rect 4426 18470 4438 18522
rect 4490 18470 34966 18522
rect 35018 18470 35030 18522
rect 35082 18470 35094 18522
rect 35146 18470 35158 18522
rect 35210 18470 38824 18522
rect 1104 18448 38824 18470
rect 11977 18411 12035 18417
rect 11977 18377 11989 18411
rect 12023 18408 12035 18411
rect 12066 18408 12072 18420
rect 12023 18380 12072 18408
rect 12023 18377 12035 18380
rect 11977 18371 12035 18377
rect 12066 18368 12072 18380
rect 12124 18368 12130 18420
rect 14458 18408 14464 18420
rect 14419 18380 14464 18408
rect 14458 18368 14464 18380
rect 14516 18368 14522 18420
rect 14734 18408 14740 18420
rect 14695 18380 14740 18408
rect 14734 18368 14740 18380
rect 14792 18408 14798 18420
rect 14792 18380 15792 18408
rect 14792 18368 14798 18380
rect 9858 18272 9864 18284
rect 9819 18244 9864 18272
rect 9858 18232 9864 18244
rect 9916 18232 9922 18284
rect 12434 18272 12440 18284
rect 12395 18244 12440 18272
rect 12434 18232 12440 18244
rect 12492 18232 12498 18284
rect 12713 18275 12771 18281
rect 12713 18241 12725 18275
rect 12759 18272 12771 18275
rect 13446 18272 13452 18284
rect 12759 18244 13452 18272
rect 12759 18241 12771 18244
rect 12713 18235 12771 18241
rect 13446 18232 13452 18244
rect 13504 18232 13510 18284
rect 10137 18207 10195 18213
rect 10137 18204 10149 18207
rect 9968 18176 10149 18204
rect 9674 18068 9680 18080
rect 9635 18040 9680 18068
rect 9674 18028 9680 18040
rect 9732 18068 9738 18080
rect 9968 18068 9996 18176
rect 10137 18173 10149 18176
rect 10183 18173 10195 18207
rect 10137 18167 10195 18173
rect 11517 18207 11575 18213
rect 11517 18173 11529 18207
rect 11563 18204 11575 18207
rect 12158 18204 12164 18216
rect 11563 18176 12164 18204
rect 11563 18173 11575 18176
rect 11517 18167 11575 18173
rect 12158 18164 12164 18176
rect 12216 18204 12222 18216
rect 15381 18207 15439 18213
rect 12216 18176 14412 18204
rect 12216 18164 12222 18176
rect 13814 18068 13820 18080
rect 9732 18040 9996 18068
rect 13775 18040 13820 18068
rect 9732 18028 9738 18040
rect 13814 18028 13820 18040
rect 13872 18028 13878 18080
rect 14384 18068 14412 18176
rect 15381 18173 15393 18207
rect 15427 18204 15439 18207
rect 15470 18204 15476 18216
rect 15427 18176 15476 18204
rect 15427 18173 15439 18176
rect 15381 18167 15439 18173
rect 15470 18164 15476 18176
rect 15528 18164 15534 18216
rect 15562 18164 15568 18216
rect 15620 18204 15626 18216
rect 15764 18213 15792 18380
rect 15930 18368 15936 18420
rect 15988 18408 15994 18420
rect 16945 18411 17003 18417
rect 16945 18408 16957 18411
rect 15988 18380 16957 18408
rect 15988 18368 15994 18380
rect 16945 18377 16957 18380
rect 16991 18377 17003 18411
rect 17310 18408 17316 18420
rect 17271 18380 17316 18408
rect 16945 18371 17003 18377
rect 17310 18368 17316 18380
rect 17368 18368 17374 18420
rect 18138 18368 18144 18420
rect 18196 18408 18202 18420
rect 18509 18411 18567 18417
rect 18509 18408 18521 18411
rect 18196 18380 18521 18408
rect 18196 18368 18202 18380
rect 18509 18377 18521 18380
rect 18555 18377 18567 18411
rect 18966 18408 18972 18420
rect 18927 18380 18972 18408
rect 18509 18371 18567 18377
rect 16298 18340 16304 18352
rect 16259 18312 16304 18340
rect 16298 18300 16304 18312
rect 16356 18300 16362 18352
rect 15749 18207 15807 18213
rect 15620 18176 15665 18204
rect 15620 18164 15626 18176
rect 15749 18173 15761 18207
rect 15795 18173 15807 18207
rect 18524 18204 18552 18371
rect 18966 18368 18972 18380
rect 19024 18368 19030 18420
rect 22557 18411 22615 18417
rect 22557 18377 22569 18411
rect 22603 18408 22615 18411
rect 22738 18408 22744 18420
rect 22603 18380 22744 18408
rect 22603 18377 22615 18380
rect 22557 18371 22615 18377
rect 22738 18368 22744 18380
rect 22796 18368 22802 18420
rect 18785 18207 18843 18213
rect 18785 18204 18797 18207
rect 18524 18176 18797 18204
rect 15749 18167 15807 18173
rect 18785 18173 18797 18176
rect 18831 18173 18843 18207
rect 18785 18167 18843 18173
rect 14918 18136 14924 18148
rect 14879 18108 14924 18136
rect 14918 18096 14924 18108
rect 14976 18096 14982 18148
rect 15580 18136 15608 18164
rect 16390 18136 16396 18148
rect 15580 18108 16396 18136
rect 16390 18096 16396 18108
rect 16448 18136 16454 18148
rect 16577 18139 16635 18145
rect 16577 18136 16589 18139
rect 16448 18108 16589 18136
rect 16448 18096 16454 18108
rect 16577 18105 16589 18108
rect 16623 18136 16635 18139
rect 17034 18136 17040 18148
rect 16623 18108 17040 18136
rect 16623 18105 16635 18108
rect 16577 18099 16635 18105
rect 17034 18096 17040 18108
rect 17092 18096 17098 18148
rect 17954 18136 17960 18148
rect 17144 18108 17960 18136
rect 17144 18068 17172 18108
rect 17954 18096 17960 18108
rect 18012 18096 18018 18148
rect 14384 18040 17172 18068
rect 17865 18071 17923 18077
rect 17865 18037 17877 18071
rect 17911 18068 17923 18071
rect 18782 18068 18788 18080
rect 17911 18040 18788 18068
rect 17911 18037 17923 18040
rect 17865 18031 17923 18037
rect 18782 18028 18788 18040
rect 18840 18028 18846 18080
rect 22094 18028 22100 18080
rect 22152 18068 22158 18080
rect 22462 18068 22468 18080
rect 22152 18040 22468 18068
rect 22152 18028 22158 18040
rect 22462 18028 22468 18040
rect 22520 18068 22526 18080
rect 22833 18071 22891 18077
rect 22833 18068 22845 18071
rect 22520 18040 22845 18068
rect 22520 18028 22526 18040
rect 22833 18037 22845 18040
rect 22879 18037 22891 18071
rect 22833 18031 22891 18037
rect 1104 17978 38824 18000
rect 1104 17926 19606 17978
rect 19658 17926 19670 17978
rect 19722 17926 19734 17978
rect 19786 17926 19798 17978
rect 19850 17926 38824 17978
rect 1104 17904 38824 17926
rect 9858 17864 9864 17876
rect 9819 17836 9864 17864
rect 9858 17824 9864 17836
rect 9916 17824 9922 17876
rect 11517 17867 11575 17873
rect 11517 17833 11529 17867
rect 11563 17864 11575 17867
rect 12342 17864 12348 17876
rect 11563 17836 12348 17864
rect 11563 17833 11575 17836
rect 11517 17827 11575 17833
rect 12342 17824 12348 17836
rect 12400 17824 12406 17876
rect 14826 17824 14832 17876
rect 14884 17864 14890 17876
rect 14921 17867 14979 17873
rect 14921 17864 14933 17867
rect 14884 17836 14933 17864
rect 14884 17824 14890 17836
rect 14921 17833 14933 17836
rect 14967 17833 14979 17867
rect 14921 17827 14979 17833
rect 18414 17824 18420 17876
rect 18472 17864 18478 17876
rect 18509 17867 18567 17873
rect 18509 17864 18521 17867
rect 18472 17836 18521 17864
rect 18472 17824 18478 17836
rect 18509 17833 18521 17836
rect 18555 17833 18567 17867
rect 18509 17827 18567 17833
rect 18969 17867 19027 17873
rect 18969 17833 18981 17867
rect 19015 17864 19027 17867
rect 19242 17864 19248 17876
rect 19015 17836 19248 17864
rect 19015 17833 19027 17836
rect 18969 17827 19027 17833
rect 19242 17824 19248 17836
rect 19300 17824 19306 17876
rect 11885 17799 11943 17805
rect 11885 17765 11897 17799
rect 11931 17796 11943 17799
rect 12802 17796 12808 17808
rect 11931 17768 12808 17796
rect 11931 17765 11943 17768
rect 11885 17759 11943 17765
rect 12802 17756 12808 17768
rect 12860 17756 12866 17808
rect 17862 17756 17868 17808
rect 17920 17796 17926 17808
rect 19061 17799 19119 17805
rect 19061 17796 19073 17799
rect 17920 17768 19073 17796
rect 17920 17756 17926 17768
rect 19061 17765 19073 17768
rect 19107 17765 19119 17799
rect 19061 17759 19119 17765
rect 12618 17728 12624 17740
rect 12579 17700 12624 17728
rect 12618 17688 12624 17700
rect 12676 17688 12682 17740
rect 11974 17660 11980 17672
rect 11935 17632 11980 17660
rect 11974 17620 11980 17632
rect 12032 17620 12038 17672
rect 12713 17663 12771 17669
rect 12713 17629 12725 17663
rect 12759 17629 12771 17663
rect 12820 17660 12848 17756
rect 12986 17728 12992 17740
rect 12899 17700 12992 17728
rect 12986 17688 12992 17700
rect 13044 17728 13050 17740
rect 13722 17728 13728 17740
rect 13044 17700 13728 17728
rect 13044 17688 13050 17700
rect 13722 17688 13728 17700
rect 13780 17688 13786 17740
rect 15378 17728 15384 17740
rect 15339 17700 15384 17728
rect 15378 17688 15384 17700
rect 15436 17688 15442 17740
rect 17034 17728 17040 17740
rect 16995 17700 17040 17728
rect 17034 17688 17040 17700
rect 17092 17688 17098 17740
rect 17494 17688 17500 17740
rect 17552 17728 17558 17740
rect 17589 17731 17647 17737
rect 17589 17728 17601 17731
rect 17552 17700 17601 17728
rect 17552 17688 17558 17700
rect 17589 17697 17601 17700
rect 17635 17697 17647 17731
rect 17589 17691 17647 17697
rect 17773 17731 17831 17737
rect 17773 17697 17785 17731
rect 17819 17728 17831 17731
rect 17880 17728 17908 17756
rect 17819 17700 17908 17728
rect 17819 17697 17831 17700
rect 17773 17691 17831 17697
rect 17954 17688 17960 17740
rect 18012 17728 18018 17740
rect 19150 17728 19156 17740
rect 18012 17700 19156 17728
rect 18012 17688 18018 17700
rect 19150 17688 19156 17700
rect 19208 17728 19214 17740
rect 19705 17731 19763 17737
rect 19705 17728 19717 17731
rect 19208 17700 19717 17728
rect 19208 17688 19214 17700
rect 19705 17697 19717 17700
rect 19751 17728 19763 17731
rect 20070 17728 20076 17740
rect 19751 17700 20076 17728
rect 19751 17697 19763 17700
rect 19705 17691 19763 17697
rect 20070 17688 20076 17700
rect 20128 17688 20134 17740
rect 12897 17663 12955 17669
rect 12897 17660 12909 17663
rect 12820 17632 12909 17660
rect 12713 17623 12771 17629
rect 12897 17629 12909 17632
rect 12943 17629 12955 17663
rect 15286 17660 15292 17672
rect 15247 17632 15292 17660
rect 12897 17623 12955 17629
rect 12158 17552 12164 17604
rect 12216 17592 12222 17604
rect 12728 17592 12756 17623
rect 15286 17620 15292 17632
rect 15344 17620 15350 17672
rect 16942 17660 16948 17672
rect 16855 17632 16948 17660
rect 16942 17620 16948 17632
rect 17000 17620 17006 17672
rect 13722 17592 13728 17604
rect 12216 17564 13728 17592
rect 12216 17552 12222 17564
rect 13722 17552 13728 17564
rect 13780 17552 13786 17604
rect 16960 17592 16988 17620
rect 18598 17592 18604 17604
rect 16960 17564 18604 17592
rect 18598 17552 18604 17564
rect 18656 17552 18662 17604
rect 9858 17484 9864 17536
rect 9916 17524 9922 17536
rect 12894 17524 12900 17536
rect 9916 17496 12900 17524
rect 9916 17484 9922 17496
rect 12894 17484 12900 17496
rect 12952 17524 12958 17536
rect 13449 17527 13507 17533
rect 13449 17524 13461 17527
rect 12952 17496 13461 17524
rect 12952 17484 12958 17496
rect 13449 17493 13461 17496
rect 13495 17493 13507 17527
rect 15562 17524 15568 17536
rect 15523 17496 15568 17524
rect 13449 17487 13507 17493
rect 15562 17484 15568 17496
rect 15620 17484 15626 17536
rect 16209 17527 16267 17533
rect 16209 17493 16221 17527
rect 16255 17524 16267 17527
rect 16482 17524 16488 17536
rect 16255 17496 16488 17524
rect 16255 17493 16267 17496
rect 16209 17487 16267 17493
rect 16482 17484 16488 17496
rect 16540 17484 16546 17536
rect 18049 17527 18107 17533
rect 18049 17493 18061 17527
rect 18095 17524 18107 17527
rect 18414 17524 18420 17536
rect 18095 17496 18420 17524
rect 18095 17493 18107 17496
rect 18049 17487 18107 17493
rect 18414 17484 18420 17496
rect 18472 17484 18478 17536
rect 1104 17434 38824 17456
rect 1104 17382 4246 17434
rect 4298 17382 4310 17434
rect 4362 17382 4374 17434
rect 4426 17382 4438 17434
rect 4490 17382 34966 17434
rect 35018 17382 35030 17434
rect 35082 17382 35094 17434
rect 35146 17382 35158 17434
rect 35210 17382 38824 17434
rect 1104 17360 38824 17382
rect 8386 17320 8392 17332
rect 8347 17292 8392 17320
rect 8386 17280 8392 17292
rect 8444 17280 8450 17332
rect 11701 17323 11759 17329
rect 11701 17289 11713 17323
rect 11747 17320 11759 17323
rect 12618 17320 12624 17332
rect 11747 17292 12624 17320
rect 11747 17289 11759 17292
rect 11701 17283 11759 17289
rect 12618 17280 12624 17292
rect 12676 17280 12682 17332
rect 12713 17323 12771 17329
rect 12713 17289 12725 17323
rect 12759 17320 12771 17323
rect 12802 17320 12808 17332
rect 12759 17292 12808 17320
rect 12759 17289 12771 17292
rect 12713 17283 12771 17289
rect 12802 17280 12808 17292
rect 12860 17280 12866 17332
rect 14461 17323 14519 17329
rect 14461 17289 14473 17323
rect 14507 17320 14519 17323
rect 14921 17323 14979 17329
rect 14921 17320 14933 17323
rect 14507 17292 14933 17320
rect 14507 17289 14519 17292
rect 14461 17283 14519 17289
rect 14921 17289 14933 17292
rect 14967 17320 14979 17323
rect 15286 17320 15292 17332
rect 14967 17292 15292 17320
rect 14967 17289 14979 17292
rect 14921 17283 14979 17289
rect 15286 17280 15292 17292
rect 15344 17280 15350 17332
rect 17494 17280 17500 17332
rect 17552 17320 17558 17332
rect 18233 17323 18291 17329
rect 18233 17320 18245 17323
rect 17552 17292 18245 17320
rect 17552 17280 17558 17292
rect 18233 17289 18245 17292
rect 18279 17289 18291 17323
rect 18598 17320 18604 17332
rect 18559 17292 18604 17320
rect 18233 17283 18291 17289
rect 18598 17280 18604 17292
rect 18656 17280 18662 17332
rect 19150 17320 19156 17332
rect 19111 17292 19156 17320
rect 19150 17280 19156 17292
rect 19208 17280 19214 17332
rect 12069 17255 12127 17261
rect 12069 17221 12081 17255
rect 12115 17252 12127 17255
rect 12158 17252 12164 17264
rect 12115 17224 12164 17252
rect 12115 17221 12127 17224
rect 12069 17215 12127 17221
rect 12158 17212 12164 17224
rect 12216 17212 12222 17264
rect 17405 17255 17463 17261
rect 17405 17221 17417 17255
rect 17451 17252 17463 17255
rect 17862 17252 17868 17264
rect 17451 17224 17868 17252
rect 17451 17221 17463 17224
rect 17405 17215 17463 17221
rect 17862 17212 17868 17224
rect 17920 17212 17926 17264
rect 12894 17184 12900 17196
rect 12855 17156 12900 17184
rect 12894 17144 12900 17156
rect 12952 17144 12958 17196
rect 13173 17187 13231 17193
rect 13173 17153 13185 17187
rect 13219 17184 13231 17187
rect 13538 17184 13544 17196
rect 13219 17156 13544 17184
rect 13219 17153 13231 17156
rect 13173 17147 13231 17153
rect 13538 17144 13544 17156
rect 13596 17144 13602 17196
rect 15289 17187 15347 17193
rect 15289 17153 15301 17187
rect 15335 17184 15347 17187
rect 15378 17184 15384 17196
rect 15335 17156 15384 17184
rect 15335 17153 15347 17156
rect 15289 17147 15347 17153
rect 15378 17144 15384 17156
rect 15436 17144 15442 17196
rect 15657 17187 15715 17193
rect 15657 17153 15669 17187
rect 15703 17184 15715 17187
rect 15703 17156 16160 17184
rect 15703 17153 15715 17156
rect 15657 17147 15715 17153
rect 8573 17119 8631 17125
rect 8573 17085 8585 17119
rect 8619 17116 8631 17119
rect 15749 17119 15807 17125
rect 8619 17088 8984 17116
rect 8619 17085 8631 17088
rect 8573 17079 8631 17085
rect 8956 16989 8984 17088
rect 15749 17085 15761 17119
rect 15795 17116 15807 17119
rect 15838 17116 15844 17128
rect 15795 17088 15844 17116
rect 15795 17085 15807 17088
rect 15749 17079 15807 17085
rect 15838 17076 15844 17088
rect 15896 17076 15902 17128
rect 15933 17119 15991 17125
rect 15933 17085 15945 17119
rect 15979 17085 15991 17119
rect 16132 17116 16160 17156
rect 16942 17144 16948 17196
rect 17000 17184 17006 17196
rect 17773 17187 17831 17193
rect 17773 17184 17785 17187
rect 17000 17156 17785 17184
rect 17000 17144 17006 17156
rect 17773 17153 17785 17156
rect 17819 17153 17831 17187
rect 17773 17147 17831 17153
rect 16390 17116 16396 17128
rect 16132 17088 16396 17116
rect 15933 17079 15991 17085
rect 15948 17048 15976 17079
rect 16390 17076 16396 17088
rect 16448 17076 16454 17128
rect 16482 17076 16488 17128
rect 16540 17116 16546 17128
rect 17494 17116 17500 17128
rect 16540 17088 17500 17116
rect 16540 17076 16546 17088
rect 17494 17076 17500 17088
rect 17552 17076 17558 17128
rect 16500 17048 16528 17076
rect 15948 17020 16528 17048
rect 17037 17051 17095 17057
rect 17037 17017 17049 17051
rect 17083 17048 17095 17051
rect 17310 17048 17316 17060
rect 17083 17020 17316 17048
rect 17083 17017 17095 17020
rect 17037 17011 17095 17017
rect 17310 17008 17316 17020
rect 17368 17008 17374 17060
rect 8941 16983 8999 16989
rect 8941 16949 8953 16983
rect 8987 16980 8999 16983
rect 9490 16980 9496 16992
rect 8987 16952 9496 16980
rect 8987 16949 8999 16952
rect 8941 16943 8999 16949
rect 9490 16940 9496 16952
rect 9548 16940 9554 16992
rect 1104 16890 38824 16912
rect 1104 16838 19606 16890
rect 19658 16838 19670 16890
rect 19722 16838 19734 16890
rect 19786 16838 19798 16890
rect 19850 16838 38824 16890
rect 1104 16816 38824 16838
rect 1394 16736 1400 16788
rect 1452 16776 1458 16788
rect 1581 16779 1639 16785
rect 1581 16776 1593 16779
rect 1452 16748 1593 16776
rect 1452 16736 1458 16748
rect 1581 16745 1593 16748
rect 1627 16745 1639 16779
rect 1581 16739 1639 16745
rect 12069 16779 12127 16785
rect 12069 16745 12081 16779
rect 12115 16776 12127 16779
rect 12986 16776 12992 16788
rect 12115 16748 12992 16776
rect 12115 16745 12127 16748
rect 12069 16739 12127 16745
rect 12986 16736 12992 16748
rect 13044 16736 13050 16788
rect 15838 16776 15844 16788
rect 15799 16748 15844 16776
rect 15838 16736 15844 16748
rect 15896 16736 15902 16788
rect 15562 16708 15568 16720
rect 13832 16680 15568 16708
rect 13832 16652 13860 16680
rect 15562 16668 15568 16680
rect 15620 16668 15626 16720
rect 25314 16708 25320 16720
rect 25275 16680 25320 16708
rect 25314 16668 25320 16680
rect 25372 16668 25378 16720
rect 12989 16643 13047 16649
rect 12989 16609 13001 16643
rect 13035 16640 13047 16643
rect 13538 16640 13544 16652
rect 13035 16612 13544 16640
rect 13035 16609 13047 16612
rect 12989 16603 13047 16609
rect 13538 16600 13544 16612
rect 13596 16640 13602 16652
rect 13814 16640 13820 16652
rect 13596 16612 13676 16640
rect 13727 16612 13820 16640
rect 13596 16600 13602 16612
rect 13648 16572 13676 16612
rect 13814 16600 13820 16612
rect 13872 16600 13878 16652
rect 14001 16643 14059 16649
rect 14001 16609 14013 16643
rect 14047 16609 14059 16643
rect 14001 16603 14059 16609
rect 14185 16643 14243 16649
rect 14185 16609 14197 16643
rect 14231 16640 14243 16643
rect 15010 16640 15016 16652
rect 14231 16612 15016 16640
rect 14231 16609 14243 16612
rect 14185 16603 14243 16609
rect 14016 16572 14044 16603
rect 14090 16572 14096 16584
rect 13648 16544 14096 16572
rect 14090 16532 14096 16544
rect 14148 16532 14154 16584
rect 13630 16504 13636 16516
rect 13591 16476 13636 16504
rect 13630 16464 13636 16476
rect 13688 16464 13694 16516
rect 13722 16464 13728 16516
rect 13780 16504 13786 16516
rect 14200 16504 14228 16603
rect 15010 16600 15016 16612
rect 15068 16600 15074 16652
rect 16209 16643 16267 16649
rect 16209 16609 16221 16643
rect 16255 16640 16267 16643
rect 16945 16643 17003 16649
rect 16945 16640 16957 16643
rect 16255 16612 16957 16640
rect 16255 16609 16267 16612
rect 16209 16603 16267 16609
rect 16945 16609 16957 16612
rect 16991 16640 17003 16643
rect 17494 16640 17500 16652
rect 16991 16612 17500 16640
rect 16991 16609 17003 16612
rect 16945 16603 17003 16609
rect 17494 16600 17500 16612
rect 17552 16600 17558 16652
rect 17678 16640 17684 16652
rect 17591 16612 17684 16640
rect 17678 16600 17684 16612
rect 17736 16640 17742 16652
rect 18322 16640 18328 16652
rect 17736 16612 18328 16640
rect 17736 16600 17742 16612
rect 18322 16600 18328 16612
rect 18380 16600 18386 16652
rect 23661 16643 23719 16649
rect 23661 16609 23673 16643
rect 23707 16640 23719 16643
rect 24302 16640 24308 16652
rect 23707 16612 24308 16640
rect 23707 16609 23719 16612
rect 23661 16603 23719 16609
rect 24302 16600 24308 16612
rect 24360 16600 24366 16652
rect 16390 16532 16396 16584
rect 16448 16572 16454 16584
rect 16758 16572 16764 16584
rect 16448 16544 16764 16572
rect 16448 16532 16454 16544
rect 16758 16532 16764 16544
rect 16816 16532 16822 16584
rect 23842 16532 23848 16584
rect 23900 16572 23906 16584
rect 23937 16575 23995 16581
rect 23937 16572 23949 16575
rect 23900 16544 23949 16572
rect 23900 16532 23906 16544
rect 23937 16541 23949 16544
rect 23983 16541 23995 16575
rect 23937 16535 23995 16541
rect 13780 16476 14228 16504
rect 13780 16464 13786 16476
rect 17954 16436 17960 16448
rect 17915 16408 17960 16436
rect 17954 16396 17960 16408
rect 18012 16396 18018 16448
rect 1104 16346 38824 16368
rect 1104 16294 4246 16346
rect 4298 16294 4310 16346
rect 4362 16294 4374 16346
rect 4426 16294 4438 16346
rect 4490 16294 34966 16346
rect 35018 16294 35030 16346
rect 35082 16294 35094 16346
rect 35146 16294 35158 16346
rect 35210 16294 38824 16346
rect 1104 16272 38824 16294
rect 2961 16235 3019 16241
rect 2961 16201 2973 16235
rect 3007 16232 3019 16235
rect 3234 16232 3240 16244
rect 3007 16204 3240 16232
rect 3007 16201 3019 16204
rect 2961 16195 3019 16201
rect 3234 16192 3240 16204
rect 3292 16192 3298 16244
rect 13814 16232 13820 16244
rect 13775 16204 13820 16232
rect 13814 16192 13820 16204
rect 13872 16192 13878 16244
rect 14090 16232 14096 16244
rect 14051 16204 14096 16232
rect 14090 16192 14096 16204
rect 14148 16192 14154 16244
rect 17221 16235 17279 16241
rect 17221 16201 17233 16235
rect 17267 16232 17279 16235
rect 17494 16232 17500 16244
rect 17267 16204 17500 16232
rect 17267 16201 17279 16204
rect 17221 16195 17279 16201
rect 17494 16192 17500 16204
rect 17552 16192 17558 16244
rect 9490 16124 9496 16176
rect 9548 16164 9554 16176
rect 10045 16167 10103 16173
rect 10045 16164 10057 16167
rect 9548 16136 10057 16164
rect 9548 16124 9554 16136
rect 10045 16133 10057 16136
rect 10091 16164 10103 16167
rect 10962 16164 10968 16176
rect 10091 16136 10968 16164
rect 10091 16133 10103 16136
rect 10045 16127 10103 16133
rect 10962 16124 10968 16136
rect 11020 16124 11026 16176
rect 13449 16167 13507 16173
rect 13449 16133 13461 16167
rect 13495 16164 13507 16167
rect 13722 16164 13728 16176
rect 13495 16136 13728 16164
rect 13495 16133 13507 16136
rect 13449 16127 13507 16133
rect 13722 16124 13728 16136
rect 13780 16124 13786 16176
rect 16853 16167 16911 16173
rect 16853 16133 16865 16167
rect 16899 16164 16911 16167
rect 17678 16164 17684 16176
rect 16899 16136 17684 16164
rect 16899 16133 16911 16136
rect 16853 16127 16911 16133
rect 17678 16124 17684 16136
rect 17736 16124 17742 16176
rect 1394 16096 1400 16108
rect 1355 16068 1400 16096
rect 1394 16056 1400 16068
rect 1452 16056 1458 16108
rect 1578 16056 1584 16108
rect 1636 16096 1642 16108
rect 1673 16099 1731 16105
rect 1673 16096 1685 16099
rect 1636 16068 1685 16096
rect 1636 16056 1642 16068
rect 1673 16065 1685 16068
rect 1719 16065 1731 16099
rect 1673 16059 1731 16065
rect 10226 16028 10232 16040
rect 10187 16000 10232 16028
rect 10226 15988 10232 16000
rect 10284 16028 10290 16040
rect 10505 16031 10563 16037
rect 10505 16028 10517 16031
rect 10284 16000 10517 16028
rect 10284 15988 10290 16000
rect 10505 15997 10517 16000
rect 10551 15997 10563 16031
rect 10505 15991 10563 15997
rect 15197 16031 15255 16037
rect 15197 15997 15209 16031
rect 15243 16028 15255 16031
rect 15654 16028 15660 16040
rect 15243 16000 15660 16028
rect 15243 15997 15255 16000
rect 15197 15991 15255 15997
rect 15654 15988 15660 16000
rect 15712 15988 15718 16040
rect 14826 15920 14832 15972
rect 14884 15960 14890 15972
rect 16390 15960 16396 15972
rect 14884 15932 16396 15960
rect 14884 15920 14890 15932
rect 16390 15920 16396 15932
rect 16448 15920 16454 15972
rect 15378 15892 15384 15904
rect 15339 15864 15384 15892
rect 15378 15852 15384 15864
rect 15436 15852 15442 15904
rect 23842 15892 23848 15904
rect 23803 15864 23848 15892
rect 23842 15852 23848 15864
rect 23900 15852 23906 15904
rect 24302 15892 24308 15904
rect 24215 15864 24308 15892
rect 24302 15852 24308 15864
rect 24360 15892 24366 15904
rect 24762 15892 24768 15904
rect 24360 15864 24768 15892
rect 24360 15852 24366 15864
rect 24762 15852 24768 15864
rect 24820 15852 24826 15904
rect 1104 15802 38824 15824
rect 1104 15750 19606 15802
rect 19658 15750 19670 15802
rect 19722 15750 19734 15802
rect 19786 15750 19798 15802
rect 19850 15750 38824 15802
rect 1104 15728 38824 15750
rect 17954 15648 17960 15700
rect 18012 15688 18018 15700
rect 18417 15691 18475 15697
rect 18417 15688 18429 15691
rect 18012 15660 18429 15688
rect 18012 15648 18018 15660
rect 18417 15657 18429 15660
rect 18463 15657 18475 15691
rect 18417 15651 18475 15657
rect 18046 15620 18052 15632
rect 18007 15592 18052 15620
rect 18046 15580 18052 15592
rect 18104 15580 18110 15632
rect 21174 15552 21180 15564
rect 21135 15524 21180 15552
rect 21174 15512 21180 15524
rect 21232 15512 21238 15564
rect 20901 15487 20959 15493
rect 20901 15453 20913 15487
rect 20947 15484 20959 15487
rect 21266 15484 21272 15496
rect 20947 15456 21272 15484
rect 20947 15453 20959 15456
rect 20901 15447 20959 15453
rect 21266 15444 21272 15456
rect 21324 15484 21330 15496
rect 22002 15484 22008 15496
rect 21324 15456 22008 15484
rect 21324 15444 21330 15456
rect 22002 15444 22008 15456
rect 22060 15444 22066 15496
rect 1578 15348 1584 15360
rect 1539 15320 1584 15348
rect 1578 15308 1584 15320
rect 1636 15308 1642 15360
rect 15838 15308 15844 15360
rect 15896 15348 15902 15360
rect 16025 15351 16083 15357
rect 16025 15348 16037 15351
rect 15896 15320 16037 15348
rect 15896 15308 15902 15320
rect 16025 15317 16037 15320
rect 16071 15317 16083 15351
rect 22462 15348 22468 15360
rect 22423 15320 22468 15348
rect 16025 15311 16083 15317
rect 22462 15308 22468 15320
rect 22520 15308 22526 15360
rect 1104 15258 38824 15280
rect 1104 15206 4246 15258
rect 4298 15206 4310 15258
rect 4362 15206 4374 15258
rect 4426 15206 4438 15258
rect 4490 15206 34966 15258
rect 35018 15206 35030 15258
rect 35082 15206 35094 15258
rect 35146 15206 35158 15258
rect 35210 15206 38824 15258
rect 1104 15184 38824 15206
rect 15194 15104 15200 15156
rect 15252 15144 15258 15156
rect 15841 15147 15899 15153
rect 15841 15144 15853 15147
rect 15252 15116 15853 15144
rect 15252 15104 15258 15116
rect 15841 15113 15853 15116
rect 15887 15144 15899 15147
rect 16850 15144 16856 15156
rect 15887 15116 16856 15144
rect 15887 15113 15899 15116
rect 15841 15107 15899 15113
rect 16850 15104 16856 15116
rect 16908 15104 16914 15156
rect 18322 15144 18328 15156
rect 18283 15116 18328 15144
rect 18322 15104 18328 15116
rect 18380 15104 18386 15156
rect 20993 15147 21051 15153
rect 20993 15113 21005 15147
rect 21039 15144 21051 15147
rect 21174 15144 21180 15156
rect 21039 15116 21180 15144
rect 21039 15113 21051 15116
rect 20993 15107 21051 15113
rect 21174 15104 21180 15116
rect 21232 15104 21238 15156
rect 16022 15036 16028 15088
rect 16080 15076 16086 15088
rect 16301 15079 16359 15085
rect 16301 15076 16313 15079
rect 16080 15048 16313 15076
rect 16080 15036 16086 15048
rect 16301 15045 16313 15048
rect 16347 15045 16359 15079
rect 18598 15076 18604 15088
rect 16301 15039 16359 15045
rect 17788 15048 18604 15076
rect 13354 14968 13360 15020
rect 13412 15008 13418 15020
rect 13541 15011 13599 15017
rect 13541 15008 13553 15011
rect 13412 14980 13553 15008
rect 13412 14968 13418 14980
rect 13541 14977 13553 14980
rect 13587 14977 13599 15011
rect 13814 15008 13820 15020
rect 13775 14980 13820 15008
rect 13541 14971 13599 14977
rect 13814 14968 13820 14980
rect 13872 14968 13878 15020
rect 15286 14968 15292 15020
rect 15344 15008 15350 15020
rect 17788 15017 17816 15048
rect 18598 15036 18604 15048
rect 18656 15076 18662 15088
rect 18656 15048 19196 15076
rect 18656 15036 18662 15048
rect 17773 15011 17831 15017
rect 17773 15008 17785 15011
rect 15344 14980 17785 15008
rect 15344 14968 15350 14980
rect 17773 14977 17785 14980
rect 17819 14977 17831 15011
rect 17773 14971 17831 14977
rect 17954 14968 17960 15020
rect 18012 15008 18018 15020
rect 18012 14980 19104 15008
rect 18012 14968 18018 14980
rect 13449 14943 13507 14949
rect 13449 14909 13461 14943
rect 13495 14940 13507 14943
rect 13832 14940 13860 14968
rect 15473 14943 15531 14949
rect 15473 14940 15485 14943
rect 13495 14912 15485 14940
rect 13495 14909 13507 14912
rect 13449 14903 13507 14909
rect 15473 14909 15485 14912
rect 15519 14909 15531 14943
rect 15473 14903 15531 14909
rect 15194 14872 15200 14884
rect 15155 14844 15200 14872
rect 15194 14832 15200 14844
rect 15252 14832 15258 14884
rect 15488 14872 15516 14903
rect 15838 14900 15844 14952
rect 15896 14940 15902 14952
rect 16485 14943 16543 14949
rect 16485 14940 16497 14943
rect 15896 14912 16497 14940
rect 15896 14900 15902 14912
rect 16485 14909 16497 14912
rect 16531 14909 16543 14943
rect 16669 14943 16727 14949
rect 16669 14940 16681 14943
rect 16485 14903 16543 14909
rect 16592 14912 16681 14940
rect 15488 14844 15976 14872
rect 15948 14804 15976 14844
rect 16592 14804 16620 14912
rect 16669 14909 16681 14912
rect 16715 14909 16727 14943
rect 16850 14940 16856 14952
rect 16811 14912 16856 14940
rect 16669 14903 16727 14909
rect 16850 14900 16856 14912
rect 16908 14900 16914 14952
rect 18046 14900 18052 14952
rect 18104 14940 18110 14952
rect 19076 14949 19104 14980
rect 19168 14949 19196 15048
rect 18509 14943 18567 14949
rect 18509 14940 18521 14943
rect 18104 14912 18521 14940
rect 18104 14900 18110 14912
rect 18509 14909 18521 14912
rect 18555 14909 18567 14943
rect 18509 14903 18567 14909
rect 18693 14943 18751 14949
rect 18693 14909 18705 14943
rect 18739 14909 18751 14943
rect 18693 14903 18751 14909
rect 19061 14943 19119 14949
rect 19061 14909 19073 14943
rect 19107 14909 19119 14943
rect 19061 14903 19119 14909
rect 19153 14943 19211 14949
rect 19153 14909 19165 14943
rect 19199 14909 19211 14943
rect 19153 14903 19211 14909
rect 17497 14875 17555 14881
rect 17497 14841 17509 14875
rect 17543 14872 17555 14875
rect 18708 14872 18736 14903
rect 18966 14872 18972 14884
rect 17543 14844 18972 14872
rect 17543 14841 17555 14844
rect 17497 14835 17555 14841
rect 18966 14832 18972 14844
rect 19024 14832 19030 14884
rect 21266 14804 21272 14816
rect 15948 14776 16620 14804
rect 21227 14776 21272 14804
rect 21266 14764 21272 14776
rect 21324 14764 21330 14816
rect 1104 14714 38824 14736
rect 1104 14662 19606 14714
rect 19658 14662 19670 14714
rect 19722 14662 19734 14714
rect 19786 14662 19798 14714
rect 19850 14662 38824 14714
rect 1104 14640 38824 14662
rect 11425 14603 11483 14609
rect 11425 14569 11437 14603
rect 11471 14600 11483 14603
rect 13354 14600 13360 14612
rect 11471 14572 13360 14600
rect 11471 14569 11483 14572
rect 11425 14563 11483 14569
rect 13354 14560 13360 14572
rect 13412 14600 13418 14612
rect 13541 14603 13599 14609
rect 13541 14600 13553 14603
rect 13412 14572 13553 14600
rect 13412 14560 13418 14572
rect 13541 14569 13553 14572
rect 13587 14569 13599 14603
rect 18966 14600 18972 14612
rect 18927 14572 18972 14600
rect 13541 14563 13599 14569
rect 18966 14560 18972 14572
rect 19024 14560 19030 14612
rect 15838 14532 15844 14544
rect 15799 14504 15844 14532
rect 15838 14492 15844 14504
rect 15896 14492 15902 14544
rect 11054 14424 11060 14476
rect 11112 14464 11118 14476
rect 11514 14464 11520 14476
rect 11112 14436 11520 14464
rect 11112 14424 11118 14436
rect 11514 14424 11520 14436
rect 11572 14464 11578 14476
rect 11609 14467 11667 14473
rect 11609 14464 11621 14467
rect 11572 14436 11621 14464
rect 11572 14424 11578 14436
rect 11609 14433 11621 14436
rect 11655 14433 11667 14467
rect 11609 14427 11667 14433
rect 15194 14424 15200 14476
rect 15252 14464 15258 14476
rect 15381 14467 15439 14473
rect 15381 14464 15393 14467
rect 15252 14436 15393 14464
rect 15252 14424 15258 14436
rect 15381 14433 15393 14436
rect 15427 14433 15439 14467
rect 15381 14427 15439 14433
rect 17865 14467 17923 14473
rect 17865 14433 17877 14467
rect 17911 14464 17923 14467
rect 17954 14464 17960 14476
rect 17911 14436 17960 14464
rect 17911 14433 17923 14436
rect 17865 14427 17923 14433
rect 17954 14424 17960 14436
rect 18012 14424 18018 14476
rect 23290 14464 23296 14476
rect 23251 14436 23296 14464
rect 23290 14424 23296 14436
rect 23348 14424 23354 14476
rect 15286 14396 15292 14408
rect 15247 14368 15292 14396
rect 15286 14356 15292 14368
rect 15344 14356 15350 14408
rect 17494 14356 17500 14408
rect 17552 14396 17558 14408
rect 17589 14399 17647 14405
rect 17589 14396 17601 14399
rect 17552 14368 17601 14396
rect 17552 14356 17558 14368
rect 17589 14365 17601 14368
rect 17635 14396 17647 14399
rect 18322 14396 18328 14408
rect 17635 14368 18328 14396
rect 17635 14365 17647 14368
rect 17589 14359 17647 14365
rect 18322 14356 18328 14368
rect 18380 14356 18386 14408
rect 22094 14220 22100 14272
rect 22152 14260 22158 14272
rect 23106 14260 23112 14272
rect 22152 14232 23112 14260
rect 22152 14220 22158 14232
rect 23106 14220 23112 14232
rect 23164 14220 23170 14272
rect 1104 14170 38824 14192
rect 1104 14118 4246 14170
rect 4298 14118 4310 14170
rect 4362 14118 4374 14170
rect 4426 14118 4438 14170
rect 4490 14118 34966 14170
rect 35018 14118 35030 14170
rect 35082 14118 35094 14170
rect 35146 14118 35158 14170
rect 35210 14118 38824 14170
rect 1104 14096 38824 14118
rect 11514 14056 11520 14068
rect 11475 14028 11520 14056
rect 11514 14016 11520 14028
rect 11572 14016 11578 14068
rect 15194 14016 15200 14068
rect 15252 14056 15258 14068
rect 15657 14059 15715 14065
rect 15657 14056 15669 14059
rect 15252 14028 15669 14056
rect 15252 14016 15258 14028
rect 15657 14025 15669 14028
rect 15703 14025 15715 14059
rect 15657 14019 15715 14025
rect 17681 14059 17739 14065
rect 17681 14025 17693 14059
rect 17727 14056 17739 14059
rect 17954 14056 17960 14068
rect 17727 14028 17960 14056
rect 17727 14025 17739 14028
rect 17681 14019 17739 14025
rect 17954 14016 17960 14028
rect 18012 14016 18018 14068
rect 18322 14056 18328 14068
rect 18283 14028 18328 14056
rect 18322 14016 18328 14028
rect 18380 14016 18386 14068
rect 23201 14059 23259 14065
rect 23201 14025 23213 14059
rect 23247 14056 23259 14059
rect 23290 14056 23296 14068
rect 23247 14028 23296 14056
rect 23247 14025 23259 14028
rect 23201 14019 23259 14025
rect 23290 14016 23296 14028
rect 23348 14016 23354 14068
rect 15286 13988 15292 14000
rect 15247 13960 15292 13988
rect 15286 13948 15292 13960
rect 15344 13948 15350 14000
rect 24946 13988 24952 14000
rect 24907 13960 24952 13988
rect 24946 13948 24952 13960
rect 25004 13948 25010 14000
rect 25130 13852 25136 13864
rect 25091 13824 25136 13852
rect 25130 13812 25136 13824
rect 25188 13852 25194 13864
rect 25409 13855 25467 13861
rect 25409 13852 25421 13855
rect 25188 13824 25421 13852
rect 25188 13812 25194 13824
rect 25409 13821 25421 13824
rect 25455 13821 25467 13855
rect 25409 13815 25467 13821
rect 1104 13626 38824 13648
rect 1104 13574 19606 13626
rect 19658 13574 19670 13626
rect 19722 13574 19734 13626
rect 19786 13574 19798 13626
rect 19850 13574 38824 13626
rect 1104 13552 38824 13574
rect 13354 13472 13360 13524
rect 13412 13512 13418 13524
rect 13633 13515 13691 13521
rect 13633 13512 13645 13515
rect 13412 13484 13645 13512
rect 13412 13472 13418 13484
rect 13633 13481 13645 13484
rect 13679 13481 13691 13515
rect 13633 13475 13691 13481
rect 21266 13472 21272 13524
rect 21324 13512 21330 13524
rect 21821 13515 21879 13521
rect 21821 13512 21833 13515
rect 21324 13484 21833 13512
rect 21324 13472 21330 13484
rect 21821 13481 21833 13484
rect 21867 13481 21879 13515
rect 21821 13475 21879 13481
rect 17862 13444 17868 13456
rect 16776 13416 17868 13444
rect 16776 13388 16804 13416
rect 17862 13404 17868 13416
rect 17920 13404 17926 13456
rect 16758 13376 16764 13388
rect 16671 13348 16764 13376
rect 16758 13336 16764 13348
rect 16816 13336 16822 13388
rect 16942 13376 16948 13388
rect 16903 13348 16948 13376
rect 16942 13336 16948 13348
rect 17000 13336 17006 13388
rect 17310 13376 17316 13388
rect 17271 13348 17316 13376
rect 17310 13336 17316 13348
rect 17368 13336 17374 13388
rect 21910 13336 21916 13388
rect 21968 13376 21974 13388
rect 22005 13379 22063 13385
rect 22005 13376 22017 13379
rect 21968 13348 22017 13376
rect 21968 13336 21974 13348
rect 22005 13345 22017 13348
rect 22051 13345 22063 13379
rect 22005 13339 22063 13345
rect 16482 13308 16488 13320
rect 16443 13280 16488 13308
rect 16482 13268 16488 13280
rect 16540 13268 16546 13320
rect 16574 13268 16580 13320
rect 16632 13308 16638 13320
rect 17221 13311 17279 13317
rect 17221 13308 17233 13311
rect 16632 13280 17233 13308
rect 16632 13268 16638 13280
rect 17221 13277 17233 13280
rect 17267 13277 17279 13311
rect 17221 13271 17279 13277
rect 1104 13082 38824 13104
rect 1104 13030 4246 13082
rect 4298 13030 4310 13082
rect 4362 13030 4374 13082
rect 4426 13030 4438 13082
rect 4490 13030 34966 13082
rect 35018 13030 35030 13082
rect 35082 13030 35094 13082
rect 35146 13030 35158 13082
rect 35210 13030 38824 13082
rect 1104 13008 38824 13030
rect 15010 12928 15016 12980
rect 15068 12968 15074 12980
rect 16393 12971 16451 12977
rect 16393 12968 16405 12971
rect 15068 12940 16405 12968
rect 15068 12928 15074 12940
rect 16393 12937 16405 12940
rect 16439 12968 16451 12971
rect 16574 12968 16580 12980
rect 16439 12940 16580 12968
rect 16439 12937 16451 12940
rect 16393 12931 16451 12937
rect 16574 12928 16580 12940
rect 16632 12928 16638 12980
rect 16942 12928 16948 12980
rect 17000 12968 17006 12980
rect 17037 12971 17095 12977
rect 17037 12968 17049 12971
rect 17000 12940 17049 12968
rect 17000 12928 17006 12940
rect 17037 12937 17049 12940
rect 17083 12968 17095 12971
rect 17126 12968 17132 12980
rect 17083 12940 17132 12968
rect 17083 12937 17095 12940
rect 17037 12931 17095 12937
rect 17126 12928 17132 12940
rect 17184 12928 17190 12980
rect 21910 12968 21916 12980
rect 21871 12940 21916 12968
rect 21910 12928 21916 12940
rect 21968 12928 21974 12980
rect 15930 12860 15936 12912
rect 15988 12900 15994 12912
rect 16025 12903 16083 12909
rect 16025 12900 16037 12903
rect 15988 12872 16037 12900
rect 15988 12860 15994 12872
rect 16025 12869 16037 12872
rect 16071 12900 16083 12903
rect 17310 12900 17316 12912
rect 16071 12872 17316 12900
rect 16071 12869 16083 12872
rect 16025 12863 16083 12869
rect 17310 12860 17316 12872
rect 17368 12860 17374 12912
rect 13541 12835 13599 12841
rect 13541 12801 13553 12835
rect 13587 12832 13599 12835
rect 13906 12832 13912 12844
rect 13587 12804 13912 12832
rect 13587 12801 13599 12804
rect 13541 12795 13599 12801
rect 13906 12792 13912 12804
rect 13964 12832 13970 12844
rect 14918 12832 14924 12844
rect 13964 12804 14924 12832
rect 13964 12792 13970 12804
rect 14918 12792 14924 12804
rect 14976 12792 14982 12844
rect 16758 12832 16764 12844
rect 16719 12804 16764 12832
rect 16758 12792 16764 12804
rect 16816 12792 16822 12844
rect 12434 12724 12440 12776
rect 12492 12764 12498 12776
rect 13354 12764 13360 12776
rect 12492 12736 13360 12764
rect 12492 12724 12498 12736
rect 13354 12724 13360 12736
rect 13412 12764 13418 12776
rect 13633 12767 13691 12773
rect 13633 12764 13645 12767
rect 13412 12736 13645 12764
rect 13412 12724 13418 12736
rect 13633 12733 13645 12736
rect 13679 12764 13691 12767
rect 14734 12764 14740 12776
rect 13679 12736 14740 12764
rect 13679 12733 13691 12736
rect 13633 12727 13691 12733
rect 14734 12724 14740 12736
rect 14792 12724 14798 12776
rect 15102 12588 15108 12640
rect 15160 12628 15166 12640
rect 15197 12631 15255 12637
rect 15197 12628 15209 12631
rect 15160 12600 15209 12628
rect 15160 12588 15166 12600
rect 15197 12597 15209 12600
rect 15243 12597 15255 12631
rect 15197 12591 15255 12597
rect 30282 12588 30288 12640
rect 30340 12628 30346 12640
rect 30466 12628 30472 12640
rect 30340 12600 30472 12628
rect 30340 12588 30346 12600
rect 30466 12588 30472 12600
rect 30524 12588 30530 12640
rect 1104 12538 38824 12560
rect 1104 12486 19606 12538
rect 19658 12486 19670 12538
rect 19722 12486 19734 12538
rect 19786 12486 19798 12538
rect 19850 12486 38824 12538
rect 1104 12464 38824 12486
rect 17126 12384 17132 12436
rect 17184 12424 17190 12436
rect 17497 12427 17555 12433
rect 17497 12424 17509 12427
rect 17184 12396 17509 12424
rect 17184 12384 17190 12396
rect 17497 12393 17509 12396
rect 17543 12393 17555 12427
rect 17497 12387 17555 12393
rect 34698 12384 34704 12436
rect 34756 12424 34762 12436
rect 35342 12424 35348 12436
rect 34756 12396 35348 12424
rect 34756 12384 34762 12396
rect 35342 12384 35348 12396
rect 35400 12384 35406 12436
rect 13170 12356 13176 12368
rect 13131 12328 13176 12356
rect 13170 12316 13176 12328
rect 13228 12316 13234 12368
rect 13998 12356 14004 12368
rect 13832 12328 14004 12356
rect 13633 12291 13691 12297
rect 13633 12257 13645 12291
rect 13679 12288 13691 12291
rect 13722 12288 13728 12300
rect 13679 12260 13728 12288
rect 13679 12257 13691 12260
rect 13633 12251 13691 12257
rect 13722 12248 13728 12260
rect 13780 12248 13786 12300
rect 13832 12297 13860 12328
rect 13998 12316 14004 12328
rect 14056 12356 14062 12368
rect 15102 12356 15108 12368
rect 14056 12328 15108 12356
rect 14056 12316 14062 12328
rect 15102 12316 15108 12328
rect 15160 12316 15166 12368
rect 18414 12316 18420 12368
rect 18472 12356 18478 12368
rect 18472 12328 19656 12356
rect 18472 12316 18478 12328
rect 13817 12291 13875 12297
rect 13817 12257 13829 12291
rect 13863 12257 13875 12291
rect 13817 12251 13875 12257
rect 13906 12248 13912 12300
rect 13964 12288 13970 12300
rect 14185 12291 14243 12297
rect 14185 12288 14197 12291
rect 13964 12260 14197 12288
rect 13964 12248 13970 12260
rect 14185 12257 14197 12260
rect 14231 12257 14243 12291
rect 14185 12251 14243 12257
rect 14369 12291 14427 12297
rect 14369 12257 14381 12291
rect 14415 12288 14427 12291
rect 15010 12288 15016 12300
rect 14415 12260 15016 12288
rect 14415 12257 14427 12260
rect 14369 12251 14427 12257
rect 12710 12180 12716 12232
rect 12768 12220 12774 12232
rect 13354 12220 13360 12232
rect 12768 12192 13360 12220
rect 12768 12180 12774 12192
rect 13354 12180 13360 12192
rect 13412 12220 13418 12232
rect 14384 12220 14412 12251
rect 15010 12248 15016 12260
rect 15068 12248 15074 12300
rect 16117 12291 16175 12297
rect 16117 12257 16129 12291
rect 16163 12288 16175 12291
rect 17494 12288 17500 12300
rect 16163 12260 17500 12288
rect 16163 12257 16175 12260
rect 16117 12251 16175 12257
rect 17494 12248 17500 12260
rect 17552 12248 17558 12300
rect 19242 12288 19248 12300
rect 19203 12260 19248 12288
rect 19242 12248 19248 12260
rect 19300 12248 19306 12300
rect 19628 12297 19656 12328
rect 19613 12291 19671 12297
rect 19613 12257 19625 12291
rect 19659 12257 19671 12291
rect 19613 12251 19671 12257
rect 16390 12220 16396 12232
rect 13412 12192 14412 12220
rect 16351 12192 16396 12220
rect 13412 12180 13418 12192
rect 16390 12180 16396 12192
rect 16448 12180 16454 12232
rect 18046 12180 18052 12232
rect 18104 12220 18110 12232
rect 18322 12220 18328 12232
rect 18104 12192 18328 12220
rect 18104 12180 18110 12192
rect 18322 12180 18328 12192
rect 18380 12220 18386 12232
rect 19061 12223 19119 12229
rect 19061 12220 19073 12223
rect 18380 12192 19073 12220
rect 18380 12180 18386 12192
rect 19061 12189 19073 12192
rect 19107 12189 19119 12223
rect 19061 12183 19119 12189
rect 19521 12223 19579 12229
rect 19521 12189 19533 12223
rect 19567 12189 19579 12223
rect 19521 12183 19579 12189
rect 18598 12112 18604 12164
rect 18656 12152 18662 12164
rect 19536 12152 19564 12183
rect 18656 12124 19564 12152
rect 18656 12112 18662 12124
rect 15286 12044 15292 12096
rect 15344 12084 15350 12096
rect 15473 12087 15531 12093
rect 15473 12084 15485 12087
rect 15344 12056 15485 12084
rect 15344 12044 15350 12056
rect 15473 12053 15485 12056
rect 15519 12084 15531 12087
rect 15746 12084 15752 12096
rect 15519 12056 15752 12084
rect 15519 12053 15531 12056
rect 15473 12047 15531 12053
rect 15746 12044 15752 12056
rect 15804 12044 15810 12096
rect 17862 12044 17868 12096
rect 17920 12084 17926 12096
rect 18414 12084 18420 12096
rect 17920 12056 18420 12084
rect 17920 12044 17926 12056
rect 18414 12044 18420 12056
rect 18472 12044 18478 12096
rect 18874 12084 18880 12096
rect 18835 12056 18880 12084
rect 18874 12044 18880 12056
rect 18932 12044 18938 12096
rect 1104 11994 38824 12016
rect 1104 11942 4246 11994
rect 4298 11942 4310 11994
rect 4362 11942 4374 11994
rect 4426 11942 4438 11994
rect 4490 11942 34966 11994
rect 35018 11942 35030 11994
rect 35082 11942 35094 11994
rect 35146 11942 35158 11994
rect 35210 11942 38824 11994
rect 1104 11920 38824 11942
rect 13265 11883 13323 11889
rect 13265 11849 13277 11883
rect 13311 11880 13323 11883
rect 13354 11880 13360 11892
rect 13311 11852 13360 11880
rect 13311 11849 13323 11852
rect 13265 11843 13323 11849
rect 13354 11840 13360 11852
rect 13412 11840 13418 11892
rect 13998 11880 14004 11892
rect 13959 11852 14004 11880
rect 13998 11840 14004 11852
rect 14056 11840 14062 11892
rect 14734 11840 14740 11892
rect 14792 11880 14798 11892
rect 14921 11883 14979 11889
rect 14921 11880 14933 11883
rect 14792 11852 14933 11880
rect 14792 11840 14798 11852
rect 14921 11849 14933 11852
rect 14967 11849 14979 11883
rect 14921 11843 14979 11849
rect 15381 11883 15439 11889
rect 15381 11849 15393 11883
rect 15427 11880 15439 11883
rect 15930 11880 15936 11892
rect 15427 11852 15936 11880
rect 15427 11849 15439 11852
rect 15381 11843 15439 11849
rect 12897 11815 12955 11821
rect 12897 11781 12909 11815
rect 12943 11812 12955 11815
rect 13906 11812 13912 11824
rect 12943 11784 13912 11812
rect 12943 11781 12955 11784
rect 12897 11775 12955 11781
rect 13906 11772 13912 11784
rect 13964 11772 13970 11824
rect 14936 11744 14964 11843
rect 15930 11840 15936 11852
rect 15988 11880 15994 11892
rect 16390 11880 16396 11892
rect 15988 11852 16396 11880
rect 15988 11840 15994 11852
rect 16390 11840 16396 11852
rect 16448 11840 16454 11892
rect 17494 11880 17500 11892
rect 17455 11852 17500 11880
rect 17494 11840 17500 11852
rect 17552 11840 17558 11892
rect 18322 11880 18328 11892
rect 18283 11852 18328 11880
rect 18322 11840 18328 11852
rect 18380 11840 18386 11892
rect 20993 11883 21051 11889
rect 20993 11849 21005 11883
rect 21039 11880 21051 11883
rect 21542 11880 21548 11892
rect 21039 11852 21548 11880
rect 21039 11849 21051 11852
rect 20993 11843 21051 11849
rect 21542 11840 21548 11852
rect 21600 11840 21606 11892
rect 15473 11747 15531 11753
rect 15473 11744 15485 11747
rect 14936 11716 15485 11744
rect 15473 11713 15485 11716
rect 15519 11713 15531 11747
rect 15473 11707 15531 11713
rect 19337 11747 19395 11753
rect 19337 11713 19349 11747
rect 19383 11744 19395 11747
rect 19383 11716 19748 11744
rect 19383 11713 19395 11716
rect 19337 11707 19395 11713
rect 15286 11636 15292 11688
rect 15344 11676 15350 11688
rect 15749 11679 15807 11685
rect 15749 11676 15761 11679
rect 15344 11648 15761 11676
rect 15344 11636 15350 11648
rect 15749 11645 15761 11648
rect 15795 11645 15807 11679
rect 19426 11676 19432 11688
rect 19387 11648 19432 11676
rect 15749 11639 15807 11645
rect 19426 11636 19432 11648
rect 19484 11636 19490 11688
rect 19720 11685 19748 11716
rect 19705 11679 19763 11685
rect 19705 11645 19717 11679
rect 19751 11676 19763 11679
rect 19978 11676 19984 11688
rect 19751 11648 19984 11676
rect 19751 11645 19763 11648
rect 19705 11639 19763 11645
rect 19978 11636 19984 11648
rect 20036 11636 20042 11688
rect 17865 11611 17923 11617
rect 17865 11577 17877 11611
rect 17911 11608 17923 11611
rect 19242 11608 19248 11620
rect 17911 11580 19248 11608
rect 17911 11577 17923 11580
rect 17865 11571 17923 11577
rect 19242 11568 19248 11580
rect 19300 11568 19306 11620
rect 13633 11543 13691 11549
rect 13633 11509 13645 11543
rect 13679 11540 13691 11543
rect 13722 11540 13728 11552
rect 13679 11512 13728 11540
rect 13679 11509 13691 11512
rect 13633 11503 13691 11509
rect 13722 11500 13728 11512
rect 13780 11500 13786 11552
rect 16206 11500 16212 11552
rect 16264 11540 16270 11552
rect 16853 11543 16911 11549
rect 16853 11540 16865 11543
rect 16264 11512 16865 11540
rect 16264 11500 16270 11512
rect 16853 11509 16865 11512
rect 16899 11509 16911 11543
rect 18598 11540 18604 11552
rect 18559 11512 18604 11540
rect 16853 11503 16911 11509
rect 18598 11500 18604 11512
rect 18656 11500 18662 11552
rect 1104 11450 38824 11472
rect 1104 11398 19606 11450
rect 19658 11398 19670 11450
rect 19722 11398 19734 11450
rect 19786 11398 19798 11450
rect 19850 11398 38824 11450
rect 1104 11376 38824 11398
rect 15286 11228 15292 11280
rect 15344 11268 15350 11280
rect 19242 11268 19248 11280
rect 15344 11240 16620 11268
rect 19203 11240 19248 11268
rect 15344 11228 15350 11240
rect 16206 11200 16212 11212
rect 16167 11172 16212 11200
rect 16206 11160 16212 11172
rect 16264 11160 16270 11212
rect 16592 11209 16620 11240
rect 19242 11228 19248 11240
rect 19300 11228 19306 11280
rect 16577 11203 16635 11209
rect 16577 11169 16589 11203
rect 16623 11169 16635 11203
rect 18598 11200 18604 11212
rect 16577 11163 16635 11169
rect 17236 11172 18604 11200
rect 13722 11092 13728 11144
rect 13780 11132 13786 11144
rect 16301 11135 16359 11141
rect 16301 11132 16313 11135
rect 13780 11104 16313 11132
rect 13780 11092 13786 11104
rect 16301 11101 16313 11104
rect 16347 11132 16359 11135
rect 16390 11132 16396 11144
rect 16347 11104 16396 11132
rect 16347 11101 16359 11104
rect 16301 11095 16359 11101
rect 16390 11092 16396 11104
rect 16448 11092 16454 11144
rect 16482 11092 16488 11144
rect 16540 11132 16546 11144
rect 17236 11132 17264 11172
rect 18598 11160 18604 11172
rect 18656 11160 18662 11212
rect 16540 11104 17264 11132
rect 16540 11092 16546 11104
rect 17494 11092 17500 11144
rect 17552 11132 17558 11144
rect 17589 11135 17647 11141
rect 17589 11132 17601 11135
rect 17552 11104 17601 11132
rect 17552 11092 17558 11104
rect 17589 11101 17601 11104
rect 17635 11101 17647 11135
rect 17862 11132 17868 11144
rect 17823 11104 17868 11132
rect 17589 11095 17647 11101
rect 17862 11092 17868 11104
rect 17920 11092 17926 11144
rect 15838 11064 15844 11076
rect 15799 11036 15844 11064
rect 15838 11024 15844 11036
rect 15896 11024 15902 11076
rect 18598 11024 18604 11076
rect 18656 11064 18662 11076
rect 19426 11064 19432 11076
rect 18656 11036 19432 11064
rect 18656 11024 18662 11036
rect 19426 11024 19432 11036
rect 19484 11064 19490 11076
rect 19521 11067 19579 11073
rect 19521 11064 19533 11067
rect 19484 11036 19533 11064
rect 19484 11024 19490 11036
rect 19521 11033 19533 11036
rect 19567 11033 19579 11067
rect 19521 11027 19579 11033
rect 1104 10906 38824 10928
rect 1104 10854 4246 10906
rect 4298 10854 4310 10906
rect 4362 10854 4374 10906
rect 4426 10854 4438 10906
rect 4490 10854 34966 10906
rect 35018 10854 35030 10906
rect 35082 10854 35094 10906
rect 35146 10854 35158 10906
rect 35210 10854 38824 10906
rect 1104 10832 38824 10854
rect 15286 10792 15292 10804
rect 15247 10764 15292 10792
rect 15286 10752 15292 10764
rect 15344 10752 15350 10804
rect 16206 10752 16212 10804
rect 16264 10792 16270 10804
rect 16301 10795 16359 10801
rect 16301 10792 16313 10795
rect 16264 10764 16313 10792
rect 16264 10752 16270 10764
rect 16301 10761 16313 10764
rect 16347 10761 16359 10795
rect 16301 10755 16359 10761
rect 17681 10795 17739 10801
rect 17681 10761 17693 10795
rect 17727 10792 17739 10795
rect 17862 10792 17868 10804
rect 17727 10764 17868 10792
rect 17727 10761 17739 10764
rect 17681 10755 17739 10761
rect 17862 10752 17868 10764
rect 17920 10752 17926 10804
rect 16025 10727 16083 10733
rect 16025 10693 16037 10727
rect 16071 10724 16083 10727
rect 16390 10724 16396 10736
rect 16071 10696 16396 10724
rect 16071 10693 16083 10696
rect 16025 10687 16083 10693
rect 16390 10684 16396 10696
rect 16448 10684 16454 10736
rect 17494 10684 17500 10736
rect 17552 10724 17558 10736
rect 18230 10724 18236 10736
rect 17552 10696 18236 10724
rect 17552 10684 17558 10696
rect 18230 10684 18236 10696
rect 18288 10724 18294 10736
rect 18598 10724 18604 10736
rect 18288 10696 18604 10724
rect 18288 10684 18294 10696
rect 18598 10684 18604 10696
rect 18656 10684 18662 10736
rect 15657 10659 15715 10665
rect 15657 10625 15669 10659
rect 15703 10656 15715 10659
rect 16482 10656 16488 10668
rect 15703 10628 16488 10656
rect 15703 10625 15715 10628
rect 15657 10619 15715 10625
rect 16482 10616 16488 10628
rect 16540 10616 16546 10668
rect 1104 10362 38824 10384
rect 1104 10310 19606 10362
rect 19658 10310 19670 10362
rect 19722 10310 19734 10362
rect 19786 10310 19798 10362
rect 19850 10310 38824 10362
rect 1104 10288 38824 10310
rect 8757 10183 8815 10189
rect 8757 10149 8769 10183
rect 8803 10180 8815 10183
rect 9398 10180 9404 10192
rect 8803 10152 9404 10180
rect 8803 10149 8815 10152
rect 8757 10143 8815 10149
rect 9398 10140 9404 10152
rect 9456 10140 9462 10192
rect 1578 10072 1584 10124
rect 1636 10112 1642 10124
rect 1765 10115 1823 10121
rect 1765 10112 1777 10115
rect 1636 10084 1777 10112
rect 1636 10072 1642 10084
rect 1765 10081 1777 10084
rect 1811 10081 1823 10115
rect 1765 10075 1823 10081
rect 2038 10072 2044 10124
rect 2096 10072 2102 10124
rect 7098 10112 7104 10124
rect 7059 10084 7104 10112
rect 7098 10072 7104 10084
rect 7156 10072 7162 10124
rect 7190 10072 7196 10124
rect 7248 10112 7254 10124
rect 7377 10115 7435 10121
rect 7377 10112 7389 10115
rect 7248 10084 7389 10112
rect 7248 10072 7254 10084
rect 7377 10081 7389 10084
rect 7423 10081 7435 10115
rect 7377 10075 7435 10081
rect 1394 10004 1400 10056
rect 1452 10044 1458 10056
rect 1489 10047 1547 10053
rect 1489 10044 1501 10047
rect 1452 10016 1501 10044
rect 1452 10004 1458 10016
rect 1489 10013 1501 10016
rect 1535 10044 1547 10047
rect 2056 10044 2084 10072
rect 3142 10044 3148 10056
rect 1535 10016 2084 10044
rect 3103 10016 3148 10044
rect 1535 10013 1547 10016
rect 1489 10007 1547 10013
rect 3142 10004 3148 10016
rect 3200 10004 3206 10056
rect 1104 9818 38824 9840
rect 1104 9766 4246 9818
rect 4298 9766 4310 9818
rect 4362 9766 4374 9818
rect 4426 9766 4438 9818
rect 4490 9766 34966 9818
rect 35018 9766 35030 9818
rect 35082 9766 35094 9818
rect 35146 9766 35158 9818
rect 35210 9766 38824 9818
rect 1104 9744 38824 9766
rect 2038 9704 2044 9716
rect 1999 9676 2044 9704
rect 2038 9664 2044 9676
rect 2096 9664 2102 9716
rect 7098 9664 7104 9716
rect 7156 9704 7162 9716
rect 7469 9707 7527 9713
rect 7469 9704 7481 9707
rect 7156 9676 7481 9704
rect 7156 9664 7162 9676
rect 7469 9673 7481 9676
rect 7515 9673 7527 9707
rect 7469 9667 7527 9673
rect 2866 9596 2872 9648
rect 2924 9636 2930 9648
rect 3326 9636 3332 9648
rect 2924 9608 3332 9636
rect 2924 9596 2930 9608
rect 3326 9596 3332 9608
rect 3384 9596 3390 9648
rect 1578 9364 1584 9376
rect 1539 9336 1584 9364
rect 1578 9324 1584 9336
rect 1636 9324 1642 9376
rect 7190 9364 7196 9376
rect 7151 9336 7196 9364
rect 7190 9324 7196 9336
rect 7248 9324 7254 9376
rect 1104 9274 38824 9296
rect 1104 9222 19606 9274
rect 19658 9222 19670 9274
rect 19722 9222 19734 9274
rect 19786 9222 19798 9274
rect 19850 9222 38824 9274
rect 1104 9200 38824 9222
rect 1104 8730 38824 8752
rect 1104 8678 4246 8730
rect 4298 8678 4310 8730
rect 4362 8678 4374 8730
rect 4426 8678 4438 8730
rect 4490 8678 34966 8730
rect 35018 8678 35030 8730
rect 35082 8678 35094 8730
rect 35146 8678 35158 8730
rect 35210 8678 38824 8730
rect 1104 8656 38824 8678
rect 1104 8186 38824 8208
rect 1104 8134 19606 8186
rect 19658 8134 19670 8186
rect 19722 8134 19734 8186
rect 19786 8134 19798 8186
rect 19850 8134 38824 8186
rect 1104 8112 38824 8134
rect 37458 7692 37464 7744
rect 37516 7732 37522 7744
rect 39574 7732 39580 7744
rect 37516 7704 39580 7732
rect 37516 7692 37522 7704
rect 39574 7692 39580 7704
rect 39632 7692 39638 7744
rect 1104 7642 38824 7664
rect 1104 7590 4246 7642
rect 4298 7590 4310 7642
rect 4362 7590 4374 7642
rect 4426 7590 4438 7642
rect 4490 7590 34966 7642
rect 35018 7590 35030 7642
rect 35082 7590 35094 7642
rect 35146 7590 35158 7642
rect 35210 7590 38824 7642
rect 1104 7568 38824 7590
rect 4614 7488 4620 7540
rect 4672 7528 4678 7540
rect 5074 7528 5080 7540
rect 4672 7500 5080 7528
rect 4672 7488 4678 7500
rect 5074 7488 5080 7500
rect 5132 7488 5138 7540
rect 37550 7488 37556 7540
rect 37608 7528 37614 7540
rect 39114 7528 39120 7540
rect 37608 7500 39120 7528
rect 37608 7488 37614 7500
rect 39114 7488 39120 7500
rect 39172 7488 39178 7540
rect 12342 7284 12348 7336
rect 12400 7324 12406 7336
rect 13446 7324 13452 7336
rect 12400 7296 13452 7324
rect 12400 7284 12406 7296
rect 13446 7284 13452 7296
rect 13504 7284 13510 7336
rect 1104 7098 38824 7120
rect 1104 7046 19606 7098
rect 19658 7046 19670 7098
rect 19722 7046 19734 7098
rect 19786 7046 19798 7098
rect 19850 7046 38824 7098
rect 1104 7024 38824 7046
rect 1104 6554 38824 6576
rect 1104 6502 4246 6554
rect 4298 6502 4310 6554
rect 4362 6502 4374 6554
rect 4426 6502 4438 6554
rect 4490 6502 34966 6554
rect 35018 6502 35030 6554
rect 35082 6502 35094 6554
rect 35146 6502 35158 6554
rect 35210 6502 38824 6554
rect 1104 6480 38824 6502
rect 35897 6307 35955 6313
rect 35897 6273 35909 6307
rect 35943 6304 35955 6307
rect 36262 6304 36268 6316
rect 35943 6276 36268 6304
rect 35943 6273 35955 6276
rect 35897 6267 35955 6273
rect 36262 6264 36268 6276
rect 36320 6264 36326 6316
rect 35986 6236 35992 6248
rect 35947 6208 35992 6236
rect 35986 6196 35992 6208
rect 36044 6196 36050 6248
rect 37366 6100 37372 6112
rect 37327 6072 37372 6100
rect 37366 6060 37372 6072
rect 37424 6060 37430 6112
rect 1104 6010 38824 6032
rect 1104 5958 19606 6010
rect 19658 5958 19670 6010
rect 19722 5958 19734 6010
rect 19786 5958 19798 6010
rect 19850 5958 38824 6010
rect 1104 5936 38824 5958
rect 35986 5692 35992 5704
rect 35947 5664 35992 5692
rect 35986 5652 35992 5664
rect 36044 5652 36050 5704
rect 1104 5466 38824 5488
rect 1104 5414 4246 5466
rect 4298 5414 4310 5466
rect 4362 5414 4374 5466
rect 4426 5414 4438 5466
rect 4490 5414 34966 5466
rect 35018 5414 35030 5466
rect 35082 5414 35094 5466
rect 35146 5414 35158 5466
rect 35210 5414 38824 5466
rect 1104 5392 38824 5414
rect 1104 4922 38824 4944
rect 1104 4870 19606 4922
rect 19658 4870 19670 4922
rect 19722 4870 19734 4922
rect 19786 4870 19798 4922
rect 19850 4870 38824 4922
rect 1104 4848 38824 4870
rect 13998 4808 14004 4820
rect 13959 4780 14004 4808
rect 13998 4768 14004 4780
rect 14056 4768 14062 4820
rect 21726 4768 21732 4820
rect 21784 4808 21790 4820
rect 22002 4808 22008 4820
rect 21784 4780 22008 4808
rect 21784 4768 21790 4780
rect 22002 4768 22008 4780
rect 22060 4768 22066 4820
rect 28994 4768 29000 4820
rect 29052 4808 29058 4820
rect 29362 4808 29368 4820
rect 29052 4780 29368 4808
rect 29052 4768 29058 4780
rect 29362 4768 29368 4780
rect 29420 4768 29426 4820
rect 33134 4768 33140 4820
rect 33192 4808 33198 4820
rect 33502 4808 33508 4820
rect 33192 4780 33508 4808
rect 33192 4768 33198 4780
rect 33502 4768 33508 4780
rect 33560 4768 33566 4820
rect 12434 4632 12440 4684
rect 12492 4672 12498 4684
rect 12492 4644 12537 4672
rect 12492 4632 12498 4644
rect 12710 4604 12716 4616
rect 12671 4576 12716 4604
rect 12710 4564 12716 4576
rect 12768 4564 12774 4616
rect 1104 4378 38824 4400
rect 1104 4326 4246 4378
rect 4298 4326 4310 4378
rect 4362 4326 4374 4378
rect 4426 4326 4438 4378
rect 4490 4326 34966 4378
rect 35018 4326 35030 4378
rect 35082 4326 35094 4378
rect 35146 4326 35158 4378
rect 35210 4326 38824 4378
rect 1104 4304 38824 4326
rect 12710 4264 12716 4276
rect 12671 4236 12716 4264
rect 12710 4224 12716 4236
rect 12768 4224 12774 4276
rect 12434 4156 12440 4208
rect 12492 4196 12498 4208
rect 12989 4199 13047 4205
rect 12989 4196 13001 4199
rect 12492 4168 13001 4196
rect 12492 4156 12498 4168
rect 12989 4165 13001 4168
rect 13035 4196 13047 4199
rect 13541 4199 13599 4205
rect 13541 4196 13553 4199
rect 13035 4168 13553 4196
rect 13035 4165 13047 4168
rect 12989 4159 13047 4165
rect 13541 4165 13553 4168
rect 13587 4165 13599 4199
rect 13541 4159 13599 4165
rect 6914 4088 6920 4140
rect 6972 4128 6978 4140
rect 8202 4128 8208 4140
rect 6972 4100 8208 4128
rect 6972 4088 6978 4100
rect 8202 4088 8208 4100
rect 8260 4088 8266 4140
rect 8386 4088 8392 4140
rect 8444 4128 8450 4140
rect 9214 4128 9220 4140
rect 8444 4100 9220 4128
rect 8444 4088 8450 4100
rect 9214 4088 9220 4100
rect 9272 4088 9278 4140
rect 10134 4088 10140 4140
rect 10192 4128 10198 4140
rect 10686 4128 10692 4140
rect 10192 4100 10692 4128
rect 10192 4088 10198 4100
rect 10686 4088 10692 4100
rect 10744 4088 10750 4140
rect 17954 4088 17960 4140
rect 18012 4128 18018 4140
rect 19150 4128 19156 4140
rect 18012 4100 19156 4128
rect 18012 4088 18018 4100
rect 19150 4088 19156 4100
rect 19208 4088 19214 4140
rect 19429 4131 19487 4137
rect 19429 4097 19441 4131
rect 19475 4128 19487 4131
rect 21177 4131 21235 4137
rect 19475 4100 19840 4128
rect 19475 4097 19487 4100
rect 19429 4091 19487 4097
rect 19812 4069 19840 4100
rect 21177 4097 21189 4131
rect 21223 4128 21235 4131
rect 21818 4128 21824 4140
rect 21223 4100 21824 4128
rect 21223 4097 21235 4100
rect 21177 4091 21235 4097
rect 21818 4088 21824 4100
rect 21876 4088 21882 4140
rect 19521 4063 19579 4069
rect 19521 4029 19533 4063
rect 19567 4029 19579 4063
rect 19521 4023 19579 4029
rect 19797 4063 19855 4069
rect 19797 4029 19809 4063
rect 19843 4060 19855 4063
rect 22738 4060 22744 4072
rect 19843 4032 22744 4060
rect 19843 4029 19855 4032
rect 19797 4023 19855 4029
rect 19426 3952 19432 4004
rect 19484 3992 19490 4004
rect 19536 3992 19564 4023
rect 22738 4020 22744 4032
rect 22796 4020 22802 4072
rect 19484 3964 19564 3992
rect 19484 3952 19490 3964
rect 11974 3884 11980 3936
rect 12032 3924 12038 3936
rect 12710 3924 12716 3936
rect 12032 3896 12716 3924
rect 12032 3884 12038 3896
rect 12710 3884 12716 3896
rect 12768 3884 12774 3936
rect 1104 3834 38824 3856
rect 1104 3782 19606 3834
rect 19658 3782 19670 3834
rect 19722 3782 19734 3834
rect 19786 3782 19798 3834
rect 19850 3782 38824 3834
rect 1104 3760 38824 3782
rect 14274 3720 14280 3732
rect 14235 3692 14280 3720
rect 14274 3680 14280 3692
rect 14332 3680 14338 3732
rect 12434 3544 12440 3596
rect 12492 3584 12498 3596
rect 12713 3587 12771 3593
rect 12713 3584 12725 3587
rect 12492 3556 12725 3584
rect 12492 3544 12498 3556
rect 12713 3553 12725 3556
rect 12759 3553 12771 3587
rect 12713 3547 12771 3553
rect 12802 3544 12808 3596
rect 12860 3584 12866 3596
rect 12989 3587 13047 3593
rect 12989 3584 13001 3587
rect 12860 3556 13001 3584
rect 12860 3544 12866 3556
rect 12989 3553 13001 3556
rect 13035 3553 13047 3587
rect 12989 3547 13047 3553
rect 14 3476 20 3528
rect 72 3516 78 3528
rect 1302 3516 1308 3528
rect 72 3488 1308 3516
rect 72 3476 78 3488
rect 1302 3476 1308 3488
rect 1360 3476 1366 3528
rect 19426 3340 19432 3392
rect 19484 3380 19490 3392
rect 19613 3383 19671 3389
rect 19613 3380 19625 3383
rect 19484 3352 19625 3380
rect 19484 3340 19490 3352
rect 19613 3349 19625 3352
rect 19659 3380 19671 3383
rect 20806 3380 20812 3392
rect 19659 3352 20812 3380
rect 19659 3349 19671 3352
rect 19613 3343 19671 3349
rect 20806 3340 20812 3352
rect 20864 3340 20870 3392
rect 1104 3290 38824 3312
rect 1104 3238 4246 3290
rect 4298 3238 4310 3290
rect 4362 3238 4374 3290
rect 4426 3238 4438 3290
rect 4490 3238 34966 3290
rect 35018 3238 35030 3290
rect 35082 3238 35094 3290
rect 35146 3238 35158 3290
rect 35210 3238 38824 3290
rect 1104 3216 38824 3238
rect 12253 3179 12311 3185
rect 12253 3145 12265 3179
rect 12299 3176 12311 3179
rect 12434 3176 12440 3188
rect 12299 3148 12440 3176
rect 12299 3145 12311 3148
rect 12253 3139 12311 3145
rect 12434 3136 12440 3148
rect 12492 3136 12498 3188
rect 14826 3136 14832 3188
rect 14884 3176 14890 3188
rect 14921 3179 14979 3185
rect 14921 3176 14933 3179
rect 14884 3148 14933 3176
rect 14884 3136 14890 3148
rect 14921 3145 14933 3148
rect 14967 3145 14979 3179
rect 14921 3139 14979 3145
rect 22281 3179 22339 3185
rect 22281 3145 22293 3179
rect 22327 3176 22339 3179
rect 22370 3176 22376 3188
rect 22327 3148 22376 3176
rect 22327 3145 22339 3148
rect 22281 3139 22339 3145
rect 22370 3136 22376 3148
rect 22428 3136 22434 3188
rect 12452 2972 12480 3136
rect 20714 3068 20720 3120
rect 20772 3068 20778 3120
rect 13449 3043 13507 3049
rect 13449 3009 13461 3043
rect 13495 3040 13507 3043
rect 13814 3040 13820 3052
rect 13495 3012 13820 3040
rect 13495 3009 13507 3012
rect 13449 3003 13507 3009
rect 13814 3000 13820 3012
rect 13872 3000 13878 3052
rect 20625 3043 20683 3049
rect 20625 3009 20637 3043
rect 20671 3040 20683 3043
rect 20732 3040 20760 3068
rect 20993 3043 21051 3049
rect 20993 3040 21005 3043
rect 20671 3012 21005 3040
rect 20671 3009 20683 3012
rect 20625 3003 20683 3009
rect 20993 3009 21005 3012
rect 21039 3009 21051 3043
rect 20993 3003 21051 3009
rect 12526 2972 12532 2984
rect 12439 2944 12532 2972
rect 12526 2932 12532 2944
rect 12584 2972 12590 2984
rect 13541 2975 13599 2981
rect 13541 2972 13553 2975
rect 12584 2944 13553 2972
rect 12584 2932 12590 2944
rect 13541 2941 13553 2944
rect 13587 2941 13599 2975
rect 13541 2935 13599 2941
rect 20717 2975 20775 2981
rect 20717 2941 20729 2975
rect 20763 2972 20775 2975
rect 20806 2972 20812 2984
rect 20763 2944 20812 2972
rect 20763 2941 20775 2944
rect 20717 2935 20775 2941
rect 20806 2932 20812 2944
rect 20864 2932 20870 2984
rect 11054 2864 11060 2916
rect 11112 2904 11118 2916
rect 12434 2904 12440 2916
rect 11112 2876 12440 2904
rect 11112 2864 11118 2876
rect 12434 2864 12440 2876
rect 12492 2864 12498 2916
rect 12802 2836 12808 2848
rect 12763 2808 12808 2836
rect 12802 2796 12808 2808
rect 12860 2796 12866 2848
rect 1104 2746 38824 2768
rect 1104 2694 19606 2746
rect 19658 2694 19670 2746
rect 19722 2694 19734 2746
rect 19786 2694 19798 2746
rect 19850 2694 38824 2746
rect 1104 2672 38824 2694
rect 12434 2592 12440 2644
rect 12492 2632 12498 2644
rect 14182 2632 14188 2644
rect 12492 2604 12537 2632
rect 14143 2604 14188 2632
rect 12492 2592 12498 2604
rect 14182 2592 14188 2604
rect 14240 2592 14246 2644
rect 20806 2632 20812 2644
rect 20767 2604 20812 2632
rect 20806 2592 20812 2604
rect 20864 2592 20870 2644
rect 28442 2632 28448 2644
rect 28403 2604 28448 2632
rect 28442 2592 28448 2604
rect 28500 2592 28506 2644
rect 12452 2496 12480 2592
rect 12897 2499 12955 2505
rect 12897 2496 12909 2499
rect 12452 2468 12909 2496
rect 12897 2465 12909 2468
rect 12943 2465 12955 2499
rect 12897 2459 12955 2465
rect 17773 2499 17831 2505
rect 17773 2465 17785 2499
rect 17819 2496 17831 2499
rect 18230 2496 18236 2508
rect 17819 2468 18236 2496
rect 17819 2465 17831 2468
rect 17773 2459 17831 2465
rect 18230 2456 18236 2468
rect 18288 2496 18294 2508
rect 18601 2499 18659 2505
rect 18601 2496 18613 2499
rect 18288 2468 18613 2496
rect 18288 2456 18294 2468
rect 18601 2465 18613 2468
rect 18647 2465 18659 2499
rect 24581 2499 24639 2505
rect 24581 2496 24593 2499
rect 18601 2459 18659 2465
rect 23768 2468 24593 2496
rect 12069 2431 12127 2437
rect 12069 2397 12081 2431
rect 12115 2428 12127 2431
rect 12526 2428 12532 2440
rect 12115 2400 12532 2428
rect 12115 2397 12127 2400
rect 12069 2391 12127 2397
rect 12526 2388 12532 2400
rect 12584 2428 12590 2440
rect 12621 2431 12679 2437
rect 12621 2428 12633 2431
rect 12584 2400 12633 2428
rect 12584 2388 12590 2400
rect 12621 2397 12633 2400
rect 12667 2397 12679 2431
rect 12621 2391 12679 2397
rect 18141 2431 18199 2437
rect 18141 2397 18153 2431
rect 18187 2428 18199 2431
rect 18877 2431 18935 2437
rect 18877 2428 18889 2431
rect 18187 2400 18889 2428
rect 18187 2397 18199 2400
rect 18141 2391 18199 2397
rect 18877 2397 18889 2400
rect 18923 2428 18935 2431
rect 18966 2428 18972 2440
rect 18923 2400 18972 2428
rect 18923 2397 18935 2400
rect 18877 2391 18935 2397
rect 18966 2388 18972 2400
rect 19024 2388 19030 2440
rect 23768 2372 23796 2468
rect 24581 2465 24593 2468
rect 24627 2465 24639 2499
rect 24581 2459 24639 2465
rect 25961 2499 26019 2505
rect 25961 2465 25973 2499
rect 26007 2496 26019 2499
rect 27614 2496 27620 2508
rect 26007 2468 27620 2496
rect 26007 2465 26019 2468
rect 25961 2459 26019 2465
rect 27614 2456 27620 2468
rect 27672 2456 27678 2508
rect 24305 2431 24363 2437
rect 24305 2428 24317 2431
rect 24228 2400 24317 2428
rect 23750 2360 23756 2372
rect 23711 2332 23756 2360
rect 23750 2320 23756 2332
rect 23808 2320 23814 2372
rect 19794 2252 19800 2304
rect 19852 2292 19858 2304
rect 19981 2295 20039 2301
rect 19981 2292 19993 2295
rect 19852 2264 19993 2292
rect 19852 2252 19858 2264
rect 19981 2261 19993 2264
rect 20027 2261 20039 2295
rect 19981 2255 20039 2261
rect 23477 2295 23535 2301
rect 23477 2261 23489 2295
rect 23523 2292 23535 2295
rect 24228 2292 24256 2400
rect 24305 2397 24317 2400
rect 24351 2428 24363 2431
rect 26142 2428 26148 2440
rect 24351 2400 26148 2428
rect 24351 2397 24363 2400
rect 24305 2391 24363 2397
rect 26142 2388 26148 2400
rect 26200 2428 26206 2440
rect 26237 2431 26295 2437
rect 26237 2428 26249 2431
rect 26200 2400 26249 2428
rect 26200 2388 26206 2400
rect 26237 2397 26249 2400
rect 26283 2428 26295 2431
rect 26888 2431 26946 2437
rect 26888 2428 26900 2431
rect 26283 2400 26900 2428
rect 26283 2397 26295 2400
rect 26237 2391 26295 2397
rect 26888 2397 26900 2400
rect 26934 2397 26946 2431
rect 27154 2428 27160 2440
rect 27067 2400 27160 2428
rect 26888 2391 26946 2397
rect 27154 2388 27160 2400
rect 27212 2428 27218 2440
rect 28534 2428 28540 2440
rect 27212 2400 28540 2428
rect 27212 2388 27218 2400
rect 28534 2388 28540 2400
rect 28592 2388 28598 2440
rect 23523 2264 24256 2292
rect 26697 2295 26755 2301
rect 23523 2261 23535 2264
rect 23477 2255 23535 2261
rect 26697 2261 26709 2295
rect 26743 2292 26755 2295
rect 27154 2292 27160 2304
rect 26743 2264 27160 2292
rect 26743 2261 26755 2264
rect 26697 2255 26755 2261
rect 27154 2252 27160 2264
rect 27212 2252 27218 2304
rect 1104 2202 38824 2224
rect 1104 2150 4246 2202
rect 4298 2150 4310 2202
rect 4362 2150 4374 2202
rect 4426 2150 4438 2202
rect 4490 2150 34966 2202
rect 35018 2150 35030 2202
rect 35082 2150 35094 2202
rect 35146 2150 35158 2202
rect 35210 2150 38824 2202
rect 1104 2128 38824 2150
rect 23474 1368 23480 1420
rect 23532 1408 23538 1420
rect 24578 1408 24584 1420
rect 23532 1380 24584 1408
rect 23532 1368 23538 1380
rect 24578 1368 24584 1380
rect 24636 1368 24642 1420
rect 474 1232 480 1284
rect 532 1272 538 1284
rect 4798 1272 4804 1284
rect 532 1244 4804 1272
rect 532 1232 538 1244
rect 4798 1232 4804 1244
rect 4856 1232 4862 1284
rect 3234 892 3240 944
rect 3292 932 3298 944
rect 3326 932 3332 944
rect 3292 904 3332 932
rect 3292 892 3298 904
rect 3326 892 3332 904
rect 3384 892 3390 944
<< via1 >>
rect 21180 77868 21232 77920
rect 24308 77868 24360 77920
rect 19606 77766 19658 77818
rect 19670 77766 19722 77818
rect 19734 77766 19786 77818
rect 19798 77766 19850 77818
rect 3976 77664 4028 77716
rect 33508 77664 33560 77716
rect 4068 77528 4120 77580
rect 24308 77571 24360 77580
rect 24308 77537 24317 77571
rect 24317 77537 24351 77571
rect 24351 77537 24360 77571
rect 24308 77528 24360 77537
rect 18052 77367 18104 77376
rect 18052 77333 18061 77367
rect 18061 77333 18095 77367
rect 18095 77333 18104 77367
rect 18052 77324 18104 77333
rect 29092 77460 29144 77512
rect 35348 77392 35400 77444
rect 24676 77324 24728 77376
rect 28080 77324 28132 77376
rect 28908 77324 28960 77376
rect 29460 77367 29512 77376
rect 29460 77333 29469 77367
rect 29469 77333 29503 77367
rect 29503 77333 29512 77367
rect 29460 77324 29512 77333
rect 4246 77222 4298 77274
rect 4310 77222 4362 77274
rect 4374 77222 4426 77274
rect 4438 77222 4490 77274
rect 34966 77222 35018 77274
rect 35030 77222 35082 77274
rect 35094 77222 35146 77274
rect 35158 77222 35210 77274
rect 24216 77120 24268 77172
rect 24400 77163 24452 77172
rect 24400 77129 24409 77163
rect 24409 77129 24443 77163
rect 24443 77129 24452 77163
rect 24400 77120 24452 77129
rect 29092 77163 29144 77172
rect 29092 77129 29101 77163
rect 29101 77129 29135 77163
rect 29135 77129 29144 77163
rect 29092 77120 29144 77129
rect 32220 77120 32272 77172
rect 24308 77052 24360 77104
rect 16120 76984 16172 77036
rect 18420 76984 18472 77036
rect 15476 76959 15528 76968
rect 15476 76925 15485 76959
rect 15485 76925 15519 76959
rect 15519 76925 15528 76959
rect 15476 76916 15528 76925
rect 17592 76916 17644 76968
rect 18052 76959 18104 76968
rect 18052 76925 18061 76959
rect 18061 76925 18095 76959
rect 18095 76925 18104 76959
rect 18052 76916 18104 76925
rect 21088 76959 21140 76968
rect 21088 76925 21097 76959
rect 21097 76925 21131 76959
rect 21131 76925 21140 76959
rect 21088 76916 21140 76925
rect 17684 76848 17736 76900
rect 19340 76780 19392 76832
rect 20904 76823 20956 76832
rect 20904 76789 20913 76823
rect 20913 76789 20947 76823
rect 20947 76789 20956 76823
rect 24676 76916 24728 76968
rect 28816 76916 28868 76968
rect 29460 76959 29512 76968
rect 29460 76925 29469 76959
rect 29469 76925 29503 76959
rect 29503 76925 29512 76959
rect 29460 76916 29512 76925
rect 20904 76780 20956 76789
rect 26976 76780 27028 76832
rect 19606 76678 19658 76730
rect 19670 76678 19722 76730
rect 19734 76678 19786 76730
rect 19798 76678 19850 76730
rect 21916 76440 21968 76492
rect 15476 76372 15528 76424
rect 17592 76415 17644 76424
rect 17592 76381 17601 76415
rect 17601 76381 17635 76415
rect 17635 76381 17644 76415
rect 17592 76372 17644 76381
rect 17776 76372 17828 76424
rect 22008 76372 22060 76424
rect 28816 76415 28868 76424
rect 28816 76381 28825 76415
rect 28825 76381 28859 76415
rect 28859 76381 28868 76415
rect 28816 76372 28868 76381
rect 29000 76372 29052 76424
rect 20536 76304 20588 76356
rect 21180 76347 21232 76356
rect 21180 76313 21189 76347
rect 21189 76313 21223 76347
rect 21223 76313 21232 76347
rect 21180 76304 21232 76313
rect 17868 76236 17920 76288
rect 22928 76279 22980 76288
rect 22928 76245 22937 76279
rect 22937 76245 22971 76279
rect 22971 76245 22980 76279
rect 22928 76236 22980 76245
rect 24124 76279 24176 76288
rect 24124 76245 24133 76279
rect 24133 76245 24167 76279
rect 24167 76245 24176 76279
rect 24676 76279 24728 76288
rect 24124 76236 24176 76245
rect 24676 76245 24685 76279
rect 24685 76245 24719 76279
rect 24719 76245 24728 76279
rect 24676 76236 24728 76245
rect 30380 76279 30432 76288
rect 30380 76245 30389 76279
rect 30389 76245 30423 76279
rect 30423 76245 30432 76279
rect 30380 76236 30432 76245
rect 4246 76134 4298 76186
rect 4310 76134 4362 76186
rect 4374 76134 4426 76186
rect 4438 76134 4490 76186
rect 34966 76134 35018 76186
rect 35030 76134 35082 76186
rect 35094 76134 35146 76186
rect 35158 76134 35210 76186
rect 22008 76032 22060 76084
rect 29000 76032 29052 76084
rect 17868 75964 17920 76016
rect 28816 75964 28868 76016
rect 17500 75896 17552 75948
rect 17592 75896 17644 75948
rect 19248 75896 19300 75948
rect 19340 75896 19392 75948
rect 112 75828 164 75880
rect 940 75828 992 75880
rect 25320 75828 25372 75880
rect 25872 75871 25924 75880
rect 25872 75837 25881 75871
rect 25881 75837 25915 75871
rect 25915 75837 25924 75871
rect 25872 75828 25924 75837
rect 27528 75803 27580 75812
rect 27528 75769 27537 75803
rect 27537 75769 27571 75803
rect 27571 75769 27580 75803
rect 27528 75760 27580 75769
rect 17776 75692 17828 75744
rect 20076 75692 20128 75744
rect 22008 75735 22060 75744
rect 22008 75701 22017 75735
rect 22017 75701 22051 75735
rect 22051 75701 22060 75735
rect 22008 75692 22060 75701
rect 19606 75590 19658 75642
rect 19670 75590 19722 75642
rect 19734 75590 19786 75642
rect 19798 75590 19850 75642
rect 29828 75463 29880 75472
rect 29828 75429 29837 75463
rect 29837 75429 29871 75463
rect 29871 75429 29880 75463
rect 29828 75420 29880 75429
rect 30380 75352 30432 75404
rect 29368 75284 29420 75336
rect 30656 75327 30708 75336
rect 30656 75293 30665 75327
rect 30665 75293 30699 75327
rect 30699 75293 30708 75327
rect 30656 75284 30708 75293
rect 19248 75148 19300 75200
rect 25964 75191 26016 75200
rect 25964 75157 25973 75191
rect 25973 75157 26007 75191
rect 26007 75157 26016 75191
rect 25964 75148 26016 75157
rect 4246 75046 4298 75098
rect 4310 75046 4362 75098
rect 4374 75046 4426 75098
rect 4438 75046 4490 75098
rect 34966 75046 35018 75098
rect 35030 75046 35082 75098
rect 35094 75046 35146 75098
rect 35158 75046 35210 75098
rect 30380 74987 30432 74996
rect 30380 74953 30389 74987
rect 30389 74953 30423 74987
rect 30423 74953 30432 74987
rect 30380 74944 30432 74953
rect 20076 74851 20128 74860
rect 20076 74817 20085 74851
rect 20085 74817 20119 74851
rect 20119 74817 20128 74851
rect 20076 74808 20128 74817
rect 9680 74740 9732 74792
rect 10876 74740 10928 74792
rect 15200 74740 15252 74792
rect 16488 74740 16540 74792
rect 19892 74740 19944 74792
rect 20536 74740 20588 74792
rect 37372 74740 37424 74792
rect 38660 74740 38712 74792
rect 2780 74604 2832 74656
rect 3884 74604 3936 74656
rect 19432 74604 19484 74656
rect 20076 74604 20128 74656
rect 20812 74604 20864 74656
rect 29368 74604 29420 74656
rect 30656 74604 30708 74656
rect 33140 74604 33192 74656
rect 34060 74604 34112 74656
rect 19606 74502 19658 74554
rect 19670 74502 19722 74554
rect 19734 74502 19786 74554
rect 19798 74502 19850 74554
rect 19892 74375 19944 74384
rect 19892 74341 19901 74375
rect 19901 74341 19935 74375
rect 19935 74341 19944 74375
rect 19892 74332 19944 74341
rect 4246 73958 4298 74010
rect 4310 73958 4362 74010
rect 4374 73958 4426 74010
rect 4438 73958 4490 74010
rect 34966 73958 35018 74010
rect 35030 73958 35082 74010
rect 35094 73958 35146 74010
rect 35158 73958 35210 74010
rect 26332 73856 26384 73908
rect 27160 73856 27212 73908
rect 19606 73414 19658 73466
rect 19670 73414 19722 73466
rect 19734 73414 19786 73466
rect 19798 73414 19850 73466
rect 19340 72972 19392 73024
rect 28816 72972 28868 73024
rect 4246 72870 4298 72922
rect 4310 72870 4362 72922
rect 4374 72870 4426 72922
rect 4438 72870 4490 72922
rect 34966 72870 35018 72922
rect 35030 72870 35082 72922
rect 35094 72870 35146 72922
rect 35158 72870 35210 72922
rect 19432 72564 19484 72616
rect 19340 72539 19392 72548
rect 19340 72505 19349 72539
rect 19349 72505 19383 72539
rect 19383 72505 19392 72539
rect 19340 72496 19392 72505
rect 21088 72471 21140 72480
rect 21088 72437 21097 72471
rect 21097 72437 21131 72471
rect 21131 72437 21140 72471
rect 21088 72428 21140 72437
rect 19606 72326 19658 72378
rect 19670 72326 19722 72378
rect 19734 72326 19786 72378
rect 19798 72326 19850 72378
rect 19524 71927 19576 71936
rect 19524 71893 19533 71927
rect 19533 71893 19567 71927
rect 19567 71893 19576 71927
rect 19524 71884 19576 71893
rect 4246 71782 4298 71834
rect 4310 71782 4362 71834
rect 4374 71782 4426 71834
rect 4438 71782 4490 71834
rect 34966 71782 35018 71834
rect 35030 71782 35082 71834
rect 35094 71782 35146 71834
rect 35158 71782 35210 71834
rect 19606 71238 19658 71290
rect 19670 71238 19722 71290
rect 19734 71238 19786 71290
rect 19798 71238 19850 71290
rect 22100 71000 22152 71052
rect 22744 71000 22796 71052
rect 23204 71000 23256 71052
rect 24308 70975 24360 70984
rect 24308 70941 24317 70975
rect 24317 70941 24351 70975
rect 24351 70941 24360 70975
rect 24308 70932 24360 70941
rect 4246 70694 4298 70746
rect 4310 70694 4362 70746
rect 4374 70694 4426 70746
rect 4438 70694 4490 70746
rect 34966 70694 35018 70746
rect 35030 70694 35082 70746
rect 35094 70694 35146 70746
rect 35158 70694 35210 70746
rect 22744 70592 22796 70644
rect 23388 70592 23440 70644
rect 23204 70456 23256 70508
rect 19606 70150 19658 70202
rect 19670 70150 19722 70202
rect 19734 70150 19786 70202
rect 19798 70150 19850 70202
rect 23480 69844 23532 69896
rect 23940 69887 23992 69896
rect 23940 69853 23949 69887
rect 23949 69853 23983 69887
rect 23983 69853 23992 69887
rect 23940 69844 23992 69853
rect 24216 69887 24268 69896
rect 24216 69853 24225 69887
rect 24225 69853 24259 69887
rect 24259 69853 24268 69887
rect 24216 69844 24268 69853
rect 24676 69708 24728 69760
rect 4246 69606 4298 69658
rect 4310 69606 4362 69658
rect 4374 69606 4426 69658
rect 4438 69606 4490 69658
rect 34966 69606 35018 69658
rect 35030 69606 35082 69658
rect 35094 69606 35146 69658
rect 35158 69606 35210 69658
rect 23940 69504 23992 69556
rect 25964 69547 26016 69556
rect 25964 69513 25973 69547
rect 25973 69513 26007 69547
rect 26007 69513 26016 69547
rect 25964 69504 26016 69513
rect 24216 69436 24268 69488
rect 25228 69232 25280 69284
rect 19606 69062 19658 69114
rect 19670 69062 19722 69114
rect 19734 69062 19786 69114
rect 19798 69062 19850 69114
rect 22836 68867 22888 68876
rect 22836 68833 22845 68867
rect 22845 68833 22879 68867
rect 22879 68833 22888 68867
rect 22836 68824 22888 68833
rect 25228 68867 25280 68876
rect 25228 68833 25237 68867
rect 25237 68833 25271 68867
rect 25271 68833 25280 68867
rect 25228 68824 25280 68833
rect 22560 68799 22612 68808
rect 22560 68765 22569 68799
rect 22569 68765 22603 68799
rect 22603 68765 22612 68799
rect 22560 68756 22612 68765
rect 22744 68756 22796 68808
rect 23940 68663 23992 68672
rect 23940 68629 23949 68663
rect 23949 68629 23983 68663
rect 23983 68629 23992 68663
rect 23940 68620 23992 68629
rect 24032 68620 24084 68672
rect 4246 68518 4298 68570
rect 4310 68518 4362 68570
rect 4374 68518 4426 68570
rect 4438 68518 4490 68570
rect 34966 68518 35018 68570
rect 35030 68518 35082 68570
rect 35094 68518 35146 68570
rect 35158 68518 35210 68570
rect 22836 68416 22888 68468
rect 24676 68280 24728 68332
rect 22560 68212 22612 68264
rect 24032 68255 24084 68264
rect 24032 68221 24041 68255
rect 24041 68221 24075 68255
rect 24075 68221 24084 68255
rect 24032 68212 24084 68221
rect 25872 68144 25924 68196
rect 19606 67974 19658 68026
rect 19670 67974 19722 68026
rect 19734 67974 19786 68026
rect 19798 67974 19850 68026
rect 19340 67872 19392 67924
rect 20904 67872 20956 67924
rect 14004 67600 14056 67652
rect 14096 67600 14148 67652
rect 24032 67600 24084 67652
rect 24492 67600 24544 67652
rect 25228 67600 25280 67652
rect 26424 67532 26476 67584
rect 4246 67430 4298 67482
rect 4310 67430 4362 67482
rect 4374 67430 4426 67482
rect 4438 67430 4490 67482
rect 34966 67430 35018 67482
rect 35030 67430 35082 67482
rect 35094 67430 35146 67482
rect 35158 67430 35210 67482
rect 26424 67371 26476 67380
rect 26424 67337 26433 67371
rect 26433 67337 26467 67371
rect 26467 67337 26476 67371
rect 26424 67328 26476 67337
rect 27068 66988 27120 67040
rect 19606 66886 19658 66938
rect 19670 66886 19722 66938
rect 19734 66886 19786 66938
rect 19798 66886 19850 66938
rect 4246 66342 4298 66394
rect 4310 66342 4362 66394
rect 4374 66342 4426 66394
rect 4438 66342 4490 66394
rect 34966 66342 35018 66394
rect 35030 66342 35082 66394
rect 35094 66342 35146 66394
rect 35158 66342 35210 66394
rect 17224 66240 17276 66292
rect 17500 66240 17552 66292
rect 17224 66104 17276 66156
rect 17592 66104 17644 66156
rect 19606 65798 19658 65850
rect 19670 65798 19722 65850
rect 19734 65798 19786 65850
rect 19798 65798 19850 65850
rect 1768 65399 1820 65408
rect 1768 65365 1777 65399
rect 1777 65365 1811 65399
rect 1811 65365 1820 65399
rect 1768 65356 1820 65365
rect 4246 65254 4298 65306
rect 4310 65254 4362 65306
rect 4374 65254 4426 65306
rect 4438 65254 4490 65306
rect 34966 65254 35018 65306
rect 35030 65254 35082 65306
rect 35094 65254 35146 65306
rect 35158 65254 35210 65306
rect 1584 65195 1636 65204
rect 1584 65161 1593 65195
rect 1593 65161 1627 65195
rect 1627 65161 1636 65195
rect 1584 65152 1636 65161
rect 1584 65016 1636 65068
rect 1768 65059 1820 65068
rect 1768 65025 1777 65059
rect 1777 65025 1811 65059
rect 1811 65025 1820 65059
rect 1768 65016 1820 65025
rect 4620 64880 4672 64932
rect 19606 64710 19658 64762
rect 19670 64710 19722 64762
rect 19734 64710 19786 64762
rect 19798 64710 19850 64762
rect 1584 64311 1636 64320
rect 1584 64277 1593 64311
rect 1593 64277 1627 64311
rect 1627 64277 1636 64311
rect 1584 64268 1636 64277
rect 4246 64166 4298 64218
rect 4310 64166 4362 64218
rect 4374 64166 4426 64218
rect 4438 64166 4490 64218
rect 34966 64166 35018 64218
rect 35030 64166 35082 64218
rect 35094 64166 35146 64218
rect 35158 64166 35210 64218
rect 1860 63971 1912 63980
rect 1860 63937 1869 63971
rect 1869 63937 1903 63971
rect 1903 63937 1912 63971
rect 1860 63928 1912 63937
rect 3884 63928 3936 63980
rect 1584 63903 1636 63912
rect 1584 63869 1593 63903
rect 1593 63869 1627 63903
rect 1627 63869 1636 63903
rect 1584 63860 1636 63869
rect 2688 63860 2740 63912
rect 4160 63903 4212 63912
rect 4160 63869 4169 63903
rect 4169 63869 4203 63903
rect 4203 63869 4212 63903
rect 4160 63860 4212 63869
rect 4252 63792 4304 63844
rect 5080 63903 5132 63912
rect 5080 63869 5089 63903
rect 5089 63869 5123 63903
rect 5123 63869 5132 63903
rect 5080 63860 5132 63869
rect 5080 63724 5132 63776
rect 19606 63622 19658 63674
rect 19670 63622 19722 63674
rect 19734 63622 19786 63674
rect 19798 63622 19850 63674
rect 1860 63520 1912 63572
rect 4252 63563 4304 63572
rect 4252 63529 4261 63563
rect 4261 63529 4295 63563
rect 4295 63529 4304 63563
rect 4252 63520 4304 63529
rect 4620 63384 4672 63436
rect 13820 63384 13872 63436
rect 20352 63384 20404 63436
rect 21640 63384 21692 63436
rect 2688 63316 2740 63368
rect 5172 63316 5224 63368
rect 21088 63359 21140 63368
rect 21088 63325 21097 63359
rect 21097 63325 21131 63359
rect 21131 63325 21140 63359
rect 21088 63316 21140 63325
rect 14004 63248 14056 63300
rect 21732 63291 21784 63300
rect 21732 63257 21741 63291
rect 21741 63257 21775 63291
rect 21775 63257 21784 63291
rect 21732 63248 21784 63257
rect 6920 63180 6972 63232
rect 18604 63180 18656 63232
rect 18880 63180 18932 63232
rect 4246 63078 4298 63130
rect 4310 63078 4362 63130
rect 4374 63078 4426 63130
rect 4438 63078 4490 63130
rect 34966 63078 35018 63130
rect 35030 63078 35082 63130
rect 35094 63078 35146 63130
rect 35158 63078 35210 63130
rect 4620 62976 4672 63028
rect 20352 63019 20404 63028
rect 20352 62985 20361 63019
rect 20361 62985 20395 63019
rect 20395 62985 20404 63019
rect 20352 62976 20404 62985
rect 18880 62840 18932 62892
rect 20076 62840 20128 62892
rect 22284 62883 22336 62892
rect 22284 62849 22293 62883
rect 22293 62849 22327 62883
rect 22327 62849 22336 62883
rect 22284 62840 22336 62849
rect 21088 62815 21140 62824
rect 18604 62704 18656 62756
rect 21088 62781 21097 62815
rect 21097 62781 21131 62815
rect 21131 62781 21140 62815
rect 21088 62772 21140 62781
rect 21456 62772 21508 62824
rect 5172 62679 5224 62688
rect 5172 62645 5181 62679
rect 5181 62645 5215 62679
rect 5215 62645 5224 62679
rect 5172 62636 5224 62645
rect 13820 62636 13872 62688
rect 21732 62772 21784 62824
rect 28724 62772 28776 62824
rect 28908 62772 28960 62824
rect 22008 62636 22060 62688
rect 19606 62534 19658 62586
rect 19670 62534 19722 62586
rect 19734 62534 19786 62586
rect 19798 62534 19850 62586
rect 18512 62296 18564 62348
rect 18880 62296 18932 62348
rect 26056 62296 26108 62348
rect 26516 62339 26568 62348
rect 26516 62305 26525 62339
rect 26525 62305 26559 62339
rect 26559 62305 26568 62339
rect 26516 62296 26568 62305
rect 26792 62339 26844 62348
rect 26792 62305 26801 62339
rect 26801 62305 26835 62339
rect 26835 62305 26844 62339
rect 26792 62296 26844 62305
rect 18420 62271 18472 62280
rect 18420 62237 18429 62271
rect 18429 62237 18463 62271
rect 18463 62237 18472 62271
rect 18420 62228 18472 62237
rect 25780 62228 25832 62280
rect 25964 62228 26016 62280
rect 19064 62203 19116 62212
rect 19064 62169 19073 62203
rect 19073 62169 19107 62203
rect 19107 62169 19116 62203
rect 19064 62160 19116 62169
rect 21180 62135 21232 62144
rect 21180 62101 21189 62135
rect 21189 62101 21223 62135
rect 21223 62101 21232 62135
rect 21180 62092 21232 62101
rect 21732 62092 21784 62144
rect 22008 62135 22060 62144
rect 22008 62101 22017 62135
rect 22017 62101 22051 62135
rect 22051 62101 22060 62135
rect 22008 62092 22060 62101
rect 27804 62092 27856 62144
rect 4246 61990 4298 62042
rect 4310 61990 4362 62042
rect 4374 61990 4426 62042
rect 4438 61990 4490 62042
rect 34966 61990 35018 62042
rect 35030 61990 35082 62042
rect 35094 61990 35146 62042
rect 35158 61990 35210 62042
rect 18420 61888 18472 61940
rect 26792 61888 26844 61940
rect 26516 61820 26568 61872
rect 13176 61591 13228 61600
rect 13176 61557 13185 61591
rect 13185 61557 13219 61591
rect 13219 61557 13228 61591
rect 13176 61548 13228 61557
rect 13912 61548 13964 61600
rect 18512 61548 18564 61600
rect 18880 61548 18932 61600
rect 20076 61548 20128 61600
rect 21916 61548 21968 61600
rect 19606 61446 19658 61498
rect 19670 61446 19722 61498
rect 19734 61446 19786 61498
rect 19798 61446 19850 61498
rect 20352 61344 20404 61396
rect 10968 61251 11020 61260
rect 10968 61217 10977 61251
rect 10977 61217 11011 61251
rect 11011 61217 11020 61251
rect 10968 61208 11020 61217
rect 19340 61208 19392 61260
rect 21916 61251 21968 61260
rect 21364 61140 21416 61192
rect 21916 61217 21925 61251
rect 21925 61217 21959 61251
rect 21959 61217 21968 61251
rect 21916 61208 21968 61217
rect 22008 61140 22060 61192
rect 20260 61072 20312 61124
rect 20720 61072 20772 61124
rect 10784 61047 10836 61056
rect 10784 61013 10793 61047
rect 10793 61013 10827 61047
rect 10827 61013 10836 61047
rect 10784 61004 10836 61013
rect 20076 61004 20128 61056
rect 22100 61004 22152 61056
rect 22560 61047 22612 61056
rect 22560 61013 22569 61047
rect 22569 61013 22603 61047
rect 22603 61013 22612 61047
rect 22560 61004 22612 61013
rect 26056 61004 26108 61056
rect 4246 60902 4298 60954
rect 4310 60902 4362 60954
rect 4374 60902 4426 60954
rect 4438 60902 4490 60954
rect 34966 60902 35018 60954
rect 35030 60902 35082 60954
rect 35094 60902 35146 60954
rect 35158 60902 35210 60954
rect 10968 60800 11020 60852
rect 18420 60800 18472 60852
rect 21364 60800 21416 60852
rect 23020 60800 23072 60852
rect 9404 60732 9456 60784
rect 20628 60775 20680 60784
rect 20628 60741 20637 60775
rect 20637 60741 20671 60775
rect 20671 60741 20680 60775
rect 20628 60732 20680 60741
rect 20076 60664 20128 60716
rect 24308 60664 24360 60716
rect 31208 60707 31260 60716
rect 31208 60673 31217 60707
rect 31217 60673 31251 60707
rect 31251 60673 31260 60707
rect 31208 60664 31260 60673
rect 37464 60664 37516 60716
rect 9496 60596 9548 60648
rect 19984 60639 20036 60648
rect 19984 60605 19993 60639
rect 19993 60605 20027 60639
rect 20027 60605 20036 60639
rect 19984 60596 20036 60605
rect 20260 60639 20312 60648
rect 20260 60605 20269 60639
rect 20269 60605 20303 60639
rect 20303 60605 20312 60639
rect 20260 60596 20312 60605
rect 20536 60596 20588 60648
rect 22100 60596 22152 60648
rect 19432 60528 19484 60580
rect 20076 60528 20128 60580
rect 21548 60528 21600 60580
rect 22376 60596 22428 60648
rect 22560 60639 22612 60648
rect 22560 60605 22569 60639
rect 22569 60605 22603 60639
rect 22603 60605 22612 60639
rect 22560 60596 22612 60605
rect 25504 60596 25556 60648
rect 26056 60596 26108 60648
rect 26240 60639 26292 60648
rect 26240 60605 26249 60639
rect 26249 60605 26283 60639
rect 26283 60605 26292 60639
rect 30932 60639 30984 60648
rect 26240 60596 26292 60605
rect 30932 60605 30941 60639
rect 30941 60605 30975 60639
rect 30975 60605 30984 60639
rect 30932 60596 30984 60605
rect 35808 60639 35860 60648
rect 35808 60605 35817 60639
rect 35817 60605 35851 60639
rect 35851 60605 35860 60639
rect 35808 60596 35860 60605
rect 26516 60528 26568 60580
rect 19340 60503 19392 60512
rect 19340 60469 19349 60503
rect 19349 60469 19383 60503
rect 19383 60469 19392 60503
rect 19340 60460 19392 60469
rect 21640 60503 21692 60512
rect 21640 60469 21649 60503
rect 21649 60469 21683 60503
rect 21683 60469 21692 60503
rect 21640 60460 21692 60469
rect 22376 60460 22428 60512
rect 32312 60503 32364 60512
rect 32312 60469 32321 60503
rect 32321 60469 32355 60503
rect 32355 60469 32364 60503
rect 32312 60460 32364 60469
rect 37372 60503 37424 60512
rect 37372 60469 37381 60503
rect 37381 60469 37415 60503
rect 37415 60469 37424 60503
rect 37372 60460 37424 60469
rect 19606 60358 19658 60410
rect 19670 60358 19722 60410
rect 19734 60358 19786 60410
rect 19798 60358 19850 60410
rect 20352 60299 20404 60308
rect 20352 60265 20361 60299
rect 20361 60265 20395 60299
rect 20395 60265 20404 60299
rect 20352 60256 20404 60265
rect 21548 60256 21600 60308
rect 24492 60299 24544 60308
rect 19248 60163 19300 60172
rect 19248 60129 19257 60163
rect 19257 60129 19291 60163
rect 19291 60129 19300 60163
rect 19248 60120 19300 60129
rect 19708 60120 19760 60172
rect 20168 60120 20220 60172
rect 24492 60265 24501 60299
rect 24501 60265 24535 60299
rect 24535 60265 24544 60299
rect 24492 60256 24544 60265
rect 25320 60299 25372 60308
rect 25320 60265 25329 60299
rect 25329 60265 25363 60299
rect 25363 60265 25372 60299
rect 25320 60256 25372 60265
rect 29552 60299 29604 60308
rect 29552 60265 29561 60299
rect 29561 60265 29595 60299
rect 29595 60265 29604 60299
rect 29552 60256 29604 60265
rect 30472 60256 30524 60308
rect 30932 60299 30984 60308
rect 30932 60265 30941 60299
rect 30941 60265 30975 60299
rect 30975 60265 30984 60299
rect 30932 60256 30984 60265
rect 22836 60163 22888 60172
rect 18052 60052 18104 60104
rect 20444 60052 20496 60104
rect 21088 60095 21140 60104
rect 21088 60061 21097 60095
rect 21097 60061 21131 60095
rect 21131 60061 21140 60095
rect 21088 60052 21140 60061
rect 20168 59984 20220 60036
rect 22836 60129 22845 60163
rect 22845 60129 22879 60163
rect 22879 60129 22888 60163
rect 22836 60120 22888 60129
rect 27804 60120 27856 60172
rect 28172 60120 28224 60172
rect 29184 60120 29236 60172
rect 21824 60095 21876 60104
rect 21824 60061 21833 60095
rect 21833 60061 21867 60095
rect 21867 60061 21876 60095
rect 21824 60052 21876 60061
rect 26608 60095 26660 60104
rect 26608 60061 26617 60095
rect 26617 60061 26651 60095
rect 26651 60061 26660 60095
rect 26608 60052 26660 60061
rect 23020 60027 23072 60036
rect 23020 59993 23029 60027
rect 23029 59993 23063 60027
rect 23063 59993 23072 60027
rect 23020 59984 23072 59993
rect 18604 59959 18656 59968
rect 18604 59925 18613 59959
rect 18613 59925 18647 59959
rect 18647 59925 18656 59959
rect 18604 59916 18656 59925
rect 19524 59959 19576 59968
rect 19524 59925 19533 59959
rect 19533 59925 19567 59959
rect 19567 59925 19576 59959
rect 19524 59916 19576 59925
rect 19892 59959 19944 59968
rect 19892 59925 19901 59959
rect 19901 59925 19935 59959
rect 19935 59925 19944 59959
rect 19892 59916 19944 59925
rect 21824 59916 21876 59968
rect 23848 59959 23900 59968
rect 23848 59925 23857 59959
rect 23857 59925 23891 59959
rect 23891 59925 23900 59959
rect 23848 59916 23900 59925
rect 24308 59916 24360 59968
rect 29920 59916 29972 59968
rect 35256 59916 35308 59968
rect 35808 59959 35860 59968
rect 35808 59925 35817 59959
rect 35817 59925 35851 59959
rect 35851 59925 35860 59959
rect 35808 59916 35860 59925
rect 4246 59814 4298 59866
rect 4310 59814 4362 59866
rect 4374 59814 4426 59866
rect 4438 59814 4490 59866
rect 34966 59814 35018 59866
rect 35030 59814 35082 59866
rect 35094 59814 35146 59866
rect 35158 59814 35210 59866
rect 17868 59755 17920 59764
rect 17868 59721 17877 59755
rect 17877 59721 17911 59755
rect 17911 59721 17920 59755
rect 17868 59712 17920 59721
rect 19892 59712 19944 59764
rect 22836 59755 22888 59764
rect 22836 59721 22845 59755
rect 22845 59721 22879 59755
rect 22879 59721 22888 59755
rect 22836 59712 22888 59721
rect 25504 59755 25556 59764
rect 25504 59721 25513 59755
rect 25513 59721 25547 59755
rect 25547 59721 25556 59755
rect 25504 59712 25556 59721
rect 19984 59644 20036 59696
rect 22192 59644 22244 59696
rect 27252 59687 27304 59696
rect 27252 59653 27261 59687
rect 27261 59653 27295 59687
rect 27295 59653 27304 59687
rect 27252 59644 27304 59653
rect 20536 59576 20588 59628
rect 20628 59619 20680 59628
rect 20628 59585 20637 59619
rect 20637 59585 20671 59619
rect 20671 59585 20680 59619
rect 20628 59576 20680 59585
rect 22744 59576 22796 59628
rect 24400 59576 24452 59628
rect 26608 59619 26660 59628
rect 26608 59585 26617 59619
rect 26617 59585 26651 59619
rect 26651 59585 26660 59619
rect 26608 59576 26660 59585
rect 30380 59619 30432 59628
rect 30380 59585 30389 59619
rect 30389 59585 30423 59619
rect 30423 59585 30432 59619
rect 30380 59576 30432 59585
rect 18604 59551 18656 59560
rect 18604 59517 18613 59551
rect 18613 59517 18647 59551
rect 18647 59517 18656 59551
rect 18604 59508 18656 59517
rect 20168 59551 20220 59560
rect 20168 59517 20177 59551
rect 20177 59517 20211 59551
rect 20211 59517 20220 59551
rect 20168 59508 20220 59517
rect 20352 59508 20404 59560
rect 21824 59551 21876 59560
rect 21824 59517 21833 59551
rect 21833 59517 21867 59551
rect 21867 59517 21876 59551
rect 21824 59508 21876 59517
rect 22376 59551 22428 59560
rect 22376 59517 22385 59551
rect 22385 59517 22419 59551
rect 22419 59517 22428 59551
rect 24216 59551 24268 59560
rect 22376 59508 22428 59517
rect 18144 59372 18196 59424
rect 19524 59440 19576 59492
rect 19708 59440 19760 59492
rect 24216 59517 24225 59551
rect 24225 59517 24259 59551
rect 24259 59517 24268 59551
rect 24216 59508 24268 59517
rect 26792 59551 26844 59560
rect 26792 59517 26801 59551
rect 26801 59517 26835 59551
rect 26835 59517 26844 59551
rect 26792 59508 26844 59517
rect 26516 59440 26568 59492
rect 29000 59508 29052 59560
rect 32312 59576 32364 59628
rect 20536 59372 20588 59424
rect 20904 59415 20956 59424
rect 20904 59381 20913 59415
rect 20913 59381 20947 59415
rect 20947 59381 20956 59415
rect 20904 59372 20956 59381
rect 23296 59415 23348 59424
rect 23296 59381 23305 59415
rect 23305 59381 23339 59415
rect 23339 59381 23348 59415
rect 23296 59372 23348 59381
rect 28172 59415 28224 59424
rect 28172 59381 28181 59415
rect 28181 59381 28215 59415
rect 28215 59381 28224 59415
rect 28172 59372 28224 59381
rect 29184 59372 29236 59424
rect 29920 59372 29972 59424
rect 19606 59270 19658 59322
rect 19670 59270 19722 59322
rect 19734 59270 19786 59322
rect 19798 59270 19850 59322
rect 1584 59211 1636 59220
rect 1584 59177 1593 59211
rect 1593 59177 1627 59211
rect 1627 59177 1636 59211
rect 1584 59168 1636 59177
rect 21548 59211 21600 59220
rect 21548 59177 21557 59211
rect 21557 59177 21591 59211
rect 21591 59177 21600 59211
rect 21548 59168 21600 59177
rect 22100 59168 22152 59220
rect 22376 59211 22428 59220
rect 22376 59177 22385 59211
rect 22385 59177 22419 59211
rect 22419 59177 22428 59211
rect 22376 59168 22428 59177
rect 19248 59143 19300 59152
rect 19248 59109 19257 59143
rect 19257 59109 19291 59143
rect 19291 59109 19300 59143
rect 19248 59100 19300 59109
rect 19984 59100 20036 59152
rect 21824 59100 21876 59152
rect 24492 59100 24544 59152
rect 26516 59143 26568 59152
rect 16580 59032 16632 59084
rect 17408 59032 17460 59084
rect 20904 59075 20956 59084
rect 20904 59041 20913 59075
rect 20913 59041 20947 59075
rect 20947 59041 20956 59075
rect 20904 59032 20956 59041
rect 23020 59075 23072 59084
rect 23020 59041 23029 59075
rect 23029 59041 23063 59075
rect 23063 59041 23072 59075
rect 23020 59032 23072 59041
rect 23296 59075 23348 59084
rect 23296 59041 23305 59075
rect 23305 59041 23339 59075
rect 23339 59041 23348 59075
rect 23296 59032 23348 59041
rect 23848 59032 23900 59084
rect 24308 59032 24360 59084
rect 26516 59109 26525 59143
rect 26525 59109 26559 59143
rect 26559 59109 26568 59143
rect 26516 59100 26568 59109
rect 26608 59100 26660 59152
rect 29092 59143 29144 59152
rect 27252 59032 27304 59084
rect 29092 59109 29101 59143
rect 29101 59109 29135 59143
rect 29135 59109 29144 59143
rect 29092 59100 29144 59109
rect 29828 59075 29880 59084
rect 29828 59041 29837 59075
rect 29837 59041 29871 59075
rect 29871 59041 29880 59075
rect 29828 59032 29880 59041
rect 35256 59032 35308 59084
rect 35440 59075 35492 59084
rect 35440 59041 35449 59075
rect 35449 59041 35483 59075
rect 35483 59041 35492 59075
rect 35440 59032 35492 59041
rect 17224 58964 17276 59016
rect 17868 58964 17920 59016
rect 18052 59007 18104 59016
rect 18052 58973 18061 59007
rect 18061 58973 18095 59007
rect 18095 58973 18104 59007
rect 18052 58964 18104 58973
rect 18972 58964 19024 59016
rect 20444 58964 20496 59016
rect 22744 58964 22796 59016
rect 25136 58964 25188 59016
rect 27068 59007 27120 59016
rect 27068 58973 27077 59007
rect 27077 58973 27111 59007
rect 27111 58973 27120 59007
rect 27068 58964 27120 58973
rect 29000 59007 29052 59016
rect 29000 58973 29009 59007
rect 29009 58973 29043 59007
rect 29043 58973 29052 59007
rect 29000 58964 29052 58973
rect 29736 58964 29788 59016
rect 19984 58896 20036 58948
rect 23388 58939 23440 58948
rect 23388 58905 23397 58939
rect 23397 58905 23431 58939
rect 23431 58905 23440 58939
rect 23388 58896 23440 58905
rect 25228 58939 25280 58948
rect 25228 58905 25237 58939
rect 25237 58905 25271 58939
rect 25271 58905 25280 58939
rect 25228 58896 25280 58905
rect 16764 58828 16816 58880
rect 17408 58828 17460 58880
rect 17776 58828 17828 58880
rect 18052 58828 18104 58880
rect 18328 58871 18380 58880
rect 18328 58837 18337 58871
rect 18337 58837 18371 58871
rect 18371 58837 18380 58871
rect 18328 58828 18380 58837
rect 19064 58828 19116 58880
rect 19892 58871 19944 58880
rect 19892 58837 19901 58871
rect 19901 58837 19935 58871
rect 19935 58837 19944 58871
rect 19892 58828 19944 58837
rect 20536 58828 20588 58880
rect 21916 58871 21968 58880
rect 21916 58837 21925 58871
rect 21925 58837 21959 58871
rect 21959 58837 21968 58871
rect 21916 58828 21968 58837
rect 24216 58828 24268 58880
rect 24584 58828 24636 58880
rect 35808 58828 35860 58880
rect 4246 58726 4298 58778
rect 4310 58726 4362 58778
rect 4374 58726 4426 58778
rect 4438 58726 4490 58778
rect 34966 58726 35018 58778
rect 35030 58726 35082 58778
rect 35094 58726 35146 58778
rect 35158 58726 35210 58778
rect 17224 58624 17276 58676
rect 19064 58667 19116 58676
rect 19064 58633 19088 58667
rect 19088 58633 19116 58667
rect 19064 58624 19116 58633
rect 19432 58624 19484 58676
rect 23020 58624 23072 58676
rect 25136 58667 25188 58676
rect 25136 58633 25145 58667
rect 25145 58633 25179 58667
rect 25179 58633 25188 58667
rect 25136 58624 25188 58633
rect 35440 58624 35492 58676
rect 19156 58599 19208 58608
rect 19156 58565 19165 58599
rect 19165 58565 19199 58599
rect 19199 58565 19208 58599
rect 19156 58556 19208 58565
rect 1584 58531 1636 58540
rect 1584 58497 1593 58531
rect 1593 58497 1627 58531
rect 1627 58497 1636 58531
rect 1584 58488 1636 58497
rect 1860 58531 1912 58540
rect 1860 58497 1869 58531
rect 1869 58497 1903 58531
rect 1903 58497 1912 58531
rect 1860 58488 1912 58497
rect 21180 58531 21232 58540
rect 16948 58463 17000 58472
rect 16948 58429 16957 58463
rect 16957 58429 16991 58463
rect 16991 58429 17000 58463
rect 16948 58420 17000 58429
rect 18972 58420 19024 58472
rect 21180 58497 21189 58531
rect 21189 58497 21223 58531
rect 21223 58497 21232 58531
rect 21180 58488 21232 58497
rect 21916 58488 21968 58540
rect 24124 58556 24176 58608
rect 27252 58556 27304 58608
rect 27712 58599 27764 58608
rect 27712 58565 27721 58599
rect 27721 58565 27755 58599
rect 27755 58565 27764 58599
rect 27712 58556 27764 58565
rect 21640 58420 21692 58472
rect 21824 58420 21876 58472
rect 24768 58531 24820 58540
rect 24768 58497 24777 58531
rect 24777 58497 24811 58531
rect 24811 58497 24820 58531
rect 24768 58488 24820 58497
rect 22376 58420 22428 58472
rect 24216 58463 24268 58472
rect 24216 58429 24225 58463
rect 24225 58429 24259 58463
rect 24259 58429 24268 58463
rect 24216 58420 24268 58429
rect 24492 58420 24544 58472
rect 19156 58352 19208 58404
rect 23020 58352 23072 58404
rect 25228 58352 25280 58404
rect 2964 58327 3016 58336
rect 2964 58293 2973 58327
rect 2973 58293 3007 58327
rect 3007 58293 3016 58327
rect 2964 58284 3016 58293
rect 16580 58284 16632 58336
rect 18144 58284 18196 58336
rect 19984 58327 20036 58336
rect 19984 58293 19993 58327
rect 19993 58293 20027 58327
rect 20027 58293 20036 58327
rect 19984 58284 20036 58293
rect 20536 58327 20588 58336
rect 20536 58293 20545 58327
rect 20545 58293 20579 58327
rect 20579 58293 20588 58327
rect 20536 58284 20588 58293
rect 22744 58284 22796 58336
rect 25320 58284 25372 58336
rect 26884 58463 26936 58472
rect 26884 58429 26893 58463
rect 26893 58429 26927 58463
rect 26927 58429 26936 58463
rect 26884 58420 26936 58429
rect 26792 58327 26844 58336
rect 26792 58293 26801 58327
rect 26801 58293 26835 58327
rect 26835 58293 26844 58327
rect 27620 58420 27672 58472
rect 29000 58420 29052 58472
rect 26792 58284 26844 58293
rect 27620 58284 27672 58336
rect 29736 58284 29788 58336
rect 35256 58284 35308 58336
rect 19606 58182 19658 58234
rect 19670 58182 19722 58234
rect 19734 58182 19786 58234
rect 19798 58182 19850 58234
rect 1860 58080 1912 58132
rect 15660 58123 15712 58132
rect 15660 58089 15669 58123
rect 15669 58089 15703 58123
rect 15703 58089 15712 58123
rect 15660 58080 15712 58089
rect 19340 58080 19392 58132
rect 24492 58080 24544 58132
rect 26608 58080 26660 58132
rect 29828 58080 29880 58132
rect 15108 57944 15160 57996
rect 20904 58055 20956 58064
rect 20904 58021 20913 58055
rect 20913 58021 20947 58055
rect 20947 58021 20956 58055
rect 20904 58012 20956 58021
rect 9128 57876 9180 57928
rect 9496 57876 9548 57928
rect 13728 57876 13780 57928
rect 13912 57876 13964 57928
rect 19156 57944 19208 57996
rect 18052 57876 18104 57928
rect 18972 57876 19024 57928
rect 20168 57919 20220 57928
rect 20168 57885 20177 57919
rect 20177 57885 20211 57919
rect 20211 57885 20220 57919
rect 23296 57944 23348 57996
rect 20168 57876 20220 57885
rect 22744 57919 22796 57928
rect 16488 57740 16540 57792
rect 16672 57783 16724 57792
rect 16672 57749 16681 57783
rect 16681 57749 16715 57783
rect 16715 57749 16724 57783
rect 16672 57740 16724 57749
rect 19064 57808 19116 57860
rect 20904 57808 20956 57860
rect 22744 57885 22753 57919
rect 22753 57885 22787 57919
rect 22787 57885 22796 57919
rect 22744 57876 22796 57885
rect 22836 57876 22888 57928
rect 28724 58012 28776 58064
rect 24032 57944 24084 57996
rect 25228 57944 25280 57996
rect 28448 57987 28500 57996
rect 28448 57953 28457 57987
rect 28457 57953 28491 57987
rect 28491 57953 28500 57987
rect 28448 57944 28500 57953
rect 28816 57944 28868 57996
rect 22468 57808 22520 57860
rect 24308 57851 24360 57860
rect 24308 57817 24317 57851
rect 24317 57817 24351 57851
rect 24351 57817 24360 57851
rect 24308 57808 24360 57817
rect 17132 57740 17184 57792
rect 17408 57783 17460 57792
rect 17408 57749 17417 57783
rect 17417 57749 17451 57783
rect 17451 57749 17460 57783
rect 17408 57740 17460 57749
rect 18972 57783 19024 57792
rect 18972 57749 18981 57783
rect 18981 57749 19015 57783
rect 19015 57749 19024 57783
rect 18972 57740 19024 57749
rect 19432 57740 19484 57792
rect 20628 57740 20680 57792
rect 21180 57783 21232 57792
rect 21180 57749 21189 57783
rect 21189 57749 21223 57783
rect 21223 57749 21232 57783
rect 21180 57740 21232 57749
rect 21364 57783 21416 57792
rect 21364 57749 21373 57783
rect 21373 57749 21407 57783
rect 21407 57749 21416 57783
rect 21364 57740 21416 57749
rect 22008 57783 22060 57792
rect 22008 57749 22017 57783
rect 22017 57749 22051 57783
rect 22051 57749 22060 57783
rect 22008 57740 22060 57749
rect 22376 57783 22428 57792
rect 22376 57749 22385 57783
rect 22385 57749 22419 57783
rect 22419 57749 22428 57783
rect 22376 57740 22428 57749
rect 23480 57740 23532 57792
rect 24216 57740 24268 57792
rect 24768 57740 24820 57792
rect 27344 57876 27396 57928
rect 28540 57876 28592 57928
rect 28632 57919 28684 57928
rect 28632 57885 28641 57919
rect 28641 57885 28675 57919
rect 28675 57885 28684 57919
rect 28632 57876 28684 57885
rect 30012 57876 30064 57928
rect 30564 57876 30616 57928
rect 26884 57740 26936 57792
rect 28356 57740 28408 57792
rect 4246 57638 4298 57690
rect 4310 57638 4362 57690
rect 4374 57638 4426 57690
rect 4438 57638 4490 57690
rect 34966 57638 35018 57690
rect 35030 57638 35082 57690
rect 35094 57638 35146 57690
rect 35158 57638 35210 57690
rect 14280 57579 14332 57588
rect 14280 57545 14289 57579
rect 14289 57545 14323 57579
rect 14323 57545 14332 57579
rect 14280 57536 14332 57545
rect 15108 57536 15160 57588
rect 17868 57579 17920 57588
rect 17868 57545 17877 57579
rect 17877 57545 17911 57579
rect 17911 57545 17920 57579
rect 17868 57536 17920 57545
rect 19064 57536 19116 57588
rect 19616 57579 19668 57588
rect 19616 57545 19625 57579
rect 19625 57545 19659 57579
rect 19659 57545 19668 57579
rect 19616 57536 19668 57545
rect 18144 57468 18196 57520
rect 19432 57511 19484 57520
rect 19432 57477 19441 57511
rect 19441 57477 19475 57511
rect 19475 57477 19484 57511
rect 21180 57536 21232 57588
rect 24124 57579 24176 57588
rect 24124 57545 24133 57579
rect 24133 57545 24167 57579
rect 24167 57545 24176 57579
rect 24124 57536 24176 57545
rect 25136 57536 25188 57588
rect 29000 57579 29052 57588
rect 19432 57468 19484 57477
rect 22008 57468 22060 57520
rect 25228 57511 25280 57520
rect 15016 57307 15068 57316
rect 15016 57273 15025 57307
rect 15025 57273 15059 57307
rect 15059 57273 15068 57307
rect 16580 57332 16632 57384
rect 18144 57375 18196 57384
rect 18144 57341 18153 57375
rect 18153 57341 18187 57375
rect 18187 57341 18196 57375
rect 18144 57332 18196 57341
rect 19432 57332 19484 57384
rect 20444 57400 20496 57452
rect 21916 57400 21968 57452
rect 20720 57375 20772 57384
rect 20720 57341 20729 57375
rect 20729 57341 20763 57375
rect 20763 57341 20772 57375
rect 20720 57332 20772 57341
rect 21364 57332 21416 57384
rect 22284 57375 22336 57384
rect 22284 57341 22293 57375
rect 22293 57341 22327 57375
rect 22327 57341 22336 57375
rect 22284 57332 22336 57341
rect 22376 57332 22428 57384
rect 25228 57477 25237 57511
rect 25237 57477 25271 57511
rect 25271 57477 25280 57511
rect 25228 57468 25280 57477
rect 15016 57264 15068 57273
rect 17408 57264 17460 57316
rect 17868 57264 17920 57316
rect 19156 57307 19208 57316
rect 19156 57273 19165 57307
rect 19165 57273 19199 57307
rect 19199 57273 19208 57307
rect 19156 57264 19208 57273
rect 22744 57332 22796 57384
rect 23572 57332 23624 57384
rect 24124 57332 24176 57384
rect 29000 57545 29009 57579
rect 29009 57545 29043 57579
rect 29043 57545 29052 57579
rect 29000 57536 29052 57545
rect 27252 57511 27304 57520
rect 27252 57477 27261 57511
rect 27261 57477 27295 57511
rect 27295 57477 27304 57511
rect 27252 57468 27304 57477
rect 27528 57400 27580 57452
rect 26700 57332 26752 57384
rect 28448 57400 28500 57452
rect 28632 57400 28684 57452
rect 28356 57375 28408 57384
rect 25596 57264 25648 57316
rect 28356 57341 28365 57375
rect 28365 57341 28399 57375
rect 28399 57341 28408 57375
rect 28356 57332 28408 57341
rect 29000 57332 29052 57384
rect 35256 57375 35308 57384
rect 35256 57341 35265 57375
rect 35265 57341 35299 57375
rect 35299 57341 35308 57375
rect 35256 57332 35308 57341
rect 35808 57332 35860 57384
rect 28724 57264 28776 57316
rect 18052 57196 18104 57248
rect 18972 57239 19024 57248
rect 18972 57205 18981 57239
rect 18981 57205 19015 57239
rect 19015 57205 19024 57239
rect 18972 57196 19024 57205
rect 19248 57196 19300 57248
rect 20444 57196 20496 57248
rect 20628 57196 20680 57248
rect 20904 57196 20956 57248
rect 23296 57196 23348 57248
rect 24308 57196 24360 57248
rect 28540 57196 28592 57248
rect 35900 57196 35952 57248
rect 19606 57094 19658 57146
rect 19670 57094 19722 57146
rect 19734 57094 19786 57146
rect 19798 57094 19850 57146
rect 19064 56992 19116 57044
rect 20168 57035 20220 57044
rect 20168 57001 20177 57035
rect 20177 57001 20211 57035
rect 20211 57001 20220 57035
rect 20168 56992 20220 57001
rect 20720 57035 20772 57044
rect 20720 57001 20729 57035
rect 20729 57001 20763 57035
rect 20763 57001 20772 57035
rect 20720 56992 20772 57001
rect 19156 56924 19208 56976
rect 19340 56924 19392 56976
rect 21456 56967 21508 56976
rect 21456 56933 21465 56967
rect 21465 56933 21499 56967
rect 21499 56933 21508 56967
rect 21456 56924 21508 56933
rect 14280 56856 14332 56908
rect 15476 56856 15528 56908
rect 16488 56856 16540 56908
rect 18328 56856 18380 56908
rect 17868 56831 17920 56840
rect 17868 56797 17877 56831
rect 17877 56797 17911 56831
rect 17911 56797 17920 56831
rect 17868 56788 17920 56797
rect 18696 56788 18748 56840
rect 18972 56788 19024 56840
rect 20444 56856 20496 56908
rect 21548 56856 21600 56908
rect 22836 57035 22888 57044
rect 22836 57001 22845 57035
rect 22845 57001 22879 57035
rect 22879 57001 22888 57035
rect 22836 56992 22888 57001
rect 26700 57035 26752 57044
rect 26700 57001 26709 57035
rect 26709 57001 26743 57035
rect 26743 57001 26752 57035
rect 26700 56992 26752 57001
rect 27344 56924 27396 56976
rect 22100 56856 22152 56908
rect 22928 56856 22980 56908
rect 23296 56899 23348 56908
rect 23296 56865 23305 56899
rect 23305 56865 23339 56899
rect 23339 56865 23348 56899
rect 23296 56856 23348 56865
rect 23480 56856 23532 56908
rect 24860 56856 24912 56908
rect 26516 56899 26568 56908
rect 26516 56865 26525 56899
rect 26525 56865 26559 56899
rect 26559 56865 26568 56899
rect 26516 56856 26568 56865
rect 27620 56856 27672 56908
rect 28264 56856 28316 56908
rect 28908 56924 28960 56976
rect 19432 56831 19484 56840
rect 19432 56797 19441 56831
rect 19441 56797 19475 56831
rect 19475 56797 19484 56831
rect 19432 56788 19484 56797
rect 22560 56788 22612 56840
rect 24400 56831 24452 56840
rect 24400 56797 24409 56831
rect 24409 56797 24443 56831
rect 24443 56797 24452 56831
rect 24400 56788 24452 56797
rect 24676 56788 24728 56840
rect 27528 56788 27580 56840
rect 28632 56788 28684 56840
rect 17500 56720 17552 56772
rect 18144 56720 18196 56772
rect 19340 56763 19392 56772
rect 19340 56729 19349 56763
rect 19349 56729 19383 56763
rect 19383 56729 19392 56763
rect 19340 56720 19392 56729
rect 21088 56720 21140 56772
rect 22008 56720 22060 56772
rect 28448 56720 28500 56772
rect 28908 56763 28960 56772
rect 28908 56729 28917 56763
rect 28917 56729 28951 56763
rect 28951 56729 28960 56763
rect 28908 56720 28960 56729
rect 14004 56695 14056 56704
rect 14004 56661 14013 56695
rect 14013 56661 14047 56695
rect 14047 56661 14056 56695
rect 14004 56652 14056 56661
rect 14464 56652 14516 56704
rect 15016 56652 15068 56704
rect 16488 56652 16540 56704
rect 19064 56652 19116 56704
rect 19524 56695 19576 56704
rect 19524 56661 19533 56695
rect 19533 56661 19567 56695
rect 19567 56661 19576 56695
rect 19524 56652 19576 56661
rect 22376 56652 22428 56704
rect 24768 56652 24820 56704
rect 25136 56695 25188 56704
rect 25136 56661 25145 56695
rect 25145 56661 25179 56695
rect 25179 56661 25188 56695
rect 25136 56652 25188 56661
rect 25504 56652 25556 56704
rect 25780 56652 25832 56704
rect 34612 56652 34664 56704
rect 35256 56695 35308 56704
rect 35256 56661 35265 56695
rect 35265 56661 35299 56695
rect 35299 56661 35308 56695
rect 35256 56652 35308 56661
rect 4246 56550 4298 56602
rect 4310 56550 4362 56602
rect 4374 56550 4426 56602
rect 4438 56550 4490 56602
rect 34966 56550 35018 56602
rect 35030 56550 35082 56602
rect 35094 56550 35146 56602
rect 35158 56550 35210 56602
rect 13268 56491 13320 56500
rect 13268 56457 13277 56491
rect 13277 56457 13311 56491
rect 13311 56457 13320 56491
rect 13268 56448 13320 56457
rect 15752 56491 15804 56500
rect 15752 56457 15761 56491
rect 15761 56457 15795 56491
rect 15795 56457 15804 56491
rect 15752 56448 15804 56457
rect 17500 56448 17552 56500
rect 17868 56491 17920 56500
rect 17868 56457 17877 56491
rect 17877 56457 17911 56491
rect 17911 56457 17920 56491
rect 17868 56448 17920 56457
rect 19432 56448 19484 56500
rect 19524 56448 19576 56500
rect 19984 56448 20036 56500
rect 21364 56491 21416 56500
rect 21364 56457 21373 56491
rect 21373 56457 21407 56491
rect 21407 56457 21416 56491
rect 21364 56448 21416 56457
rect 21456 56448 21508 56500
rect 23296 56491 23348 56500
rect 23296 56457 23305 56491
rect 23305 56457 23339 56491
rect 23339 56457 23348 56491
rect 23296 56448 23348 56457
rect 27344 56448 27396 56500
rect 27528 56491 27580 56500
rect 27528 56457 27537 56491
rect 27537 56457 27571 56491
rect 27571 56457 27580 56491
rect 27528 56448 27580 56457
rect 18052 56380 18104 56432
rect 18972 56380 19024 56432
rect 19156 56380 19208 56432
rect 19616 56380 19668 56432
rect 20260 56380 20312 56432
rect 14188 56355 14240 56364
rect 14188 56321 14197 56355
rect 14197 56321 14231 56355
rect 14231 56321 14240 56355
rect 14188 56312 14240 56321
rect 19340 56312 19392 56364
rect 20904 56380 20956 56432
rect 21916 56380 21968 56432
rect 21456 56355 21508 56364
rect 13268 56244 13320 56296
rect 14004 56244 14056 56296
rect 14280 56176 14332 56228
rect 13544 56151 13596 56160
rect 13544 56117 13553 56151
rect 13553 56117 13587 56151
rect 13587 56117 13596 56151
rect 13544 56108 13596 56117
rect 17224 56108 17276 56160
rect 18328 56176 18380 56228
rect 20168 56244 20220 56296
rect 21456 56321 21465 56355
rect 21465 56321 21499 56355
rect 21499 56321 21508 56355
rect 21456 56312 21508 56321
rect 24952 56312 25004 56364
rect 26056 56355 26108 56364
rect 26056 56321 26065 56355
rect 26065 56321 26099 56355
rect 26099 56321 26108 56355
rect 26056 56312 26108 56321
rect 28356 56355 28408 56364
rect 28356 56321 28365 56355
rect 28365 56321 28399 56355
rect 28399 56321 28408 56355
rect 28356 56312 28408 56321
rect 21916 56244 21968 56296
rect 22284 56244 22336 56296
rect 23664 56287 23716 56296
rect 23664 56253 23673 56287
rect 23673 56253 23707 56287
rect 23707 56253 23716 56287
rect 23664 56244 23716 56253
rect 25136 56287 25188 56296
rect 25136 56253 25145 56287
rect 25145 56253 25179 56287
rect 25179 56253 25188 56287
rect 25136 56244 25188 56253
rect 25320 56244 25372 56296
rect 25780 56244 25832 56296
rect 27804 56287 27856 56296
rect 27804 56253 27813 56287
rect 27813 56253 27847 56287
rect 27847 56253 27856 56287
rect 27804 56244 27856 56253
rect 20904 56219 20956 56228
rect 20904 56185 20913 56219
rect 20913 56185 20947 56219
rect 20947 56185 20956 56219
rect 20904 56176 20956 56185
rect 21364 56176 21416 56228
rect 26332 56176 26384 56228
rect 17592 56108 17644 56160
rect 19340 56151 19392 56160
rect 19340 56117 19349 56151
rect 19349 56117 19383 56151
rect 19383 56117 19392 56151
rect 19340 56108 19392 56117
rect 19432 56108 19484 56160
rect 22100 56108 22152 56160
rect 22560 56151 22612 56160
rect 22560 56117 22569 56151
rect 22569 56117 22603 56151
rect 22603 56117 22612 56151
rect 22560 56108 22612 56117
rect 23480 56108 23532 56160
rect 23848 56151 23900 56160
rect 23848 56117 23857 56151
rect 23857 56117 23891 56151
rect 23891 56117 23900 56151
rect 23848 56108 23900 56117
rect 24492 56151 24544 56160
rect 24492 56117 24501 56151
rect 24501 56117 24535 56151
rect 24535 56117 24544 56151
rect 24492 56108 24544 56117
rect 24768 56108 24820 56160
rect 26516 56151 26568 56160
rect 26516 56117 26525 56151
rect 26525 56117 26559 56151
rect 26559 56117 26568 56151
rect 26516 56108 26568 56117
rect 28356 56108 28408 56160
rect 19606 56006 19658 56058
rect 19670 56006 19722 56058
rect 19734 56006 19786 56058
rect 19798 56006 19850 56058
rect 14372 55947 14424 55956
rect 14372 55913 14381 55947
rect 14381 55913 14415 55947
rect 14415 55913 14424 55947
rect 14372 55904 14424 55913
rect 17500 55947 17552 55956
rect 17500 55913 17509 55947
rect 17509 55913 17543 55947
rect 17543 55913 17552 55947
rect 17500 55904 17552 55913
rect 18696 55947 18748 55956
rect 18696 55913 18705 55947
rect 18705 55913 18739 55947
rect 18739 55913 18748 55947
rect 18696 55904 18748 55913
rect 19064 55947 19116 55956
rect 19064 55913 19073 55947
rect 19073 55913 19107 55947
rect 19107 55913 19116 55947
rect 19064 55904 19116 55913
rect 20260 55947 20312 55956
rect 20260 55913 20269 55947
rect 20269 55913 20303 55947
rect 20303 55913 20312 55947
rect 20260 55904 20312 55913
rect 22836 55904 22888 55956
rect 24492 55904 24544 55956
rect 27068 55904 27120 55956
rect 28540 55947 28592 55956
rect 28540 55913 28549 55947
rect 28549 55913 28583 55947
rect 28583 55913 28592 55947
rect 28540 55904 28592 55913
rect 12716 55836 12768 55888
rect 15016 55836 15068 55888
rect 19984 55879 20036 55888
rect 19984 55845 19993 55879
rect 19993 55845 20027 55879
rect 20027 55845 20036 55879
rect 19984 55836 20036 55845
rect 12256 55768 12308 55820
rect 13176 55811 13228 55820
rect 13176 55777 13185 55811
rect 13185 55777 13219 55811
rect 13219 55777 13228 55811
rect 13176 55768 13228 55777
rect 14832 55768 14884 55820
rect 16856 55811 16908 55820
rect 16856 55777 16865 55811
rect 16865 55777 16899 55811
rect 16899 55777 16908 55811
rect 16856 55768 16908 55777
rect 18328 55811 18380 55820
rect 18328 55777 18337 55811
rect 18337 55777 18371 55811
rect 18371 55777 18380 55811
rect 18328 55768 18380 55777
rect 19064 55768 19116 55820
rect 20720 55768 20772 55820
rect 21088 55811 21140 55820
rect 21088 55777 21097 55811
rect 21097 55777 21131 55811
rect 21131 55777 21140 55811
rect 21088 55768 21140 55777
rect 22928 55811 22980 55820
rect 22928 55777 22937 55811
rect 22937 55777 22971 55811
rect 22971 55777 22980 55811
rect 22928 55768 22980 55777
rect 23112 55768 23164 55820
rect 23940 55768 23992 55820
rect 24952 55811 25004 55820
rect 24952 55777 24961 55811
rect 24961 55777 24995 55811
rect 24995 55777 25004 55811
rect 24952 55768 25004 55777
rect 13636 55700 13688 55752
rect 15476 55743 15528 55752
rect 15476 55709 15485 55743
rect 15485 55709 15519 55743
rect 15519 55709 15528 55743
rect 15476 55700 15528 55709
rect 16948 55700 17000 55752
rect 17224 55743 17276 55752
rect 17224 55709 17233 55743
rect 17233 55709 17267 55743
rect 17267 55709 17276 55743
rect 17224 55700 17276 55709
rect 18420 55743 18472 55752
rect 18420 55709 18429 55743
rect 18429 55709 18463 55743
rect 18463 55709 18472 55743
rect 18420 55700 18472 55709
rect 12440 55564 12492 55616
rect 13452 55564 13504 55616
rect 13912 55564 13964 55616
rect 15016 55564 15068 55616
rect 15660 55632 15712 55684
rect 16028 55675 16080 55684
rect 16028 55641 16037 55675
rect 16037 55641 16071 55675
rect 16071 55641 16080 55675
rect 16028 55632 16080 55641
rect 19156 55632 19208 55684
rect 19340 55700 19392 55752
rect 21180 55700 21232 55752
rect 22468 55700 22520 55752
rect 16488 55564 16540 55616
rect 20260 55632 20312 55684
rect 25596 55768 25648 55820
rect 28264 55811 28316 55820
rect 26516 55700 26568 55752
rect 28264 55777 28273 55811
rect 28273 55777 28307 55811
rect 28307 55777 28316 55811
rect 28264 55768 28316 55777
rect 33232 55768 33284 55820
rect 34428 55768 34480 55820
rect 33600 55700 33652 55752
rect 34612 55700 34664 55752
rect 19524 55607 19576 55616
rect 19524 55573 19533 55607
rect 19533 55573 19567 55607
rect 19567 55573 19576 55607
rect 20720 55607 20772 55616
rect 19524 55564 19576 55573
rect 20720 55573 20729 55607
rect 20729 55573 20763 55607
rect 20763 55573 20772 55607
rect 20720 55564 20772 55573
rect 20996 55564 21048 55616
rect 22560 55564 22612 55616
rect 23296 55564 23348 55616
rect 23664 55607 23716 55616
rect 23664 55573 23673 55607
rect 23673 55573 23707 55607
rect 23707 55573 23716 55607
rect 23664 55564 23716 55573
rect 24860 55564 24912 55616
rect 25780 55564 25832 55616
rect 27804 55564 27856 55616
rect 32680 55564 32732 55616
rect 4246 55462 4298 55514
rect 4310 55462 4362 55514
rect 4374 55462 4426 55514
rect 4438 55462 4490 55514
rect 34966 55462 35018 55514
rect 35030 55462 35082 55514
rect 35094 55462 35146 55514
rect 35158 55462 35210 55514
rect 12256 55403 12308 55412
rect 12256 55369 12265 55403
rect 12265 55369 12299 55403
rect 12299 55369 12308 55403
rect 12256 55360 12308 55369
rect 12716 55403 12768 55412
rect 12716 55369 12725 55403
rect 12725 55369 12759 55403
rect 12759 55369 12768 55403
rect 12716 55360 12768 55369
rect 13912 55360 13964 55412
rect 14648 55360 14700 55412
rect 15476 55360 15528 55412
rect 16764 55360 16816 55412
rect 16948 55360 17000 55412
rect 20168 55360 20220 55412
rect 22836 55360 22888 55412
rect 24952 55360 25004 55412
rect 33232 55403 33284 55412
rect 33232 55369 33241 55403
rect 33241 55369 33275 55403
rect 33275 55369 33284 55403
rect 33232 55360 33284 55369
rect 12348 55224 12400 55276
rect 12532 55224 12584 55276
rect 15016 55335 15068 55344
rect 15016 55301 15040 55335
rect 15040 55301 15068 55335
rect 15016 55292 15068 55301
rect 13176 55224 13228 55276
rect 14464 55224 14516 55276
rect 14188 55156 14240 55208
rect 15108 55156 15160 55208
rect 15292 55156 15344 55208
rect 15936 55156 15988 55208
rect 24216 55292 24268 55344
rect 26516 55292 26568 55344
rect 17868 55224 17920 55276
rect 20260 55224 20312 55276
rect 20720 55224 20772 55276
rect 21088 55224 21140 55276
rect 26240 55224 26292 55276
rect 19064 55156 19116 55208
rect 19616 55199 19668 55208
rect 19616 55165 19625 55199
rect 19625 55165 19659 55199
rect 19659 55165 19668 55199
rect 19616 55156 19668 55165
rect 21180 55199 21232 55208
rect 21180 55165 21189 55199
rect 21189 55165 21223 55199
rect 21223 55165 21232 55199
rect 21180 55156 21232 55165
rect 23664 55199 23716 55208
rect 14832 55131 14884 55140
rect 14832 55097 14841 55131
rect 14841 55097 14875 55131
rect 14875 55097 14884 55131
rect 14832 55088 14884 55097
rect 16120 55088 16172 55140
rect 18052 55131 18104 55140
rect 15200 55020 15252 55072
rect 18052 55097 18061 55131
rect 18061 55097 18095 55131
rect 18095 55097 18104 55131
rect 18052 55088 18104 55097
rect 21088 55088 21140 55140
rect 23664 55165 23673 55199
rect 23673 55165 23707 55199
rect 23707 55165 23716 55199
rect 23664 55156 23716 55165
rect 23848 55156 23900 55208
rect 24492 55199 24544 55208
rect 24492 55165 24501 55199
rect 24501 55165 24535 55199
rect 24535 55165 24544 55199
rect 24492 55156 24544 55165
rect 28264 55224 28316 55276
rect 31576 55267 31628 55276
rect 31576 55233 31585 55267
rect 31585 55233 31619 55267
rect 31619 55233 31628 55267
rect 31576 55224 31628 55233
rect 27988 55199 28040 55208
rect 26608 55088 26660 55140
rect 27988 55165 27997 55199
rect 27997 55165 28031 55199
rect 28031 55165 28040 55199
rect 27988 55156 28040 55165
rect 31760 55156 31812 55208
rect 33600 55267 33652 55276
rect 33600 55233 33609 55267
rect 33609 55233 33643 55267
rect 33643 55233 33652 55267
rect 33600 55224 33652 55233
rect 32680 55199 32732 55208
rect 32680 55165 32689 55199
rect 32689 55165 32723 55199
rect 32723 55165 32732 55199
rect 32680 55156 32732 55165
rect 31944 55131 31996 55140
rect 31944 55097 31953 55131
rect 31953 55097 31987 55131
rect 31987 55097 31996 55131
rect 31944 55088 31996 55097
rect 16580 55063 16632 55072
rect 16580 55029 16589 55063
rect 16589 55029 16623 55063
rect 16623 55029 16632 55063
rect 16580 55020 16632 55029
rect 17500 55063 17552 55072
rect 17500 55029 17509 55063
rect 17509 55029 17543 55063
rect 17543 55029 17552 55063
rect 17500 55020 17552 55029
rect 19340 55063 19392 55072
rect 19340 55029 19349 55063
rect 19349 55029 19383 55063
rect 19383 55029 19392 55063
rect 19340 55020 19392 55029
rect 19432 55020 19484 55072
rect 20444 55063 20496 55072
rect 20444 55029 20453 55063
rect 20453 55029 20487 55063
rect 20487 55029 20496 55063
rect 20444 55020 20496 55029
rect 21640 55020 21692 55072
rect 23940 55020 23992 55072
rect 26332 55020 26384 55072
rect 26792 55020 26844 55072
rect 19606 54918 19658 54970
rect 19670 54918 19722 54970
rect 19734 54918 19786 54970
rect 19798 54918 19850 54970
rect 13636 54859 13688 54868
rect 13636 54825 13645 54859
rect 13645 54825 13679 54859
rect 13679 54825 13688 54859
rect 13636 54816 13688 54825
rect 15476 54816 15528 54868
rect 15660 54816 15712 54868
rect 16580 54816 16632 54868
rect 17592 54859 17644 54868
rect 17592 54825 17601 54859
rect 17601 54825 17635 54859
rect 17635 54825 17644 54859
rect 17592 54816 17644 54825
rect 19064 54816 19116 54868
rect 21916 54816 21968 54868
rect 23848 54816 23900 54868
rect 23940 54859 23992 54868
rect 23940 54825 23949 54859
rect 23949 54825 23983 54859
rect 23983 54825 23992 54859
rect 23940 54816 23992 54825
rect 14832 54748 14884 54800
rect 18052 54748 18104 54800
rect 13176 54723 13228 54732
rect 13176 54689 13185 54723
rect 13185 54689 13219 54723
rect 13219 54689 13228 54723
rect 13176 54680 13228 54689
rect 13360 54680 13412 54732
rect 14188 54723 14240 54732
rect 14188 54689 14197 54723
rect 14197 54689 14231 54723
rect 14231 54689 14240 54723
rect 14188 54680 14240 54689
rect 17224 54680 17276 54732
rect 19248 54748 19300 54800
rect 19432 54791 19484 54800
rect 19432 54757 19441 54791
rect 19441 54757 19475 54791
rect 19475 54757 19484 54791
rect 19432 54748 19484 54757
rect 20628 54748 20680 54800
rect 19340 54723 19392 54732
rect 19340 54689 19349 54723
rect 19349 54689 19383 54723
rect 19383 54689 19392 54723
rect 19340 54680 19392 54689
rect 19616 54680 19668 54732
rect 20168 54680 20220 54732
rect 21456 54680 21508 54732
rect 21640 54680 21692 54732
rect 22836 54748 22888 54800
rect 24308 54748 24360 54800
rect 25136 54748 25188 54800
rect 22744 54723 22796 54732
rect 22744 54689 22753 54723
rect 22753 54689 22787 54723
rect 22787 54689 22796 54723
rect 22744 54680 22796 54689
rect 23940 54680 23992 54732
rect 25044 54723 25096 54732
rect 25044 54689 25053 54723
rect 25053 54689 25087 54723
rect 25087 54689 25096 54723
rect 25044 54680 25096 54689
rect 26240 54748 26292 54800
rect 25964 54680 26016 54732
rect 28080 54816 28132 54868
rect 29000 54680 29052 54732
rect 15292 54612 15344 54664
rect 16856 54612 16908 54664
rect 18788 54612 18840 54664
rect 22284 54612 22336 54664
rect 22468 54612 22520 54664
rect 23112 54655 23164 54664
rect 23112 54621 23121 54655
rect 23121 54621 23155 54655
rect 23155 54621 23164 54655
rect 23112 54612 23164 54621
rect 25504 54655 25556 54664
rect 14372 54587 14424 54596
rect 14372 54553 14381 54587
rect 14381 54553 14415 54587
rect 14415 54553 14424 54587
rect 14372 54544 14424 54553
rect 16028 54587 16080 54596
rect 16028 54553 16037 54587
rect 16037 54553 16071 54587
rect 16071 54553 16080 54587
rect 16028 54544 16080 54553
rect 16580 54544 16632 54596
rect 17500 54544 17552 54596
rect 18512 54544 18564 54596
rect 20260 54544 20312 54596
rect 25504 54621 25513 54655
rect 25513 54621 25547 54655
rect 25547 54621 25556 54655
rect 25504 54612 25556 54621
rect 27528 54612 27580 54664
rect 28816 54612 28868 54664
rect 25412 54544 25464 54596
rect 13360 54519 13412 54528
rect 13360 54485 13369 54519
rect 13369 54485 13403 54519
rect 13403 54485 13412 54519
rect 13360 54476 13412 54485
rect 15016 54476 15068 54528
rect 15844 54476 15896 54528
rect 16488 54476 16540 54528
rect 20720 54476 20772 54528
rect 21088 54519 21140 54528
rect 21088 54485 21097 54519
rect 21097 54485 21131 54519
rect 21131 54485 21140 54519
rect 21088 54476 21140 54485
rect 24492 54519 24544 54528
rect 24492 54485 24501 54519
rect 24501 54485 24535 54519
rect 24535 54485 24544 54519
rect 24492 54476 24544 54485
rect 25780 54476 25832 54528
rect 26884 54476 26936 54528
rect 29092 54476 29144 54528
rect 31760 54519 31812 54528
rect 31760 54485 31769 54519
rect 31769 54485 31803 54519
rect 31803 54485 31812 54519
rect 31760 54476 31812 54485
rect 4246 54374 4298 54426
rect 4310 54374 4362 54426
rect 4374 54374 4426 54426
rect 4438 54374 4490 54426
rect 34966 54374 35018 54426
rect 35030 54374 35082 54426
rect 35094 54374 35146 54426
rect 35158 54374 35210 54426
rect 13176 54315 13228 54324
rect 13176 54281 13185 54315
rect 13185 54281 13219 54315
rect 13219 54281 13228 54315
rect 13176 54272 13228 54281
rect 14188 54272 14240 54324
rect 16856 54315 16908 54324
rect 16856 54281 16865 54315
rect 16865 54281 16899 54315
rect 16899 54281 16908 54315
rect 16856 54272 16908 54281
rect 17592 54315 17644 54324
rect 17592 54281 17601 54315
rect 17601 54281 17635 54315
rect 17635 54281 17644 54315
rect 17592 54272 17644 54281
rect 18052 54272 18104 54324
rect 19340 54272 19392 54324
rect 22008 54272 22060 54324
rect 22192 54272 22244 54324
rect 15844 54204 15896 54256
rect 17776 54204 17828 54256
rect 19616 54247 19668 54256
rect 19616 54213 19625 54247
rect 19625 54213 19659 54247
rect 19659 54213 19668 54247
rect 19616 54204 19668 54213
rect 14004 54136 14056 54188
rect 14464 54136 14516 54188
rect 17224 54136 17276 54188
rect 19432 54136 19484 54188
rect 20628 54136 20680 54188
rect 21180 54136 21232 54188
rect 21456 54136 21508 54188
rect 22376 54136 22428 54188
rect 12440 54068 12492 54120
rect 14372 54068 14424 54120
rect 14832 54000 14884 54052
rect 14740 53975 14792 53984
rect 14740 53941 14749 53975
rect 14749 53941 14783 53975
rect 14783 53941 14792 53975
rect 18604 54111 18656 54120
rect 18604 54077 18613 54111
rect 18613 54077 18647 54111
rect 18647 54077 18656 54111
rect 18604 54068 18656 54077
rect 18788 54111 18840 54120
rect 18788 54077 18797 54111
rect 18797 54077 18831 54111
rect 18831 54077 18840 54111
rect 18788 54068 18840 54077
rect 21640 54068 21692 54120
rect 22008 54068 22060 54120
rect 22560 54111 22612 54120
rect 14740 53932 14792 53941
rect 19616 54000 19668 54052
rect 20076 54000 20128 54052
rect 20720 54000 20772 54052
rect 21088 54000 21140 54052
rect 19340 53932 19392 53984
rect 20260 53932 20312 53984
rect 20444 53975 20496 53984
rect 20444 53941 20453 53975
rect 20453 53941 20487 53975
rect 20487 53941 20496 53975
rect 21916 54000 21968 54052
rect 22560 54077 22569 54111
rect 22569 54077 22603 54111
rect 22603 54077 22612 54111
rect 23848 54272 23900 54324
rect 24308 54315 24360 54324
rect 24308 54281 24317 54315
rect 24317 54281 24351 54315
rect 24351 54281 24360 54315
rect 24308 54272 24360 54281
rect 27896 54315 27948 54324
rect 27896 54281 27905 54315
rect 27905 54281 27939 54315
rect 27939 54281 27948 54315
rect 27896 54272 27948 54281
rect 28816 54272 28868 54324
rect 29000 54272 29052 54324
rect 29552 54272 29604 54324
rect 30288 54272 30340 54324
rect 23940 54204 23992 54256
rect 24768 54204 24820 54256
rect 25412 54136 25464 54188
rect 25596 54179 25648 54188
rect 25596 54145 25605 54179
rect 25605 54145 25639 54179
rect 25639 54145 25648 54179
rect 25596 54136 25648 54145
rect 26240 54136 26292 54188
rect 22560 54068 22612 54077
rect 24952 54068 25004 54120
rect 25044 54068 25096 54120
rect 25504 54111 25556 54120
rect 25504 54077 25513 54111
rect 25513 54077 25547 54111
rect 25547 54077 25556 54111
rect 25504 54068 25556 54077
rect 26700 54068 26752 54120
rect 26792 54111 26844 54120
rect 26792 54077 26801 54111
rect 26801 54077 26835 54111
rect 26835 54077 26844 54111
rect 26792 54068 26844 54077
rect 27896 54068 27948 54120
rect 22376 54000 22428 54052
rect 24492 54043 24544 54052
rect 24492 54009 24501 54043
rect 24501 54009 24535 54043
rect 24535 54009 24544 54043
rect 24492 54000 24544 54009
rect 26240 54000 26292 54052
rect 26884 54043 26936 54052
rect 20444 53932 20496 53941
rect 22836 53932 22888 53984
rect 25964 53975 26016 53984
rect 25964 53941 25973 53975
rect 25973 53941 26007 53975
rect 26007 53941 26016 53975
rect 25964 53932 26016 53941
rect 26332 53975 26384 53984
rect 26332 53941 26341 53975
rect 26341 53941 26375 53975
rect 26375 53941 26384 53975
rect 26332 53932 26384 53941
rect 26884 54009 26893 54043
rect 26893 54009 26927 54043
rect 26927 54009 26936 54043
rect 26884 54000 26936 54009
rect 19606 53830 19658 53882
rect 19670 53830 19722 53882
rect 19734 53830 19786 53882
rect 19798 53830 19850 53882
rect 14464 53728 14516 53780
rect 14648 53728 14700 53780
rect 16396 53728 16448 53780
rect 17592 53728 17644 53780
rect 19340 53728 19392 53780
rect 19984 53728 20036 53780
rect 20444 53728 20496 53780
rect 20628 53771 20680 53780
rect 20628 53737 20637 53771
rect 20637 53737 20671 53771
rect 20671 53737 20680 53771
rect 20628 53728 20680 53737
rect 22376 53728 22428 53780
rect 22928 53728 22980 53780
rect 15108 53703 15160 53712
rect 15108 53669 15117 53703
rect 15117 53669 15151 53703
rect 15151 53669 15160 53703
rect 15108 53660 15160 53669
rect 15660 53660 15712 53712
rect 15936 53703 15988 53712
rect 15936 53669 15945 53703
rect 15945 53669 15979 53703
rect 15979 53669 15988 53703
rect 15936 53660 15988 53669
rect 16304 53703 16356 53712
rect 16304 53669 16313 53703
rect 16313 53669 16347 53703
rect 16347 53669 16356 53703
rect 16304 53660 16356 53669
rect 16580 53703 16632 53712
rect 16580 53669 16589 53703
rect 16589 53669 16623 53703
rect 16623 53669 16632 53703
rect 16580 53660 16632 53669
rect 16948 53660 17000 53712
rect 14280 53592 14332 53644
rect 14372 53592 14424 53644
rect 16764 53592 16816 53644
rect 16856 53592 16908 53644
rect 17500 53635 17552 53644
rect 17500 53601 17509 53635
rect 17509 53601 17543 53635
rect 17543 53601 17552 53635
rect 17500 53592 17552 53601
rect 18604 53660 18656 53712
rect 19616 53703 19668 53712
rect 19616 53669 19625 53703
rect 19625 53669 19659 53703
rect 19659 53669 19668 53703
rect 19616 53660 19668 53669
rect 20720 53660 20772 53712
rect 21548 53703 21600 53712
rect 21548 53669 21557 53703
rect 21557 53669 21591 53703
rect 21591 53669 21600 53703
rect 21548 53660 21600 53669
rect 23572 53660 23624 53712
rect 18972 53592 19024 53644
rect 21640 53635 21692 53644
rect 21640 53601 21649 53635
rect 21649 53601 21683 53635
rect 21683 53601 21692 53635
rect 21640 53592 21692 53601
rect 22376 53592 22428 53644
rect 23848 53592 23900 53644
rect 24124 53635 24176 53644
rect 24124 53601 24133 53635
rect 24133 53601 24167 53635
rect 24167 53601 24176 53635
rect 24124 53592 24176 53601
rect 24492 53635 24544 53644
rect 24492 53601 24501 53635
rect 24501 53601 24535 53635
rect 24535 53601 24544 53635
rect 24492 53592 24544 53601
rect 24676 53592 24728 53644
rect 27344 53635 27396 53644
rect 27344 53601 27353 53635
rect 27353 53601 27387 53635
rect 27387 53601 27396 53635
rect 27344 53592 27396 53601
rect 27528 53635 27580 53644
rect 27528 53601 27537 53635
rect 27537 53601 27571 53635
rect 27571 53601 27580 53635
rect 27528 53592 27580 53601
rect 28172 53635 28224 53644
rect 28172 53601 28181 53635
rect 28181 53601 28215 53635
rect 28215 53601 28224 53635
rect 28172 53592 28224 53601
rect 19432 53524 19484 53576
rect 20352 53524 20404 53576
rect 21364 53524 21416 53576
rect 14924 53456 14976 53508
rect 17960 53499 18012 53508
rect 17960 53465 17969 53499
rect 17969 53465 18003 53499
rect 18003 53465 18012 53499
rect 17960 53456 18012 53465
rect 19064 53499 19116 53508
rect 14740 53431 14792 53440
rect 14740 53397 14749 53431
rect 14749 53397 14783 53431
rect 14783 53397 14792 53431
rect 14740 53388 14792 53397
rect 15660 53388 15712 53440
rect 19064 53465 19073 53499
rect 19073 53465 19107 53499
rect 19107 53465 19116 53499
rect 19064 53456 19116 53465
rect 18604 53431 18656 53440
rect 18604 53397 18613 53431
rect 18613 53397 18647 53431
rect 18647 53397 18656 53431
rect 18604 53388 18656 53397
rect 23296 53524 23348 53576
rect 26332 53524 26384 53576
rect 23848 53456 23900 53508
rect 24400 53499 24452 53508
rect 24400 53465 24409 53499
rect 24409 53465 24443 53499
rect 24443 53465 24452 53499
rect 24400 53456 24452 53465
rect 25228 53456 25280 53508
rect 27160 53499 27212 53508
rect 27160 53465 27169 53499
rect 27169 53465 27203 53499
rect 27203 53465 27212 53499
rect 27160 53456 27212 53465
rect 23296 53388 23348 53440
rect 24952 53431 25004 53440
rect 24952 53397 24961 53431
rect 24961 53397 24995 53431
rect 24995 53397 25004 53431
rect 24952 53388 25004 53397
rect 25504 53388 25556 53440
rect 26240 53431 26292 53440
rect 26240 53397 26249 53431
rect 26249 53397 26283 53431
rect 26283 53397 26292 53431
rect 26240 53388 26292 53397
rect 26700 53431 26752 53440
rect 26700 53397 26709 53431
rect 26709 53397 26743 53431
rect 26743 53397 26752 53431
rect 26700 53388 26752 53397
rect 4246 53286 4298 53338
rect 4310 53286 4362 53338
rect 4374 53286 4426 53338
rect 4438 53286 4490 53338
rect 34966 53286 35018 53338
rect 35030 53286 35082 53338
rect 35094 53286 35146 53338
rect 35158 53286 35210 53338
rect 13820 53184 13872 53236
rect 15844 53184 15896 53236
rect 16580 53184 16632 53236
rect 16856 53184 16908 53236
rect 17408 53184 17460 53236
rect 18604 53184 18656 53236
rect 19524 53227 19576 53236
rect 19524 53193 19533 53227
rect 19533 53193 19567 53227
rect 19567 53193 19576 53227
rect 19524 53184 19576 53193
rect 22560 53184 22612 53236
rect 23480 53227 23532 53236
rect 23480 53193 23489 53227
rect 23489 53193 23523 53227
rect 23523 53193 23532 53227
rect 23480 53184 23532 53193
rect 24768 53227 24820 53236
rect 24768 53193 24777 53227
rect 24777 53193 24811 53227
rect 24811 53193 24820 53227
rect 24768 53184 24820 53193
rect 29552 53227 29604 53236
rect 29552 53193 29561 53227
rect 29561 53193 29595 53227
rect 29595 53193 29604 53227
rect 29552 53184 29604 53193
rect 14280 53159 14332 53168
rect 14280 53125 14289 53159
rect 14289 53125 14323 53159
rect 14323 53125 14332 53159
rect 14280 53116 14332 53125
rect 14648 53116 14700 53168
rect 18236 53116 18288 53168
rect 19984 53159 20036 53168
rect 19984 53125 19993 53159
rect 19993 53125 20027 53159
rect 20027 53125 20036 53159
rect 19984 53116 20036 53125
rect 20260 53116 20312 53168
rect 21824 53116 21876 53168
rect 15660 53048 15712 53100
rect 16764 53091 16816 53100
rect 16764 53057 16773 53091
rect 16773 53057 16807 53091
rect 16807 53057 16816 53091
rect 16764 53048 16816 53057
rect 15292 53023 15344 53032
rect 15292 52989 15301 53023
rect 15301 52989 15335 53023
rect 15335 52989 15344 53023
rect 15292 52980 15344 52989
rect 15936 52980 15988 53032
rect 16396 53023 16448 53032
rect 16396 52989 16405 53023
rect 16405 52989 16439 53023
rect 16439 52989 16448 53023
rect 16396 52980 16448 52989
rect 17776 52980 17828 53032
rect 18144 53023 18196 53032
rect 18144 52989 18153 53023
rect 18153 52989 18187 53023
rect 18187 52989 18196 53023
rect 18144 52980 18196 52989
rect 18512 53023 18564 53032
rect 18512 52989 18521 53023
rect 18521 52989 18555 53023
rect 18555 52989 18564 53023
rect 18512 52980 18564 52989
rect 18972 53023 19024 53032
rect 18972 52989 18981 53023
rect 18981 52989 19015 53023
rect 19015 52989 19024 53023
rect 18972 52980 19024 52989
rect 20720 53048 20772 53100
rect 23756 53159 23808 53168
rect 23756 53125 23765 53159
rect 23765 53125 23799 53159
rect 23799 53125 23808 53159
rect 23756 53116 23808 53125
rect 23940 53116 23992 53168
rect 20536 52980 20588 53032
rect 21364 53023 21416 53032
rect 21364 52989 21373 53023
rect 21373 52989 21407 53023
rect 21407 52989 21416 53023
rect 21364 52980 21416 52989
rect 22284 53023 22336 53032
rect 15476 52844 15528 52896
rect 22284 52989 22293 53023
rect 22293 52989 22327 53023
rect 22327 52989 22336 53023
rect 22284 52980 22336 52989
rect 25596 53048 25648 53100
rect 22376 52912 22428 52964
rect 17868 52844 17920 52896
rect 18788 52844 18840 52896
rect 22928 52844 22980 52896
rect 25228 53023 25280 53032
rect 25228 52989 25237 53023
rect 25237 52989 25271 53023
rect 25271 52989 25280 53023
rect 25228 52980 25280 52989
rect 23940 52844 23992 52896
rect 24768 52844 24820 52896
rect 26240 52980 26292 53032
rect 26516 52980 26568 53032
rect 27160 52980 27212 53032
rect 25780 52912 25832 52964
rect 26792 52912 26844 52964
rect 26240 52844 26292 52896
rect 26332 52844 26384 52896
rect 27160 52887 27212 52896
rect 27160 52853 27169 52887
rect 27169 52853 27203 52887
rect 27203 52853 27212 52887
rect 27160 52844 27212 52853
rect 27344 52844 27396 52896
rect 19606 52742 19658 52794
rect 19670 52742 19722 52794
rect 19734 52742 19786 52794
rect 19798 52742 19850 52794
rect 14740 52683 14792 52692
rect 14740 52649 14749 52683
rect 14749 52649 14783 52683
rect 14783 52649 14792 52683
rect 14740 52640 14792 52649
rect 16580 52640 16632 52692
rect 18328 52683 18380 52692
rect 18328 52649 18337 52683
rect 18337 52649 18371 52683
rect 18371 52649 18380 52683
rect 18328 52640 18380 52649
rect 20628 52640 20680 52692
rect 21640 52683 21692 52692
rect 21640 52649 21649 52683
rect 21649 52649 21683 52683
rect 21683 52649 21692 52683
rect 21640 52640 21692 52649
rect 23112 52640 23164 52692
rect 23756 52683 23808 52692
rect 15476 52572 15528 52624
rect 16212 52615 16264 52624
rect 16212 52581 16221 52615
rect 16221 52581 16255 52615
rect 16255 52581 16264 52615
rect 16212 52572 16264 52581
rect 16948 52572 17000 52624
rect 20444 52572 20496 52624
rect 20996 52572 21048 52624
rect 22100 52572 22152 52624
rect 9956 52504 10008 52556
rect 10784 52504 10836 52556
rect 15660 52547 15712 52556
rect 15660 52513 15669 52547
rect 15669 52513 15703 52547
rect 15703 52513 15712 52547
rect 15660 52504 15712 52513
rect 15752 52547 15804 52556
rect 15752 52513 15761 52547
rect 15761 52513 15795 52547
rect 15795 52513 15804 52547
rect 15752 52504 15804 52513
rect 11888 52479 11940 52488
rect 11888 52445 11897 52479
rect 11897 52445 11931 52479
rect 11931 52445 11940 52479
rect 11888 52436 11940 52445
rect 15200 52436 15252 52488
rect 16764 52504 16816 52556
rect 17960 52504 18012 52556
rect 18696 52504 18748 52556
rect 19432 52547 19484 52556
rect 19432 52513 19441 52547
rect 19441 52513 19475 52547
rect 19475 52513 19484 52547
rect 19432 52504 19484 52513
rect 19892 52504 19944 52556
rect 20536 52504 20588 52556
rect 20904 52547 20956 52556
rect 20904 52513 20913 52547
rect 20913 52513 20947 52547
rect 20947 52513 20956 52547
rect 20904 52504 20956 52513
rect 22192 52504 22244 52556
rect 17592 52479 17644 52488
rect 17592 52445 17601 52479
rect 17601 52445 17635 52479
rect 17635 52445 17644 52479
rect 17592 52436 17644 52445
rect 17776 52436 17828 52488
rect 18972 52368 19024 52420
rect 19984 52436 20036 52488
rect 20260 52436 20312 52488
rect 20720 52436 20772 52488
rect 23756 52649 23765 52683
rect 23765 52649 23799 52683
rect 23799 52649 23808 52683
rect 23756 52640 23808 52649
rect 23940 52640 23992 52692
rect 25780 52640 25832 52692
rect 29092 52683 29144 52692
rect 24952 52615 25004 52624
rect 24952 52581 24961 52615
rect 24961 52581 24995 52615
rect 24995 52581 25004 52615
rect 24952 52572 25004 52581
rect 27436 52615 27488 52624
rect 27436 52581 27445 52615
rect 27445 52581 27479 52615
rect 27479 52581 27488 52615
rect 27436 52572 27488 52581
rect 24676 52547 24728 52556
rect 24676 52513 24685 52547
rect 24685 52513 24719 52547
rect 24719 52513 24728 52547
rect 24676 52504 24728 52513
rect 25780 52504 25832 52556
rect 27528 52504 27580 52556
rect 29092 52649 29101 52683
rect 29101 52649 29135 52683
rect 29135 52649 29144 52683
rect 29092 52640 29144 52649
rect 29460 52547 29512 52556
rect 29460 52513 29469 52547
rect 29469 52513 29503 52547
rect 29503 52513 29512 52547
rect 29460 52504 29512 52513
rect 29552 52504 29604 52556
rect 24492 52436 24544 52488
rect 19340 52368 19392 52420
rect 16948 52300 17000 52352
rect 18144 52300 18196 52352
rect 18788 52300 18840 52352
rect 22100 52343 22152 52352
rect 22100 52309 22109 52343
rect 22109 52309 22143 52343
rect 22143 52309 22152 52343
rect 22836 52368 22888 52420
rect 27160 52436 27212 52488
rect 28264 52479 28316 52488
rect 24952 52368 25004 52420
rect 28264 52445 28273 52479
rect 28273 52445 28307 52479
rect 28307 52445 28316 52479
rect 28264 52436 28316 52445
rect 30288 52436 30340 52488
rect 30748 52479 30800 52488
rect 30748 52445 30757 52479
rect 30757 52445 30791 52479
rect 30791 52445 30800 52479
rect 30748 52436 30800 52445
rect 34704 52436 34756 52488
rect 35808 52436 35860 52488
rect 28356 52368 28408 52420
rect 22100 52300 22152 52309
rect 26240 52300 26292 52352
rect 26792 52343 26844 52352
rect 26792 52309 26801 52343
rect 26801 52309 26835 52343
rect 26835 52309 26844 52343
rect 26792 52300 26844 52309
rect 26884 52300 26936 52352
rect 4246 52198 4298 52250
rect 4310 52198 4362 52250
rect 4374 52198 4426 52250
rect 4438 52198 4490 52250
rect 34966 52198 35018 52250
rect 35030 52198 35082 52250
rect 35094 52198 35146 52250
rect 35158 52198 35210 52250
rect 9956 52096 10008 52148
rect 10784 52096 10836 52148
rect 15200 52096 15252 52148
rect 15660 52096 15712 52148
rect 18696 52096 18748 52148
rect 19064 52139 19116 52148
rect 19064 52105 19073 52139
rect 19073 52105 19107 52139
rect 19107 52105 19116 52139
rect 19064 52096 19116 52105
rect 20904 52096 20956 52148
rect 23112 52096 23164 52148
rect 23296 52096 23348 52148
rect 25136 52139 25188 52148
rect 25136 52105 25145 52139
rect 25145 52105 25179 52139
rect 25179 52105 25188 52139
rect 25136 52096 25188 52105
rect 25504 52139 25556 52148
rect 25504 52105 25513 52139
rect 25513 52105 25547 52139
rect 25547 52105 25556 52139
rect 25504 52096 25556 52105
rect 27712 52139 27764 52148
rect 27712 52105 27721 52139
rect 27721 52105 27755 52139
rect 27755 52105 27764 52139
rect 27712 52096 27764 52105
rect 28264 52096 28316 52148
rect 29460 52096 29512 52148
rect 17960 52028 18012 52080
rect 22284 52071 22336 52080
rect 22284 52037 22293 52071
rect 22293 52037 22327 52071
rect 22327 52037 22336 52071
rect 22284 52028 22336 52037
rect 23940 52028 23992 52080
rect 16120 52003 16172 52012
rect 16120 51969 16129 52003
rect 16129 51969 16163 52003
rect 16163 51969 16172 52003
rect 16120 51960 16172 51969
rect 16672 52003 16724 52012
rect 16672 51969 16681 52003
rect 16681 51969 16715 52003
rect 16715 51969 16724 52003
rect 16672 51960 16724 51969
rect 18328 51960 18380 52012
rect 24124 51960 24176 52012
rect 24860 51960 24912 52012
rect 27620 52028 27672 52080
rect 27344 52003 27396 52012
rect 16948 51935 17000 51944
rect 16948 51901 16957 51935
rect 16957 51901 16991 51935
rect 16991 51901 17000 51935
rect 16948 51892 17000 51901
rect 17776 51892 17828 51944
rect 18604 51892 18656 51944
rect 19156 51892 19208 51944
rect 19984 51892 20036 51944
rect 20260 51935 20312 51944
rect 20260 51901 20269 51935
rect 20269 51901 20303 51935
rect 20303 51901 20312 51935
rect 20260 51892 20312 51901
rect 20444 51935 20496 51944
rect 20444 51901 20453 51935
rect 20453 51901 20487 51935
rect 20487 51901 20496 51935
rect 20444 51892 20496 51901
rect 21548 51935 21600 51944
rect 21548 51901 21557 51935
rect 21557 51901 21591 51935
rect 21591 51901 21600 51935
rect 21548 51892 21600 51901
rect 22376 51935 22428 51944
rect 22376 51901 22385 51935
rect 22385 51901 22419 51935
rect 22419 51901 22428 51935
rect 22376 51892 22428 51901
rect 22560 51935 22612 51944
rect 22560 51901 22569 51935
rect 22569 51901 22603 51935
rect 22603 51901 22612 51935
rect 22560 51892 22612 51901
rect 23480 51935 23532 51944
rect 23480 51901 23489 51935
rect 23489 51901 23523 51935
rect 23523 51901 23532 51935
rect 23480 51892 23532 51901
rect 27344 51969 27353 52003
rect 27353 51969 27387 52003
rect 27387 51969 27396 52003
rect 27344 51960 27396 51969
rect 30564 52003 30616 52012
rect 30564 51969 30573 52003
rect 30573 51969 30607 52003
rect 30607 51969 30616 52003
rect 30564 51960 30616 51969
rect 26792 51935 26844 51944
rect 17868 51867 17920 51876
rect 17868 51833 17877 51867
rect 17877 51833 17911 51867
rect 17911 51833 17920 51867
rect 18420 51867 18472 51876
rect 17868 51824 17920 51833
rect 18420 51833 18429 51867
rect 18429 51833 18463 51867
rect 18463 51833 18472 51867
rect 18420 51824 18472 51833
rect 19248 51824 19300 51876
rect 15752 51756 15804 51808
rect 18972 51756 19024 51808
rect 21640 51824 21692 51876
rect 23296 51824 23348 51876
rect 26792 51901 26801 51935
rect 26801 51901 26835 51935
rect 26835 51901 26844 51935
rect 26792 51892 26844 51901
rect 26884 51935 26936 51944
rect 26884 51901 26893 51935
rect 26893 51901 26927 51935
rect 26927 51901 26936 51935
rect 26884 51892 26936 51901
rect 28080 51892 28132 51944
rect 29092 51935 29144 51944
rect 29092 51901 29101 51935
rect 29101 51901 29135 51935
rect 29135 51901 29144 51935
rect 29092 51892 29144 51901
rect 30288 51935 30340 51944
rect 30288 51901 30297 51935
rect 30297 51901 30331 51935
rect 30331 51901 30340 51935
rect 30288 51892 30340 51901
rect 21456 51799 21508 51808
rect 21456 51765 21465 51799
rect 21465 51765 21499 51799
rect 21499 51765 21508 51799
rect 21456 51756 21508 51765
rect 22192 51756 22244 51808
rect 24676 51799 24728 51808
rect 24676 51765 24685 51799
rect 24685 51765 24719 51799
rect 24719 51765 24728 51799
rect 24676 51756 24728 51765
rect 25780 51824 25832 51876
rect 25320 51756 25372 51808
rect 26240 51756 26292 51808
rect 27528 51824 27580 51876
rect 28264 51756 28316 51808
rect 29000 51756 29052 51808
rect 31760 51756 31812 51808
rect 19606 51654 19658 51706
rect 19670 51654 19722 51706
rect 19734 51654 19786 51706
rect 19798 51654 19850 51706
rect 15108 51595 15160 51604
rect 15108 51561 15117 51595
rect 15117 51561 15151 51595
rect 15151 51561 15160 51595
rect 15108 51552 15160 51561
rect 15476 51595 15528 51604
rect 15476 51561 15485 51595
rect 15485 51561 15519 51595
rect 15519 51561 15528 51595
rect 15476 51552 15528 51561
rect 18604 51552 18656 51604
rect 18788 51595 18840 51604
rect 18788 51561 18797 51595
rect 18797 51561 18831 51595
rect 18831 51561 18840 51595
rect 18788 51552 18840 51561
rect 20260 51595 20312 51604
rect 20260 51561 20269 51595
rect 20269 51561 20303 51595
rect 20303 51561 20312 51595
rect 20260 51552 20312 51561
rect 20536 51552 20588 51604
rect 21364 51595 21416 51604
rect 21364 51561 21373 51595
rect 21373 51561 21407 51595
rect 21407 51561 21416 51595
rect 21364 51552 21416 51561
rect 21824 51595 21876 51604
rect 21824 51561 21833 51595
rect 21833 51561 21867 51595
rect 21867 51561 21876 51595
rect 21824 51552 21876 51561
rect 22008 51552 22060 51604
rect 23296 51595 23348 51604
rect 23296 51561 23305 51595
rect 23305 51561 23339 51595
rect 23339 51561 23348 51595
rect 23296 51552 23348 51561
rect 24860 51552 24912 51604
rect 26884 51552 26936 51604
rect 27988 51552 28040 51604
rect 30288 51552 30340 51604
rect 30656 51595 30708 51604
rect 30656 51561 30665 51595
rect 30665 51561 30699 51595
rect 30699 51561 30708 51595
rect 30656 51552 30708 51561
rect 14924 51484 14976 51536
rect 17776 51484 17828 51536
rect 20076 51484 20128 51536
rect 21180 51484 21232 51536
rect 16028 51459 16080 51468
rect 16028 51425 16037 51459
rect 16037 51425 16071 51459
rect 16071 51425 16080 51459
rect 16028 51416 16080 51425
rect 17408 51459 17460 51468
rect 17408 51425 17417 51459
rect 17417 51425 17451 51459
rect 17451 51425 17460 51459
rect 17408 51416 17460 51425
rect 17868 51459 17920 51468
rect 17868 51425 17877 51459
rect 17877 51425 17911 51459
rect 17911 51425 17920 51459
rect 17868 51416 17920 51425
rect 20904 51459 20956 51468
rect 16580 51348 16632 51400
rect 17500 51348 17552 51400
rect 18972 51391 19024 51400
rect 18972 51357 18981 51391
rect 18981 51357 19015 51391
rect 19015 51357 19024 51391
rect 18972 51348 19024 51357
rect 19524 51391 19576 51400
rect 19524 51357 19533 51391
rect 19533 51357 19567 51391
rect 19567 51357 19576 51391
rect 19524 51348 19576 51357
rect 17960 51323 18012 51332
rect 17960 51289 17969 51323
rect 17969 51289 18003 51323
rect 18003 51289 18012 51323
rect 17960 51280 18012 51289
rect 19800 51280 19852 51332
rect 20904 51425 20913 51459
rect 20913 51425 20947 51459
rect 20947 51425 20956 51459
rect 20904 51416 20956 51425
rect 22376 51484 22428 51536
rect 22560 51484 22612 51536
rect 27252 51527 27304 51536
rect 27252 51493 27261 51527
rect 27261 51493 27295 51527
rect 27295 51493 27304 51527
rect 27252 51484 27304 51493
rect 29092 51484 29144 51536
rect 21732 51416 21784 51468
rect 19984 51391 20036 51400
rect 19984 51357 19993 51391
rect 19993 51357 20027 51391
rect 20027 51357 20036 51391
rect 19984 51348 20036 51357
rect 21364 51348 21416 51400
rect 22008 51416 22060 51468
rect 23940 51459 23992 51468
rect 22100 51348 22152 51400
rect 23940 51425 23949 51459
rect 23949 51425 23983 51459
rect 23983 51425 23992 51459
rect 23940 51416 23992 51425
rect 23112 51348 23164 51400
rect 24308 51416 24360 51468
rect 24952 51459 25004 51468
rect 24952 51425 24961 51459
rect 24961 51425 24995 51459
rect 24995 51425 25004 51459
rect 24952 51416 25004 51425
rect 25044 51416 25096 51468
rect 25320 51416 25372 51468
rect 26976 51459 27028 51468
rect 22284 51280 22336 51332
rect 14740 51255 14792 51264
rect 14740 51221 14749 51255
rect 14749 51221 14783 51255
rect 14783 51221 14792 51255
rect 14740 51212 14792 51221
rect 16212 51255 16264 51264
rect 16212 51221 16221 51255
rect 16221 51221 16255 51255
rect 16255 51221 16264 51255
rect 16212 51212 16264 51221
rect 21732 51212 21784 51264
rect 24768 51348 24820 51400
rect 26976 51425 26985 51459
rect 26985 51425 27019 51459
rect 27019 51425 27028 51459
rect 26976 51416 27028 51425
rect 26884 51348 26936 51400
rect 28356 51391 28408 51400
rect 28356 51357 28365 51391
rect 28365 51357 28399 51391
rect 28399 51357 28408 51391
rect 28356 51348 28408 51357
rect 28448 51391 28500 51400
rect 28448 51357 28457 51391
rect 28457 51357 28491 51391
rect 28491 51357 28500 51391
rect 28448 51348 28500 51357
rect 29552 51416 29604 51468
rect 30196 51459 30248 51468
rect 30196 51425 30205 51459
rect 30205 51425 30239 51459
rect 30239 51425 30248 51459
rect 30196 51416 30248 51425
rect 31392 51459 31444 51468
rect 31392 51425 31401 51459
rect 31401 51425 31435 51459
rect 31435 51425 31444 51459
rect 31392 51416 31444 51425
rect 33692 51416 33744 51468
rect 30288 51280 30340 51332
rect 26332 51212 26384 51264
rect 27528 51255 27580 51264
rect 27528 51221 27537 51255
rect 27537 51221 27571 51255
rect 27571 51221 27580 51255
rect 27528 51212 27580 51221
rect 28908 51212 28960 51264
rect 29552 51212 29604 51264
rect 30104 51255 30156 51264
rect 30104 51221 30113 51255
rect 30113 51221 30147 51255
rect 30147 51221 30156 51255
rect 30104 51212 30156 51221
rect 30380 51255 30432 51264
rect 30380 51221 30389 51255
rect 30389 51221 30423 51255
rect 30423 51221 30432 51255
rect 30380 51212 30432 51221
rect 31484 51212 31536 51264
rect 33600 51212 33652 51264
rect 34152 51212 34204 51264
rect 4246 51110 4298 51162
rect 4310 51110 4362 51162
rect 4374 51110 4426 51162
rect 4438 51110 4490 51162
rect 34966 51110 35018 51162
rect 35030 51110 35082 51162
rect 35094 51110 35146 51162
rect 35158 51110 35210 51162
rect 15016 51008 15068 51060
rect 16028 51051 16080 51060
rect 16028 51017 16037 51051
rect 16037 51017 16071 51051
rect 16071 51017 16080 51051
rect 16028 51008 16080 51017
rect 18604 51008 18656 51060
rect 19800 51051 19852 51060
rect 19800 51017 19809 51051
rect 19809 51017 19843 51051
rect 19843 51017 19852 51051
rect 19800 51008 19852 51017
rect 20352 51051 20404 51060
rect 20352 51017 20361 51051
rect 20361 51017 20395 51051
rect 20395 51017 20404 51051
rect 20352 51008 20404 51017
rect 22008 51051 22060 51060
rect 22008 51017 22017 51051
rect 22017 51017 22051 51051
rect 22051 51017 22060 51051
rect 22008 51008 22060 51017
rect 22284 51051 22336 51060
rect 22284 51017 22293 51051
rect 22293 51017 22327 51051
rect 22327 51017 22336 51051
rect 22284 51008 22336 51017
rect 23388 51008 23440 51060
rect 16212 50940 16264 50992
rect 18880 50983 18932 50992
rect 16580 50872 16632 50924
rect 18880 50949 18889 50983
rect 18889 50949 18923 50983
rect 18923 50949 18932 50983
rect 18880 50940 18932 50949
rect 24308 51008 24360 51060
rect 24860 51051 24912 51060
rect 24860 51017 24869 51051
rect 24869 51017 24903 51051
rect 24903 51017 24912 51051
rect 24860 51008 24912 51017
rect 28080 51008 28132 51060
rect 28356 51008 28408 51060
rect 30196 51008 30248 51060
rect 31392 51008 31444 51060
rect 15108 50847 15160 50856
rect 15108 50813 15117 50847
rect 15117 50813 15151 50847
rect 15151 50813 15160 50847
rect 15108 50804 15160 50813
rect 16672 50847 16724 50856
rect 16672 50813 16681 50847
rect 16681 50813 16715 50847
rect 16715 50813 16724 50847
rect 16672 50804 16724 50813
rect 17224 50872 17276 50924
rect 17868 50872 17920 50924
rect 17316 50736 17368 50788
rect 17500 50779 17552 50788
rect 17500 50745 17509 50779
rect 17509 50745 17543 50779
rect 17543 50745 17552 50779
rect 17500 50736 17552 50745
rect 18788 50804 18840 50856
rect 19248 50804 19300 50856
rect 20720 50804 20772 50856
rect 21640 50872 21692 50924
rect 22008 50872 22060 50924
rect 21364 50847 21416 50856
rect 18236 50736 18288 50788
rect 20444 50736 20496 50788
rect 21364 50813 21373 50847
rect 21373 50813 21407 50847
rect 21407 50813 21416 50847
rect 21364 50804 21416 50813
rect 24768 50940 24820 50992
rect 27620 50940 27672 50992
rect 27344 50872 27396 50924
rect 28724 50872 28776 50924
rect 30012 50872 30064 50924
rect 30564 50872 30616 50924
rect 17960 50668 18012 50720
rect 18144 50668 18196 50720
rect 19984 50668 20036 50720
rect 20352 50668 20404 50720
rect 20904 50668 20956 50720
rect 21180 50668 21232 50720
rect 22008 50668 22060 50720
rect 24860 50804 24912 50856
rect 25504 50804 25556 50856
rect 27068 50804 27120 50856
rect 26424 50736 26476 50788
rect 27988 50736 28040 50788
rect 28172 50779 28224 50788
rect 28172 50745 28181 50779
rect 28181 50745 28215 50779
rect 28215 50745 28224 50779
rect 28172 50736 28224 50745
rect 30840 50847 30892 50856
rect 30840 50813 30849 50847
rect 30849 50813 30883 50847
rect 30883 50813 30892 50847
rect 30840 50804 30892 50813
rect 33692 50847 33744 50856
rect 33692 50813 33701 50847
rect 33701 50813 33735 50847
rect 33735 50813 33744 50847
rect 33692 50804 33744 50813
rect 24308 50668 24360 50720
rect 26884 50711 26936 50720
rect 26884 50677 26893 50711
rect 26893 50677 26927 50711
rect 26927 50677 26936 50711
rect 26884 50668 26936 50677
rect 27528 50668 27580 50720
rect 27804 50668 27856 50720
rect 28356 50668 28408 50720
rect 29000 50711 29052 50720
rect 29000 50677 29009 50711
rect 29009 50677 29043 50711
rect 29043 50677 29052 50711
rect 29000 50668 29052 50677
rect 29460 50668 29512 50720
rect 29736 50668 29788 50720
rect 30932 50668 30984 50720
rect 31024 50711 31076 50720
rect 31024 50677 31033 50711
rect 31033 50677 31067 50711
rect 31067 50677 31076 50711
rect 31024 50668 31076 50677
rect 34796 50668 34848 50720
rect 35440 50668 35492 50720
rect 19606 50566 19658 50618
rect 19670 50566 19722 50618
rect 19734 50566 19786 50618
rect 19798 50566 19850 50618
rect 17868 50464 17920 50516
rect 21364 50464 21416 50516
rect 23940 50464 23992 50516
rect 26976 50464 27028 50516
rect 27528 50464 27580 50516
rect 28172 50464 28224 50516
rect 30472 50464 30524 50516
rect 18512 50396 18564 50448
rect 21088 50396 21140 50448
rect 14832 50124 14884 50176
rect 15660 50328 15712 50380
rect 17960 50328 18012 50380
rect 18972 50328 19024 50380
rect 20628 50328 20680 50380
rect 21732 50371 21784 50380
rect 21732 50337 21741 50371
rect 21741 50337 21775 50371
rect 21775 50337 21784 50371
rect 21732 50328 21784 50337
rect 22284 50371 22336 50380
rect 22284 50337 22293 50371
rect 22293 50337 22327 50371
rect 22327 50337 22336 50371
rect 22284 50328 22336 50337
rect 22652 50371 22704 50380
rect 22652 50337 22661 50371
rect 22661 50337 22695 50371
rect 22695 50337 22704 50371
rect 22652 50328 22704 50337
rect 15292 50303 15344 50312
rect 15292 50269 15301 50303
rect 15301 50269 15335 50303
rect 15335 50269 15344 50303
rect 15292 50260 15344 50269
rect 17408 50260 17460 50312
rect 18052 50260 18104 50312
rect 19340 50260 19392 50312
rect 20168 50260 20220 50312
rect 22192 50192 22244 50244
rect 22928 50396 22980 50448
rect 27068 50396 27120 50448
rect 27712 50396 27764 50448
rect 24124 50328 24176 50380
rect 24492 50371 24544 50380
rect 24492 50337 24501 50371
rect 24501 50337 24535 50371
rect 24535 50337 24544 50371
rect 24492 50328 24544 50337
rect 27252 50328 27304 50380
rect 28356 50371 28408 50380
rect 28356 50337 28365 50371
rect 28365 50337 28399 50371
rect 28399 50337 28408 50371
rect 28356 50328 28408 50337
rect 29092 50328 29144 50380
rect 31484 50371 31536 50380
rect 31484 50337 31493 50371
rect 31493 50337 31527 50371
rect 31527 50337 31536 50371
rect 31484 50328 31536 50337
rect 23664 50303 23716 50312
rect 23664 50269 23673 50303
rect 23673 50269 23707 50303
rect 23707 50269 23716 50303
rect 23664 50260 23716 50269
rect 23848 50260 23900 50312
rect 28264 50260 28316 50312
rect 29552 50303 29604 50312
rect 29552 50269 29561 50303
rect 29561 50269 29595 50303
rect 29595 50269 29604 50303
rect 29552 50260 29604 50269
rect 29736 50260 29788 50312
rect 27804 50192 27856 50244
rect 28540 50192 28592 50244
rect 15200 50124 15252 50176
rect 16304 50124 16356 50176
rect 22468 50124 22520 50176
rect 25320 50124 25372 50176
rect 25596 50124 25648 50176
rect 28908 50167 28960 50176
rect 28908 50133 28917 50167
rect 28917 50133 28951 50167
rect 28951 50133 28960 50167
rect 28908 50124 28960 50133
rect 29276 50167 29328 50176
rect 29276 50133 29285 50167
rect 29285 50133 29319 50167
rect 29319 50133 29328 50167
rect 29276 50124 29328 50133
rect 4246 50022 4298 50074
rect 4310 50022 4362 50074
rect 4374 50022 4426 50074
rect 4438 50022 4490 50074
rect 34966 50022 35018 50074
rect 35030 50022 35082 50074
rect 35094 50022 35146 50074
rect 35158 50022 35210 50074
rect 17224 49920 17276 49972
rect 17316 49920 17368 49972
rect 15200 49852 15252 49904
rect 15660 49852 15712 49904
rect 15384 49827 15436 49836
rect 15384 49793 15393 49827
rect 15393 49793 15427 49827
rect 15427 49793 15436 49827
rect 15384 49784 15436 49793
rect 13820 49716 13872 49768
rect 15660 49716 15712 49768
rect 18236 49920 18288 49972
rect 18144 49852 18196 49904
rect 19340 49920 19392 49972
rect 16304 49759 16356 49768
rect 16304 49725 16313 49759
rect 16313 49725 16347 49759
rect 16347 49725 16356 49759
rect 16304 49716 16356 49725
rect 18236 49759 18288 49768
rect 18236 49725 18245 49759
rect 18245 49725 18279 49759
rect 18279 49725 18288 49759
rect 18236 49716 18288 49725
rect 18604 49759 18656 49768
rect 18604 49725 18613 49759
rect 18613 49725 18647 49759
rect 18647 49725 18656 49759
rect 18604 49716 18656 49725
rect 21732 49920 21784 49972
rect 22560 49920 22612 49972
rect 22928 49920 22980 49972
rect 24124 49920 24176 49972
rect 28356 49963 28408 49972
rect 28356 49929 28365 49963
rect 28365 49929 28399 49963
rect 28399 49929 28408 49963
rect 28356 49920 28408 49929
rect 29552 49920 29604 49972
rect 30656 49920 30708 49972
rect 31944 49920 31996 49972
rect 32220 49963 32272 49972
rect 32220 49929 32229 49963
rect 32229 49929 32263 49963
rect 32263 49929 32272 49963
rect 32220 49920 32272 49929
rect 21088 49852 21140 49904
rect 20076 49759 20128 49768
rect 20076 49725 20085 49759
rect 20085 49725 20119 49759
rect 20119 49725 20128 49759
rect 20076 49716 20128 49725
rect 20260 49648 20312 49700
rect 21088 49759 21140 49768
rect 21088 49725 21097 49759
rect 21097 49725 21131 49759
rect 21131 49725 21140 49759
rect 21088 49716 21140 49725
rect 22192 49759 22244 49768
rect 22192 49725 22201 49759
rect 22201 49725 22235 49759
rect 22235 49725 22244 49759
rect 22192 49716 22244 49725
rect 23940 49852 23992 49904
rect 24308 49852 24360 49904
rect 23480 49827 23532 49836
rect 23480 49793 23489 49827
rect 23489 49793 23523 49827
rect 23523 49793 23532 49827
rect 23480 49784 23532 49793
rect 23388 49716 23440 49768
rect 23940 49759 23992 49768
rect 23940 49725 23949 49759
rect 23949 49725 23983 49759
rect 23983 49725 23992 49759
rect 25136 49784 25188 49836
rect 26240 49852 26292 49904
rect 26332 49852 26384 49904
rect 25964 49784 26016 49836
rect 26976 49784 27028 49836
rect 23940 49716 23992 49725
rect 25596 49716 25648 49768
rect 27528 49759 27580 49768
rect 22284 49648 22336 49700
rect 25228 49648 25280 49700
rect 25504 49648 25556 49700
rect 27528 49725 27537 49759
rect 27537 49725 27571 49759
rect 27571 49725 27580 49759
rect 27528 49716 27580 49725
rect 27804 49716 27856 49768
rect 27896 49759 27948 49768
rect 27896 49725 27905 49759
rect 27905 49725 27939 49759
rect 27939 49725 27948 49759
rect 27896 49716 27948 49725
rect 28632 49716 28684 49768
rect 29828 49852 29880 49904
rect 30104 49784 30156 49836
rect 30564 49784 30616 49836
rect 31208 49827 31260 49836
rect 31208 49793 31217 49827
rect 31217 49793 31251 49827
rect 31251 49793 31260 49827
rect 31208 49784 31260 49793
rect 29092 49759 29144 49768
rect 29092 49725 29101 49759
rect 29101 49725 29135 49759
rect 29135 49725 29144 49759
rect 29092 49716 29144 49725
rect 29276 49716 29328 49768
rect 29828 49716 29880 49768
rect 31024 49759 31076 49768
rect 26332 49648 26384 49700
rect 31024 49725 31033 49759
rect 31033 49725 31067 49759
rect 31067 49725 31076 49759
rect 31024 49716 31076 49725
rect 30380 49648 30432 49700
rect 22192 49623 22244 49632
rect 22192 49589 22201 49623
rect 22201 49589 22235 49623
rect 22235 49589 22244 49623
rect 22192 49580 22244 49589
rect 23756 49580 23808 49632
rect 25596 49623 25648 49632
rect 25596 49589 25605 49623
rect 25605 49589 25639 49623
rect 25639 49589 25648 49623
rect 25596 49580 25648 49589
rect 25964 49580 26016 49632
rect 19606 49478 19658 49530
rect 19670 49478 19722 49530
rect 19734 49478 19786 49530
rect 19798 49478 19850 49530
rect 17868 49376 17920 49428
rect 19432 49376 19484 49428
rect 20260 49419 20312 49428
rect 20260 49385 20269 49419
rect 20269 49385 20303 49419
rect 20303 49385 20312 49419
rect 20260 49376 20312 49385
rect 20720 49419 20772 49428
rect 20720 49385 20729 49419
rect 20729 49385 20763 49419
rect 20763 49385 20772 49419
rect 20720 49376 20772 49385
rect 21548 49376 21600 49428
rect 22560 49376 22612 49428
rect 24032 49376 24084 49428
rect 24768 49376 24820 49428
rect 25044 49376 25096 49428
rect 25596 49376 25648 49428
rect 26700 49376 26752 49428
rect 27252 49376 27304 49428
rect 29736 49376 29788 49428
rect 30380 49376 30432 49428
rect 31668 49376 31720 49428
rect 13268 49351 13320 49360
rect 13268 49317 13277 49351
rect 13277 49317 13311 49351
rect 13311 49317 13320 49351
rect 13268 49308 13320 49317
rect 13728 49283 13780 49292
rect 13728 49249 13737 49283
rect 13737 49249 13771 49283
rect 13771 49249 13780 49283
rect 13728 49240 13780 49249
rect 13544 49172 13596 49224
rect 14004 49240 14056 49292
rect 15016 49308 15068 49360
rect 13268 49104 13320 49156
rect 15292 49240 15344 49292
rect 15476 49240 15528 49292
rect 17408 49240 17460 49292
rect 17868 49172 17920 49224
rect 18604 49172 18656 49224
rect 18972 49240 19024 49292
rect 20628 49240 20680 49292
rect 22284 49283 22336 49292
rect 22284 49249 22293 49283
rect 22293 49249 22327 49283
rect 22327 49249 22336 49283
rect 22284 49240 22336 49249
rect 22652 49283 22704 49292
rect 22652 49249 22661 49283
rect 22661 49249 22695 49283
rect 22695 49249 22704 49283
rect 22652 49240 22704 49249
rect 23572 49240 23624 49292
rect 24032 49283 24084 49292
rect 24032 49249 24041 49283
rect 24041 49249 24075 49283
rect 24075 49249 24084 49283
rect 24032 49240 24084 49249
rect 26792 49308 26844 49360
rect 27528 49351 27580 49360
rect 27528 49317 27537 49351
rect 27537 49317 27571 49351
rect 27571 49317 27580 49351
rect 27528 49308 27580 49317
rect 29276 49308 29328 49360
rect 26700 49283 26752 49292
rect 26700 49249 26709 49283
rect 26709 49249 26743 49283
rect 26743 49249 26752 49283
rect 26700 49240 26752 49249
rect 28724 49240 28776 49292
rect 28816 49283 28868 49292
rect 28816 49249 28825 49283
rect 28825 49249 28859 49283
rect 28859 49249 28868 49283
rect 29920 49283 29972 49292
rect 28816 49240 28868 49249
rect 29920 49249 29929 49283
rect 29929 49249 29963 49283
rect 29963 49249 29972 49283
rect 29920 49240 29972 49249
rect 19708 49172 19760 49224
rect 24768 49215 24820 49224
rect 24768 49181 24777 49215
rect 24777 49181 24811 49215
rect 24811 49181 24820 49215
rect 24768 49172 24820 49181
rect 27068 49215 27120 49224
rect 27068 49181 27077 49215
rect 27077 49181 27111 49215
rect 27111 49181 27120 49215
rect 27068 49172 27120 49181
rect 27988 49172 28040 49224
rect 29460 49172 29512 49224
rect 18696 49147 18748 49156
rect 18696 49113 18705 49147
rect 18705 49113 18739 49147
rect 18739 49113 18748 49147
rect 18696 49104 18748 49113
rect 22376 49104 22428 49156
rect 14832 49036 14884 49088
rect 17776 49036 17828 49088
rect 23848 49036 23900 49088
rect 25964 49036 26016 49088
rect 26240 49079 26292 49088
rect 26240 49045 26249 49079
rect 26249 49045 26283 49079
rect 26283 49045 26292 49079
rect 26240 49036 26292 49045
rect 31208 49079 31260 49088
rect 31208 49045 31217 49079
rect 31217 49045 31251 49079
rect 31251 49045 31260 49079
rect 31208 49036 31260 49045
rect 4246 48934 4298 48986
rect 4310 48934 4362 48986
rect 4374 48934 4426 48986
rect 4438 48934 4490 48986
rect 34966 48934 35018 48986
rect 35030 48934 35082 48986
rect 35094 48934 35146 48986
rect 35158 48934 35210 48986
rect 14004 48832 14056 48884
rect 15292 48832 15344 48884
rect 17408 48875 17460 48884
rect 17408 48841 17417 48875
rect 17417 48841 17451 48875
rect 17451 48841 17460 48875
rect 17408 48832 17460 48841
rect 17868 48875 17920 48884
rect 17868 48841 17877 48875
rect 17877 48841 17911 48875
rect 17911 48841 17920 48875
rect 17868 48832 17920 48841
rect 18236 48875 18288 48884
rect 18236 48841 18245 48875
rect 18245 48841 18279 48875
rect 18279 48841 18288 48875
rect 18236 48832 18288 48841
rect 15384 48807 15436 48816
rect 15384 48773 15393 48807
rect 15393 48773 15427 48807
rect 15427 48773 15436 48807
rect 15384 48764 15436 48773
rect 13268 48671 13320 48680
rect 13268 48637 13277 48671
rect 13277 48637 13311 48671
rect 13311 48637 13320 48671
rect 13268 48628 13320 48637
rect 13544 48671 13596 48680
rect 13544 48637 13553 48671
rect 13553 48637 13587 48671
rect 13587 48637 13596 48671
rect 13544 48628 13596 48637
rect 20076 48832 20128 48884
rect 20628 48832 20680 48884
rect 20996 48875 21048 48884
rect 20996 48841 21005 48875
rect 21005 48841 21039 48875
rect 21039 48841 21048 48875
rect 20996 48832 21048 48841
rect 24952 48832 25004 48884
rect 25412 48832 25464 48884
rect 26700 48832 26752 48884
rect 28724 48875 28776 48884
rect 28724 48841 28733 48875
rect 28733 48841 28767 48875
rect 28767 48841 28776 48875
rect 28724 48832 28776 48841
rect 29920 48832 29972 48884
rect 30748 48832 30800 48884
rect 31208 48832 31260 48884
rect 31392 48875 31444 48884
rect 31392 48841 31401 48875
rect 31401 48841 31435 48875
rect 31435 48841 31444 48875
rect 31392 48832 31444 48841
rect 23572 48764 23624 48816
rect 27620 48764 27672 48816
rect 19248 48739 19300 48748
rect 19248 48705 19257 48739
rect 19257 48705 19291 48739
rect 19291 48705 19300 48739
rect 19248 48696 19300 48705
rect 19524 48696 19576 48748
rect 19432 48671 19484 48680
rect 19432 48637 19441 48671
rect 19441 48637 19475 48671
rect 19475 48637 19484 48671
rect 19432 48628 19484 48637
rect 19984 48671 20036 48680
rect 19984 48637 19993 48671
rect 19993 48637 20027 48671
rect 20027 48637 20036 48671
rect 19984 48628 20036 48637
rect 20352 48628 20404 48680
rect 22100 48696 22152 48748
rect 22376 48696 22428 48748
rect 23020 48696 23072 48748
rect 22560 48671 22612 48680
rect 22560 48637 22569 48671
rect 22569 48637 22603 48671
rect 22603 48637 22612 48671
rect 22560 48628 22612 48637
rect 22744 48671 22796 48680
rect 22744 48637 22753 48671
rect 22753 48637 22787 48671
rect 22787 48637 22796 48671
rect 22744 48628 22796 48637
rect 14648 48535 14700 48544
rect 14648 48501 14657 48535
rect 14657 48501 14691 48535
rect 14691 48501 14700 48535
rect 14648 48492 14700 48501
rect 17224 48492 17276 48544
rect 20904 48535 20956 48544
rect 20904 48501 20913 48535
rect 20913 48501 20947 48535
rect 20947 48501 20956 48535
rect 20904 48492 20956 48501
rect 22284 48492 22336 48544
rect 22560 48492 22612 48544
rect 24124 48492 24176 48544
rect 26240 48696 26292 48748
rect 25044 48628 25096 48680
rect 29460 48739 29512 48748
rect 29460 48705 29469 48739
rect 29469 48705 29503 48739
rect 29503 48705 29512 48739
rect 29460 48696 29512 48705
rect 30288 48739 30340 48748
rect 30288 48705 30297 48739
rect 30297 48705 30331 48739
rect 30331 48705 30340 48739
rect 30288 48696 30340 48705
rect 27160 48671 27212 48680
rect 24952 48492 25004 48544
rect 25228 48560 25280 48612
rect 26332 48560 26384 48612
rect 27160 48637 27169 48671
rect 27169 48637 27203 48671
rect 27203 48637 27212 48671
rect 27160 48628 27212 48637
rect 28172 48671 28224 48680
rect 28172 48637 28181 48671
rect 28181 48637 28215 48671
rect 28215 48637 28224 48671
rect 28172 48628 28224 48637
rect 29828 48628 29880 48680
rect 31208 48671 31260 48680
rect 31208 48637 31217 48671
rect 31217 48637 31251 48671
rect 31251 48637 31260 48671
rect 31208 48628 31260 48637
rect 25780 48492 25832 48544
rect 25964 48492 26016 48544
rect 26792 48492 26844 48544
rect 27436 48492 27488 48544
rect 27988 48535 28040 48544
rect 27988 48501 27997 48535
rect 27997 48501 28031 48535
rect 28031 48501 28040 48535
rect 27988 48492 28040 48501
rect 28540 48492 28592 48544
rect 28816 48492 28868 48544
rect 29276 48492 29328 48544
rect 30656 48535 30708 48544
rect 30656 48501 30665 48535
rect 30665 48501 30699 48535
rect 30699 48501 30708 48535
rect 30656 48492 30708 48501
rect 19606 48390 19658 48442
rect 19670 48390 19722 48442
rect 19734 48390 19786 48442
rect 19798 48390 19850 48442
rect 9128 48288 9180 48340
rect 9404 48288 9456 48340
rect 13544 48288 13596 48340
rect 15476 48288 15528 48340
rect 17224 48288 17276 48340
rect 18972 48288 19024 48340
rect 22652 48288 22704 48340
rect 11612 48263 11664 48272
rect 11612 48229 11621 48263
rect 11621 48229 11655 48263
rect 11655 48229 11664 48263
rect 11612 48220 11664 48229
rect 15108 48263 15160 48272
rect 15108 48229 15117 48263
rect 15117 48229 15151 48263
rect 15151 48229 15160 48263
rect 15108 48220 15160 48229
rect 18420 48263 18472 48272
rect 18420 48229 18429 48263
rect 18429 48229 18463 48263
rect 18463 48229 18472 48263
rect 18420 48220 18472 48229
rect 18604 48220 18656 48272
rect 19984 48220 20036 48272
rect 20444 48220 20496 48272
rect 22376 48263 22428 48272
rect 22376 48229 22385 48263
rect 22385 48229 22419 48263
rect 22419 48229 22428 48263
rect 22376 48220 22428 48229
rect 23020 48263 23072 48272
rect 23020 48229 23029 48263
rect 23029 48229 23063 48263
rect 23063 48229 23072 48263
rect 23020 48220 23072 48229
rect 25044 48288 25096 48340
rect 25596 48331 25648 48340
rect 25596 48297 25605 48331
rect 25605 48297 25639 48331
rect 25639 48297 25648 48331
rect 28172 48331 28224 48340
rect 25596 48288 25648 48297
rect 28172 48297 28181 48331
rect 28181 48297 28215 48331
rect 28215 48297 28224 48331
rect 28172 48288 28224 48297
rect 28724 48288 28776 48340
rect 29460 48331 29512 48340
rect 29460 48297 29469 48331
rect 29469 48297 29503 48331
rect 29503 48297 29512 48331
rect 29460 48288 29512 48297
rect 29828 48331 29880 48340
rect 29828 48297 29837 48331
rect 29837 48297 29871 48331
rect 29871 48297 29880 48331
rect 29828 48288 29880 48297
rect 23572 48220 23624 48272
rect 24124 48220 24176 48272
rect 10968 48152 11020 48204
rect 12256 48195 12308 48204
rect 12256 48161 12265 48195
rect 12265 48161 12299 48195
rect 12299 48161 12308 48195
rect 12256 48152 12308 48161
rect 12808 48195 12860 48204
rect 12164 48127 12216 48136
rect 12164 48093 12173 48127
rect 12173 48093 12207 48127
rect 12207 48093 12216 48127
rect 12164 48084 12216 48093
rect 11428 47991 11480 48000
rect 11428 47957 11437 47991
rect 11437 47957 11471 47991
rect 11471 47957 11480 47991
rect 12808 48161 12817 48195
rect 12817 48161 12851 48195
rect 12851 48161 12860 48195
rect 12808 48152 12860 48161
rect 14280 48152 14332 48204
rect 14648 48152 14700 48204
rect 15844 48152 15896 48204
rect 16120 48195 16172 48204
rect 14004 48084 14056 48136
rect 16120 48161 16129 48195
rect 16129 48161 16163 48195
rect 16163 48161 16172 48195
rect 16120 48152 16172 48161
rect 19064 48195 19116 48204
rect 19064 48161 19073 48195
rect 19073 48161 19107 48195
rect 19107 48161 19116 48195
rect 19064 48152 19116 48161
rect 19432 48195 19484 48204
rect 19432 48161 19441 48195
rect 19441 48161 19475 48195
rect 19475 48161 19484 48195
rect 19432 48152 19484 48161
rect 21180 48195 21232 48204
rect 21180 48161 21189 48195
rect 21189 48161 21223 48195
rect 21223 48161 21232 48195
rect 21180 48152 21232 48161
rect 21456 48195 21508 48204
rect 21456 48161 21465 48195
rect 21465 48161 21499 48195
rect 21499 48161 21508 48195
rect 21456 48152 21508 48161
rect 22560 48195 22612 48204
rect 22560 48161 22569 48195
rect 22569 48161 22603 48195
rect 22603 48161 22612 48195
rect 22560 48152 22612 48161
rect 23848 48195 23900 48204
rect 23848 48161 23857 48195
rect 23857 48161 23891 48195
rect 23891 48161 23900 48195
rect 23848 48152 23900 48161
rect 13728 48016 13780 48068
rect 16672 48084 16724 48136
rect 19984 48127 20036 48136
rect 19984 48093 19993 48127
rect 19993 48093 20027 48127
rect 20027 48093 20036 48127
rect 19984 48084 20036 48093
rect 20720 48084 20772 48136
rect 15568 48059 15620 48068
rect 15568 48025 15577 48059
rect 15577 48025 15611 48059
rect 15611 48025 15620 48059
rect 15568 48016 15620 48025
rect 19892 48016 19944 48068
rect 20260 48016 20312 48068
rect 21088 48016 21140 48068
rect 23388 48084 23440 48136
rect 24492 48152 24544 48204
rect 26424 48220 26476 48272
rect 26608 48220 26660 48272
rect 27620 48220 27672 48272
rect 28448 48220 28500 48272
rect 26792 48152 26844 48204
rect 27068 48152 27120 48204
rect 27528 48152 27580 48204
rect 27804 48195 27856 48204
rect 27804 48161 27813 48195
rect 27813 48161 27847 48195
rect 27847 48161 27856 48195
rect 27804 48152 27856 48161
rect 28540 48195 28592 48204
rect 28540 48161 28549 48195
rect 28549 48161 28583 48195
rect 28583 48161 28592 48195
rect 28540 48152 28592 48161
rect 29552 48195 29604 48204
rect 29552 48161 29561 48195
rect 29561 48161 29595 48195
rect 29595 48161 29604 48195
rect 29552 48152 29604 48161
rect 29920 48195 29972 48204
rect 29920 48161 29929 48195
rect 29929 48161 29963 48195
rect 29963 48161 29972 48195
rect 29920 48152 29972 48161
rect 30380 48152 30432 48204
rect 24308 48084 24360 48136
rect 24676 48127 24728 48136
rect 24676 48093 24685 48127
rect 24685 48093 24719 48127
rect 24719 48093 24728 48127
rect 24676 48084 24728 48093
rect 31392 48084 31444 48136
rect 23664 48016 23716 48068
rect 28080 48016 28132 48068
rect 28908 48016 28960 48068
rect 29092 48016 29144 48068
rect 29460 48016 29512 48068
rect 29644 48016 29696 48068
rect 11428 47948 11480 47957
rect 14648 47991 14700 48000
rect 14648 47957 14657 47991
rect 14657 47957 14691 47991
rect 14691 47957 14700 47991
rect 14648 47948 14700 47957
rect 24032 47948 24084 48000
rect 26240 47991 26292 48000
rect 26240 47957 26249 47991
rect 26249 47957 26283 47991
rect 26283 47957 26292 47991
rect 26240 47948 26292 47957
rect 29000 47948 29052 48000
rect 30840 47948 30892 48000
rect 4246 47846 4298 47898
rect 4310 47846 4362 47898
rect 4374 47846 4426 47898
rect 4438 47846 4490 47898
rect 34966 47846 35018 47898
rect 35030 47846 35082 47898
rect 35094 47846 35146 47898
rect 35158 47846 35210 47898
rect 10968 47787 11020 47796
rect 10968 47753 10977 47787
rect 10977 47753 11011 47787
rect 11011 47753 11020 47787
rect 10968 47744 11020 47753
rect 12808 47744 12860 47796
rect 13176 47744 13228 47796
rect 13820 47744 13872 47796
rect 14280 47787 14332 47796
rect 14280 47753 14289 47787
rect 14289 47753 14323 47787
rect 14323 47753 14332 47787
rect 14280 47744 14332 47753
rect 16672 47787 16724 47796
rect 16672 47753 16681 47787
rect 16681 47753 16715 47787
rect 16715 47753 16724 47787
rect 16672 47744 16724 47753
rect 18604 47787 18656 47796
rect 18604 47753 18613 47787
rect 18613 47753 18647 47787
rect 18647 47753 18656 47787
rect 18604 47744 18656 47753
rect 19064 47744 19116 47796
rect 19432 47744 19484 47796
rect 20076 47744 20128 47796
rect 21180 47744 21232 47796
rect 22744 47744 22796 47796
rect 23388 47744 23440 47796
rect 27068 47744 27120 47796
rect 29092 47787 29144 47796
rect 29092 47753 29101 47787
rect 29101 47753 29135 47787
rect 29135 47753 29144 47787
rect 29092 47744 29144 47753
rect 31116 47787 31168 47796
rect 31116 47753 31125 47787
rect 31125 47753 31159 47787
rect 31159 47753 31168 47787
rect 31116 47744 31168 47753
rect 12164 47719 12216 47728
rect 12164 47685 12173 47719
rect 12173 47685 12207 47719
rect 12207 47685 12216 47719
rect 12164 47676 12216 47685
rect 12624 47608 12676 47660
rect 23940 47676 23992 47728
rect 15108 47608 15160 47660
rect 22008 47608 22060 47660
rect 23664 47608 23716 47660
rect 24952 47608 25004 47660
rect 26332 47608 26384 47660
rect 29276 47676 29328 47728
rect 32404 47719 32456 47728
rect 32404 47685 32413 47719
rect 32413 47685 32447 47719
rect 32447 47685 32456 47719
rect 32404 47676 32456 47685
rect 12992 47583 13044 47592
rect 12992 47549 13001 47583
rect 13001 47549 13035 47583
rect 13035 47549 13044 47583
rect 12992 47540 13044 47549
rect 13268 47540 13320 47592
rect 13452 47583 13504 47592
rect 13452 47549 13461 47583
rect 13461 47549 13495 47583
rect 13495 47549 13504 47583
rect 14648 47583 14700 47592
rect 13452 47540 13504 47549
rect 14648 47549 14657 47583
rect 14657 47549 14691 47583
rect 14691 47549 14700 47583
rect 14648 47540 14700 47549
rect 15292 47540 15344 47592
rect 16120 47540 16172 47592
rect 16856 47583 16908 47592
rect 14004 47404 14056 47456
rect 15752 47447 15804 47456
rect 15752 47413 15761 47447
rect 15761 47413 15795 47447
rect 15795 47413 15804 47447
rect 15752 47404 15804 47413
rect 16856 47549 16865 47583
rect 16865 47549 16899 47583
rect 16899 47549 16908 47583
rect 16856 47540 16908 47549
rect 21088 47583 21140 47592
rect 21088 47549 21097 47583
rect 21097 47549 21131 47583
rect 21131 47549 21140 47583
rect 21088 47540 21140 47549
rect 21640 47540 21692 47592
rect 23388 47540 23440 47592
rect 24032 47540 24084 47592
rect 24492 47583 24544 47592
rect 24492 47549 24501 47583
rect 24501 47549 24535 47583
rect 24535 47549 24544 47583
rect 24492 47540 24544 47549
rect 24676 47583 24728 47592
rect 24676 47549 24685 47583
rect 24685 47549 24719 47583
rect 24719 47549 24728 47583
rect 24676 47540 24728 47549
rect 25596 47540 25648 47592
rect 27712 47583 27764 47592
rect 27712 47549 27721 47583
rect 27721 47549 27755 47583
rect 27755 47549 27764 47583
rect 27712 47540 27764 47549
rect 27804 47540 27856 47592
rect 27988 47540 28040 47592
rect 23572 47472 23624 47524
rect 25320 47472 25372 47524
rect 25964 47472 26016 47524
rect 27528 47472 27580 47524
rect 29092 47540 29144 47592
rect 29920 47608 29972 47660
rect 29828 47540 29880 47592
rect 30840 47583 30892 47592
rect 30840 47549 30849 47583
rect 30849 47549 30883 47583
rect 30883 47549 30892 47583
rect 30840 47540 30892 47549
rect 30932 47583 30984 47592
rect 30932 47549 30941 47583
rect 30941 47549 30975 47583
rect 30975 47549 30984 47583
rect 30932 47540 30984 47549
rect 30380 47515 30432 47524
rect 30380 47481 30389 47515
rect 30389 47481 30423 47515
rect 30423 47481 30432 47515
rect 30380 47472 30432 47481
rect 31024 47472 31076 47524
rect 20076 47404 20128 47456
rect 25596 47404 25648 47456
rect 26792 47404 26844 47456
rect 28540 47447 28592 47456
rect 28540 47413 28549 47447
rect 28549 47413 28583 47447
rect 28583 47413 28592 47447
rect 28540 47404 28592 47413
rect 29368 47447 29420 47456
rect 29368 47413 29377 47447
rect 29377 47413 29411 47447
rect 29411 47413 29420 47447
rect 29368 47404 29420 47413
rect 30656 47447 30708 47456
rect 30656 47413 30665 47447
rect 30665 47413 30699 47447
rect 30699 47413 30708 47447
rect 30656 47404 30708 47413
rect 19606 47302 19658 47354
rect 19670 47302 19722 47354
rect 19734 47302 19786 47354
rect 19798 47302 19850 47354
rect 12256 47200 12308 47252
rect 13452 47200 13504 47252
rect 19432 47200 19484 47252
rect 21180 47243 21232 47252
rect 21180 47209 21189 47243
rect 21189 47209 21223 47243
rect 21223 47209 21232 47243
rect 21180 47200 21232 47209
rect 21456 47243 21508 47252
rect 21456 47209 21465 47243
rect 21465 47209 21499 47243
rect 21499 47209 21508 47243
rect 21456 47200 21508 47209
rect 22560 47200 22612 47252
rect 23756 47200 23808 47252
rect 24124 47200 24176 47252
rect 25412 47243 25464 47252
rect 25412 47209 25421 47243
rect 25421 47209 25455 47243
rect 25455 47209 25464 47243
rect 25412 47200 25464 47209
rect 25780 47243 25832 47252
rect 25780 47209 25789 47243
rect 25789 47209 25823 47243
rect 25823 47209 25832 47243
rect 25780 47200 25832 47209
rect 27068 47200 27120 47252
rect 28448 47243 28500 47252
rect 28448 47209 28457 47243
rect 28457 47209 28491 47243
rect 28491 47209 28500 47243
rect 28448 47200 28500 47209
rect 29828 47243 29880 47252
rect 29828 47209 29837 47243
rect 29837 47209 29871 47243
rect 29871 47209 29880 47243
rect 29828 47200 29880 47209
rect 30196 47243 30248 47252
rect 30196 47209 30205 47243
rect 30205 47209 30239 47243
rect 30239 47209 30248 47243
rect 30196 47200 30248 47209
rect 31392 47243 31444 47252
rect 31392 47209 31401 47243
rect 31401 47209 31435 47243
rect 31435 47209 31444 47243
rect 31392 47200 31444 47209
rect 12992 47132 13044 47184
rect 15844 47175 15896 47184
rect 15844 47141 15853 47175
rect 15853 47141 15887 47175
rect 15887 47141 15896 47175
rect 15844 47132 15896 47141
rect 11428 47064 11480 47116
rect 13912 47107 13964 47116
rect 13912 47073 13921 47107
rect 13921 47073 13955 47107
rect 13955 47073 13964 47107
rect 13912 47064 13964 47073
rect 15752 47064 15804 47116
rect 17316 47064 17368 47116
rect 19892 47064 19944 47116
rect 11704 46996 11756 47048
rect 14004 46996 14056 47048
rect 16948 47039 17000 47048
rect 16948 47005 16957 47039
rect 16957 47005 16991 47039
rect 16991 47005 17000 47039
rect 16948 46996 17000 47005
rect 23020 47132 23072 47184
rect 23848 47132 23900 47184
rect 24216 47132 24268 47184
rect 20352 46971 20404 46980
rect 20352 46937 20361 46971
rect 20361 46937 20395 46971
rect 20395 46937 20404 46971
rect 20352 46928 20404 46937
rect 21916 46971 21968 46980
rect 21916 46937 21925 46971
rect 21925 46937 21959 46971
rect 21959 46937 21968 46971
rect 21916 46928 21968 46937
rect 1400 46860 1452 46912
rect 14924 46903 14976 46912
rect 14924 46869 14933 46903
rect 14933 46869 14967 46903
rect 14967 46869 14976 46903
rect 14924 46860 14976 46869
rect 22100 47064 22152 47116
rect 23664 46996 23716 47048
rect 24308 46996 24360 47048
rect 22192 46928 22244 46980
rect 23572 46928 23624 46980
rect 25596 47132 25648 47184
rect 26884 47132 26936 47184
rect 28540 47132 28592 47184
rect 30748 47175 30800 47184
rect 30748 47141 30757 47175
rect 30757 47141 30791 47175
rect 30791 47141 30800 47175
rect 30748 47132 30800 47141
rect 31852 47132 31904 47184
rect 25228 47107 25280 47116
rect 25228 47073 25237 47107
rect 25237 47073 25271 47107
rect 25271 47073 25280 47107
rect 25228 47064 25280 47073
rect 27160 47107 27212 47116
rect 27160 47073 27169 47107
rect 27169 47073 27203 47107
rect 27203 47073 27212 47107
rect 27160 47064 27212 47073
rect 27528 47107 27580 47116
rect 27528 47073 27537 47107
rect 27537 47073 27571 47107
rect 27571 47073 27580 47107
rect 27528 47064 27580 47073
rect 29000 47107 29052 47116
rect 29000 47073 29009 47107
rect 29009 47073 29043 47107
rect 29043 47073 29052 47107
rect 29000 47064 29052 47073
rect 29276 47064 29328 47116
rect 26884 46996 26936 47048
rect 27436 46996 27488 47048
rect 27712 46996 27764 47048
rect 28908 46996 28960 47048
rect 29092 46996 29144 47048
rect 29920 47064 29972 47116
rect 30564 47107 30616 47116
rect 30564 47073 30573 47107
rect 30573 47073 30607 47107
rect 30607 47073 30616 47107
rect 30564 47064 30616 47073
rect 31024 47064 31076 47116
rect 32128 47107 32180 47116
rect 32128 47073 32137 47107
rect 32137 47073 32171 47107
rect 32171 47073 32180 47107
rect 32128 47064 32180 47073
rect 30380 47039 30432 47048
rect 30380 47005 30389 47039
rect 30389 47005 30423 47039
rect 30423 47005 30432 47039
rect 30380 46996 30432 47005
rect 31116 47039 31168 47048
rect 31116 47005 31125 47039
rect 31125 47005 31159 47039
rect 31159 47005 31168 47039
rect 31116 46996 31168 47005
rect 28816 46971 28868 46980
rect 22284 46860 22336 46912
rect 22744 46860 22796 46912
rect 28816 46937 28825 46971
rect 28825 46937 28859 46971
rect 28859 46937 28868 46971
rect 28816 46928 28868 46937
rect 24032 46860 24084 46912
rect 29644 46860 29696 46912
rect 4246 46758 4298 46810
rect 4310 46758 4362 46810
rect 4374 46758 4426 46810
rect 4438 46758 4490 46810
rect 34966 46758 35018 46810
rect 35030 46758 35082 46810
rect 35094 46758 35146 46810
rect 35158 46758 35210 46810
rect 11704 46699 11756 46708
rect 11704 46665 11713 46699
rect 11713 46665 11747 46699
rect 11747 46665 11756 46699
rect 11704 46656 11756 46665
rect 13912 46656 13964 46708
rect 19892 46699 19944 46708
rect 19892 46665 19901 46699
rect 19901 46665 19935 46699
rect 19935 46665 19944 46699
rect 19892 46656 19944 46665
rect 20904 46656 20956 46708
rect 22008 46656 22060 46708
rect 25228 46699 25280 46708
rect 25228 46665 25237 46699
rect 25237 46665 25271 46699
rect 25271 46665 25280 46699
rect 25228 46656 25280 46665
rect 27160 46656 27212 46708
rect 29092 46699 29144 46708
rect 29092 46665 29101 46699
rect 29101 46665 29135 46699
rect 29135 46665 29144 46699
rect 29092 46656 29144 46665
rect 29552 46656 29604 46708
rect 32128 46699 32180 46708
rect 22192 46588 22244 46640
rect 1676 46563 1728 46572
rect 1676 46529 1685 46563
rect 1685 46529 1719 46563
rect 1719 46529 1728 46563
rect 1676 46520 1728 46529
rect 12716 46563 12768 46572
rect 12716 46529 12725 46563
rect 12725 46529 12759 46563
rect 12759 46529 12768 46563
rect 12716 46520 12768 46529
rect 13452 46520 13504 46572
rect 14556 46520 14608 46572
rect 22468 46563 22520 46572
rect 22468 46529 22477 46563
rect 22477 46529 22511 46563
rect 22511 46529 22520 46563
rect 22468 46520 22520 46529
rect 28172 46588 28224 46640
rect 28632 46588 28684 46640
rect 24676 46563 24728 46572
rect 1400 46495 1452 46504
rect 1400 46461 1409 46495
rect 1409 46461 1443 46495
rect 1443 46461 1452 46495
rect 1400 46452 1452 46461
rect 11704 46452 11756 46504
rect 12440 46495 12492 46504
rect 12440 46461 12449 46495
rect 12449 46461 12483 46495
rect 12483 46461 12492 46495
rect 12440 46452 12492 46461
rect 15016 46452 15068 46504
rect 15568 46495 15620 46504
rect 15568 46461 15577 46495
rect 15577 46461 15611 46495
rect 15611 46461 15620 46495
rect 15568 46452 15620 46461
rect 15660 46452 15712 46504
rect 20996 46495 21048 46504
rect 20996 46461 21005 46495
rect 21005 46461 21039 46495
rect 21039 46461 21048 46495
rect 20996 46452 21048 46461
rect 21916 46452 21968 46504
rect 22100 46495 22152 46504
rect 22100 46461 22109 46495
rect 22109 46461 22143 46495
rect 22143 46461 22152 46495
rect 22100 46452 22152 46461
rect 22928 46452 22980 46504
rect 24676 46529 24685 46563
rect 24685 46529 24719 46563
rect 24719 46529 24728 46563
rect 24676 46520 24728 46529
rect 26516 46520 26568 46572
rect 32128 46665 32137 46699
rect 32137 46665 32171 46699
rect 32171 46665 32180 46699
rect 32128 46656 32180 46665
rect 31852 46588 31904 46640
rect 24032 46452 24084 46504
rect 24860 46452 24912 46504
rect 26608 46452 26660 46504
rect 27068 46452 27120 46504
rect 28172 46495 28224 46504
rect 3056 46427 3108 46436
rect 3056 46393 3065 46427
rect 3065 46393 3099 46427
rect 3099 46393 3108 46427
rect 3056 46384 3108 46393
rect 16948 46384 17000 46436
rect 17500 46384 17552 46436
rect 26424 46384 26476 46436
rect 28172 46461 28181 46495
rect 28181 46461 28215 46495
rect 28215 46461 28224 46495
rect 28172 46452 28224 46461
rect 11428 46359 11480 46368
rect 11428 46325 11437 46359
rect 11437 46325 11471 46359
rect 11471 46325 11480 46359
rect 11428 46316 11480 46325
rect 12348 46316 12400 46368
rect 12716 46316 12768 46368
rect 14004 46316 14056 46368
rect 17316 46316 17368 46368
rect 25780 46316 25832 46368
rect 27804 46316 27856 46368
rect 28080 46316 28132 46368
rect 31944 46520 31996 46572
rect 29552 46452 29604 46504
rect 28908 46316 28960 46368
rect 31208 46359 31260 46368
rect 31208 46325 31217 46359
rect 31217 46325 31251 46359
rect 31251 46325 31260 46359
rect 31208 46316 31260 46325
rect 31760 46359 31812 46368
rect 31760 46325 31769 46359
rect 31769 46325 31803 46359
rect 31803 46325 31812 46359
rect 31760 46316 31812 46325
rect 19606 46214 19658 46266
rect 19670 46214 19722 46266
rect 19734 46214 19786 46266
rect 19798 46214 19850 46266
rect 1676 46155 1728 46164
rect 1676 46121 1685 46155
rect 1685 46121 1719 46155
rect 1719 46121 1728 46155
rect 1676 46112 1728 46121
rect 8852 46155 8904 46164
rect 8852 46121 8861 46155
rect 8861 46121 8895 46155
rect 8895 46121 8904 46155
rect 8852 46112 8904 46121
rect 9680 46112 9732 46164
rect 12440 46112 12492 46164
rect 13360 46155 13412 46164
rect 13360 46121 13369 46155
rect 13369 46121 13403 46155
rect 13403 46121 13412 46155
rect 13360 46112 13412 46121
rect 13912 46112 13964 46164
rect 15752 46112 15804 46164
rect 22100 46112 22152 46164
rect 22376 46112 22428 46164
rect 23664 46155 23716 46164
rect 23664 46121 23673 46155
rect 23673 46121 23707 46155
rect 23707 46121 23716 46155
rect 23664 46112 23716 46121
rect 25964 46112 26016 46164
rect 27252 46112 27304 46164
rect 27436 46112 27488 46164
rect 28632 46155 28684 46164
rect 14924 46044 14976 46096
rect 22928 46044 22980 46096
rect 28632 46121 28641 46155
rect 28641 46121 28675 46155
rect 28675 46121 28684 46155
rect 28632 46112 28684 46121
rect 29276 46112 29328 46164
rect 29460 46112 29512 46164
rect 30380 46155 30432 46164
rect 30380 46121 30389 46155
rect 30389 46121 30423 46155
rect 30423 46121 30432 46155
rect 30380 46112 30432 46121
rect 30564 46112 30616 46164
rect 30932 46112 30984 46164
rect 31760 46112 31812 46164
rect 28540 46044 28592 46096
rect 29184 46044 29236 46096
rect 12808 46019 12860 46028
rect 12808 45985 12817 46019
rect 12817 45985 12851 46019
rect 12851 45985 12860 46019
rect 12808 45976 12860 45985
rect 14740 45976 14792 46028
rect 21180 45976 21232 46028
rect 22284 45976 22336 46028
rect 22744 46019 22796 46028
rect 14004 45908 14056 45960
rect 22744 45985 22753 46019
rect 22753 45985 22787 46019
rect 22787 45985 22796 46019
rect 22744 45976 22796 45985
rect 24860 46019 24912 46028
rect 24860 45985 24869 46019
rect 24869 45985 24903 46019
rect 24903 45985 24912 46019
rect 24860 45976 24912 45985
rect 27528 46019 27580 46028
rect 27528 45985 27537 46019
rect 27537 45985 27571 46019
rect 27571 45985 27580 46019
rect 27528 45976 27580 45985
rect 27620 45976 27672 46028
rect 28356 45976 28408 46028
rect 29092 45976 29144 46028
rect 31024 45976 31076 46028
rect 32128 46019 32180 46028
rect 32128 45985 32137 46019
rect 32137 45985 32171 46019
rect 32171 45985 32180 46019
rect 32128 45976 32180 45985
rect 32220 46019 32272 46028
rect 32220 45985 32229 46019
rect 32229 45985 32263 46019
rect 32263 45985 32272 46019
rect 32220 45976 32272 45985
rect 22928 45951 22980 45960
rect 21640 45883 21692 45892
rect 21640 45849 21649 45883
rect 21649 45849 21683 45883
rect 21683 45849 21692 45883
rect 21640 45840 21692 45849
rect 13268 45772 13320 45824
rect 15660 45772 15712 45824
rect 22376 45840 22428 45892
rect 22928 45917 22937 45951
rect 22937 45917 22971 45951
rect 22971 45917 22980 45951
rect 22928 45908 22980 45917
rect 24032 45951 24084 45960
rect 24032 45917 24041 45951
rect 24041 45917 24075 45951
rect 24075 45917 24084 45951
rect 24032 45908 24084 45917
rect 23388 45840 23440 45892
rect 24308 45840 24360 45892
rect 24676 45908 24728 45960
rect 23480 45772 23532 45824
rect 25412 45815 25464 45824
rect 25412 45781 25421 45815
rect 25421 45781 25455 45815
rect 25455 45781 25464 45815
rect 25412 45772 25464 45781
rect 26424 45772 26476 45824
rect 30472 45772 30524 45824
rect 31392 45772 31444 45824
rect 32404 45815 32456 45824
rect 32404 45781 32413 45815
rect 32413 45781 32447 45815
rect 32447 45781 32456 45815
rect 32404 45772 32456 45781
rect 4246 45670 4298 45722
rect 4310 45670 4362 45722
rect 4374 45670 4426 45722
rect 4438 45670 4490 45722
rect 34966 45670 35018 45722
rect 35030 45670 35082 45722
rect 35094 45670 35146 45722
rect 35158 45670 35210 45722
rect 14740 45611 14792 45620
rect 14740 45577 14749 45611
rect 14749 45577 14783 45611
rect 14783 45577 14792 45611
rect 14740 45568 14792 45577
rect 8760 45500 8812 45552
rect 9864 45475 9916 45484
rect 9864 45441 9873 45475
rect 9873 45441 9907 45475
rect 9907 45441 9916 45475
rect 9864 45432 9916 45441
rect 13360 45475 13412 45484
rect 13360 45441 13369 45475
rect 13369 45441 13403 45475
rect 13403 45441 13412 45475
rect 13360 45432 13412 45441
rect 9128 45364 9180 45416
rect 9680 45364 9732 45416
rect 13452 45364 13504 45416
rect 22928 45568 22980 45620
rect 23388 45568 23440 45620
rect 23480 45500 23532 45552
rect 24676 45500 24728 45552
rect 23940 45432 23992 45484
rect 25964 45568 26016 45620
rect 26516 45568 26568 45620
rect 27620 45611 27672 45620
rect 27620 45577 27629 45611
rect 27629 45577 27663 45611
rect 27663 45577 27672 45611
rect 27620 45568 27672 45577
rect 28172 45568 28224 45620
rect 31024 45568 31076 45620
rect 32128 45611 32180 45620
rect 32128 45577 32137 45611
rect 32137 45577 32171 45611
rect 32171 45577 32180 45611
rect 32128 45568 32180 45577
rect 32220 45568 32272 45620
rect 28080 45543 28132 45552
rect 28080 45509 28089 45543
rect 28089 45509 28123 45543
rect 28123 45509 28132 45543
rect 28080 45500 28132 45509
rect 29092 45543 29144 45552
rect 29092 45509 29101 45543
rect 29101 45509 29135 45543
rect 29135 45509 29144 45543
rect 29092 45500 29144 45509
rect 29460 45500 29512 45552
rect 29736 45500 29788 45552
rect 25412 45432 25464 45484
rect 26608 45432 26660 45484
rect 25044 45364 25096 45416
rect 26516 45364 26568 45416
rect 26792 45407 26844 45416
rect 26792 45373 26801 45407
rect 26801 45373 26835 45407
rect 26835 45373 26844 45407
rect 26792 45364 26844 45373
rect 26884 45407 26936 45416
rect 26884 45373 26893 45407
rect 26893 45373 26927 45407
rect 26927 45373 26936 45407
rect 27988 45432 28040 45484
rect 29000 45432 29052 45484
rect 26884 45364 26936 45373
rect 27344 45407 27396 45416
rect 27344 45373 27353 45407
rect 27353 45373 27387 45407
rect 27387 45373 27396 45407
rect 27344 45364 27396 45373
rect 8576 45296 8628 45348
rect 22468 45296 22520 45348
rect 12808 45271 12860 45280
rect 12808 45237 12817 45271
rect 12817 45237 12851 45271
rect 12851 45237 12860 45271
rect 12808 45228 12860 45237
rect 14004 45228 14056 45280
rect 21180 45228 21232 45280
rect 22744 45228 22796 45280
rect 24124 45296 24176 45348
rect 28172 45407 28224 45416
rect 28172 45373 28181 45407
rect 28181 45373 28215 45407
rect 28215 45373 28224 45407
rect 28172 45364 28224 45373
rect 28908 45364 28960 45416
rect 30196 45364 30248 45416
rect 31484 45364 31536 45416
rect 29276 45339 29328 45348
rect 29276 45305 29285 45339
rect 29285 45305 29319 45339
rect 29319 45305 29328 45339
rect 29276 45296 29328 45305
rect 24860 45228 24912 45280
rect 27988 45228 28040 45280
rect 28448 45228 28500 45280
rect 29184 45228 29236 45280
rect 29736 45296 29788 45348
rect 30932 45296 30984 45348
rect 31392 45296 31444 45348
rect 31576 45339 31628 45348
rect 31576 45305 31585 45339
rect 31585 45305 31619 45339
rect 31619 45305 31628 45339
rect 31576 45296 31628 45305
rect 19606 45126 19658 45178
rect 19670 45126 19722 45178
rect 19734 45126 19786 45178
rect 19798 45126 19850 45178
rect 8760 45024 8812 45076
rect 13360 45024 13412 45076
rect 14740 45024 14792 45076
rect 22468 45067 22520 45076
rect 22468 45033 22477 45067
rect 22477 45033 22511 45067
rect 22511 45033 22520 45067
rect 22468 45024 22520 45033
rect 22744 45067 22796 45076
rect 22744 45033 22753 45067
rect 22753 45033 22787 45067
rect 22787 45033 22796 45067
rect 22744 45024 22796 45033
rect 23020 45024 23072 45076
rect 23756 45067 23808 45076
rect 23756 45033 23765 45067
rect 23765 45033 23799 45067
rect 23799 45033 23808 45067
rect 23756 45024 23808 45033
rect 24308 44999 24360 45008
rect 24308 44965 24317 44999
rect 24317 44965 24351 44999
rect 24351 44965 24360 44999
rect 24308 44956 24360 44965
rect 1768 44931 1820 44940
rect 1768 44897 1777 44931
rect 1777 44897 1811 44931
rect 1811 44897 1820 44931
rect 1768 44888 1820 44897
rect 13728 44931 13780 44940
rect 13728 44897 13737 44931
rect 13737 44897 13771 44931
rect 13771 44897 13780 44931
rect 13728 44888 13780 44897
rect 14096 44888 14148 44940
rect 23848 44931 23900 44940
rect 1400 44820 1452 44872
rect 1952 44820 2004 44872
rect 13084 44752 13136 44804
rect 13452 44795 13504 44804
rect 13452 44761 13461 44795
rect 13461 44761 13495 44795
rect 13495 44761 13504 44795
rect 13452 44752 13504 44761
rect 14464 44752 14516 44804
rect 3056 44727 3108 44736
rect 3056 44693 3065 44727
rect 3065 44693 3099 44727
rect 3099 44693 3108 44727
rect 3056 44684 3108 44693
rect 12900 44727 12952 44736
rect 12900 44693 12909 44727
rect 12909 44693 12943 44727
rect 12943 44693 12952 44727
rect 12900 44684 12952 44693
rect 14004 44727 14056 44736
rect 14004 44693 14013 44727
rect 14013 44693 14047 44727
rect 14047 44693 14056 44727
rect 14004 44684 14056 44693
rect 15108 44684 15160 44736
rect 23848 44897 23857 44931
rect 23857 44897 23891 44931
rect 23891 44897 23900 44931
rect 23848 44888 23900 44897
rect 24676 44888 24728 44940
rect 24952 44888 25004 44940
rect 26332 45024 26384 45076
rect 27436 45067 27488 45076
rect 27436 45033 27445 45067
rect 27445 45033 27479 45067
rect 27479 45033 27488 45067
rect 27436 45024 27488 45033
rect 28356 45024 28408 45076
rect 28540 45024 28592 45076
rect 27620 44888 27672 44940
rect 28540 44931 28592 44940
rect 28540 44897 28549 44931
rect 28549 44897 28583 44931
rect 28583 44897 28592 44931
rect 28540 44888 28592 44897
rect 29920 45024 29972 45076
rect 30472 45024 30524 45076
rect 30840 45024 30892 45076
rect 31484 45067 31536 45076
rect 31484 45033 31493 45067
rect 31493 45033 31527 45067
rect 31527 45033 31536 45067
rect 31484 45024 31536 45033
rect 29552 44931 29604 44940
rect 29552 44897 29561 44931
rect 29561 44897 29595 44931
rect 29595 44897 29604 44931
rect 29552 44888 29604 44897
rect 26700 44820 26752 44872
rect 28632 44820 28684 44872
rect 29828 44863 29880 44872
rect 29828 44829 29837 44863
rect 29837 44829 29871 44863
rect 29871 44829 29880 44863
rect 29828 44820 29880 44829
rect 26884 44752 26936 44804
rect 27712 44752 27764 44804
rect 28080 44752 28132 44804
rect 22376 44684 22428 44736
rect 25228 44684 25280 44736
rect 25780 44684 25832 44736
rect 25964 44727 26016 44736
rect 25964 44693 25973 44727
rect 25973 44693 26007 44727
rect 26007 44693 26016 44727
rect 25964 44684 26016 44693
rect 26792 44684 26844 44736
rect 27252 44684 27304 44736
rect 27804 44684 27856 44736
rect 31852 44727 31904 44736
rect 31852 44693 31861 44727
rect 31861 44693 31895 44727
rect 31895 44693 31904 44727
rect 31852 44684 31904 44693
rect 4246 44582 4298 44634
rect 4310 44582 4362 44634
rect 4374 44582 4426 44634
rect 4438 44582 4490 44634
rect 34966 44582 35018 44634
rect 35030 44582 35082 44634
rect 35094 44582 35146 44634
rect 35158 44582 35210 44634
rect 1768 44480 1820 44532
rect 8116 44523 8168 44532
rect 8116 44489 8125 44523
rect 8125 44489 8159 44523
rect 8159 44489 8168 44523
rect 8116 44480 8168 44489
rect 13728 44480 13780 44532
rect 15936 44523 15988 44532
rect 13820 44412 13872 44464
rect 14096 44412 14148 44464
rect 15936 44489 15945 44523
rect 15945 44489 15979 44523
rect 15979 44489 15988 44523
rect 15936 44480 15988 44489
rect 24676 44480 24728 44532
rect 26700 44480 26752 44532
rect 26884 44480 26936 44532
rect 28632 44480 28684 44532
rect 28908 44480 28960 44532
rect 31116 44523 31168 44532
rect 31116 44489 31125 44523
rect 31125 44489 31159 44523
rect 31159 44489 31168 44523
rect 31116 44480 31168 44489
rect 37648 44523 37700 44532
rect 37648 44489 37657 44523
rect 37657 44489 37691 44523
rect 37691 44489 37700 44523
rect 37648 44480 37700 44489
rect 16580 44412 16632 44464
rect 12532 44387 12584 44396
rect 12532 44353 12541 44387
rect 12541 44353 12575 44387
rect 12575 44353 12584 44387
rect 12532 44344 12584 44353
rect 12900 44387 12952 44396
rect 12900 44353 12909 44387
rect 12909 44353 12943 44387
rect 12943 44353 12952 44387
rect 12900 44344 12952 44353
rect 25964 44344 26016 44396
rect 2044 44319 2096 44328
rect 2044 44285 2053 44319
rect 2053 44285 2087 44319
rect 2087 44285 2096 44319
rect 2044 44276 2096 44285
rect 8300 44319 8352 44328
rect 8300 44285 8309 44319
rect 8309 44285 8343 44319
rect 8343 44285 8352 44319
rect 8300 44276 8352 44285
rect 12256 44276 12308 44328
rect 13084 44319 13136 44328
rect 13084 44285 13093 44319
rect 13093 44285 13127 44319
rect 13127 44285 13136 44319
rect 13084 44276 13136 44285
rect 10968 44208 11020 44260
rect 12532 44208 12584 44260
rect 11796 44140 11848 44192
rect 12808 44140 12860 44192
rect 15936 44276 15988 44328
rect 23848 44276 23900 44328
rect 24032 44319 24084 44328
rect 24032 44285 24041 44319
rect 24041 44285 24075 44319
rect 24075 44285 24084 44319
rect 24032 44276 24084 44285
rect 24216 44319 24268 44328
rect 24216 44285 24225 44319
rect 24225 44285 24259 44319
rect 24259 44285 24268 44319
rect 24216 44276 24268 44285
rect 26148 44276 26200 44328
rect 26608 44344 26660 44396
rect 27528 44344 27580 44396
rect 26424 44319 26476 44328
rect 26424 44285 26433 44319
rect 26433 44285 26467 44319
rect 26467 44285 26476 44319
rect 27896 44412 27948 44464
rect 27988 44412 28040 44464
rect 27712 44344 27764 44396
rect 30840 44387 30892 44396
rect 30840 44353 30849 44387
rect 30849 44353 30883 44387
rect 30883 44353 30892 44387
rect 30840 44344 30892 44353
rect 26424 44276 26476 44285
rect 28908 44276 28960 44328
rect 29092 44319 29144 44328
rect 29092 44285 29101 44319
rect 29101 44285 29135 44319
rect 29135 44285 29144 44319
rect 29092 44276 29144 44285
rect 29920 44276 29972 44328
rect 30748 44319 30800 44328
rect 30748 44285 30757 44319
rect 30757 44285 30791 44319
rect 30791 44285 30800 44319
rect 30748 44276 30800 44285
rect 34152 44276 34204 44328
rect 36084 44319 36136 44328
rect 36084 44285 36093 44319
rect 36093 44285 36127 44319
rect 36127 44285 36136 44319
rect 36084 44276 36136 44285
rect 36360 44319 36412 44328
rect 36360 44285 36369 44319
rect 36369 44285 36403 44319
rect 36403 44285 36412 44319
rect 36360 44276 36412 44285
rect 24952 44208 25004 44260
rect 25504 44208 25556 44260
rect 27344 44251 27396 44260
rect 27344 44217 27353 44251
rect 27353 44217 27387 44251
rect 27387 44217 27396 44251
rect 27344 44208 27396 44217
rect 27620 44208 27672 44260
rect 22376 44183 22428 44192
rect 22376 44149 22385 44183
rect 22385 44149 22419 44183
rect 22419 44149 22428 44183
rect 22376 44140 22428 44149
rect 29828 44208 29880 44260
rect 31116 44208 31168 44260
rect 19606 44038 19658 44090
rect 19670 44038 19722 44090
rect 19734 44038 19786 44090
rect 19798 44038 19850 44090
rect 8300 43979 8352 43988
rect 8300 43945 8309 43979
rect 8309 43945 8343 43979
rect 8343 43945 8352 43979
rect 8300 43936 8352 43945
rect 12532 43979 12584 43988
rect 12532 43945 12541 43979
rect 12541 43945 12575 43979
rect 12575 43945 12584 43979
rect 12532 43936 12584 43945
rect 11336 43800 11388 43852
rect 13084 43800 13136 43852
rect 13360 43936 13412 43988
rect 17316 43936 17368 43988
rect 15384 43843 15436 43852
rect 15384 43809 15393 43843
rect 15393 43809 15427 43843
rect 15427 43809 15436 43843
rect 15384 43800 15436 43809
rect 16580 43800 16632 43852
rect 17776 43800 17828 43852
rect 24308 43936 24360 43988
rect 24860 43936 24912 43988
rect 25964 43979 26016 43988
rect 25964 43945 25973 43979
rect 25973 43945 26007 43979
rect 26007 43945 26016 43979
rect 25964 43936 26016 43945
rect 26332 43979 26384 43988
rect 26332 43945 26341 43979
rect 26341 43945 26375 43979
rect 26375 43945 26384 43979
rect 26332 43936 26384 43945
rect 26608 43979 26660 43988
rect 26608 43945 26617 43979
rect 26617 43945 26651 43979
rect 26651 43945 26660 43979
rect 26608 43936 26660 43945
rect 27988 43979 28040 43988
rect 27988 43945 27997 43979
rect 27997 43945 28031 43979
rect 28031 43945 28040 43979
rect 27988 43936 28040 43945
rect 29368 43936 29420 43988
rect 36084 43979 36136 43988
rect 36084 43945 36093 43979
rect 36093 43945 36127 43979
rect 36127 43945 36136 43979
rect 36084 43936 36136 43945
rect 28908 43868 28960 43920
rect 20904 43843 20956 43852
rect 20904 43809 20913 43843
rect 20913 43809 20947 43843
rect 20947 43809 20956 43843
rect 20904 43800 20956 43809
rect 23848 43800 23900 43852
rect 24216 43843 24268 43852
rect 24216 43809 24225 43843
rect 24225 43809 24259 43843
rect 24259 43809 24268 43843
rect 24216 43800 24268 43809
rect 25228 43843 25280 43852
rect 25228 43809 25237 43843
rect 25237 43809 25271 43843
rect 25271 43809 25280 43843
rect 25228 43800 25280 43809
rect 25596 43800 25648 43852
rect 26516 43843 26568 43852
rect 26516 43809 26525 43843
rect 26525 43809 26559 43843
rect 26559 43809 26568 43843
rect 26516 43800 26568 43809
rect 27344 43800 27396 43852
rect 27528 43800 27580 43852
rect 27988 43800 28040 43852
rect 28356 43843 28408 43852
rect 28356 43809 28365 43843
rect 28365 43809 28399 43843
rect 28399 43809 28408 43843
rect 28356 43800 28408 43809
rect 29000 43800 29052 43852
rect 29460 43800 29512 43852
rect 29920 43800 29972 43852
rect 11152 43732 11204 43784
rect 12256 43732 12308 43784
rect 15292 43775 15344 43784
rect 15292 43741 15301 43775
rect 15301 43741 15335 43775
rect 15335 43741 15344 43775
rect 15292 43732 15344 43741
rect 21180 43775 21232 43784
rect 21180 43741 21189 43775
rect 21189 43741 21223 43775
rect 21223 43741 21232 43775
rect 21180 43732 21232 43741
rect 28632 43732 28684 43784
rect 29276 43775 29328 43784
rect 29276 43741 29285 43775
rect 29285 43741 29319 43775
rect 29319 43741 29328 43775
rect 29276 43732 29328 43741
rect 29552 43732 29604 43784
rect 23572 43707 23624 43716
rect 23572 43673 23581 43707
rect 23581 43673 23615 43707
rect 23615 43673 23624 43707
rect 23572 43664 23624 43673
rect 25044 43664 25096 43716
rect 27436 43664 27488 43716
rect 29920 43664 29972 43716
rect 15108 43596 15160 43648
rect 22008 43596 22060 43648
rect 30380 43639 30432 43648
rect 30380 43605 30389 43639
rect 30389 43605 30423 43639
rect 30423 43605 30432 43639
rect 30380 43596 30432 43605
rect 4246 43494 4298 43546
rect 4310 43494 4362 43546
rect 4374 43494 4426 43546
rect 4438 43494 4490 43546
rect 34966 43494 35018 43546
rect 35030 43494 35082 43546
rect 35094 43494 35146 43546
rect 35158 43494 35210 43546
rect 11152 43392 11204 43444
rect 11336 43435 11388 43444
rect 11336 43401 11345 43435
rect 11345 43401 11379 43435
rect 11379 43401 11388 43435
rect 11336 43392 11388 43401
rect 15292 43435 15344 43444
rect 15292 43401 15301 43435
rect 15301 43401 15335 43435
rect 15335 43401 15344 43435
rect 15292 43392 15344 43401
rect 17776 43435 17828 43444
rect 17776 43401 17785 43435
rect 17785 43401 17819 43435
rect 17819 43401 17828 43435
rect 17776 43392 17828 43401
rect 21180 43392 21232 43444
rect 27896 43435 27948 43444
rect 27896 43401 27905 43435
rect 27905 43401 27939 43435
rect 27939 43401 27948 43435
rect 27896 43392 27948 43401
rect 28080 43392 28132 43444
rect 20904 43324 20956 43376
rect 21364 43324 21416 43376
rect 28356 43392 28408 43444
rect 29184 43392 29236 43444
rect 29920 43392 29972 43444
rect 29276 43324 29328 43376
rect 13084 43299 13136 43308
rect 13084 43265 13093 43299
rect 13093 43265 13127 43299
rect 13127 43265 13136 43299
rect 13084 43256 13136 43265
rect 15384 43256 15436 43308
rect 24492 43256 24544 43308
rect 24676 43256 24728 43308
rect 25504 43299 25556 43308
rect 25504 43265 25513 43299
rect 25513 43265 25547 43299
rect 25547 43265 25556 43299
rect 25504 43256 25556 43265
rect 26700 43256 26752 43308
rect 27436 43299 27488 43308
rect 27436 43265 27445 43299
rect 27445 43265 27479 43299
rect 27479 43265 27488 43299
rect 27436 43256 27488 43265
rect 29368 43299 29420 43308
rect 29368 43265 29377 43299
rect 29377 43265 29411 43299
rect 29411 43265 29420 43299
rect 29368 43256 29420 43265
rect 30380 43324 30432 43376
rect 12624 43052 12676 43104
rect 14096 43188 14148 43240
rect 25136 43188 25188 43240
rect 26332 43188 26384 43240
rect 27160 43188 27212 43240
rect 29736 43188 29788 43240
rect 24676 43163 24728 43172
rect 24676 43129 24685 43163
rect 24685 43129 24719 43163
rect 24719 43129 24728 43163
rect 24676 43120 24728 43129
rect 27068 43120 27120 43172
rect 29460 43163 29512 43172
rect 29460 43129 29469 43163
rect 29469 43129 29503 43163
rect 29503 43129 29512 43163
rect 29460 43120 29512 43129
rect 23848 43095 23900 43104
rect 23848 43061 23857 43095
rect 23857 43061 23891 43095
rect 23891 43061 23900 43095
rect 23848 43052 23900 43061
rect 26516 43052 26568 43104
rect 19606 42950 19658 43002
rect 19670 42950 19722 43002
rect 19734 42950 19786 43002
rect 19798 42950 19850 43002
rect 14096 42891 14148 42900
rect 14096 42857 14105 42891
rect 14105 42857 14139 42891
rect 14139 42857 14148 42891
rect 14096 42848 14148 42857
rect 14740 42848 14792 42900
rect 24492 42891 24544 42900
rect 24492 42857 24501 42891
rect 24501 42857 24535 42891
rect 24535 42857 24544 42891
rect 24492 42848 24544 42857
rect 25136 42848 25188 42900
rect 27344 42848 27396 42900
rect 29000 42848 29052 42900
rect 29092 42848 29144 42900
rect 29736 42848 29788 42900
rect 26608 42780 26660 42832
rect 12900 42755 12952 42764
rect 12900 42721 12909 42755
rect 12909 42721 12943 42755
rect 12943 42721 12952 42755
rect 12900 42712 12952 42721
rect 13084 42755 13136 42764
rect 13084 42721 13093 42755
rect 13093 42721 13127 42755
rect 13127 42721 13136 42755
rect 13084 42712 13136 42721
rect 13360 42712 13412 42764
rect 14096 42712 14148 42764
rect 14832 42712 14884 42764
rect 20904 42755 20956 42764
rect 20904 42721 20913 42755
rect 20913 42721 20947 42755
rect 20947 42721 20956 42755
rect 20904 42712 20956 42721
rect 20996 42712 21048 42764
rect 22008 42712 22060 42764
rect 24124 42755 24176 42764
rect 24124 42721 24133 42755
rect 24133 42721 24167 42755
rect 24167 42721 24176 42755
rect 24124 42712 24176 42721
rect 25780 42712 25832 42764
rect 26976 42712 27028 42764
rect 27252 42755 27304 42764
rect 27252 42721 27261 42755
rect 27261 42721 27295 42755
rect 27295 42721 27304 42755
rect 27252 42712 27304 42721
rect 27620 42755 27672 42764
rect 27620 42721 27629 42755
rect 27629 42721 27663 42755
rect 27663 42721 27672 42755
rect 27620 42712 27672 42721
rect 29000 42712 29052 42764
rect 29460 42755 29512 42764
rect 29460 42721 29469 42755
rect 29469 42721 29503 42755
rect 29503 42721 29512 42755
rect 29460 42712 29512 42721
rect 34152 42712 34204 42764
rect 27528 42644 27580 42696
rect 28540 42644 28592 42696
rect 28724 42687 28776 42696
rect 28724 42653 28733 42687
rect 28733 42653 28767 42687
rect 28767 42653 28776 42687
rect 28724 42644 28776 42653
rect 29276 42644 29328 42696
rect 34060 42687 34112 42696
rect 34060 42653 34069 42687
rect 34069 42653 34103 42687
rect 34103 42653 34112 42687
rect 34060 42644 34112 42653
rect 35164 42687 35216 42696
rect 35164 42653 35173 42687
rect 35173 42653 35207 42687
rect 35207 42653 35216 42687
rect 35164 42644 35216 42653
rect 12716 42619 12768 42628
rect 12716 42585 12725 42619
rect 12725 42585 12759 42619
rect 12759 42585 12768 42619
rect 12716 42576 12768 42585
rect 19708 42508 19760 42560
rect 25228 42551 25280 42560
rect 25228 42517 25237 42551
rect 25237 42517 25271 42551
rect 25271 42517 25280 42551
rect 25228 42508 25280 42517
rect 25964 42508 26016 42560
rect 4246 42406 4298 42458
rect 4310 42406 4362 42458
rect 4374 42406 4426 42458
rect 4438 42406 4490 42458
rect 34966 42406 35018 42458
rect 35030 42406 35082 42458
rect 35094 42406 35146 42458
rect 35158 42406 35210 42458
rect 12716 42304 12768 42356
rect 12992 42304 13044 42356
rect 20996 42347 21048 42356
rect 20996 42313 21005 42347
rect 21005 42313 21039 42347
rect 21039 42313 21048 42347
rect 20996 42304 21048 42313
rect 26976 42347 27028 42356
rect 12164 42236 12216 42288
rect 13360 42236 13412 42288
rect 14372 42279 14424 42288
rect 14372 42245 14381 42279
rect 14381 42245 14415 42279
rect 14415 42245 14424 42279
rect 14372 42236 14424 42245
rect 20904 42236 20956 42288
rect 25688 42236 25740 42288
rect 12992 42211 13044 42220
rect 12992 42177 13001 42211
rect 13001 42177 13035 42211
rect 13035 42177 13044 42211
rect 12992 42168 13044 42177
rect 13728 42168 13780 42220
rect 14188 42100 14240 42152
rect 15108 42168 15160 42220
rect 26976 42313 26985 42347
rect 26985 42313 27019 42347
rect 27019 42313 27028 42347
rect 26976 42304 27028 42313
rect 27528 42304 27580 42356
rect 28080 42347 28132 42356
rect 28080 42313 28089 42347
rect 28089 42313 28123 42347
rect 28123 42313 28132 42347
rect 28080 42304 28132 42313
rect 29000 42347 29052 42356
rect 29000 42313 29009 42347
rect 29009 42313 29043 42347
rect 29043 42313 29052 42347
rect 29000 42304 29052 42313
rect 29460 42347 29512 42356
rect 29460 42313 29469 42347
rect 29469 42313 29503 42347
rect 29503 42313 29512 42347
rect 29460 42304 29512 42313
rect 34152 42347 34204 42356
rect 34152 42313 34161 42347
rect 34161 42313 34195 42347
rect 34195 42313 34204 42347
rect 34152 42304 34204 42313
rect 34612 42304 34664 42356
rect 27988 42236 28040 42288
rect 29276 42236 29328 42288
rect 26700 42168 26752 42220
rect 14740 42143 14792 42152
rect 14740 42109 14749 42143
rect 14749 42109 14783 42143
rect 14783 42109 14792 42143
rect 14740 42100 14792 42109
rect 12900 41964 12952 42016
rect 14556 41964 14608 42016
rect 15016 42100 15068 42152
rect 19708 42143 19760 42152
rect 19708 42109 19717 42143
rect 19717 42109 19751 42143
rect 19751 42109 19760 42143
rect 19708 42100 19760 42109
rect 19064 42007 19116 42016
rect 19064 41973 19073 42007
rect 19073 41973 19107 42007
rect 19107 41973 19116 42007
rect 19064 41964 19116 41973
rect 19340 42007 19392 42016
rect 19340 41973 19349 42007
rect 19349 41973 19383 42007
rect 19383 41973 19392 42007
rect 20444 42032 20496 42084
rect 24124 42100 24176 42152
rect 25688 42143 25740 42152
rect 25688 42109 25697 42143
rect 25697 42109 25731 42143
rect 25731 42109 25740 42143
rect 25688 42100 25740 42109
rect 25964 42100 26016 42152
rect 28080 42100 28132 42152
rect 24308 42007 24360 42016
rect 19340 41964 19392 41973
rect 24308 41973 24317 42007
rect 24317 41973 24351 42007
rect 24351 41973 24360 42007
rect 24308 41964 24360 41973
rect 28172 42032 28224 42084
rect 26608 41964 26660 42016
rect 28080 41964 28132 42016
rect 28264 41964 28316 42016
rect 34060 41964 34112 42016
rect 19606 41862 19658 41914
rect 19670 41862 19722 41914
rect 19734 41862 19786 41914
rect 19798 41862 19850 41914
rect 12440 41760 12492 41812
rect 13084 41760 13136 41812
rect 14188 41803 14240 41812
rect 14188 41769 14197 41803
rect 14197 41769 14231 41803
rect 14231 41769 14240 41803
rect 14188 41760 14240 41769
rect 20904 41760 20956 41812
rect 24216 41760 24268 41812
rect 25688 41760 25740 41812
rect 27160 41760 27212 41812
rect 5724 41735 5776 41744
rect 5724 41701 5733 41735
rect 5733 41701 5767 41735
rect 5767 41701 5776 41735
rect 5724 41692 5776 41701
rect 12900 41692 12952 41744
rect 4160 41624 4212 41676
rect 13452 41624 13504 41676
rect 19892 41667 19944 41676
rect 19892 41633 19901 41667
rect 19901 41633 19935 41667
rect 19935 41633 19944 41667
rect 19892 41624 19944 41633
rect 23572 41624 23624 41676
rect 3976 41556 4028 41608
rect 10324 41599 10376 41608
rect 10324 41565 10333 41599
rect 10333 41565 10367 41599
rect 10367 41565 10376 41599
rect 10324 41556 10376 41565
rect 10508 41556 10560 41608
rect 12624 41556 12676 41608
rect 12900 41556 12952 41608
rect 13084 41599 13136 41608
rect 13084 41565 13093 41599
rect 13093 41565 13127 41599
rect 13127 41565 13136 41599
rect 13084 41556 13136 41565
rect 19064 41556 19116 41608
rect 19524 41556 19576 41608
rect 23756 41599 23808 41608
rect 23756 41565 23765 41599
rect 23765 41565 23799 41599
rect 23799 41565 23808 41599
rect 23756 41556 23808 41565
rect 27252 41599 27304 41608
rect 27252 41565 27261 41599
rect 27261 41565 27295 41599
rect 27295 41565 27304 41599
rect 27252 41556 27304 41565
rect 27528 41599 27580 41608
rect 27528 41565 27537 41599
rect 27537 41565 27571 41599
rect 27571 41565 27580 41599
rect 27528 41556 27580 41565
rect 30196 41556 30248 41608
rect 11612 41420 11664 41472
rect 19432 41420 19484 41472
rect 24860 41463 24912 41472
rect 24860 41429 24869 41463
rect 24869 41429 24903 41463
rect 24903 41429 24912 41463
rect 24860 41420 24912 41429
rect 29460 41420 29512 41472
rect 30012 41420 30064 41472
rect 4246 41318 4298 41370
rect 4310 41318 4362 41370
rect 4374 41318 4426 41370
rect 4438 41318 4490 41370
rect 34966 41318 35018 41370
rect 35030 41318 35082 41370
rect 35094 41318 35146 41370
rect 35158 41318 35210 41370
rect 10508 41216 10560 41268
rect 23756 41216 23808 41268
rect 27528 41216 27580 41268
rect 27712 41259 27764 41268
rect 27712 41225 27721 41259
rect 27721 41225 27755 41259
rect 27755 41225 27764 41259
rect 27712 41216 27764 41225
rect 29184 41216 29236 41268
rect 34704 41216 34756 41268
rect 19892 41148 19944 41200
rect 23572 41148 23624 41200
rect 34888 41148 34940 41200
rect 30012 41080 30064 41132
rect 3976 40944 4028 40996
rect 13084 40944 13136 40996
rect 13820 40944 13872 40996
rect 19340 41012 19392 41064
rect 19892 41012 19944 41064
rect 20904 41012 20956 41064
rect 21180 41012 21232 41064
rect 21364 41055 21416 41064
rect 21364 41021 21373 41055
rect 21373 41021 21407 41055
rect 21407 41021 21416 41055
rect 21364 41012 21416 41021
rect 30196 41055 30248 41064
rect 30196 41021 30205 41055
rect 30205 41021 30239 41055
rect 30239 41021 30248 41055
rect 30196 41012 30248 41021
rect 19524 40944 19576 40996
rect 29644 40944 29696 40996
rect 4068 40919 4120 40928
rect 4068 40885 4077 40919
rect 4077 40885 4111 40919
rect 4111 40885 4120 40919
rect 4068 40876 4120 40885
rect 10324 40876 10376 40928
rect 11336 40876 11388 40928
rect 13452 40919 13504 40928
rect 13452 40885 13461 40919
rect 13461 40885 13495 40919
rect 13495 40885 13504 40919
rect 13452 40876 13504 40885
rect 18236 40919 18288 40928
rect 18236 40885 18245 40919
rect 18245 40885 18279 40919
rect 18279 40885 18288 40919
rect 18236 40876 18288 40885
rect 18972 40919 19024 40928
rect 18972 40885 18981 40919
rect 18981 40885 19015 40919
rect 19015 40885 19024 40919
rect 18972 40876 19024 40885
rect 20260 40876 20312 40928
rect 22468 40919 22520 40928
rect 22468 40885 22477 40919
rect 22477 40885 22511 40919
rect 22511 40885 22520 40919
rect 22468 40876 22520 40885
rect 19606 40774 19658 40826
rect 19670 40774 19722 40826
rect 19734 40774 19786 40826
rect 19798 40774 19850 40826
rect 20720 40672 20772 40724
rect 21180 40672 21232 40724
rect 23480 40715 23532 40724
rect 2412 40647 2464 40656
rect 2412 40613 2421 40647
rect 2421 40613 2455 40647
rect 2455 40613 2464 40647
rect 2412 40604 2464 40613
rect 4068 40604 4120 40656
rect 13452 40604 13504 40656
rect 13820 40579 13872 40588
rect 2228 40468 2280 40520
rect 13820 40545 13829 40579
rect 13829 40545 13863 40579
rect 13863 40545 13872 40579
rect 13820 40536 13872 40545
rect 15936 40579 15988 40588
rect 15936 40545 15945 40579
rect 15945 40545 15979 40579
rect 15979 40545 15988 40579
rect 15936 40536 15988 40545
rect 17868 40536 17920 40588
rect 18972 40579 19024 40588
rect 18972 40545 18981 40579
rect 18981 40545 19015 40579
rect 19015 40545 19024 40579
rect 18972 40536 19024 40545
rect 19340 40579 19392 40588
rect 19340 40545 19349 40579
rect 19349 40545 19383 40579
rect 19383 40545 19392 40579
rect 19340 40536 19392 40545
rect 19708 40579 19760 40588
rect 19708 40545 19717 40579
rect 19717 40545 19751 40579
rect 19751 40545 19760 40579
rect 19708 40536 19760 40545
rect 19984 40579 20036 40588
rect 19984 40545 19993 40579
rect 19993 40545 20027 40579
rect 20027 40545 20036 40579
rect 19984 40536 20036 40545
rect 20076 40579 20128 40588
rect 20076 40545 20085 40579
rect 20085 40545 20119 40579
rect 20119 40545 20128 40579
rect 20076 40536 20128 40545
rect 20260 40579 20312 40588
rect 20260 40545 20269 40579
rect 20269 40545 20303 40579
rect 20303 40545 20312 40579
rect 20260 40536 20312 40545
rect 21088 40536 21140 40588
rect 23480 40681 23489 40715
rect 23489 40681 23523 40715
rect 23523 40681 23532 40715
rect 23480 40672 23532 40681
rect 23388 40536 23440 40588
rect 34888 40536 34940 40588
rect 35532 40536 35584 40588
rect 11336 40511 11388 40520
rect 11336 40477 11345 40511
rect 11345 40477 11379 40511
rect 11379 40477 11388 40511
rect 11336 40468 11388 40477
rect 11612 40511 11664 40520
rect 11612 40477 11621 40511
rect 11621 40477 11655 40511
rect 11655 40477 11664 40511
rect 11612 40468 11664 40477
rect 17776 40511 17828 40520
rect 17776 40477 17785 40511
rect 17785 40477 17819 40511
rect 17819 40477 17828 40511
rect 17776 40468 17828 40477
rect 34612 40468 34664 40520
rect 35440 40468 35492 40520
rect 19708 40400 19760 40452
rect 20260 40400 20312 40452
rect 1952 40332 2004 40384
rect 14004 40375 14056 40384
rect 14004 40341 14013 40375
rect 14013 40341 14047 40375
rect 14047 40341 14056 40375
rect 14004 40332 14056 40341
rect 15200 40332 15252 40384
rect 19340 40332 19392 40384
rect 21364 40375 21416 40384
rect 21364 40341 21373 40375
rect 21373 40341 21407 40375
rect 21407 40341 21416 40375
rect 21364 40332 21416 40341
rect 25688 40375 25740 40384
rect 25688 40341 25697 40375
rect 25697 40341 25731 40375
rect 25731 40341 25740 40375
rect 25688 40332 25740 40341
rect 28448 40332 28500 40384
rect 30012 40332 30064 40384
rect 35716 40332 35768 40384
rect 4246 40230 4298 40282
rect 4310 40230 4362 40282
rect 4374 40230 4426 40282
rect 4438 40230 4490 40282
rect 34966 40230 35018 40282
rect 35030 40230 35082 40282
rect 35094 40230 35146 40282
rect 35158 40230 35210 40282
rect 17132 40171 17184 40180
rect 17132 40137 17141 40171
rect 17141 40137 17175 40171
rect 17175 40137 17184 40171
rect 17132 40128 17184 40137
rect 17868 40128 17920 40180
rect 23388 40128 23440 40180
rect 35440 40171 35492 40180
rect 35440 40137 35449 40171
rect 35449 40137 35483 40171
rect 35483 40137 35492 40171
rect 35440 40128 35492 40137
rect 9680 40060 9732 40112
rect 11336 40060 11388 40112
rect 35532 40060 35584 40112
rect 1952 39992 2004 40044
rect 20076 39992 20128 40044
rect 21364 40035 21416 40044
rect 21364 40001 21373 40035
rect 21373 40001 21407 40035
rect 21407 40001 21416 40035
rect 21364 39992 21416 40001
rect 25688 39992 25740 40044
rect 26516 39992 26568 40044
rect 1676 39924 1728 39976
rect 13084 39967 13136 39976
rect 13084 39933 13093 39967
rect 13093 39933 13127 39967
rect 13127 39933 13136 39967
rect 13084 39924 13136 39933
rect 15936 39967 15988 39976
rect 15936 39933 15945 39967
rect 15945 39933 15979 39967
rect 15979 39933 15988 39967
rect 16488 39967 16540 39976
rect 15936 39924 15988 39933
rect 16488 39933 16497 39967
rect 16497 39933 16531 39967
rect 16531 39933 16540 39967
rect 16488 39924 16540 39933
rect 17868 39967 17920 39976
rect 17868 39933 17877 39967
rect 17877 39933 17911 39967
rect 17911 39933 17920 39967
rect 17868 39924 17920 39933
rect 21180 39924 21232 39976
rect 23572 39924 23624 39976
rect 25136 39967 25188 39976
rect 25136 39933 25145 39967
rect 25145 39933 25179 39967
rect 25179 39933 25188 39967
rect 25136 39924 25188 39933
rect 4068 39856 4120 39908
rect 11612 39788 11664 39840
rect 12440 39788 12492 39840
rect 13452 39788 13504 39840
rect 13820 39788 13872 39840
rect 15476 39788 15528 39840
rect 15936 39788 15988 39840
rect 18604 39831 18656 39840
rect 18604 39797 18613 39831
rect 18613 39797 18647 39831
rect 18647 39797 18656 39831
rect 20352 39856 20404 39908
rect 20536 39899 20588 39908
rect 20536 39865 20545 39899
rect 20545 39865 20579 39899
rect 20579 39865 20588 39899
rect 20536 39856 20588 39865
rect 25780 39856 25832 39908
rect 18604 39788 18656 39797
rect 20996 39788 21048 39840
rect 26884 39924 26936 39976
rect 19606 39686 19658 39738
rect 19670 39686 19722 39738
rect 19734 39686 19786 39738
rect 19798 39686 19850 39738
rect 2412 39584 2464 39636
rect 19064 39627 19116 39636
rect 19064 39593 19073 39627
rect 19073 39593 19107 39627
rect 19107 39593 19116 39627
rect 19064 39584 19116 39593
rect 21088 39627 21140 39636
rect 21088 39593 21097 39627
rect 21097 39593 21131 39627
rect 21131 39593 21140 39627
rect 21088 39584 21140 39593
rect 21364 39584 21416 39636
rect 25136 39627 25188 39636
rect 25136 39593 25145 39627
rect 25145 39593 25179 39627
rect 25179 39593 25188 39627
rect 25136 39584 25188 39593
rect 1584 39559 1636 39568
rect 1584 39525 1593 39559
rect 1593 39525 1627 39559
rect 1627 39525 1636 39559
rect 1584 39516 1636 39525
rect 19984 39559 20036 39568
rect 19984 39525 19993 39559
rect 19993 39525 20027 39559
rect 20027 39525 20036 39559
rect 19984 39516 20036 39525
rect 26516 39559 26568 39568
rect 26516 39525 26525 39559
rect 26525 39525 26559 39559
rect 26559 39525 26568 39559
rect 26516 39516 26568 39525
rect 15568 39491 15620 39500
rect 15568 39457 15577 39491
rect 15577 39457 15611 39491
rect 15611 39457 15620 39491
rect 15568 39448 15620 39457
rect 16580 39448 16632 39500
rect 18236 39491 18288 39500
rect 18236 39457 18245 39491
rect 18245 39457 18279 39491
rect 18279 39457 18288 39491
rect 18236 39448 18288 39457
rect 19892 39491 19944 39500
rect 19892 39457 19901 39491
rect 19901 39457 19935 39491
rect 19935 39457 19944 39491
rect 19892 39448 19944 39457
rect 21180 39448 21232 39500
rect 25044 39491 25096 39500
rect 25044 39457 25053 39491
rect 25053 39457 25087 39491
rect 25087 39457 25096 39491
rect 25044 39448 25096 39457
rect 26608 39491 26660 39500
rect 26608 39457 26617 39491
rect 26617 39457 26651 39491
rect 26651 39457 26660 39491
rect 26608 39448 26660 39457
rect 35716 39448 35768 39500
rect 14188 39380 14240 39432
rect 16028 39423 16080 39432
rect 15108 39312 15160 39364
rect 16028 39389 16037 39423
rect 16037 39389 16071 39423
rect 16071 39389 16080 39423
rect 16028 39380 16080 39389
rect 16120 39380 16172 39432
rect 17776 39423 17828 39432
rect 17776 39389 17785 39423
rect 17785 39389 17819 39423
rect 17819 39389 17828 39423
rect 17776 39380 17828 39389
rect 16212 39312 16264 39364
rect 18052 39312 18104 39364
rect 21732 39380 21784 39432
rect 34704 39423 34756 39432
rect 34704 39389 34713 39423
rect 34713 39389 34747 39423
rect 34747 39389 34756 39423
rect 34704 39380 34756 39389
rect 2228 39244 2280 39296
rect 14280 39244 14332 39296
rect 15016 39287 15068 39296
rect 15016 39253 15025 39287
rect 15025 39253 15059 39287
rect 15059 39253 15068 39287
rect 15016 39244 15068 39253
rect 16304 39287 16356 39296
rect 16304 39253 16313 39287
rect 16313 39253 16347 39287
rect 16347 39253 16356 39287
rect 16304 39244 16356 39253
rect 16580 39244 16632 39296
rect 20260 39244 20312 39296
rect 22468 39244 22520 39296
rect 4246 39142 4298 39194
rect 4310 39142 4362 39194
rect 4374 39142 4426 39194
rect 4438 39142 4490 39194
rect 34966 39142 35018 39194
rect 35030 39142 35082 39194
rect 35094 39142 35146 39194
rect 35158 39142 35210 39194
rect 9404 39083 9456 39092
rect 9404 39049 9413 39083
rect 9413 39049 9447 39083
rect 9447 39049 9456 39083
rect 9404 39040 9456 39049
rect 15568 39040 15620 39092
rect 16764 39083 16816 39092
rect 1676 38947 1728 38956
rect 1676 38913 1685 38947
rect 1685 38913 1719 38947
rect 1719 38913 1728 38947
rect 1676 38904 1728 38913
rect 2412 38904 2464 38956
rect 16764 39049 16773 39083
rect 16773 39049 16807 39083
rect 16807 39049 16816 39083
rect 16764 39040 16816 39049
rect 17776 39083 17828 39092
rect 17776 39049 17785 39083
rect 17785 39049 17819 39083
rect 17819 39049 17828 39083
rect 17776 39040 17828 39049
rect 19340 39083 19392 39092
rect 19340 39049 19349 39083
rect 19349 39049 19383 39083
rect 19383 39049 19392 39083
rect 19340 39040 19392 39049
rect 20996 39083 21048 39092
rect 20996 39049 21005 39083
rect 21005 39049 21039 39083
rect 21039 39049 21048 39083
rect 20996 39040 21048 39049
rect 22468 39040 22520 39092
rect 26608 39040 26660 39092
rect 29460 39040 29512 39092
rect 18052 38947 18104 38956
rect 1952 38836 2004 38888
rect 9404 38836 9456 38888
rect 9680 38836 9732 38888
rect 13912 38836 13964 38888
rect 14280 38879 14332 38888
rect 14280 38845 14289 38879
rect 14289 38845 14323 38879
rect 14323 38845 14332 38879
rect 14280 38836 14332 38845
rect 14924 38836 14976 38888
rect 15108 38879 15160 38888
rect 15108 38845 15117 38879
rect 15117 38845 15151 38879
rect 15151 38845 15160 38879
rect 15108 38836 15160 38845
rect 18052 38913 18061 38947
rect 18061 38913 18095 38947
rect 18095 38913 18104 38947
rect 18052 38904 18104 38913
rect 18420 38904 18472 38956
rect 19984 38972 20036 39024
rect 19064 38947 19116 38956
rect 19064 38913 19073 38947
rect 19073 38913 19107 38947
rect 19107 38913 19116 38947
rect 19064 38904 19116 38913
rect 16120 38836 16172 38888
rect 16304 38836 16356 38888
rect 16488 38879 16540 38888
rect 16488 38845 16497 38879
rect 16497 38845 16531 38879
rect 16531 38845 16540 38879
rect 16488 38836 16540 38845
rect 16580 38879 16632 38888
rect 16580 38845 16589 38879
rect 16589 38845 16623 38879
rect 16623 38845 16632 38879
rect 16580 38836 16632 38845
rect 19156 38836 19208 38888
rect 20076 38836 20128 38888
rect 27252 38972 27304 39024
rect 20260 38947 20312 38956
rect 20260 38913 20269 38947
rect 20269 38913 20303 38947
rect 20303 38913 20312 38947
rect 20260 38904 20312 38913
rect 25136 38904 25188 38956
rect 26056 38904 26108 38956
rect 26516 38904 26568 38956
rect 27160 38904 27212 38956
rect 35716 39040 35768 39092
rect 25412 38879 25464 38888
rect 25412 38845 25421 38879
rect 25421 38845 25455 38879
rect 25455 38845 25464 38879
rect 25412 38836 25464 38845
rect 25780 38879 25832 38888
rect 25780 38845 25789 38879
rect 25789 38845 25823 38879
rect 25823 38845 25832 38879
rect 25780 38836 25832 38845
rect 26884 38836 26936 38888
rect 28080 38836 28132 38888
rect 29552 38836 29604 38888
rect 29920 38879 29972 38888
rect 29920 38845 29929 38879
rect 29929 38845 29963 38879
rect 29963 38845 29972 38879
rect 29920 38836 29972 38845
rect 19892 38811 19944 38820
rect 19892 38777 19901 38811
rect 19901 38777 19935 38811
rect 19935 38777 19944 38811
rect 19892 38768 19944 38777
rect 20996 38768 21048 38820
rect 21732 38768 21784 38820
rect 22468 38768 22520 38820
rect 26792 38811 26844 38820
rect 26792 38777 26801 38811
rect 26801 38777 26835 38811
rect 26835 38777 26844 38811
rect 26792 38768 26844 38777
rect 2780 38743 2832 38752
rect 2780 38709 2789 38743
rect 2789 38709 2823 38743
rect 2823 38709 2832 38743
rect 11152 38743 11204 38752
rect 2780 38700 2832 38709
rect 11152 38709 11161 38743
rect 11161 38709 11195 38743
rect 11195 38709 11204 38743
rect 11152 38700 11204 38709
rect 13084 38700 13136 38752
rect 16212 38700 16264 38752
rect 21640 38743 21692 38752
rect 21640 38709 21649 38743
rect 21649 38709 21683 38743
rect 21683 38709 21692 38743
rect 21640 38700 21692 38709
rect 30472 38700 30524 38752
rect 19606 38598 19658 38650
rect 19670 38598 19722 38650
rect 19734 38598 19786 38650
rect 19798 38598 19850 38650
rect 1676 38539 1728 38548
rect 1676 38505 1685 38539
rect 1685 38505 1719 38539
rect 1719 38505 1728 38539
rect 1676 38496 1728 38505
rect 1952 38539 2004 38548
rect 1952 38505 1961 38539
rect 1961 38505 1995 38539
rect 1995 38505 2004 38539
rect 1952 38496 2004 38505
rect 13728 38496 13780 38548
rect 13912 38496 13964 38548
rect 15936 38539 15988 38548
rect 15936 38505 15945 38539
rect 15945 38505 15979 38539
rect 15979 38505 15988 38539
rect 15936 38496 15988 38505
rect 19340 38496 19392 38548
rect 19984 38539 20036 38548
rect 19984 38505 19993 38539
rect 19993 38505 20027 38539
rect 20027 38505 20036 38539
rect 19984 38496 20036 38505
rect 20996 38496 21048 38548
rect 21180 38496 21232 38548
rect 25044 38496 25096 38548
rect 26884 38539 26936 38548
rect 26884 38505 26893 38539
rect 26893 38505 26927 38539
rect 26927 38505 26936 38539
rect 26884 38496 26936 38505
rect 27160 38539 27212 38548
rect 27160 38505 27169 38539
rect 27169 38505 27203 38539
rect 27203 38505 27212 38539
rect 27160 38496 27212 38505
rect 29920 38539 29972 38548
rect 29920 38505 29929 38539
rect 29929 38505 29963 38539
rect 29963 38505 29972 38539
rect 29920 38496 29972 38505
rect 12164 38428 12216 38480
rect 18052 38428 18104 38480
rect 25320 38428 25372 38480
rect 11796 38403 11848 38412
rect 11796 38369 11805 38403
rect 11805 38369 11839 38403
rect 11839 38369 11848 38403
rect 11796 38360 11848 38369
rect 11980 38403 12032 38412
rect 11980 38369 11989 38403
rect 11989 38369 12023 38403
rect 12023 38369 12032 38403
rect 11980 38360 12032 38369
rect 12256 38360 12308 38412
rect 12624 38360 12676 38412
rect 14096 38360 14148 38412
rect 14372 38403 14424 38412
rect 14372 38369 14381 38403
rect 14381 38369 14415 38403
rect 14415 38369 14424 38403
rect 14372 38360 14424 38369
rect 16028 38403 16080 38412
rect 16028 38369 16037 38403
rect 16037 38369 16071 38403
rect 16071 38369 16080 38403
rect 16028 38360 16080 38369
rect 16120 38360 16172 38412
rect 19064 38403 19116 38412
rect 11336 38335 11388 38344
rect 11336 38301 11345 38335
rect 11345 38301 11379 38335
rect 11379 38301 11388 38335
rect 11336 38292 11388 38301
rect 13360 38335 13412 38344
rect 13360 38301 13369 38335
rect 13369 38301 13403 38335
rect 13403 38301 13412 38335
rect 13360 38292 13412 38301
rect 13912 38335 13964 38344
rect 13912 38301 13921 38335
rect 13921 38301 13955 38335
rect 13955 38301 13964 38335
rect 19064 38369 19073 38403
rect 19073 38369 19107 38403
rect 19107 38369 19116 38403
rect 19064 38360 19116 38369
rect 19156 38360 19208 38412
rect 20444 38360 20496 38412
rect 20996 38403 21048 38412
rect 20996 38369 21005 38403
rect 21005 38369 21039 38403
rect 21039 38369 21048 38403
rect 20996 38360 21048 38369
rect 24308 38360 24360 38412
rect 13912 38292 13964 38301
rect 17408 38292 17460 38344
rect 17868 38292 17920 38344
rect 16856 38267 16908 38276
rect 16856 38233 16865 38267
rect 16865 38233 16899 38267
rect 16899 38233 16908 38267
rect 16856 38224 16908 38233
rect 18236 38224 18288 38276
rect 21088 38292 21140 38344
rect 24492 38335 24544 38344
rect 24492 38301 24501 38335
rect 24501 38301 24535 38335
rect 24535 38301 24544 38335
rect 24492 38292 24544 38301
rect 28080 38360 28132 38412
rect 25504 38292 25556 38344
rect 28356 38292 28408 38344
rect 11060 38156 11112 38208
rect 12256 38156 12308 38208
rect 12532 38156 12584 38208
rect 14740 38199 14792 38208
rect 14740 38165 14749 38199
rect 14749 38165 14783 38199
rect 14783 38165 14792 38199
rect 14740 38156 14792 38165
rect 15108 38199 15160 38208
rect 15108 38165 15117 38199
rect 15117 38165 15151 38199
rect 15151 38165 15160 38199
rect 15108 38156 15160 38165
rect 15292 38156 15344 38208
rect 18788 38156 18840 38208
rect 24124 38199 24176 38208
rect 24124 38165 24133 38199
rect 24133 38165 24167 38199
rect 24167 38165 24176 38199
rect 24124 38156 24176 38165
rect 27712 38156 27764 38208
rect 4246 38054 4298 38106
rect 4310 38054 4362 38106
rect 4374 38054 4426 38106
rect 4438 38054 4490 38106
rect 34966 38054 35018 38106
rect 35030 38054 35082 38106
rect 35094 38054 35146 38106
rect 35158 38054 35210 38106
rect 12624 37952 12676 38004
rect 13636 37995 13688 38004
rect 13636 37961 13645 37995
rect 13645 37961 13679 37995
rect 13679 37961 13688 37995
rect 13636 37952 13688 37961
rect 13912 37952 13964 38004
rect 16028 37952 16080 38004
rect 17408 37995 17460 38004
rect 17408 37961 17417 37995
rect 17417 37961 17451 37995
rect 17451 37961 17460 37995
rect 17408 37952 17460 37961
rect 17868 37995 17920 38004
rect 17868 37961 17877 37995
rect 17877 37961 17911 37995
rect 17911 37961 17920 37995
rect 17868 37952 17920 37961
rect 19800 37995 19852 38004
rect 19800 37961 19809 37995
rect 19809 37961 19843 37995
rect 19843 37961 19852 37995
rect 19800 37952 19852 37961
rect 24308 37952 24360 38004
rect 25504 37952 25556 38004
rect 11796 37884 11848 37936
rect 17132 37884 17184 37936
rect 12532 37859 12584 37868
rect 12532 37825 12541 37859
rect 12541 37825 12575 37859
rect 12575 37825 12584 37859
rect 12532 37816 12584 37825
rect 14280 37816 14332 37868
rect 11980 37680 12032 37732
rect 13544 37748 13596 37800
rect 15936 37816 15988 37868
rect 16580 37791 16632 37800
rect 16580 37757 16589 37791
rect 16589 37757 16623 37791
rect 16623 37757 16632 37791
rect 16580 37748 16632 37757
rect 16948 37791 17000 37800
rect 16948 37757 16957 37791
rect 16957 37757 16991 37791
rect 16991 37757 17000 37791
rect 16948 37748 17000 37757
rect 17132 37791 17184 37800
rect 17132 37757 17141 37791
rect 17141 37757 17175 37791
rect 17175 37757 17184 37791
rect 17132 37748 17184 37757
rect 18236 37791 18288 37800
rect 18236 37757 18245 37791
rect 18245 37757 18279 37791
rect 18279 37757 18288 37791
rect 18236 37748 18288 37757
rect 18420 37748 18472 37800
rect 18788 37791 18840 37800
rect 18788 37757 18797 37791
rect 18797 37757 18831 37791
rect 18831 37757 18840 37791
rect 18788 37748 18840 37757
rect 18880 37791 18932 37800
rect 18880 37757 18889 37791
rect 18889 37757 18923 37791
rect 18923 37757 18932 37791
rect 18880 37748 18932 37757
rect 19064 37748 19116 37800
rect 20076 37748 20128 37800
rect 28080 37952 28132 38004
rect 28356 37952 28408 38004
rect 29552 37952 29604 38004
rect 21548 37816 21600 37868
rect 27252 37816 27304 37868
rect 20812 37791 20864 37800
rect 15936 37723 15988 37732
rect 15936 37689 15945 37723
rect 15945 37689 15979 37723
rect 15979 37689 15988 37723
rect 15936 37680 15988 37689
rect 19984 37723 20036 37732
rect 19984 37689 19993 37723
rect 19993 37689 20027 37723
rect 20027 37689 20036 37723
rect 19984 37680 20036 37689
rect 20352 37680 20404 37732
rect 20812 37757 20821 37791
rect 20821 37757 20855 37791
rect 20855 37757 20864 37791
rect 20812 37748 20864 37757
rect 25412 37791 25464 37800
rect 25412 37757 25421 37791
rect 25421 37757 25455 37791
rect 25455 37757 25464 37791
rect 25412 37748 25464 37757
rect 25688 37791 25740 37800
rect 25688 37757 25697 37791
rect 25697 37757 25731 37791
rect 25731 37757 25740 37791
rect 25688 37748 25740 37757
rect 26792 37748 26844 37800
rect 27712 37791 27764 37800
rect 27712 37757 27721 37791
rect 27721 37757 27755 37791
rect 27755 37757 27764 37791
rect 27712 37748 27764 37757
rect 25964 37723 26016 37732
rect 25964 37689 25973 37723
rect 25973 37689 26007 37723
rect 26007 37689 26016 37723
rect 25964 37680 26016 37689
rect 12808 37612 12860 37664
rect 13268 37612 13320 37664
rect 16856 37612 16908 37664
rect 17960 37612 18012 37664
rect 19156 37612 19208 37664
rect 20444 37612 20496 37664
rect 21088 37612 21140 37664
rect 26884 37612 26936 37664
rect 19606 37510 19658 37562
rect 19670 37510 19722 37562
rect 19734 37510 19786 37562
rect 19798 37510 19850 37562
rect 11980 37408 12032 37460
rect 13544 37408 13596 37460
rect 18052 37408 18104 37460
rect 18420 37451 18472 37460
rect 18420 37417 18429 37451
rect 18429 37417 18463 37451
rect 18463 37417 18472 37451
rect 18420 37408 18472 37417
rect 18512 37408 18564 37460
rect 20352 37408 20404 37460
rect 20812 37408 20864 37460
rect 25688 37408 25740 37460
rect 27252 37408 27304 37460
rect 33508 37451 33560 37460
rect 33508 37417 33517 37451
rect 33517 37417 33551 37451
rect 33551 37417 33560 37451
rect 33508 37408 33560 37417
rect 14740 37340 14792 37392
rect 15752 37340 15804 37392
rect 17960 37340 18012 37392
rect 9404 37272 9456 37324
rect 11060 37315 11112 37324
rect 11060 37281 11069 37315
rect 11069 37281 11103 37315
rect 11103 37281 11112 37315
rect 11060 37272 11112 37281
rect 13728 37315 13780 37324
rect 11888 37204 11940 37256
rect 13728 37281 13737 37315
rect 13737 37281 13771 37315
rect 13771 37281 13780 37315
rect 13728 37272 13780 37281
rect 14280 37272 14332 37324
rect 15384 37272 15436 37324
rect 16120 37315 16172 37324
rect 16120 37281 16129 37315
rect 16129 37281 16163 37315
rect 16163 37281 16172 37315
rect 16120 37272 16172 37281
rect 16948 37315 17000 37324
rect 16948 37281 16957 37315
rect 16957 37281 16991 37315
rect 16991 37281 17000 37315
rect 16948 37272 17000 37281
rect 17316 37315 17368 37324
rect 17316 37281 17325 37315
rect 17325 37281 17359 37315
rect 17359 37281 17368 37315
rect 17316 37272 17368 37281
rect 18236 37272 18288 37324
rect 19984 37340 20036 37392
rect 18972 37315 19024 37324
rect 18972 37281 18981 37315
rect 18981 37281 19015 37315
rect 19015 37281 19024 37315
rect 18972 37272 19024 37281
rect 19156 37315 19208 37324
rect 19156 37281 19165 37315
rect 19165 37281 19199 37315
rect 19199 37281 19208 37315
rect 19156 37272 19208 37281
rect 23848 37272 23900 37324
rect 24952 37272 25004 37324
rect 27436 37315 27488 37324
rect 27436 37281 27445 37315
rect 27445 37281 27479 37315
rect 27479 37281 27488 37315
rect 27436 37272 27488 37281
rect 32220 37272 32272 37324
rect 13360 37204 13412 37256
rect 14832 37204 14884 37256
rect 16856 37247 16908 37256
rect 16856 37213 16865 37247
rect 16865 37213 16899 37247
rect 16899 37213 16908 37247
rect 16856 37204 16908 37213
rect 17132 37204 17184 37256
rect 23112 37247 23164 37256
rect 23112 37213 23121 37247
rect 23121 37213 23155 37247
rect 23155 37213 23164 37247
rect 23112 37204 23164 37213
rect 23296 37204 23348 37256
rect 32496 37204 32548 37256
rect 11796 37136 11848 37188
rect 14372 37136 14424 37188
rect 16212 37136 16264 37188
rect 17592 37136 17644 37188
rect 12808 37111 12860 37120
rect 12808 37077 12817 37111
rect 12817 37077 12851 37111
rect 12851 37077 12860 37111
rect 12808 37068 12860 37077
rect 14740 37111 14792 37120
rect 14740 37077 14749 37111
rect 14749 37077 14783 37111
rect 14783 37077 14792 37111
rect 14740 37068 14792 37077
rect 15660 37068 15712 37120
rect 24216 37068 24268 37120
rect 4246 36966 4298 37018
rect 4310 36966 4362 37018
rect 4374 36966 4426 37018
rect 4438 36966 4490 37018
rect 34966 36966 35018 37018
rect 35030 36966 35082 37018
rect 35094 36966 35146 37018
rect 35158 36966 35210 37018
rect 11060 36864 11112 36916
rect 12716 36864 12768 36916
rect 13176 36864 13228 36916
rect 14464 36864 14516 36916
rect 14740 36864 14792 36916
rect 15384 36864 15436 36916
rect 16028 36864 16080 36916
rect 17132 36864 17184 36916
rect 11428 36796 11480 36848
rect 15108 36796 15160 36848
rect 11796 36728 11848 36780
rect 10140 36524 10192 36576
rect 12624 36703 12676 36712
rect 12624 36669 12633 36703
rect 12633 36669 12667 36703
rect 12667 36669 12676 36703
rect 12624 36660 12676 36669
rect 12808 36728 12860 36780
rect 14648 36728 14700 36780
rect 13360 36660 13412 36712
rect 14924 36703 14976 36712
rect 14924 36669 14933 36703
rect 14933 36669 14967 36703
rect 14967 36669 14976 36703
rect 14924 36660 14976 36669
rect 15200 36703 15252 36712
rect 15200 36669 15209 36703
rect 15209 36669 15243 36703
rect 15243 36669 15252 36703
rect 15200 36660 15252 36669
rect 15660 36703 15712 36712
rect 13636 36592 13688 36644
rect 14464 36592 14516 36644
rect 15016 36592 15068 36644
rect 15660 36669 15669 36703
rect 15669 36669 15703 36703
rect 15703 36669 15712 36703
rect 15660 36660 15712 36669
rect 17776 36864 17828 36916
rect 19984 36864 20036 36916
rect 20260 36864 20312 36916
rect 21640 36907 21692 36916
rect 21640 36873 21649 36907
rect 21649 36873 21683 36907
rect 21683 36873 21692 36907
rect 21640 36864 21692 36873
rect 23296 36864 23348 36916
rect 26792 36907 26844 36916
rect 26792 36873 26801 36907
rect 26801 36873 26835 36907
rect 26835 36873 26844 36907
rect 26792 36864 26844 36873
rect 27436 36907 27488 36916
rect 27436 36873 27445 36907
rect 27445 36873 27479 36907
rect 27479 36873 27488 36907
rect 27436 36864 27488 36873
rect 32496 36907 32548 36916
rect 32496 36873 32505 36907
rect 32505 36873 32539 36907
rect 32539 36873 32548 36907
rect 32496 36864 32548 36873
rect 18236 36703 18288 36712
rect 18236 36669 18245 36703
rect 18245 36669 18279 36703
rect 18279 36669 18288 36703
rect 18236 36660 18288 36669
rect 10600 36567 10652 36576
rect 10600 36533 10609 36567
rect 10609 36533 10643 36567
rect 10643 36533 10652 36567
rect 10600 36524 10652 36533
rect 17408 36592 17460 36644
rect 17592 36592 17644 36644
rect 18880 36660 18932 36712
rect 25412 36703 25464 36712
rect 18512 36524 18564 36576
rect 19064 36524 19116 36576
rect 25412 36669 25421 36703
rect 25421 36669 25455 36703
rect 25455 36669 25464 36703
rect 25412 36660 25464 36669
rect 25688 36703 25740 36712
rect 25688 36669 25697 36703
rect 25697 36669 25731 36703
rect 25731 36669 25740 36703
rect 25688 36660 25740 36669
rect 19984 36524 20036 36576
rect 20904 36567 20956 36576
rect 20904 36533 20913 36567
rect 20913 36533 20947 36567
rect 20947 36533 20956 36567
rect 20904 36524 20956 36533
rect 21180 36524 21232 36576
rect 23112 36524 23164 36576
rect 23296 36524 23348 36576
rect 32128 36567 32180 36576
rect 32128 36533 32137 36567
rect 32137 36533 32171 36567
rect 32171 36533 32180 36567
rect 32128 36524 32180 36533
rect 19606 36422 19658 36474
rect 19670 36422 19722 36474
rect 19734 36422 19786 36474
rect 19798 36422 19850 36474
rect 10968 36363 11020 36372
rect 10968 36329 10977 36363
rect 10977 36329 11011 36363
rect 11011 36329 11020 36363
rect 10968 36320 11020 36329
rect 11888 36320 11940 36372
rect 12256 36320 12308 36372
rect 14832 36363 14884 36372
rect 14832 36329 14841 36363
rect 14841 36329 14875 36363
rect 14875 36329 14884 36363
rect 14832 36320 14884 36329
rect 15384 36320 15436 36372
rect 16672 36320 16724 36372
rect 17868 36320 17920 36372
rect 18236 36320 18288 36372
rect 18972 36363 19024 36372
rect 18972 36329 18981 36363
rect 18981 36329 19015 36363
rect 19015 36329 19024 36363
rect 18972 36320 19024 36329
rect 23848 36320 23900 36372
rect 29552 36363 29604 36372
rect 29552 36329 29561 36363
rect 29561 36329 29595 36363
rect 29595 36329 29604 36363
rect 29552 36320 29604 36329
rect 15844 36252 15896 36304
rect 17224 36252 17276 36304
rect 17684 36252 17736 36304
rect 18328 36295 18380 36304
rect 18328 36261 18337 36295
rect 18337 36261 18371 36295
rect 18371 36261 18380 36295
rect 18328 36252 18380 36261
rect 11060 36227 11112 36236
rect 11060 36193 11069 36227
rect 11069 36193 11103 36227
rect 11103 36193 11112 36227
rect 11060 36184 11112 36193
rect 11428 36184 11480 36236
rect 12164 36184 12216 36236
rect 12808 36227 12860 36236
rect 12808 36193 12817 36227
rect 12817 36193 12851 36227
rect 12851 36193 12860 36227
rect 12808 36184 12860 36193
rect 12992 36227 13044 36236
rect 12992 36193 13001 36227
rect 13001 36193 13035 36227
rect 13035 36193 13044 36227
rect 12992 36184 13044 36193
rect 15752 36227 15804 36236
rect 15752 36193 15761 36227
rect 15761 36193 15795 36227
rect 15795 36193 15804 36227
rect 15752 36184 15804 36193
rect 15936 36227 15988 36236
rect 15936 36193 15945 36227
rect 15945 36193 15979 36227
rect 15979 36193 15988 36227
rect 15936 36184 15988 36193
rect 16672 36227 16724 36236
rect 14924 36116 14976 36168
rect 16672 36193 16681 36227
rect 16681 36193 16715 36227
rect 16715 36193 16724 36227
rect 16672 36184 16724 36193
rect 17408 36184 17460 36236
rect 16304 36116 16356 36168
rect 17868 36227 17920 36236
rect 17868 36193 17877 36227
rect 17877 36193 17911 36227
rect 17911 36193 17920 36227
rect 17868 36184 17920 36193
rect 18880 36184 18932 36236
rect 19340 36227 19392 36236
rect 19340 36193 19349 36227
rect 19349 36193 19383 36227
rect 19383 36193 19392 36227
rect 19340 36184 19392 36193
rect 21180 36184 21232 36236
rect 23388 36227 23440 36236
rect 23388 36193 23397 36227
rect 23397 36193 23431 36227
rect 23431 36193 23440 36227
rect 23388 36184 23440 36193
rect 28264 36184 28316 36236
rect 23296 36116 23348 36168
rect 25412 36159 25464 36168
rect 25412 36125 25421 36159
rect 25421 36125 25455 36159
rect 25455 36125 25464 36159
rect 25412 36116 25464 36125
rect 28448 36159 28500 36168
rect 28448 36125 28457 36159
rect 28457 36125 28491 36159
rect 28491 36125 28500 36159
rect 28448 36116 28500 36125
rect 16764 36048 16816 36100
rect 17684 36048 17736 36100
rect 19248 36048 19300 36100
rect 11428 35980 11480 36032
rect 11980 36023 12032 36032
rect 11980 35989 11989 36023
rect 11989 35989 12023 36023
rect 12023 35989 12032 36023
rect 11980 35980 12032 35989
rect 14924 35980 14976 36032
rect 16948 35980 17000 36032
rect 18236 35980 18288 36032
rect 19156 35980 19208 36032
rect 19432 35980 19484 36032
rect 21088 36023 21140 36032
rect 21088 35989 21097 36023
rect 21097 35989 21131 36023
rect 21131 35989 21140 36023
rect 21088 35980 21140 35989
rect 21180 35980 21232 36032
rect 24216 35980 24268 36032
rect 4246 35878 4298 35930
rect 4310 35878 4362 35930
rect 4374 35878 4426 35930
rect 4438 35878 4490 35930
rect 34966 35878 35018 35930
rect 35030 35878 35082 35930
rect 35094 35878 35146 35930
rect 35158 35878 35210 35930
rect 10784 35819 10836 35828
rect 10784 35785 10793 35819
rect 10793 35785 10827 35819
rect 10827 35785 10836 35819
rect 10784 35776 10836 35785
rect 11060 35819 11112 35828
rect 11060 35785 11069 35819
rect 11069 35785 11103 35819
rect 11103 35785 11112 35819
rect 11060 35776 11112 35785
rect 11428 35776 11480 35828
rect 12164 35776 12216 35828
rect 12624 35776 12676 35828
rect 13360 35776 13412 35828
rect 14096 35776 14148 35828
rect 16028 35819 16080 35828
rect 16028 35785 16037 35819
rect 16037 35785 16071 35819
rect 16071 35785 16080 35819
rect 16028 35776 16080 35785
rect 16488 35819 16540 35828
rect 16488 35785 16497 35819
rect 16497 35785 16531 35819
rect 16531 35785 16540 35819
rect 16488 35776 16540 35785
rect 16672 35819 16724 35828
rect 16672 35785 16681 35819
rect 16681 35785 16715 35819
rect 16715 35785 16724 35819
rect 16672 35776 16724 35785
rect 16764 35776 16816 35828
rect 17408 35776 17460 35828
rect 17960 35776 18012 35828
rect 23388 35776 23440 35828
rect 28264 35776 28316 35828
rect 13268 35708 13320 35760
rect 13912 35708 13964 35760
rect 15844 35708 15896 35760
rect 10968 35640 11020 35692
rect 11060 35640 11112 35692
rect 14096 35640 14148 35692
rect 15292 35683 15344 35692
rect 15292 35649 15301 35683
rect 15301 35649 15335 35683
rect 15335 35649 15344 35683
rect 15292 35640 15344 35649
rect 13268 35572 13320 35624
rect 14372 35615 14424 35624
rect 14372 35581 14381 35615
rect 14381 35581 14415 35615
rect 14415 35581 14424 35615
rect 14372 35572 14424 35581
rect 14464 35572 14516 35624
rect 14924 35572 14976 35624
rect 12532 35547 12584 35556
rect 12532 35513 12541 35547
rect 12541 35513 12575 35547
rect 12575 35513 12584 35547
rect 12532 35504 12584 35513
rect 13912 35547 13964 35556
rect 13912 35513 13921 35547
rect 13921 35513 13955 35547
rect 13955 35513 13964 35547
rect 13912 35504 13964 35513
rect 15200 35504 15252 35556
rect 17960 35640 18012 35692
rect 19432 35640 19484 35692
rect 23296 35640 23348 35692
rect 18328 35615 18380 35624
rect 18328 35581 18337 35615
rect 18337 35581 18371 35615
rect 18371 35581 18380 35615
rect 18328 35572 18380 35581
rect 19248 35572 19300 35624
rect 21180 35615 21232 35624
rect 10140 35436 10192 35488
rect 19892 35504 19944 35556
rect 21180 35581 21189 35615
rect 21189 35581 21223 35615
rect 21223 35581 21232 35615
rect 21180 35572 21232 35581
rect 20628 35504 20680 35556
rect 22560 35547 22612 35556
rect 22560 35513 22569 35547
rect 22569 35513 22603 35547
rect 22603 35513 22612 35547
rect 22560 35504 22612 35513
rect 28448 35504 28500 35556
rect 28816 35504 28868 35556
rect 18880 35436 18932 35488
rect 23940 35479 23992 35488
rect 23940 35445 23949 35479
rect 23949 35445 23983 35479
rect 23983 35445 23992 35479
rect 23940 35436 23992 35445
rect 19606 35334 19658 35386
rect 19670 35334 19722 35386
rect 19734 35334 19786 35386
rect 19798 35334 19850 35386
rect 1676 35232 1728 35284
rect 1952 35232 2004 35284
rect 11336 35275 11388 35284
rect 11336 35241 11345 35275
rect 11345 35241 11379 35275
rect 11379 35241 11388 35275
rect 11336 35232 11388 35241
rect 11704 35275 11756 35284
rect 11704 35241 11713 35275
rect 11713 35241 11747 35275
rect 11747 35241 11756 35275
rect 11704 35232 11756 35241
rect 12532 35232 12584 35284
rect 13728 35232 13780 35284
rect 17592 35232 17644 35284
rect 17960 35232 18012 35284
rect 19340 35232 19392 35284
rect 21272 35232 21324 35284
rect 22652 35232 22704 35284
rect 23388 35232 23440 35284
rect 11888 35139 11940 35148
rect 11888 35105 11897 35139
rect 11897 35105 11931 35139
rect 11931 35105 11940 35139
rect 11888 35096 11940 35105
rect 12256 35164 12308 35216
rect 12992 35164 13044 35216
rect 13544 35164 13596 35216
rect 14464 35164 14516 35216
rect 17684 35207 17736 35216
rect 17684 35173 17693 35207
rect 17693 35173 17727 35207
rect 17727 35173 17736 35207
rect 17684 35164 17736 35173
rect 18052 35207 18104 35216
rect 18052 35173 18061 35207
rect 18061 35173 18095 35207
rect 18095 35173 18104 35207
rect 18052 35164 18104 35173
rect 19432 35207 19484 35216
rect 19432 35173 19441 35207
rect 19441 35173 19475 35207
rect 19475 35173 19484 35207
rect 19432 35164 19484 35173
rect 13820 35139 13872 35148
rect 13820 35105 13829 35139
rect 13829 35105 13863 35139
rect 13863 35105 13872 35139
rect 13820 35096 13872 35105
rect 14188 35139 14240 35148
rect 14188 35105 14197 35139
rect 14197 35105 14231 35139
rect 14231 35105 14240 35139
rect 15936 35139 15988 35148
rect 14188 35096 14240 35105
rect 11612 35028 11664 35080
rect 9404 34935 9456 34944
rect 9404 34901 9413 34935
rect 9413 34901 9447 34935
rect 9447 34901 9456 34935
rect 9404 34892 9456 34901
rect 12256 34892 12308 34944
rect 13360 34960 13412 35012
rect 14648 35028 14700 35080
rect 15936 35105 15945 35139
rect 15945 35105 15979 35139
rect 15979 35105 15988 35139
rect 15936 35096 15988 35105
rect 16028 35139 16080 35148
rect 16028 35105 16037 35139
rect 16037 35105 16071 35139
rect 16071 35105 16080 35139
rect 16028 35096 16080 35105
rect 18880 35139 18932 35148
rect 16396 35071 16448 35080
rect 16396 35037 16405 35071
rect 16405 35037 16439 35071
rect 16439 35037 16448 35071
rect 16396 35028 16448 35037
rect 17408 35028 17460 35080
rect 16028 34960 16080 35012
rect 13728 34892 13780 34944
rect 14464 34892 14516 34944
rect 14924 34892 14976 34944
rect 17132 34935 17184 34944
rect 17132 34901 17141 34935
rect 17141 34901 17175 34935
rect 17175 34901 17184 34935
rect 18880 35105 18889 35139
rect 18889 35105 18923 35139
rect 18923 35105 18932 35139
rect 18880 35096 18932 35105
rect 17960 35028 18012 35080
rect 19156 35096 19208 35148
rect 19340 35096 19392 35148
rect 21088 35096 21140 35148
rect 23480 35164 23532 35216
rect 22560 35096 22612 35148
rect 22652 35028 22704 35080
rect 19340 34960 19392 35012
rect 20076 35003 20128 35012
rect 20076 34969 20085 35003
rect 20085 34969 20119 35003
rect 20119 34969 20128 35003
rect 20076 34960 20128 34969
rect 20352 34960 20404 35012
rect 27896 35028 27948 35080
rect 23296 34960 23348 35012
rect 23940 34960 23992 35012
rect 18696 34935 18748 34944
rect 17132 34892 17184 34901
rect 18696 34901 18705 34935
rect 18705 34901 18739 34935
rect 18739 34901 18748 34935
rect 18696 34892 18748 34901
rect 19616 34892 19668 34944
rect 22836 34892 22888 34944
rect 23848 34935 23900 34944
rect 23848 34901 23857 34935
rect 23857 34901 23891 34935
rect 23891 34901 23900 34935
rect 23848 34892 23900 34901
rect 4246 34790 4298 34842
rect 4310 34790 4362 34842
rect 4374 34790 4426 34842
rect 4438 34790 4490 34842
rect 34966 34790 35018 34842
rect 35030 34790 35082 34842
rect 35094 34790 35146 34842
rect 35158 34790 35210 34842
rect 3056 34731 3108 34740
rect 3056 34697 3065 34731
rect 3065 34697 3099 34731
rect 3099 34697 3108 34731
rect 3056 34688 3108 34697
rect 8944 34731 8996 34740
rect 8944 34697 8953 34731
rect 8953 34697 8987 34731
rect 8987 34697 8996 34731
rect 8944 34688 8996 34697
rect 9220 34731 9272 34740
rect 9220 34697 9229 34731
rect 9229 34697 9263 34731
rect 9263 34697 9272 34731
rect 9220 34688 9272 34697
rect 11612 34688 11664 34740
rect 13360 34731 13412 34740
rect 13360 34697 13369 34731
rect 13369 34697 13403 34731
rect 13403 34697 13412 34731
rect 13360 34688 13412 34697
rect 14096 34688 14148 34740
rect 14832 34688 14884 34740
rect 16028 34688 16080 34740
rect 16580 34688 16632 34740
rect 18328 34688 18380 34740
rect 19892 34731 19944 34740
rect 19892 34697 19901 34731
rect 19901 34697 19935 34731
rect 19935 34697 19944 34731
rect 19892 34688 19944 34697
rect 21088 34688 21140 34740
rect 22560 34688 22612 34740
rect 24216 34688 24268 34740
rect 24676 34731 24728 34740
rect 24676 34697 24685 34731
rect 24685 34697 24719 34731
rect 24719 34697 24728 34731
rect 24676 34688 24728 34697
rect 28172 34688 28224 34740
rect 1676 34595 1728 34604
rect 1676 34561 1685 34595
rect 1685 34561 1719 34595
rect 1719 34561 1728 34595
rect 1676 34552 1728 34561
rect 14924 34620 14976 34672
rect 16396 34663 16448 34672
rect 11980 34552 12032 34604
rect 12808 34552 12860 34604
rect 15936 34552 15988 34604
rect 16396 34629 16405 34663
rect 16405 34629 16439 34663
rect 16439 34629 16448 34663
rect 16396 34620 16448 34629
rect 18696 34620 18748 34672
rect 20812 34663 20864 34672
rect 20812 34629 20821 34663
rect 20821 34629 20855 34663
rect 20855 34629 20864 34663
rect 20812 34620 20864 34629
rect 20996 34620 21048 34672
rect 1952 34527 2004 34536
rect 1952 34493 1961 34527
rect 1961 34493 1995 34527
rect 1995 34493 2004 34527
rect 1952 34484 2004 34493
rect 9220 34484 9272 34536
rect 9404 34527 9456 34536
rect 9404 34493 9413 34527
rect 9413 34493 9447 34527
rect 9447 34493 9456 34527
rect 9404 34484 9456 34493
rect 12992 34527 13044 34536
rect 10876 34416 10928 34468
rect 12992 34493 13001 34527
rect 13001 34493 13035 34527
rect 13035 34493 13044 34527
rect 12992 34484 13044 34493
rect 12624 34416 12676 34468
rect 14464 34527 14516 34536
rect 14464 34493 14473 34527
rect 14473 34493 14507 34527
rect 14507 34493 14516 34527
rect 14464 34484 14516 34493
rect 14096 34416 14148 34468
rect 14832 34484 14884 34536
rect 15200 34527 15252 34536
rect 15200 34493 15209 34527
rect 15209 34493 15243 34527
rect 15243 34493 15252 34527
rect 15200 34484 15252 34493
rect 16212 34484 16264 34536
rect 17592 34484 17644 34536
rect 18880 34484 18932 34536
rect 19616 34527 19668 34536
rect 19616 34493 19625 34527
rect 19625 34493 19659 34527
rect 19659 34493 19668 34527
rect 19616 34484 19668 34493
rect 20352 34484 20404 34536
rect 26700 34552 26752 34604
rect 30656 34595 30708 34604
rect 21088 34484 21140 34536
rect 22560 34527 22612 34536
rect 22560 34493 22569 34527
rect 22569 34493 22603 34527
rect 22603 34493 22612 34527
rect 22560 34484 22612 34493
rect 23480 34484 23532 34536
rect 24492 34484 24544 34536
rect 26240 34527 26292 34536
rect 26240 34493 26249 34527
rect 26249 34493 26283 34527
rect 26283 34493 26292 34527
rect 26240 34484 26292 34493
rect 28264 34484 28316 34536
rect 29276 34527 29328 34536
rect 29276 34493 29285 34527
rect 29285 34493 29319 34527
rect 29319 34493 29328 34527
rect 29276 34484 29328 34493
rect 30656 34561 30665 34595
rect 30665 34561 30699 34595
rect 30699 34561 30708 34595
rect 30656 34552 30708 34561
rect 29828 34484 29880 34536
rect 8484 34348 8536 34400
rect 12072 34348 12124 34400
rect 13728 34348 13780 34400
rect 16304 34416 16356 34468
rect 19432 34416 19484 34468
rect 21364 34416 21416 34468
rect 22652 34416 22704 34468
rect 24860 34416 24912 34468
rect 20352 34348 20404 34400
rect 22100 34348 22152 34400
rect 24032 34348 24084 34400
rect 19606 34246 19658 34298
rect 19670 34246 19722 34298
rect 19734 34246 19786 34298
rect 19798 34246 19850 34298
rect 10600 34187 10652 34196
rect 10600 34153 10609 34187
rect 10609 34153 10643 34187
rect 10643 34153 10652 34187
rect 10600 34144 10652 34153
rect 10968 34144 11020 34196
rect 11060 34076 11112 34128
rect 12256 34076 12308 34128
rect 12440 34187 12492 34196
rect 12440 34153 12449 34187
rect 12449 34153 12483 34187
rect 12483 34153 12492 34187
rect 12440 34144 12492 34153
rect 16948 34144 17000 34196
rect 18696 34144 18748 34196
rect 7564 34008 7616 34060
rect 11152 34051 11204 34060
rect 11152 34017 11161 34051
rect 11161 34017 11195 34051
rect 11195 34017 11204 34051
rect 11152 34008 11204 34017
rect 13360 34051 13412 34060
rect 13360 34017 13369 34051
rect 13369 34017 13403 34051
rect 13403 34017 13412 34051
rect 13360 34008 13412 34017
rect 14188 34008 14240 34060
rect 16212 34051 16264 34060
rect 16212 34017 16221 34051
rect 16221 34017 16255 34051
rect 16255 34017 16264 34051
rect 16212 34008 16264 34017
rect 11888 33983 11940 33992
rect 11888 33949 11897 33983
rect 11897 33949 11931 33983
rect 11931 33949 11940 33983
rect 11888 33940 11940 33949
rect 12532 33940 12584 33992
rect 12808 33983 12860 33992
rect 12808 33949 12817 33983
rect 12817 33949 12851 33983
rect 12851 33949 12860 33983
rect 12808 33940 12860 33949
rect 13912 33940 13964 33992
rect 16856 34076 16908 34128
rect 17960 34119 18012 34128
rect 17960 34085 17969 34119
rect 17969 34085 18003 34119
rect 18003 34085 18012 34119
rect 17960 34076 18012 34085
rect 18328 34119 18380 34128
rect 18328 34085 18337 34119
rect 18337 34085 18371 34119
rect 18371 34085 18380 34119
rect 18328 34076 18380 34085
rect 19248 34076 19300 34128
rect 20260 34076 20312 34128
rect 20720 34144 20772 34196
rect 24124 34187 24176 34196
rect 24124 34153 24133 34187
rect 24133 34153 24167 34187
rect 24167 34153 24176 34187
rect 24124 34144 24176 34153
rect 25044 34187 25096 34196
rect 25044 34153 25053 34187
rect 25053 34153 25087 34187
rect 25087 34153 25096 34187
rect 25044 34144 25096 34153
rect 29276 34187 29328 34196
rect 29276 34153 29285 34187
rect 29285 34153 29319 34187
rect 29319 34153 29328 34187
rect 29276 34144 29328 34153
rect 22100 34076 22152 34128
rect 18236 34008 18288 34060
rect 20352 34008 20404 34060
rect 20904 34051 20956 34060
rect 20904 34017 20913 34051
rect 20913 34017 20947 34051
rect 20947 34017 20956 34051
rect 20904 34008 20956 34017
rect 20996 34008 21048 34060
rect 23296 34008 23348 34060
rect 27620 34051 27672 34060
rect 27620 34017 27629 34051
rect 27629 34017 27663 34051
rect 27663 34017 27672 34051
rect 27620 34008 27672 34017
rect 32404 34051 32456 34060
rect 32404 34017 32413 34051
rect 32413 34017 32447 34051
rect 32447 34017 32456 34051
rect 32404 34008 32456 34017
rect 16580 33940 16632 33992
rect 17684 33940 17736 33992
rect 17868 33872 17920 33924
rect 1952 33804 2004 33856
rect 8116 33847 8168 33856
rect 8116 33813 8125 33847
rect 8125 33813 8159 33847
rect 8159 33813 8168 33847
rect 8116 33804 8168 33813
rect 8484 33847 8536 33856
rect 8484 33813 8493 33847
rect 8493 33813 8527 33847
rect 8527 33813 8536 33847
rect 8484 33804 8536 33813
rect 9220 33804 9272 33856
rect 9588 33804 9640 33856
rect 9956 33847 10008 33856
rect 9956 33813 9965 33847
rect 9965 33813 9999 33847
rect 9999 33813 10008 33847
rect 9956 33804 10008 33813
rect 12624 33804 12676 33856
rect 14096 33804 14148 33856
rect 14280 33847 14332 33856
rect 14280 33813 14289 33847
rect 14289 33813 14323 33847
rect 14323 33813 14332 33847
rect 14280 33804 14332 33813
rect 15568 33847 15620 33856
rect 15568 33813 15577 33847
rect 15577 33813 15611 33847
rect 15611 33813 15620 33847
rect 15568 33804 15620 33813
rect 15936 33847 15988 33856
rect 15936 33813 15945 33847
rect 15945 33813 15979 33847
rect 15979 33813 15988 33847
rect 15936 33804 15988 33813
rect 17408 33847 17460 33856
rect 17408 33813 17417 33847
rect 17417 33813 17451 33847
rect 17451 33813 17460 33847
rect 17408 33804 17460 33813
rect 18052 33804 18104 33856
rect 19156 33847 19208 33856
rect 19156 33813 19165 33847
rect 19165 33813 19199 33847
rect 19199 33813 19208 33847
rect 20628 33940 20680 33992
rect 23020 33983 23072 33992
rect 23020 33949 23029 33983
rect 23029 33949 23063 33983
rect 23063 33949 23072 33983
rect 23020 33940 23072 33949
rect 28264 33940 28316 33992
rect 32496 33940 32548 33992
rect 21548 33872 21600 33924
rect 23756 33872 23808 33924
rect 26332 33872 26384 33924
rect 19156 33804 19208 33813
rect 19340 33804 19392 33856
rect 20720 33847 20772 33856
rect 20720 33813 20729 33847
rect 20729 33813 20763 33847
rect 20763 33813 20772 33847
rect 20720 33804 20772 33813
rect 21272 33804 21324 33856
rect 22468 33847 22520 33856
rect 22468 33813 22477 33847
rect 22477 33813 22511 33847
rect 22511 33813 22520 33847
rect 22468 33804 22520 33813
rect 24676 33847 24728 33856
rect 24676 33813 24685 33847
rect 24685 33813 24719 33847
rect 24719 33813 24728 33847
rect 24676 33804 24728 33813
rect 26240 33847 26292 33856
rect 26240 33813 26249 33847
rect 26249 33813 26283 33847
rect 26283 33813 26292 33847
rect 26240 33804 26292 33813
rect 27712 33804 27764 33856
rect 33508 33847 33560 33856
rect 33508 33813 33517 33847
rect 33517 33813 33551 33847
rect 33551 33813 33560 33847
rect 33508 33804 33560 33813
rect 4246 33702 4298 33754
rect 4310 33702 4362 33754
rect 4374 33702 4426 33754
rect 4438 33702 4490 33754
rect 34966 33702 35018 33754
rect 35030 33702 35082 33754
rect 35094 33702 35146 33754
rect 35158 33702 35210 33754
rect 5448 33600 5500 33652
rect 7564 33643 7616 33652
rect 7564 33609 7573 33643
rect 7573 33609 7607 33643
rect 7607 33609 7616 33643
rect 7564 33600 7616 33609
rect 9404 33643 9456 33652
rect 9404 33609 9413 33643
rect 9413 33609 9447 33643
rect 9447 33609 9456 33643
rect 9404 33600 9456 33609
rect 10048 33643 10100 33652
rect 10048 33609 10057 33643
rect 10057 33609 10091 33643
rect 10091 33609 10100 33643
rect 10048 33600 10100 33609
rect 14188 33600 14240 33652
rect 15016 33600 15068 33652
rect 15660 33600 15712 33652
rect 16856 33643 16908 33652
rect 16856 33609 16865 33643
rect 16865 33609 16899 33643
rect 16899 33609 16908 33643
rect 16856 33600 16908 33609
rect 18236 33600 18288 33652
rect 19432 33600 19484 33652
rect 20904 33600 20956 33652
rect 22008 33600 22060 33652
rect 24768 33600 24820 33652
rect 25596 33643 25648 33652
rect 25596 33609 25605 33643
rect 25605 33609 25639 33643
rect 25639 33609 25648 33643
rect 25596 33600 25648 33609
rect 27620 33600 27672 33652
rect 28264 33600 28316 33652
rect 32404 33600 32456 33652
rect 32496 33643 32548 33652
rect 32496 33609 32505 33643
rect 32505 33609 32539 33643
rect 32539 33609 32548 33643
rect 32496 33600 32548 33609
rect 20076 33532 20128 33584
rect 11520 33507 11572 33516
rect 7932 33328 7984 33380
rect 9588 33396 9640 33448
rect 10508 33439 10560 33448
rect 10508 33405 10517 33439
rect 10517 33405 10551 33439
rect 10551 33405 10560 33439
rect 10508 33396 10560 33405
rect 10784 33396 10836 33448
rect 11060 33439 11112 33448
rect 11060 33405 11069 33439
rect 11069 33405 11103 33439
rect 11103 33405 11112 33439
rect 11060 33396 11112 33405
rect 11520 33473 11529 33507
rect 11529 33473 11563 33507
rect 11563 33473 11572 33507
rect 11520 33464 11572 33473
rect 12532 33464 12584 33516
rect 10048 33328 10100 33380
rect 11612 33396 11664 33448
rect 13820 33464 13872 33516
rect 14372 33464 14424 33516
rect 15200 33464 15252 33516
rect 19616 33507 19668 33516
rect 13268 33439 13320 33448
rect 12440 33328 12492 33380
rect 13268 33405 13277 33439
rect 13277 33405 13311 33439
rect 13311 33405 13320 33439
rect 13268 33396 13320 33405
rect 13544 33328 13596 33380
rect 8484 33260 8536 33312
rect 9956 33260 10008 33312
rect 11980 33260 12032 33312
rect 12072 33260 12124 33312
rect 14648 33396 14700 33448
rect 14832 33439 14884 33448
rect 14832 33405 14841 33439
rect 14841 33405 14875 33439
rect 14875 33405 14884 33439
rect 14832 33396 14884 33405
rect 15016 33439 15068 33448
rect 15016 33405 15025 33439
rect 15025 33405 15059 33439
rect 15059 33405 15068 33439
rect 15016 33396 15068 33405
rect 16580 33439 16632 33448
rect 15476 33328 15528 33380
rect 16580 33405 16589 33439
rect 16589 33405 16623 33439
rect 16623 33405 16632 33439
rect 16580 33396 16632 33405
rect 19616 33473 19625 33507
rect 19625 33473 19659 33507
rect 19659 33473 19668 33507
rect 19616 33464 19668 33473
rect 19984 33464 20036 33516
rect 21732 33464 21784 33516
rect 16948 33396 17000 33448
rect 15660 33328 15712 33380
rect 16856 33328 16908 33380
rect 17684 33328 17736 33380
rect 18696 33396 18748 33448
rect 19432 33396 19484 33448
rect 20904 33439 20956 33448
rect 20904 33405 20913 33439
rect 20913 33405 20947 33439
rect 20947 33405 20956 33439
rect 20904 33396 20956 33405
rect 21364 33396 21416 33448
rect 13912 33260 13964 33312
rect 14096 33260 14148 33312
rect 14372 33260 14424 33312
rect 15200 33260 15252 33312
rect 16212 33260 16264 33312
rect 16396 33303 16448 33312
rect 16396 33269 16405 33303
rect 16405 33269 16439 33303
rect 16439 33269 16448 33303
rect 16396 33260 16448 33269
rect 16580 33260 16632 33312
rect 18236 33303 18288 33312
rect 18236 33269 18245 33303
rect 18245 33269 18279 33303
rect 18279 33269 18288 33303
rect 18236 33260 18288 33269
rect 18788 33371 18840 33380
rect 18788 33337 18797 33371
rect 18797 33337 18831 33371
rect 18831 33337 18840 33371
rect 18788 33328 18840 33337
rect 19156 33328 19208 33380
rect 20260 33328 20312 33380
rect 21640 33328 21692 33380
rect 23756 33396 23808 33448
rect 24124 33439 24176 33448
rect 24124 33405 24133 33439
rect 24133 33405 24167 33439
rect 24167 33405 24176 33439
rect 24124 33396 24176 33405
rect 24492 33396 24544 33448
rect 24676 33439 24728 33448
rect 24676 33405 24685 33439
rect 24685 33405 24719 33439
rect 24719 33405 24728 33439
rect 24676 33396 24728 33405
rect 24860 33439 24912 33448
rect 24860 33405 24869 33439
rect 24869 33405 24903 33439
rect 24903 33405 24912 33439
rect 24860 33396 24912 33405
rect 25504 33396 25556 33448
rect 23020 33328 23072 33380
rect 25320 33328 25372 33380
rect 20352 33260 20404 33312
rect 21272 33260 21324 33312
rect 21456 33303 21508 33312
rect 21456 33269 21465 33303
rect 21465 33269 21499 33303
rect 21499 33269 21508 33303
rect 21456 33260 21508 33269
rect 22008 33260 22060 33312
rect 23112 33303 23164 33312
rect 23112 33269 23121 33303
rect 23121 33269 23155 33303
rect 23155 33269 23164 33303
rect 23112 33260 23164 33269
rect 23296 33303 23348 33312
rect 23296 33269 23305 33303
rect 23305 33269 23339 33303
rect 23339 33269 23348 33303
rect 23296 33260 23348 33269
rect 23756 33260 23808 33312
rect 26240 33303 26292 33312
rect 26240 33269 26249 33303
rect 26249 33269 26283 33303
rect 26283 33269 26292 33303
rect 26240 33260 26292 33269
rect 29276 33260 29328 33312
rect 32496 33260 32548 33312
rect 19606 33158 19658 33210
rect 19670 33158 19722 33210
rect 19734 33158 19786 33210
rect 19798 33158 19850 33210
rect 8116 33099 8168 33108
rect 8116 33065 8125 33099
rect 8125 33065 8159 33099
rect 8159 33065 8168 33099
rect 8116 33056 8168 33065
rect 8760 33099 8812 33108
rect 8760 33065 8769 33099
rect 8769 33065 8803 33099
rect 8803 33065 8812 33099
rect 8760 33056 8812 33065
rect 9588 33056 9640 33108
rect 11060 33099 11112 33108
rect 11060 33065 11069 33099
rect 11069 33065 11103 33099
rect 11103 33065 11112 33099
rect 15476 33099 15528 33108
rect 11060 33056 11112 33065
rect 9036 32988 9088 33040
rect 13084 32988 13136 33040
rect 13544 32988 13596 33040
rect 13912 32988 13964 33040
rect 8576 32963 8628 32972
rect 8576 32929 8585 32963
rect 8585 32929 8619 32963
rect 8619 32929 8628 32963
rect 8576 32920 8628 32929
rect 10968 32920 11020 32972
rect 12164 32963 12216 32972
rect 12164 32929 12173 32963
rect 12173 32929 12207 32963
rect 12207 32929 12216 32963
rect 12164 32920 12216 32929
rect 12992 32920 13044 32972
rect 15476 33065 15485 33099
rect 15485 33065 15519 33099
rect 15519 33065 15528 33099
rect 15476 33056 15528 33065
rect 17684 33056 17736 33108
rect 18604 33099 18656 33108
rect 18604 33065 18613 33099
rect 18613 33065 18647 33099
rect 18647 33065 18656 33099
rect 18604 33056 18656 33065
rect 20260 33056 20312 33108
rect 16580 33031 16632 33040
rect 16580 32997 16589 33031
rect 16589 32997 16623 33031
rect 16623 32997 16632 33031
rect 16580 32988 16632 32997
rect 16764 33031 16816 33040
rect 16764 32997 16773 33031
rect 16773 32997 16807 33031
rect 16807 32997 16816 33031
rect 16764 32988 16816 32997
rect 9220 32852 9272 32904
rect 9680 32895 9732 32904
rect 9680 32861 9689 32895
rect 9689 32861 9723 32895
rect 9723 32861 9732 32895
rect 9680 32852 9732 32861
rect 9864 32852 9916 32904
rect 11520 32852 11572 32904
rect 12624 32827 12676 32836
rect 12624 32793 12633 32827
rect 12633 32793 12667 32827
rect 12667 32793 12676 32827
rect 12624 32784 12676 32793
rect 12716 32784 12768 32836
rect 15660 32920 15712 32972
rect 16396 32963 16448 32972
rect 16396 32929 16405 32963
rect 16405 32929 16439 32963
rect 16439 32929 16448 32963
rect 16396 32920 16448 32929
rect 16948 32920 17000 32972
rect 17776 32988 17828 33040
rect 21732 33056 21784 33108
rect 26240 33056 26292 33108
rect 22008 32988 22060 33040
rect 17960 32963 18012 32972
rect 17960 32929 17969 32963
rect 17969 32929 18003 32963
rect 18003 32929 18012 32963
rect 17960 32920 18012 32929
rect 19432 32920 19484 32972
rect 15384 32852 15436 32904
rect 16028 32784 16080 32836
rect 17592 32852 17644 32904
rect 17776 32852 17828 32904
rect 18328 32895 18380 32904
rect 18328 32861 18337 32895
rect 18337 32861 18371 32895
rect 18371 32861 18380 32895
rect 18328 32852 18380 32861
rect 20352 32852 20404 32904
rect 20812 32852 20864 32904
rect 18788 32784 18840 32836
rect 19616 32784 19668 32836
rect 20536 32784 20588 32836
rect 11336 32716 11388 32768
rect 11704 32759 11756 32768
rect 11704 32725 11713 32759
rect 11713 32725 11747 32759
rect 11747 32725 11756 32759
rect 11704 32716 11756 32725
rect 12072 32759 12124 32768
rect 12072 32725 12081 32759
rect 12081 32725 12115 32759
rect 12115 32725 12124 32759
rect 12072 32716 12124 32725
rect 12256 32716 12308 32768
rect 12808 32716 12860 32768
rect 13360 32716 13412 32768
rect 13820 32716 13872 32768
rect 14464 32716 14516 32768
rect 15016 32759 15068 32768
rect 15016 32725 15025 32759
rect 15025 32725 15059 32759
rect 15059 32725 15068 32759
rect 15016 32716 15068 32725
rect 15752 32716 15804 32768
rect 16304 32716 16356 32768
rect 16672 32716 16724 32768
rect 17868 32716 17920 32768
rect 18328 32716 18380 32768
rect 18880 32716 18932 32768
rect 19064 32716 19116 32768
rect 19432 32716 19484 32768
rect 20720 32759 20772 32768
rect 20720 32725 20729 32759
rect 20729 32725 20763 32759
rect 20763 32725 20772 32759
rect 22928 32920 22980 32972
rect 24216 32963 24268 32972
rect 24216 32929 24225 32963
rect 24225 32929 24259 32963
rect 24259 32929 24268 32963
rect 24216 32920 24268 32929
rect 27344 32920 27396 32972
rect 28264 32920 28316 32972
rect 28448 32920 28500 32972
rect 28908 32963 28960 32972
rect 28908 32929 28917 32963
rect 28917 32929 28951 32963
rect 28951 32929 28960 32963
rect 28908 32920 28960 32929
rect 21640 32895 21692 32904
rect 21640 32861 21649 32895
rect 21649 32861 21683 32895
rect 21683 32861 21692 32895
rect 21640 32852 21692 32861
rect 22100 32852 22152 32904
rect 22468 32895 22520 32904
rect 22468 32861 22477 32895
rect 22477 32861 22511 32895
rect 22511 32861 22520 32895
rect 22468 32852 22520 32861
rect 23664 32895 23716 32904
rect 23664 32861 23673 32895
rect 23673 32861 23707 32895
rect 23707 32861 23716 32895
rect 23664 32852 23716 32861
rect 23756 32852 23808 32904
rect 25320 32895 25372 32904
rect 25320 32861 25329 32895
rect 25329 32861 25363 32895
rect 25363 32861 25372 32895
rect 25320 32852 25372 32861
rect 22652 32784 22704 32836
rect 24952 32784 25004 32836
rect 28172 32784 28224 32836
rect 20720 32716 20772 32725
rect 22560 32716 22612 32768
rect 23296 32759 23348 32768
rect 23296 32725 23305 32759
rect 23305 32725 23339 32759
rect 23339 32725 23348 32759
rect 23296 32716 23348 32725
rect 30012 32759 30064 32768
rect 30012 32725 30021 32759
rect 30021 32725 30055 32759
rect 30055 32725 30064 32759
rect 30012 32716 30064 32725
rect 4246 32614 4298 32666
rect 4310 32614 4362 32666
rect 4374 32614 4426 32666
rect 4438 32614 4490 32666
rect 34966 32614 35018 32666
rect 35030 32614 35082 32666
rect 35094 32614 35146 32666
rect 35158 32614 35210 32666
rect 1676 32512 1728 32564
rect 5448 32555 5500 32564
rect 5448 32521 5457 32555
rect 5457 32521 5491 32555
rect 5491 32521 5500 32555
rect 5448 32512 5500 32521
rect 7748 32555 7800 32564
rect 7748 32521 7757 32555
rect 7757 32521 7791 32555
rect 7791 32521 7800 32555
rect 7748 32512 7800 32521
rect 5448 32308 5500 32360
rect 9220 32512 9272 32564
rect 9864 32512 9916 32564
rect 11888 32555 11940 32564
rect 11888 32521 11897 32555
rect 11897 32521 11931 32555
rect 11931 32521 11940 32555
rect 11888 32512 11940 32521
rect 12164 32555 12216 32564
rect 12164 32521 12173 32555
rect 12173 32521 12207 32555
rect 12207 32521 12216 32555
rect 12164 32512 12216 32521
rect 15384 32555 15436 32564
rect 15384 32521 15393 32555
rect 15393 32521 15427 32555
rect 15427 32521 15436 32555
rect 15384 32512 15436 32521
rect 16028 32512 16080 32564
rect 16764 32512 16816 32564
rect 13084 32487 13136 32496
rect 9312 32376 9364 32428
rect 10968 32419 11020 32428
rect 10968 32385 10987 32419
rect 10987 32385 11020 32419
rect 11520 32419 11572 32428
rect 10968 32376 11020 32385
rect 11520 32385 11529 32419
rect 11529 32385 11563 32419
rect 11563 32385 11572 32419
rect 11520 32376 11572 32385
rect 9036 32308 9088 32360
rect 9680 32351 9732 32360
rect 9680 32317 9689 32351
rect 9689 32317 9723 32351
rect 9723 32317 9732 32351
rect 11060 32351 11112 32360
rect 9680 32308 9732 32317
rect 11060 32317 11069 32351
rect 11069 32317 11103 32351
rect 11103 32317 11112 32351
rect 11060 32308 11112 32317
rect 11888 32308 11940 32360
rect 13084 32453 13093 32487
rect 13093 32453 13127 32487
rect 13127 32453 13136 32487
rect 13084 32444 13136 32453
rect 14372 32444 14424 32496
rect 15292 32444 15344 32496
rect 16212 32487 16264 32496
rect 16212 32453 16221 32487
rect 16221 32453 16255 32487
rect 16255 32453 16264 32487
rect 16212 32444 16264 32453
rect 13544 32376 13596 32428
rect 12624 32308 12676 32360
rect 13820 32308 13872 32360
rect 15844 32376 15896 32428
rect 16304 32419 16356 32428
rect 16304 32385 16313 32419
rect 16313 32385 16347 32419
rect 16347 32385 16356 32419
rect 16304 32376 16356 32385
rect 10140 32283 10192 32292
rect 10140 32249 10149 32283
rect 10149 32249 10183 32283
rect 10183 32249 10192 32283
rect 10140 32240 10192 32249
rect 10876 32283 10928 32292
rect 10876 32249 10885 32283
rect 10885 32249 10919 32283
rect 10919 32249 10928 32283
rect 10876 32240 10928 32249
rect 12440 32240 12492 32292
rect 14372 32351 14424 32360
rect 14372 32317 14381 32351
rect 14381 32317 14415 32351
rect 14415 32317 14424 32351
rect 14648 32351 14700 32360
rect 14372 32308 14424 32317
rect 14648 32317 14657 32351
rect 14657 32317 14691 32351
rect 14691 32317 14700 32351
rect 14648 32308 14700 32317
rect 14832 32308 14884 32360
rect 7564 32172 7616 32224
rect 8116 32215 8168 32224
rect 8116 32181 8125 32215
rect 8125 32181 8159 32215
rect 8159 32181 8168 32215
rect 8116 32172 8168 32181
rect 13084 32172 13136 32224
rect 13452 32172 13504 32224
rect 13820 32172 13872 32224
rect 16580 32308 16632 32360
rect 15844 32240 15896 32292
rect 17316 32512 17368 32564
rect 17316 32376 17368 32428
rect 17592 32308 17644 32360
rect 18420 32308 18472 32360
rect 18880 32444 18932 32496
rect 19892 32512 19944 32564
rect 20076 32512 20128 32564
rect 21088 32512 21140 32564
rect 22100 32512 22152 32564
rect 19892 32376 19944 32428
rect 21732 32444 21784 32496
rect 23296 32444 23348 32496
rect 17960 32240 18012 32292
rect 19248 32308 19300 32360
rect 20812 32308 20864 32360
rect 21088 32376 21140 32428
rect 21456 32376 21508 32428
rect 22008 32376 22060 32428
rect 24860 32512 24912 32564
rect 25596 32555 25648 32564
rect 25596 32521 25605 32555
rect 25605 32521 25639 32555
rect 25639 32521 25648 32555
rect 25596 32512 25648 32521
rect 26332 32512 26384 32564
rect 28448 32555 28500 32564
rect 25780 32444 25832 32496
rect 24124 32376 24176 32428
rect 19064 32240 19116 32292
rect 19616 32240 19668 32292
rect 20996 32240 21048 32292
rect 21180 32240 21232 32292
rect 16580 32215 16632 32224
rect 16580 32181 16589 32215
rect 16589 32181 16623 32215
rect 16623 32181 16632 32215
rect 16580 32172 16632 32181
rect 17408 32172 17460 32224
rect 17592 32172 17644 32224
rect 18420 32172 18472 32224
rect 20904 32172 20956 32224
rect 21548 32172 21600 32224
rect 22560 32308 22612 32360
rect 23664 32351 23716 32360
rect 23664 32317 23673 32351
rect 23673 32317 23707 32351
rect 23707 32317 23716 32351
rect 23664 32308 23716 32317
rect 23940 32351 23992 32360
rect 23940 32317 23949 32351
rect 23949 32317 23983 32351
rect 23983 32317 23992 32351
rect 23940 32308 23992 32317
rect 26424 32308 26476 32360
rect 27160 32308 27212 32360
rect 28448 32521 28457 32555
rect 28457 32521 28491 32555
rect 28491 32521 28500 32555
rect 28448 32512 28500 32521
rect 28908 32555 28960 32564
rect 28908 32521 28917 32555
rect 28917 32521 28951 32555
rect 28951 32521 28960 32555
rect 28908 32512 28960 32521
rect 29184 32444 29236 32496
rect 22468 32240 22520 32292
rect 22928 32172 22980 32224
rect 26240 32240 26292 32292
rect 25688 32172 25740 32224
rect 26332 32215 26384 32224
rect 26332 32181 26341 32215
rect 26341 32181 26375 32215
rect 26375 32181 26384 32215
rect 26332 32172 26384 32181
rect 26424 32172 26476 32224
rect 19606 32070 19658 32122
rect 19670 32070 19722 32122
rect 19734 32070 19786 32122
rect 19798 32070 19850 32122
rect 6920 31968 6972 32020
rect 7840 31968 7892 32020
rect 9036 31968 9088 32020
rect 10140 31968 10192 32020
rect 10600 31968 10652 32020
rect 12992 31968 13044 32020
rect 13268 32011 13320 32020
rect 13268 31977 13277 32011
rect 13277 31977 13311 32011
rect 13311 31977 13320 32011
rect 13268 31968 13320 31977
rect 7288 31900 7340 31952
rect 8576 31875 8628 31884
rect 8576 31841 8585 31875
rect 8585 31841 8619 31875
rect 8619 31841 8628 31875
rect 8576 31832 8628 31841
rect 10232 31900 10284 31952
rect 12716 31900 12768 31952
rect 14464 31968 14516 32020
rect 14648 32011 14700 32020
rect 14648 31977 14657 32011
rect 14657 31977 14691 32011
rect 14691 31977 14700 32011
rect 14648 31968 14700 31977
rect 15752 31968 15804 32020
rect 16028 31968 16080 32020
rect 16120 31968 16172 32020
rect 16672 31968 16724 32020
rect 18972 32011 19024 32020
rect 13820 31943 13872 31952
rect 13820 31909 13829 31943
rect 13829 31909 13863 31943
rect 13863 31909 13872 31943
rect 13820 31900 13872 31909
rect 11152 31832 11204 31884
rect 13912 31875 13964 31884
rect 13912 31841 13921 31875
rect 13921 31841 13955 31875
rect 13955 31841 13964 31875
rect 13912 31832 13964 31841
rect 7656 31764 7708 31816
rect 8024 31764 8076 31816
rect 8944 31764 8996 31816
rect 9772 31764 9824 31816
rect 9864 31764 9916 31816
rect 10784 31807 10836 31816
rect 10784 31773 10793 31807
rect 10793 31773 10827 31807
rect 10827 31773 10836 31807
rect 10784 31764 10836 31773
rect 10968 31764 11020 31816
rect 13544 31764 13596 31816
rect 8760 31739 8812 31748
rect 8760 31705 8769 31739
rect 8769 31705 8803 31739
rect 8803 31705 8812 31739
rect 8760 31696 8812 31705
rect 9496 31739 9548 31748
rect 9496 31705 9505 31739
rect 9505 31705 9539 31739
rect 9539 31705 9548 31739
rect 9496 31696 9548 31705
rect 12256 31696 12308 31748
rect 12440 31696 12492 31748
rect 12532 31696 12584 31748
rect 12808 31696 12860 31748
rect 14372 31875 14424 31884
rect 14372 31841 14381 31875
rect 14381 31841 14415 31875
rect 14415 31841 14424 31875
rect 14372 31832 14424 31841
rect 14648 31832 14700 31884
rect 14924 31832 14976 31884
rect 15844 31900 15896 31952
rect 15752 31875 15804 31884
rect 15752 31841 15761 31875
rect 15761 31841 15795 31875
rect 15795 31841 15804 31875
rect 15752 31832 15804 31841
rect 16120 31875 16172 31884
rect 16120 31841 16129 31875
rect 16129 31841 16163 31875
rect 16163 31841 16172 31875
rect 16120 31832 16172 31841
rect 16396 31900 16448 31952
rect 16764 31832 16816 31884
rect 18328 31875 18380 31884
rect 18328 31841 18337 31875
rect 18337 31841 18371 31875
rect 18371 31841 18380 31875
rect 18328 31832 18380 31841
rect 18972 31977 18981 32011
rect 18981 31977 19015 32011
rect 19015 31977 19024 32011
rect 18972 31968 19024 31977
rect 20260 31968 20312 32020
rect 20812 31968 20864 32020
rect 21272 31968 21324 32020
rect 21548 31968 21600 32020
rect 23296 32011 23348 32020
rect 23296 31977 23305 32011
rect 23305 31977 23339 32011
rect 23339 31977 23348 32011
rect 23296 31968 23348 31977
rect 19616 31900 19668 31952
rect 19892 31900 19944 31952
rect 20536 31900 20588 31952
rect 22836 31943 22888 31952
rect 22836 31909 22845 31943
rect 22845 31909 22879 31943
rect 22879 31909 22888 31943
rect 22836 31900 22888 31909
rect 24216 31968 24268 32020
rect 24860 32011 24912 32020
rect 24860 31977 24869 32011
rect 24869 31977 24903 32011
rect 24903 31977 24912 32011
rect 24860 31968 24912 31977
rect 25044 31968 25096 32020
rect 27712 31968 27764 32020
rect 24124 31900 24176 31952
rect 25596 31900 25648 31952
rect 16580 31764 16632 31816
rect 17960 31764 18012 31816
rect 20260 31832 20312 31884
rect 20444 31832 20496 31884
rect 21364 31875 21416 31884
rect 21364 31841 21373 31875
rect 21373 31841 21407 31875
rect 21407 31841 21416 31875
rect 21364 31832 21416 31841
rect 21456 31832 21508 31884
rect 22468 31875 22520 31884
rect 18880 31764 18932 31816
rect 19340 31764 19392 31816
rect 20720 31764 20772 31816
rect 21640 31764 21692 31816
rect 22468 31841 22477 31875
rect 22477 31841 22511 31875
rect 22511 31841 22520 31875
rect 22468 31832 22520 31841
rect 23112 31832 23164 31884
rect 24768 31832 24820 31884
rect 24952 31875 25004 31884
rect 24952 31841 24961 31875
rect 24961 31841 24995 31875
rect 24995 31841 25004 31875
rect 24952 31832 25004 31841
rect 26792 31832 26844 31884
rect 28080 31900 28132 31952
rect 28724 31900 28776 31952
rect 29184 31875 29236 31884
rect 29184 31841 29193 31875
rect 29193 31841 29227 31875
rect 29227 31841 29236 31875
rect 29184 31832 29236 31841
rect 29460 31875 29512 31884
rect 29460 31841 29469 31875
rect 29469 31841 29503 31875
rect 29503 31841 29512 31875
rect 29460 31832 29512 31841
rect 19892 31696 19944 31748
rect 23296 31764 23348 31816
rect 24308 31764 24360 31816
rect 23940 31696 23992 31748
rect 7564 31628 7616 31680
rect 11152 31628 11204 31680
rect 11520 31628 11572 31680
rect 11796 31628 11848 31680
rect 13452 31628 13504 31680
rect 16672 31628 16724 31680
rect 19340 31628 19392 31680
rect 20812 31628 20864 31680
rect 21272 31628 21324 31680
rect 25136 31764 25188 31816
rect 27344 31764 27396 31816
rect 27620 31764 27672 31816
rect 30564 31807 30616 31816
rect 30564 31773 30573 31807
rect 30573 31773 30607 31807
rect 30607 31773 30616 31807
rect 30564 31764 30616 31773
rect 25780 31739 25832 31748
rect 25780 31705 25789 31739
rect 25789 31705 25823 31739
rect 25823 31705 25832 31739
rect 25780 31696 25832 31705
rect 27712 31628 27764 31680
rect 4246 31526 4298 31578
rect 4310 31526 4362 31578
rect 4374 31526 4426 31578
rect 4438 31526 4490 31578
rect 34966 31526 35018 31578
rect 35030 31526 35082 31578
rect 35094 31526 35146 31578
rect 35158 31526 35210 31578
rect 8484 31424 8536 31476
rect 8760 31424 8812 31476
rect 11888 31467 11940 31476
rect 11888 31433 11897 31467
rect 11897 31433 11931 31467
rect 11931 31433 11940 31467
rect 11888 31424 11940 31433
rect 12440 31424 12492 31476
rect 13268 31424 13320 31476
rect 13820 31467 13872 31476
rect 13820 31433 13829 31467
rect 13829 31433 13863 31467
rect 13863 31433 13872 31467
rect 13820 31424 13872 31433
rect 15844 31467 15896 31476
rect 15844 31433 15853 31467
rect 15853 31433 15887 31467
rect 15887 31433 15896 31467
rect 15844 31424 15896 31433
rect 19340 31424 19392 31476
rect 10876 31356 10928 31408
rect 7564 31331 7616 31340
rect 7564 31297 7573 31331
rect 7573 31297 7607 31331
rect 7607 31297 7616 31331
rect 7564 31288 7616 31297
rect 7840 31331 7892 31340
rect 7840 31297 7849 31331
rect 7849 31297 7883 31331
rect 7883 31297 7892 31331
rect 7840 31288 7892 31297
rect 10968 31288 11020 31340
rect 11060 31288 11112 31340
rect 11520 31288 11572 31340
rect 13544 31356 13596 31408
rect 15292 31356 15344 31408
rect 16304 31356 16356 31408
rect 14464 31288 14516 31340
rect 15476 31331 15528 31340
rect 15476 31297 15485 31331
rect 15485 31297 15519 31331
rect 15519 31297 15528 31331
rect 15476 31288 15528 31297
rect 17684 31356 17736 31408
rect 16580 31288 16632 31340
rect 19064 31288 19116 31340
rect 19340 31288 19392 31340
rect 10508 31152 10560 31204
rect 11980 31220 12032 31272
rect 12900 31263 12952 31272
rect 12900 31229 12909 31263
rect 12909 31229 12943 31263
rect 12943 31229 12952 31263
rect 12900 31220 12952 31229
rect 13268 31263 13320 31272
rect 13268 31229 13277 31263
rect 13277 31229 13311 31263
rect 13311 31229 13320 31263
rect 13268 31220 13320 31229
rect 13452 31220 13504 31272
rect 14372 31220 14424 31272
rect 15016 31220 15068 31272
rect 7012 31127 7064 31136
rect 7012 31093 7021 31127
rect 7021 31093 7055 31127
rect 7055 31093 7064 31127
rect 7012 31084 7064 31093
rect 7472 31127 7524 31136
rect 7472 31093 7481 31127
rect 7481 31093 7515 31127
rect 7515 31093 7524 31127
rect 7472 31084 7524 31093
rect 9036 31084 9088 31136
rect 9588 31127 9640 31136
rect 9588 31093 9597 31127
rect 9597 31093 9631 31127
rect 9631 31093 9640 31127
rect 9588 31084 9640 31093
rect 9956 31127 10008 31136
rect 9956 31093 9965 31127
rect 9965 31093 9999 31127
rect 9999 31093 10008 31127
rect 9956 31084 10008 31093
rect 10232 31084 10284 31136
rect 10968 31127 11020 31136
rect 10968 31093 10977 31127
rect 10977 31093 11011 31127
rect 11011 31093 11020 31127
rect 10968 31084 11020 31093
rect 11888 31152 11940 31204
rect 15292 31152 15344 31204
rect 15844 31152 15896 31204
rect 17316 31220 17368 31272
rect 17592 31220 17644 31272
rect 19892 31288 19944 31340
rect 16764 31195 16816 31204
rect 16764 31161 16773 31195
rect 16773 31161 16807 31195
rect 16807 31161 16816 31195
rect 16764 31152 16816 31161
rect 17224 31152 17276 31204
rect 18052 31195 18104 31204
rect 18052 31161 18061 31195
rect 18061 31161 18095 31195
rect 18095 31161 18104 31195
rect 18052 31152 18104 31161
rect 18604 31152 18656 31204
rect 21456 31424 21508 31476
rect 23112 31467 23164 31476
rect 23112 31433 23121 31467
rect 23121 31433 23155 31467
rect 23155 31433 23164 31467
rect 23112 31424 23164 31433
rect 24492 31424 24544 31476
rect 24952 31424 25004 31476
rect 26056 31467 26108 31476
rect 26056 31433 26065 31467
rect 26065 31433 26099 31467
rect 26099 31433 26108 31467
rect 26056 31424 26108 31433
rect 26792 31467 26844 31476
rect 26792 31433 26801 31467
rect 26801 31433 26835 31467
rect 26835 31433 26844 31467
rect 26792 31424 26844 31433
rect 26976 31424 27028 31476
rect 27436 31467 27488 31476
rect 27436 31433 27445 31467
rect 27445 31433 27479 31467
rect 27479 31433 27488 31467
rect 27436 31424 27488 31433
rect 28080 31467 28132 31476
rect 28080 31433 28089 31467
rect 28089 31433 28123 31467
rect 28123 31433 28132 31467
rect 28080 31424 28132 31433
rect 29460 31467 29512 31476
rect 29460 31433 29469 31467
rect 29469 31433 29503 31467
rect 29503 31433 29512 31467
rect 29460 31424 29512 31433
rect 24032 31356 24084 31408
rect 21640 31288 21692 31340
rect 22008 31288 22060 31340
rect 23940 31288 23992 31340
rect 21456 31220 21508 31272
rect 23480 31220 23532 31272
rect 25780 31288 25832 31340
rect 28448 31331 28500 31340
rect 12256 31127 12308 31136
rect 12256 31093 12265 31127
rect 12265 31093 12299 31127
rect 12299 31093 12308 31127
rect 12256 31084 12308 31093
rect 13268 31084 13320 31136
rect 16580 31127 16632 31136
rect 16580 31093 16589 31127
rect 16589 31093 16623 31127
rect 16623 31093 16632 31127
rect 16580 31084 16632 31093
rect 17960 31084 18012 31136
rect 19432 31084 19484 31136
rect 20352 31195 20404 31204
rect 20352 31161 20361 31195
rect 20361 31161 20395 31195
rect 20395 31161 20404 31195
rect 20352 31152 20404 31161
rect 22652 31152 22704 31204
rect 22836 31152 22888 31204
rect 23756 31152 23808 31204
rect 25320 31220 25372 31272
rect 28448 31297 28457 31331
rect 28457 31297 28491 31331
rect 28491 31297 28500 31331
rect 28448 31288 28500 31297
rect 26240 31263 26292 31272
rect 26240 31229 26249 31263
rect 26249 31229 26283 31263
rect 26283 31229 26292 31263
rect 26240 31220 26292 31229
rect 27252 31263 27304 31272
rect 27252 31229 27261 31263
rect 27261 31229 27295 31263
rect 27295 31229 27304 31263
rect 27252 31220 27304 31229
rect 24492 31152 24544 31204
rect 24768 31152 24820 31204
rect 26332 31152 26384 31204
rect 21456 31127 21508 31136
rect 21456 31093 21465 31127
rect 21465 31093 21499 31127
rect 21499 31093 21508 31127
rect 21456 31084 21508 31093
rect 21640 31084 21692 31136
rect 22468 31084 22520 31136
rect 23112 31084 23164 31136
rect 23388 31084 23440 31136
rect 24952 31084 25004 31136
rect 25412 31127 25464 31136
rect 25412 31093 25421 31127
rect 25421 31093 25455 31127
rect 25455 31093 25464 31127
rect 25412 31084 25464 31093
rect 26792 31084 26844 31136
rect 28724 31084 28776 31136
rect 29184 31084 29236 31136
rect 29460 31084 29512 31136
rect 19606 30982 19658 31034
rect 19670 30982 19722 31034
rect 19734 30982 19786 31034
rect 19798 30982 19850 31034
rect 7012 30880 7064 30932
rect 7748 30923 7800 30932
rect 7748 30889 7757 30923
rect 7757 30889 7791 30923
rect 7791 30889 7800 30923
rect 7748 30880 7800 30889
rect 8576 30880 8628 30932
rect 9588 30880 9640 30932
rect 10784 30880 10836 30932
rect 11244 30923 11296 30932
rect 11244 30889 11253 30923
rect 11253 30889 11287 30923
rect 11287 30889 11296 30923
rect 11244 30880 11296 30889
rect 11520 30880 11572 30932
rect 11704 30880 11756 30932
rect 12440 30880 12492 30932
rect 13728 30880 13780 30932
rect 7564 30787 7616 30796
rect 7564 30753 7573 30787
rect 7573 30753 7607 30787
rect 7607 30753 7616 30787
rect 7564 30744 7616 30753
rect 9128 30744 9180 30796
rect 8116 30676 8168 30728
rect 8208 30608 8260 30660
rect 9128 30608 9180 30660
rect 10876 30744 10928 30796
rect 12532 30812 12584 30864
rect 15200 30880 15252 30932
rect 16212 30880 16264 30932
rect 11796 30787 11848 30796
rect 11796 30753 11805 30787
rect 11805 30753 11839 30787
rect 11839 30753 11848 30787
rect 11796 30744 11848 30753
rect 11980 30744 12032 30796
rect 12624 30744 12676 30796
rect 14188 30812 14240 30864
rect 14924 30812 14976 30864
rect 16304 30855 16356 30864
rect 16304 30821 16313 30855
rect 16313 30821 16347 30855
rect 16347 30821 16356 30855
rect 16304 30812 16356 30821
rect 16856 30812 16908 30864
rect 18328 30880 18380 30932
rect 18696 30880 18748 30932
rect 19248 30923 19300 30932
rect 19248 30889 19257 30923
rect 19257 30889 19291 30923
rect 19291 30889 19300 30923
rect 19248 30880 19300 30889
rect 20720 30923 20772 30932
rect 20720 30889 20729 30923
rect 20729 30889 20763 30923
rect 20763 30889 20772 30923
rect 20720 30880 20772 30889
rect 21088 30880 21140 30932
rect 21364 30880 21416 30932
rect 22928 30923 22980 30932
rect 22928 30889 22937 30923
rect 22937 30889 22971 30923
rect 22971 30889 22980 30923
rect 22928 30880 22980 30889
rect 23664 30880 23716 30932
rect 23940 30880 23992 30932
rect 20352 30812 20404 30864
rect 21272 30855 21324 30864
rect 21272 30821 21281 30855
rect 21281 30821 21315 30855
rect 21315 30821 21324 30855
rect 21272 30812 21324 30821
rect 21732 30812 21784 30864
rect 23112 30812 23164 30864
rect 24860 30880 24912 30932
rect 11704 30676 11756 30728
rect 12900 30676 12952 30728
rect 13728 30676 13780 30728
rect 10232 30608 10284 30660
rect 8300 30540 8352 30592
rect 8484 30583 8536 30592
rect 8484 30549 8493 30583
rect 8493 30549 8527 30583
rect 8527 30549 8536 30583
rect 8484 30540 8536 30549
rect 9312 30540 9364 30592
rect 10968 30540 11020 30592
rect 12808 30608 12860 30660
rect 13084 30608 13136 30660
rect 14464 30744 14516 30796
rect 14832 30744 14884 30796
rect 16212 30744 16264 30796
rect 16764 30744 16816 30796
rect 17132 30744 17184 30796
rect 17960 30744 18012 30796
rect 15108 30676 15160 30728
rect 18236 30676 18288 30728
rect 18604 30744 18656 30796
rect 19984 30676 20036 30728
rect 16948 30608 17000 30660
rect 21364 30744 21416 30796
rect 22284 30744 22336 30796
rect 22836 30744 22888 30796
rect 24492 30744 24544 30796
rect 24860 30744 24912 30796
rect 20720 30676 20772 30728
rect 22008 30676 22060 30728
rect 24676 30676 24728 30728
rect 27344 30676 27396 30728
rect 27528 30676 27580 30728
rect 20352 30651 20404 30660
rect 20352 30617 20361 30651
rect 20361 30617 20395 30651
rect 20395 30617 20404 30651
rect 20352 30608 20404 30617
rect 22560 30651 22612 30660
rect 22560 30617 22569 30651
rect 22569 30617 22603 30651
rect 22603 30617 22612 30651
rect 22560 30608 22612 30617
rect 24308 30651 24360 30660
rect 24308 30617 24317 30651
rect 24317 30617 24351 30651
rect 24351 30617 24360 30651
rect 24308 30608 24360 30617
rect 24492 30608 24544 30660
rect 13452 30540 13504 30592
rect 15752 30583 15804 30592
rect 15752 30549 15761 30583
rect 15761 30549 15795 30583
rect 15795 30549 15804 30583
rect 15752 30540 15804 30549
rect 16212 30583 16264 30592
rect 16212 30549 16221 30583
rect 16221 30549 16255 30583
rect 16255 30549 16264 30583
rect 16212 30540 16264 30549
rect 16580 30540 16632 30592
rect 18788 30540 18840 30592
rect 19340 30540 19392 30592
rect 22468 30540 22520 30592
rect 23756 30540 23808 30592
rect 24216 30540 24268 30592
rect 24952 30540 25004 30592
rect 25412 30540 25464 30592
rect 26424 30540 26476 30592
rect 28172 30540 28224 30592
rect 28540 30583 28592 30592
rect 28540 30549 28549 30583
rect 28549 30549 28583 30583
rect 28583 30549 28592 30583
rect 28540 30540 28592 30549
rect 4246 30438 4298 30490
rect 4310 30438 4362 30490
rect 4374 30438 4426 30490
rect 4438 30438 4490 30490
rect 34966 30438 35018 30490
rect 35030 30438 35082 30490
rect 35094 30438 35146 30490
rect 35158 30438 35210 30490
rect 7564 30379 7616 30388
rect 7564 30345 7573 30379
rect 7573 30345 7607 30379
rect 7607 30345 7616 30379
rect 7564 30336 7616 30345
rect 9128 30379 9180 30388
rect 9128 30345 9137 30379
rect 9137 30345 9171 30379
rect 9171 30345 9180 30379
rect 9128 30336 9180 30345
rect 9680 30336 9732 30388
rect 9956 30379 10008 30388
rect 9956 30345 9965 30379
rect 9965 30345 9999 30379
rect 9999 30345 10008 30379
rect 9956 30336 10008 30345
rect 11244 30336 11296 30388
rect 12072 30336 12124 30388
rect 12624 30336 12676 30388
rect 14188 30379 14240 30388
rect 14188 30345 14197 30379
rect 14197 30345 14231 30379
rect 14231 30345 14240 30379
rect 14188 30336 14240 30345
rect 16304 30379 16356 30388
rect 16304 30345 16313 30379
rect 16313 30345 16347 30379
rect 16347 30345 16356 30379
rect 16304 30336 16356 30345
rect 9588 30268 9640 30320
rect 11336 30268 11388 30320
rect 12716 30311 12768 30320
rect 12716 30277 12725 30311
rect 12725 30277 12759 30311
rect 12759 30277 12768 30311
rect 12716 30268 12768 30277
rect 7656 30243 7708 30252
rect 7656 30209 7665 30243
rect 7665 30209 7699 30243
rect 7699 30209 7708 30243
rect 7656 30200 7708 30209
rect 8116 30243 8168 30252
rect 8116 30209 8125 30243
rect 8125 30209 8159 30243
rect 8159 30209 8168 30243
rect 8116 30200 8168 30209
rect 8208 30200 8260 30252
rect 10600 30200 10652 30252
rect 13728 30268 13780 30320
rect 8300 30175 8352 30184
rect 8300 30141 8309 30175
rect 8309 30141 8343 30175
rect 8343 30141 8352 30175
rect 8300 30132 8352 30141
rect 8484 30132 8536 30184
rect 9220 30064 9272 30116
rect 10784 30107 10836 30116
rect 10784 30073 10793 30107
rect 10793 30073 10827 30107
rect 10827 30073 10836 30107
rect 13268 30200 13320 30252
rect 13820 30200 13872 30252
rect 14648 30200 14700 30252
rect 14832 30268 14884 30320
rect 15568 30268 15620 30320
rect 17408 30268 17460 30320
rect 17592 30268 17644 30320
rect 18236 30336 18288 30388
rect 20444 30336 20496 30388
rect 21180 30336 21232 30388
rect 21364 30336 21416 30388
rect 19064 30311 19116 30320
rect 12900 30132 12952 30184
rect 13084 30175 13136 30184
rect 13084 30141 13093 30175
rect 13093 30141 13127 30175
rect 13127 30141 13136 30175
rect 13084 30132 13136 30141
rect 14188 30132 14240 30184
rect 15016 30132 15068 30184
rect 10784 30064 10836 30073
rect 7472 29996 7524 30048
rect 9680 30039 9732 30048
rect 9680 30005 9689 30039
rect 9689 30005 9723 30039
rect 9723 30005 9732 30039
rect 9680 29996 9732 30005
rect 10324 30039 10376 30048
rect 10324 30005 10333 30039
rect 10333 30005 10367 30039
rect 10367 30005 10376 30039
rect 10324 29996 10376 30005
rect 10968 30039 11020 30048
rect 10968 30005 10977 30039
rect 10977 30005 11011 30039
rect 11011 30005 11020 30039
rect 10968 29996 11020 30005
rect 11336 30064 11388 30116
rect 11980 30064 12032 30116
rect 13728 30064 13780 30116
rect 13912 30064 13964 30116
rect 16396 30200 16448 30252
rect 17776 30200 17828 30252
rect 18052 30243 18104 30252
rect 18052 30209 18061 30243
rect 18061 30209 18095 30243
rect 18095 30209 18104 30243
rect 18052 30200 18104 30209
rect 19064 30277 19073 30311
rect 19073 30277 19107 30311
rect 19107 30277 19116 30311
rect 19064 30268 19116 30277
rect 20076 30268 20128 30320
rect 19984 30243 20036 30252
rect 19984 30209 19993 30243
rect 19993 30209 20027 30243
rect 20027 30209 20036 30243
rect 19984 30200 20036 30209
rect 20720 30268 20772 30320
rect 21272 30268 21324 30320
rect 22008 30311 22060 30320
rect 22008 30277 22017 30311
rect 22017 30277 22051 30311
rect 22051 30277 22060 30311
rect 22008 30268 22060 30277
rect 22560 30336 22612 30388
rect 23848 30268 23900 30320
rect 25872 30336 25924 30388
rect 27528 30336 27580 30388
rect 26608 30311 26660 30320
rect 26608 30277 26617 30311
rect 26617 30277 26651 30311
rect 26651 30277 26660 30311
rect 26608 30268 26660 30277
rect 27620 30268 27672 30320
rect 22192 30200 22244 30252
rect 24768 30200 24820 30252
rect 15292 30064 15344 30116
rect 15660 30064 15712 30116
rect 17040 30064 17092 30116
rect 17132 30064 17184 30116
rect 17868 30064 17920 30116
rect 18972 30132 19024 30184
rect 20076 30132 20128 30184
rect 18420 30107 18472 30116
rect 18420 30073 18429 30107
rect 18429 30073 18463 30107
rect 18463 30073 18472 30107
rect 18420 30064 18472 30073
rect 18788 30107 18840 30116
rect 18788 30073 18797 30107
rect 18797 30073 18831 30107
rect 18831 30073 18840 30107
rect 18788 30064 18840 30073
rect 20444 30132 20496 30184
rect 21180 30175 21232 30184
rect 21180 30141 21189 30175
rect 21189 30141 21223 30175
rect 21223 30141 21232 30175
rect 21180 30132 21232 30141
rect 11244 29996 11296 30048
rect 13084 29996 13136 30048
rect 13360 29996 13412 30048
rect 13820 29996 13872 30048
rect 14648 29996 14700 30048
rect 15016 30039 15068 30048
rect 15016 30005 15025 30039
rect 15025 30005 15059 30039
rect 15059 30005 15068 30039
rect 15016 29996 15068 30005
rect 15476 29996 15528 30048
rect 16212 29996 16264 30048
rect 16672 30039 16724 30048
rect 16672 30005 16681 30039
rect 16681 30005 16715 30039
rect 16715 30005 16724 30039
rect 18328 30039 18380 30048
rect 16672 29996 16724 30005
rect 18328 30005 18337 30039
rect 18337 30005 18371 30039
rect 18371 30005 18380 30039
rect 18328 29996 18380 30005
rect 18880 29996 18932 30048
rect 19248 29996 19300 30048
rect 20720 30064 20772 30116
rect 21732 30132 21784 30184
rect 23388 30132 23440 30184
rect 23940 30175 23992 30184
rect 23940 30141 23949 30175
rect 23949 30141 23983 30175
rect 23983 30141 23992 30175
rect 23940 30132 23992 30141
rect 22192 30064 22244 30116
rect 22836 30064 22888 30116
rect 24032 30064 24084 30116
rect 24216 30132 24268 30184
rect 26608 30132 26660 30184
rect 24492 30064 24544 30116
rect 20812 29996 20864 30048
rect 22560 29996 22612 30048
rect 23664 29996 23716 30048
rect 24124 29996 24176 30048
rect 24676 30039 24728 30048
rect 24676 30005 24685 30039
rect 24685 30005 24719 30039
rect 24719 30005 24728 30039
rect 24676 29996 24728 30005
rect 24952 29996 25004 30048
rect 25320 30064 25372 30116
rect 25872 30064 25924 30116
rect 25504 30039 25556 30048
rect 25504 30005 25513 30039
rect 25513 30005 25547 30039
rect 25547 30005 25556 30039
rect 25504 29996 25556 30005
rect 26240 30039 26292 30048
rect 26240 30005 26249 30039
rect 26249 30005 26283 30039
rect 26283 30005 26292 30039
rect 26240 29996 26292 30005
rect 27344 30107 27396 30116
rect 27344 30073 27353 30107
rect 27353 30073 27387 30107
rect 27387 30073 27396 30107
rect 27344 30064 27396 30073
rect 28080 30107 28132 30116
rect 28080 30073 28089 30107
rect 28089 30073 28123 30107
rect 28123 30073 28132 30107
rect 28080 30064 28132 30073
rect 28724 29996 28776 30048
rect 29460 30039 29512 30048
rect 29460 30005 29469 30039
rect 29469 30005 29503 30039
rect 29503 30005 29512 30039
rect 29460 29996 29512 30005
rect 19606 29894 19658 29946
rect 19670 29894 19722 29946
rect 19734 29894 19786 29946
rect 19798 29894 19850 29946
rect 1676 29792 1728 29844
rect 2872 29792 2924 29844
rect 6736 29835 6788 29844
rect 6736 29801 6745 29835
rect 6745 29801 6779 29835
rect 6779 29801 6788 29835
rect 6736 29792 6788 29801
rect 9496 29835 9548 29844
rect 9496 29801 9505 29835
rect 9505 29801 9539 29835
rect 9539 29801 9548 29835
rect 9496 29792 9548 29801
rect 10876 29792 10928 29844
rect 11060 29792 11112 29844
rect 11244 29792 11296 29844
rect 11888 29792 11940 29844
rect 12072 29792 12124 29844
rect 13268 29835 13320 29844
rect 8484 29767 8536 29776
rect 8484 29733 8493 29767
rect 8493 29733 8527 29767
rect 8527 29733 8536 29767
rect 8484 29724 8536 29733
rect 13268 29801 13277 29835
rect 13277 29801 13311 29835
rect 13311 29801 13320 29835
rect 13268 29792 13320 29801
rect 14832 29835 14884 29844
rect 14832 29801 14841 29835
rect 14841 29801 14875 29835
rect 14875 29801 14884 29835
rect 14832 29792 14884 29801
rect 15476 29835 15528 29844
rect 15476 29801 15485 29835
rect 15485 29801 15519 29835
rect 15519 29801 15528 29835
rect 15476 29792 15528 29801
rect 15660 29792 15712 29844
rect 16396 29792 16448 29844
rect 16672 29792 16724 29844
rect 17868 29792 17920 29844
rect 18696 29792 18748 29844
rect 20076 29792 20128 29844
rect 20720 29792 20772 29844
rect 20996 29792 21048 29844
rect 21640 29792 21692 29844
rect 22284 29835 22336 29844
rect 22284 29801 22293 29835
rect 22293 29801 22327 29835
rect 22327 29801 22336 29835
rect 22284 29792 22336 29801
rect 23756 29792 23808 29844
rect 24308 29792 24360 29844
rect 24860 29792 24912 29844
rect 25688 29792 25740 29844
rect 7196 29656 7248 29708
rect 8116 29656 8168 29708
rect 9128 29699 9180 29708
rect 9128 29665 9137 29699
rect 9137 29665 9171 29699
rect 9171 29665 9180 29699
rect 9128 29656 9180 29665
rect 9772 29699 9824 29708
rect 9772 29665 9781 29699
rect 9781 29665 9815 29699
rect 9815 29665 9824 29699
rect 9772 29656 9824 29665
rect 11060 29656 11112 29708
rect 11244 29656 11296 29708
rect 12624 29724 12676 29776
rect 15016 29724 15068 29776
rect 16304 29724 16356 29776
rect 16580 29767 16632 29776
rect 16580 29733 16589 29767
rect 16589 29733 16623 29767
rect 16623 29733 16632 29767
rect 16580 29724 16632 29733
rect 18420 29724 18472 29776
rect 20444 29724 20496 29776
rect 21548 29724 21600 29776
rect 1676 29631 1728 29640
rect 1676 29597 1685 29631
rect 1685 29597 1719 29631
rect 1719 29597 1728 29631
rect 1676 29588 1728 29597
rect 6644 29588 6696 29640
rect 11704 29588 11756 29640
rect 10968 29563 11020 29572
rect 10968 29529 10977 29563
rect 10977 29529 11011 29563
rect 11011 29529 11020 29563
rect 10968 29520 11020 29529
rect 13728 29656 13780 29708
rect 14096 29656 14148 29708
rect 15200 29656 15252 29708
rect 18052 29699 18104 29708
rect 13360 29631 13412 29640
rect 13360 29597 13369 29631
rect 13369 29597 13403 29631
rect 13403 29597 13412 29631
rect 13360 29588 13412 29597
rect 14004 29588 14056 29640
rect 10876 29452 10928 29504
rect 11704 29495 11756 29504
rect 11704 29461 11713 29495
rect 11713 29461 11747 29495
rect 11747 29461 11756 29495
rect 11704 29452 11756 29461
rect 11888 29520 11940 29572
rect 12900 29520 12952 29572
rect 14096 29520 14148 29572
rect 15660 29588 15712 29640
rect 18052 29665 18061 29699
rect 18061 29665 18095 29699
rect 18095 29665 18104 29699
rect 18052 29656 18104 29665
rect 19524 29699 19576 29708
rect 19524 29665 19533 29699
rect 19533 29665 19567 29699
rect 19567 29665 19576 29699
rect 19524 29656 19576 29665
rect 22008 29656 22060 29708
rect 22100 29656 22152 29708
rect 23388 29724 23440 29776
rect 23480 29724 23532 29776
rect 24768 29767 24820 29776
rect 23112 29656 23164 29708
rect 24768 29733 24777 29767
rect 24777 29733 24811 29767
rect 24811 29733 24820 29767
rect 24768 29724 24820 29733
rect 25320 29767 25372 29776
rect 25320 29733 25329 29767
rect 25329 29733 25363 29767
rect 25363 29733 25372 29767
rect 27712 29792 27764 29844
rect 27896 29792 27948 29844
rect 25320 29724 25372 29733
rect 26332 29724 26384 29776
rect 25688 29656 25740 29708
rect 25872 29656 25924 29708
rect 26516 29699 26568 29708
rect 26516 29665 26525 29699
rect 26525 29665 26559 29699
rect 26559 29665 26568 29699
rect 26516 29656 26568 29665
rect 26976 29724 27028 29776
rect 27252 29767 27304 29776
rect 27252 29733 27261 29767
rect 27261 29733 27295 29767
rect 27295 29733 27304 29767
rect 27252 29724 27304 29733
rect 27896 29656 27948 29708
rect 16948 29631 17000 29640
rect 16948 29597 16957 29631
rect 16957 29597 16991 29631
rect 16991 29597 17000 29631
rect 16948 29588 17000 29597
rect 17776 29631 17828 29640
rect 17776 29597 17785 29631
rect 17785 29597 17819 29631
rect 17819 29597 17828 29631
rect 17776 29588 17828 29597
rect 19064 29588 19116 29640
rect 19708 29588 19760 29640
rect 21180 29588 21232 29640
rect 21364 29588 21416 29640
rect 21732 29588 21784 29640
rect 27620 29588 27672 29640
rect 20444 29520 20496 29572
rect 12440 29452 12492 29504
rect 12808 29495 12860 29504
rect 12808 29461 12817 29495
rect 12817 29461 12851 29495
rect 12851 29461 12860 29495
rect 12808 29452 12860 29461
rect 13268 29452 13320 29504
rect 15752 29452 15804 29504
rect 18788 29452 18840 29504
rect 20628 29495 20680 29504
rect 20628 29461 20637 29495
rect 20637 29461 20671 29495
rect 20671 29461 20680 29495
rect 20628 29452 20680 29461
rect 21180 29452 21232 29504
rect 21548 29452 21600 29504
rect 22468 29452 22520 29504
rect 22928 29495 22980 29504
rect 22928 29461 22937 29495
rect 22937 29461 22971 29495
rect 22971 29461 22980 29495
rect 22928 29452 22980 29461
rect 23940 29520 23992 29572
rect 26608 29520 26660 29572
rect 27252 29520 27304 29572
rect 26332 29452 26384 29504
rect 26976 29452 27028 29504
rect 28264 29452 28316 29504
rect 28724 29495 28776 29504
rect 28724 29461 28733 29495
rect 28733 29461 28767 29495
rect 28767 29461 28776 29495
rect 28724 29452 28776 29461
rect 4246 29350 4298 29402
rect 4310 29350 4362 29402
rect 4374 29350 4426 29402
rect 4438 29350 4490 29402
rect 34966 29350 35018 29402
rect 35030 29350 35082 29402
rect 35094 29350 35146 29402
rect 35158 29350 35210 29402
rect 1768 29248 1820 29300
rect 2780 29248 2832 29300
rect 6644 29291 6696 29300
rect 6644 29257 6653 29291
rect 6653 29257 6687 29291
rect 6687 29257 6696 29291
rect 6644 29248 6696 29257
rect 7012 29248 7064 29300
rect 7196 29248 7248 29300
rect 7288 29180 7340 29232
rect 6644 29044 6696 29096
rect 6920 29044 6972 29096
rect 7472 29112 7524 29164
rect 7840 29044 7892 29096
rect 8024 29044 8076 29096
rect 8484 29248 8536 29300
rect 9220 29248 9272 29300
rect 9312 29248 9364 29300
rect 9772 29291 9824 29300
rect 9772 29257 9781 29291
rect 9781 29257 9815 29291
rect 9815 29257 9824 29291
rect 9772 29248 9824 29257
rect 10232 29291 10284 29300
rect 10232 29257 10241 29291
rect 10241 29257 10275 29291
rect 10275 29257 10284 29291
rect 10232 29248 10284 29257
rect 10508 29291 10560 29300
rect 10508 29257 10517 29291
rect 10517 29257 10551 29291
rect 10551 29257 10560 29291
rect 10508 29248 10560 29257
rect 11888 29291 11940 29300
rect 11888 29257 11897 29291
rect 11897 29257 11931 29291
rect 11931 29257 11940 29291
rect 11888 29248 11940 29257
rect 12256 29291 12308 29300
rect 12256 29257 12265 29291
rect 12265 29257 12299 29291
rect 12299 29257 12308 29291
rect 12256 29248 12308 29257
rect 12440 29248 12492 29300
rect 15292 29248 15344 29300
rect 15476 29248 15528 29300
rect 15752 29248 15804 29300
rect 16672 29248 16724 29300
rect 17040 29248 17092 29300
rect 7380 28976 7432 29028
rect 8300 28976 8352 29028
rect 8484 28976 8536 29028
rect 8576 28976 8628 29028
rect 9588 29180 9640 29232
rect 12164 29180 12216 29232
rect 13728 29180 13780 29232
rect 8760 29112 8812 29164
rect 10600 29112 10652 29164
rect 9220 29044 9272 29096
rect 10324 29087 10376 29096
rect 10324 29053 10333 29087
rect 10333 29053 10367 29087
rect 10367 29053 10376 29087
rect 10876 29087 10928 29096
rect 10324 29044 10376 29053
rect 10876 29053 10885 29087
rect 10885 29053 10919 29087
rect 10919 29053 10928 29087
rect 10876 29044 10928 29053
rect 12256 29044 12308 29096
rect 13360 29112 13412 29164
rect 13820 29087 13872 29096
rect 11060 28976 11112 29028
rect 12992 28976 13044 29028
rect 13820 29053 13829 29087
rect 13829 29053 13863 29087
rect 13863 29053 13872 29087
rect 13820 29044 13872 29053
rect 14372 29180 14424 29232
rect 15660 29180 15712 29232
rect 14188 29112 14240 29164
rect 15016 29112 15068 29164
rect 15752 29112 15804 29164
rect 15936 29112 15988 29164
rect 14096 29044 14148 29096
rect 14372 29087 14424 29096
rect 14372 29053 14381 29087
rect 14381 29053 14415 29087
rect 14415 29053 14424 29087
rect 14372 29044 14424 29053
rect 15108 29044 15160 29096
rect 17132 29180 17184 29232
rect 17408 29248 17460 29300
rect 17776 29248 17828 29300
rect 19156 29248 19208 29300
rect 19708 29291 19760 29300
rect 19708 29257 19717 29291
rect 19717 29257 19751 29291
rect 19751 29257 19760 29291
rect 19708 29248 19760 29257
rect 19800 29248 19852 29300
rect 16580 29112 16632 29164
rect 18052 29112 18104 29164
rect 16672 29087 16724 29096
rect 16672 29053 16681 29087
rect 16681 29053 16715 29087
rect 16715 29053 16724 29087
rect 16672 29044 16724 29053
rect 18788 29044 18840 29096
rect 13912 28976 13964 29028
rect 14188 28976 14240 29028
rect 14648 28976 14700 29028
rect 16212 28976 16264 29028
rect 17132 29019 17184 29028
rect 1676 28951 1728 28960
rect 1676 28917 1685 28951
rect 1685 28917 1719 28951
rect 1719 28917 1728 28951
rect 1676 28908 1728 28917
rect 7656 28908 7708 28960
rect 8392 28908 8444 28960
rect 8668 28951 8720 28960
rect 8668 28917 8677 28951
rect 8677 28917 8711 28951
rect 8711 28917 8720 28951
rect 8668 28908 8720 28917
rect 12440 28908 12492 28960
rect 13544 28908 13596 28960
rect 15936 28908 15988 28960
rect 17132 28985 17141 29019
rect 17141 28985 17175 29019
rect 17175 28985 17184 29019
rect 17132 28976 17184 28985
rect 18420 29019 18472 29028
rect 18420 28985 18429 29019
rect 18429 28985 18463 29019
rect 18463 28985 18472 29019
rect 18420 28976 18472 28985
rect 18604 29019 18656 29028
rect 18604 28985 18613 29019
rect 18613 28985 18647 29019
rect 18647 28985 18656 29019
rect 18604 28976 18656 28985
rect 19156 29112 19208 29164
rect 20904 29248 20956 29300
rect 23112 29291 23164 29300
rect 20996 29180 21048 29232
rect 21548 29180 21600 29232
rect 23112 29257 23121 29291
rect 23121 29257 23155 29291
rect 23155 29257 23164 29291
rect 23112 29248 23164 29257
rect 23480 29291 23532 29300
rect 23480 29257 23489 29291
rect 23489 29257 23523 29291
rect 23523 29257 23532 29291
rect 23480 29248 23532 29257
rect 21916 29155 21968 29164
rect 21916 29121 21925 29155
rect 21925 29121 21959 29155
rect 21959 29121 21968 29155
rect 21916 29112 21968 29121
rect 18052 28908 18104 28960
rect 18696 28908 18748 28960
rect 19156 28976 19208 29028
rect 20628 29044 20680 29096
rect 21088 29019 21140 29028
rect 21088 28985 21097 29019
rect 21097 28985 21131 29019
rect 21131 28985 21140 29019
rect 21088 28976 21140 28985
rect 22652 29112 22704 29164
rect 23480 29112 23532 29164
rect 23848 29112 23900 29164
rect 22468 29044 22520 29096
rect 23756 29044 23808 29096
rect 25320 29248 25372 29300
rect 25872 29248 25924 29300
rect 26516 29248 26568 29300
rect 27068 29180 27120 29232
rect 26240 29155 26292 29164
rect 26240 29121 26249 29155
rect 26249 29121 26283 29155
rect 26283 29121 26292 29155
rect 26240 29112 26292 29121
rect 28356 29248 28408 29300
rect 28724 29248 28776 29300
rect 27896 29180 27948 29232
rect 28172 29180 28224 29232
rect 26792 29044 26844 29096
rect 28080 29087 28132 29096
rect 22652 29019 22704 29028
rect 22652 28985 22661 29019
rect 22661 28985 22695 29019
rect 22695 28985 22704 29019
rect 22652 28976 22704 28985
rect 25320 29019 25372 29028
rect 25320 28985 25329 29019
rect 25329 28985 25363 29019
rect 25363 28985 25372 29019
rect 25320 28976 25372 28985
rect 26332 29019 26384 29028
rect 26332 28985 26341 29019
rect 26341 28985 26375 29019
rect 26375 28985 26384 29019
rect 26332 28976 26384 28985
rect 28080 29053 28089 29087
rect 28089 29053 28123 29087
rect 28123 29053 28132 29087
rect 28080 29044 28132 29053
rect 20444 28908 20496 28960
rect 22100 28951 22152 28960
rect 22100 28917 22109 28951
rect 22109 28917 22143 28951
rect 22143 28917 22152 28951
rect 22100 28908 22152 28917
rect 26056 28908 26108 28960
rect 27436 28976 27488 29028
rect 28724 28976 28776 29028
rect 29000 29019 29052 29028
rect 29000 28985 29009 29019
rect 29009 28985 29043 29019
rect 29043 28985 29052 29019
rect 29000 28976 29052 28985
rect 19606 28806 19658 28858
rect 19670 28806 19722 28858
rect 19734 28806 19786 28858
rect 19798 28806 19850 28858
rect 8024 28704 8076 28756
rect 8484 28704 8536 28756
rect 8944 28704 8996 28756
rect 10600 28747 10652 28756
rect 10600 28713 10609 28747
rect 10609 28713 10643 28747
rect 10643 28713 10652 28747
rect 10600 28704 10652 28713
rect 11796 28747 11848 28756
rect 11796 28713 11805 28747
rect 11805 28713 11839 28747
rect 11839 28713 11848 28747
rect 11796 28704 11848 28713
rect 12348 28747 12400 28756
rect 12348 28713 12357 28747
rect 12357 28713 12391 28747
rect 12391 28713 12400 28747
rect 12348 28704 12400 28713
rect 12900 28704 12952 28756
rect 7564 28679 7616 28688
rect 7564 28645 7573 28679
rect 7573 28645 7607 28679
rect 7607 28645 7616 28679
rect 7564 28636 7616 28645
rect 9128 28679 9180 28688
rect 9128 28645 9137 28679
rect 9137 28645 9171 28679
rect 9171 28645 9180 28679
rect 9128 28636 9180 28645
rect 12256 28636 12308 28688
rect 12808 28636 12860 28688
rect 13452 28704 13504 28756
rect 14004 28704 14056 28756
rect 15108 28704 15160 28756
rect 16304 28704 16356 28756
rect 18696 28704 18748 28756
rect 18880 28704 18932 28756
rect 20444 28704 20496 28756
rect 8024 28568 8076 28620
rect 8668 28568 8720 28620
rect 8944 28568 8996 28620
rect 9772 28568 9824 28620
rect 10784 28611 10836 28620
rect 10784 28577 10793 28611
rect 10793 28577 10827 28611
rect 10827 28577 10836 28611
rect 10784 28568 10836 28577
rect 12992 28568 13044 28620
rect 14372 28636 14424 28688
rect 18972 28636 19024 28688
rect 19984 28679 20036 28688
rect 19984 28645 19993 28679
rect 19993 28645 20027 28679
rect 20027 28645 20036 28679
rect 21180 28704 21232 28756
rect 21916 28747 21968 28756
rect 21916 28713 21925 28747
rect 21925 28713 21959 28747
rect 21959 28713 21968 28747
rect 21916 28704 21968 28713
rect 22468 28704 22520 28756
rect 23112 28704 23164 28756
rect 23664 28704 23716 28756
rect 23940 28747 23992 28756
rect 23940 28713 23949 28747
rect 23949 28713 23983 28747
rect 23983 28713 23992 28747
rect 23940 28704 23992 28713
rect 24860 28704 24912 28756
rect 25596 28704 25648 28756
rect 26056 28704 26108 28756
rect 26240 28747 26292 28756
rect 26240 28713 26249 28747
rect 26249 28713 26283 28747
rect 26283 28713 26292 28747
rect 26240 28704 26292 28713
rect 20720 28679 20772 28688
rect 19984 28636 20036 28645
rect 20720 28645 20729 28679
rect 20729 28645 20763 28679
rect 20763 28645 20772 28679
rect 20720 28636 20772 28645
rect 20904 28636 20956 28688
rect 21456 28636 21508 28688
rect 22100 28636 22152 28688
rect 14464 28568 14516 28620
rect 15200 28568 15252 28620
rect 16764 28568 16816 28620
rect 17776 28568 17828 28620
rect 18328 28568 18380 28620
rect 18880 28568 18932 28620
rect 21180 28611 21232 28620
rect 21180 28577 21189 28611
rect 21189 28577 21223 28611
rect 21223 28577 21232 28611
rect 23388 28636 23440 28688
rect 27344 28704 27396 28756
rect 27712 28704 27764 28756
rect 28908 28704 28960 28756
rect 29000 28747 29052 28756
rect 29000 28713 29009 28747
rect 29009 28713 29043 28747
rect 29043 28713 29052 28747
rect 29000 28704 29052 28713
rect 26608 28636 26660 28688
rect 26792 28636 26844 28688
rect 21180 28568 21232 28577
rect 23112 28568 23164 28620
rect 24216 28611 24268 28620
rect 24216 28577 24225 28611
rect 24225 28577 24259 28611
rect 24259 28577 24268 28611
rect 24216 28568 24268 28577
rect 28172 28568 28224 28620
rect 32036 28568 32088 28620
rect 32496 28568 32548 28620
rect 7840 28500 7892 28552
rect 8392 28500 8444 28552
rect 12808 28543 12860 28552
rect 12808 28509 12817 28543
rect 12817 28509 12851 28543
rect 12851 28509 12860 28543
rect 12808 28500 12860 28509
rect 13452 28500 13504 28552
rect 14648 28500 14700 28552
rect 13728 28432 13780 28484
rect 14004 28432 14056 28484
rect 15936 28500 15988 28552
rect 18604 28500 18656 28552
rect 18972 28500 19024 28552
rect 19340 28500 19392 28552
rect 19800 28432 19852 28484
rect 20444 28500 20496 28552
rect 21272 28500 21324 28552
rect 21640 28543 21692 28552
rect 21640 28509 21649 28543
rect 21649 28509 21683 28543
rect 21683 28509 21692 28543
rect 21640 28500 21692 28509
rect 21916 28500 21968 28552
rect 22560 28500 22612 28552
rect 26792 28500 26844 28552
rect 32772 28500 32824 28552
rect 22008 28432 22060 28484
rect 26516 28432 26568 28484
rect 27344 28432 27396 28484
rect 27620 28432 27672 28484
rect 6920 28407 6972 28416
rect 6920 28373 6929 28407
rect 6929 28373 6963 28407
rect 6963 28373 6972 28407
rect 6920 28364 6972 28373
rect 7288 28407 7340 28416
rect 7288 28373 7297 28407
rect 7297 28373 7331 28407
rect 7331 28373 7340 28407
rect 7288 28364 7340 28373
rect 11060 28364 11112 28416
rect 13912 28364 13964 28416
rect 15476 28364 15528 28416
rect 16672 28407 16724 28416
rect 16672 28373 16681 28407
rect 16681 28373 16715 28407
rect 16715 28373 16724 28407
rect 16672 28364 16724 28373
rect 17592 28407 17644 28416
rect 17592 28373 17601 28407
rect 17601 28373 17635 28407
rect 17635 28373 17644 28407
rect 17592 28364 17644 28373
rect 17960 28407 18012 28416
rect 17960 28373 17969 28407
rect 17969 28373 18003 28407
rect 18003 28373 18012 28407
rect 17960 28364 18012 28373
rect 18604 28364 18656 28416
rect 21272 28364 21324 28416
rect 23940 28364 23992 28416
rect 24308 28407 24360 28416
rect 24308 28373 24317 28407
rect 24317 28373 24351 28407
rect 24351 28373 24360 28407
rect 24308 28364 24360 28373
rect 24768 28364 24820 28416
rect 25044 28364 25096 28416
rect 25596 28364 25648 28416
rect 25872 28364 25924 28416
rect 27160 28407 27212 28416
rect 27160 28373 27169 28407
rect 27169 28373 27203 28407
rect 27203 28373 27212 28407
rect 27160 28364 27212 28373
rect 28540 28407 28592 28416
rect 28540 28373 28549 28407
rect 28549 28373 28583 28407
rect 28583 28373 28592 28407
rect 28540 28364 28592 28373
rect 33784 28407 33836 28416
rect 33784 28373 33793 28407
rect 33793 28373 33827 28407
rect 33827 28373 33836 28407
rect 33784 28364 33836 28373
rect 4246 28262 4298 28314
rect 4310 28262 4362 28314
rect 4374 28262 4426 28314
rect 4438 28262 4490 28314
rect 34966 28262 35018 28314
rect 35030 28262 35082 28314
rect 35094 28262 35146 28314
rect 35158 28262 35210 28314
rect 1676 28203 1728 28212
rect 1676 28169 1685 28203
rect 1685 28169 1719 28203
rect 1719 28169 1728 28203
rect 1676 28160 1728 28169
rect 2228 28203 2280 28212
rect 2228 28169 2237 28203
rect 2237 28169 2271 28203
rect 2271 28169 2280 28203
rect 2228 28160 2280 28169
rect 8668 28160 8720 28212
rect 9496 28203 9548 28212
rect 9496 28169 9505 28203
rect 9505 28169 9539 28203
rect 9539 28169 9548 28203
rect 9496 28160 9548 28169
rect 10324 28160 10376 28212
rect 10508 28203 10560 28212
rect 10508 28169 10517 28203
rect 10517 28169 10551 28203
rect 10551 28169 10560 28203
rect 10508 28160 10560 28169
rect 10784 28203 10836 28212
rect 10784 28169 10793 28203
rect 10793 28169 10827 28203
rect 10827 28169 10836 28203
rect 10784 28160 10836 28169
rect 12440 28160 12492 28212
rect 14740 28160 14792 28212
rect 15108 28160 15160 28212
rect 17776 28203 17828 28212
rect 17776 28169 17785 28203
rect 17785 28169 17819 28203
rect 17819 28169 17828 28203
rect 17776 28160 17828 28169
rect 18236 28160 18288 28212
rect 18880 28203 18932 28212
rect 18880 28169 18889 28203
rect 18889 28169 18923 28203
rect 18923 28169 18932 28203
rect 18880 28160 18932 28169
rect 19800 28160 19852 28212
rect 20628 28160 20680 28212
rect 20996 28160 21048 28212
rect 21916 28160 21968 28212
rect 23940 28203 23992 28212
rect 23940 28169 23949 28203
rect 23949 28169 23983 28203
rect 23983 28169 23992 28203
rect 23940 28160 23992 28169
rect 25872 28203 25924 28212
rect 25872 28169 25881 28203
rect 25881 28169 25915 28203
rect 25915 28169 25924 28203
rect 25872 28160 25924 28169
rect 26608 28160 26660 28212
rect 27436 28160 27488 28212
rect 28172 28160 28224 28212
rect 29184 28160 29236 28212
rect 30012 28160 30064 28212
rect 32496 28203 32548 28212
rect 32496 28169 32505 28203
rect 32505 28169 32539 28203
rect 32539 28169 32548 28203
rect 32496 28160 32548 28169
rect 32772 28203 32824 28212
rect 32772 28169 32781 28203
rect 32781 28169 32815 28203
rect 32815 28169 32824 28203
rect 32772 28160 32824 28169
rect 8576 28092 8628 28144
rect 11612 28135 11664 28144
rect 11612 28101 11621 28135
rect 11621 28101 11655 28135
rect 11655 28101 11664 28135
rect 11612 28092 11664 28101
rect 14188 28092 14240 28144
rect 8484 28024 8536 28076
rect 9128 28067 9180 28076
rect 9128 28033 9137 28067
rect 9137 28033 9171 28067
rect 9171 28033 9180 28067
rect 9128 28024 9180 28033
rect 9588 28024 9640 28076
rect 1584 27999 1636 28008
rect 1584 27965 1593 27999
rect 1593 27965 1627 27999
rect 1627 27965 1636 27999
rect 1584 27956 1636 27965
rect 8944 27956 8996 28008
rect 10968 28024 11020 28076
rect 13176 28024 13228 28076
rect 13544 28024 13596 28076
rect 14004 28024 14056 28076
rect 7288 27931 7340 27940
rect 7288 27897 7297 27931
rect 7297 27897 7331 27931
rect 7331 27897 7340 27931
rect 7288 27888 7340 27897
rect 8392 27888 8444 27940
rect 8024 27863 8076 27872
rect 8024 27829 8033 27863
rect 8033 27829 8067 27863
rect 8067 27829 8076 27863
rect 8024 27820 8076 27829
rect 9864 27863 9916 27872
rect 9864 27829 9873 27863
rect 9873 27829 9907 27863
rect 9907 27829 9916 27863
rect 9864 27820 9916 27829
rect 12164 27956 12216 28008
rect 13728 27956 13780 28008
rect 15108 28024 15160 28076
rect 14004 27888 14056 27940
rect 14648 27956 14700 28008
rect 14464 27888 14516 27940
rect 14832 27956 14884 28008
rect 11336 27820 11388 27872
rect 11428 27820 11480 27872
rect 12440 27820 12492 27872
rect 12900 27820 12952 27872
rect 13452 27820 13504 27872
rect 14188 27820 14240 27872
rect 16764 28092 16816 28144
rect 17960 28092 18012 28144
rect 16120 28024 16172 28076
rect 16304 28067 16356 28076
rect 16304 28033 16313 28067
rect 16313 28033 16347 28067
rect 16347 28033 16356 28067
rect 16304 28024 16356 28033
rect 17224 28024 17276 28076
rect 16672 27956 16724 28008
rect 15936 27820 15988 27872
rect 18880 27956 18932 28008
rect 20260 28024 20312 28076
rect 20812 28092 20864 28144
rect 23112 28135 23164 28144
rect 23112 28101 23121 28135
rect 23121 28101 23155 28135
rect 23155 28101 23164 28135
rect 23112 28092 23164 28101
rect 24032 28092 24084 28144
rect 19800 27999 19852 28008
rect 19800 27965 19809 27999
rect 19809 27965 19843 27999
rect 19843 27965 19852 27999
rect 19800 27956 19852 27965
rect 20996 28024 21048 28076
rect 21732 28024 21784 28076
rect 23296 28024 23348 28076
rect 20812 27956 20864 28008
rect 23112 27956 23164 28008
rect 24676 27999 24728 28008
rect 20904 27888 20956 27940
rect 21732 27888 21784 27940
rect 17040 27863 17092 27872
rect 17040 27829 17049 27863
rect 17049 27829 17083 27863
rect 17083 27829 17092 27863
rect 17040 27820 17092 27829
rect 20076 27820 20128 27872
rect 20260 27820 20312 27872
rect 20444 27820 20496 27872
rect 20812 27820 20864 27872
rect 21180 27820 21232 27872
rect 21916 27863 21968 27872
rect 21916 27829 21925 27863
rect 21925 27829 21959 27863
rect 21959 27829 21968 27863
rect 21916 27820 21968 27829
rect 22192 27888 22244 27940
rect 22928 27888 22980 27940
rect 23940 27888 23992 27940
rect 24676 27965 24685 27999
rect 24685 27965 24719 27999
rect 24719 27965 24728 27999
rect 24676 27956 24728 27965
rect 24860 27999 24912 28008
rect 24860 27965 24869 27999
rect 24869 27965 24903 27999
rect 24903 27965 24912 27999
rect 24860 27956 24912 27965
rect 25596 28024 25648 28076
rect 27068 28024 27120 28076
rect 29276 27999 29328 28008
rect 29276 27965 29285 27999
rect 29285 27965 29319 27999
rect 29319 27965 29328 27999
rect 29276 27956 29328 27965
rect 22468 27820 22520 27872
rect 25044 27820 25096 27872
rect 26516 27863 26568 27872
rect 26516 27829 26525 27863
rect 26525 27829 26559 27863
rect 26559 27829 26568 27863
rect 26516 27820 26568 27829
rect 29460 27863 29512 27872
rect 29460 27829 29469 27863
rect 29469 27829 29503 27863
rect 29503 27829 29512 27863
rect 29460 27820 29512 27829
rect 19606 27718 19658 27770
rect 19670 27718 19722 27770
rect 19734 27718 19786 27770
rect 19798 27718 19850 27770
rect 8300 27616 8352 27668
rect 10784 27659 10836 27668
rect 10784 27625 10793 27659
rect 10793 27625 10827 27659
rect 10827 27625 10836 27659
rect 10784 27616 10836 27625
rect 12440 27659 12492 27668
rect 12440 27625 12449 27659
rect 12449 27625 12483 27659
rect 12483 27625 12492 27659
rect 12440 27616 12492 27625
rect 13360 27616 13412 27668
rect 14096 27616 14148 27668
rect 17316 27616 17368 27668
rect 10508 27591 10560 27600
rect 10508 27557 10517 27591
rect 10517 27557 10551 27591
rect 10551 27557 10560 27591
rect 10508 27548 10560 27557
rect 12992 27591 13044 27600
rect 6000 27480 6052 27532
rect 6828 27480 6880 27532
rect 10600 27523 10652 27532
rect 10600 27489 10609 27523
rect 10609 27489 10643 27523
rect 10643 27489 10652 27523
rect 10600 27480 10652 27489
rect 11704 27523 11756 27532
rect 11704 27489 11713 27523
rect 11713 27489 11747 27523
rect 11747 27489 11756 27523
rect 11704 27480 11756 27489
rect 12624 27480 12676 27532
rect 12992 27557 13001 27591
rect 13001 27557 13035 27591
rect 13035 27557 13044 27591
rect 12992 27548 13044 27557
rect 14924 27548 14976 27600
rect 15108 27548 15160 27600
rect 16856 27548 16908 27600
rect 17408 27591 17460 27600
rect 17408 27557 17417 27591
rect 17417 27557 17451 27591
rect 17451 27557 17460 27591
rect 17408 27548 17460 27557
rect 18328 27616 18380 27668
rect 18604 27616 18656 27668
rect 20260 27616 20312 27668
rect 20352 27616 20404 27668
rect 17776 27591 17828 27600
rect 17776 27557 17785 27591
rect 17785 27557 17819 27591
rect 17819 27557 17828 27591
rect 17776 27548 17828 27557
rect 18052 27548 18104 27600
rect 13728 27480 13780 27532
rect 13820 27523 13872 27532
rect 13820 27489 13829 27523
rect 13829 27489 13863 27523
rect 13863 27489 13872 27523
rect 13820 27480 13872 27489
rect 7104 27412 7156 27464
rect 7472 27412 7524 27464
rect 9128 27412 9180 27464
rect 10140 27455 10192 27464
rect 10140 27421 10149 27455
rect 10149 27421 10183 27455
rect 10183 27421 10192 27455
rect 10140 27412 10192 27421
rect 12256 27412 12308 27464
rect 13544 27455 13596 27464
rect 13544 27421 13553 27455
rect 13553 27421 13587 27455
rect 13587 27421 13596 27455
rect 13544 27412 13596 27421
rect 1584 27319 1636 27328
rect 1584 27285 1593 27319
rect 1593 27285 1627 27319
rect 1627 27285 1636 27319
rect 1584 27276 1636 27285
rect 8300 27319 8352 27328
rect 8300 27285 8309 27319
rect 8309 27285 8343 27319
rect 8343 27285 8352 27319
rect 8300 27276 8352 27285
rect 8392 27276 8444 27328
rect 8944 27276 8996 27328
rect 11888 27319 11940 27328
rect 11888 27285 11897 27319
rect 11897 27285 11931 27319
rect 11931 27285 11940 27319
rect 11888 27276 11940 27285
rect 13544 27276 13596 27328
rect 14740 27480 14792 27532
rect 15844 27523 15896 27532
rect 15844 27489 15853 27523
rect 15853 27489 15887 27523
rect 15887 27489 15896 27523
rect 15844 27480 15896 27489
rect 14464 27455 14516 27464
rect 14464 27421 14473 27455
rect 14473 27421 14507 27455
rect 14507 27421 14516 27455
rect 14464 27412 14516 27421
rect 16120 27523 16172 27532
rect 16120 27489 16129 27523
rect 16129 27489 16163 27523
rect 16163 27489 16172 27523
rect 16120 27480 16172 27489
rect 17592 27523 17644 27532
rect 16212 27412 16264 27464
rect 16304 27412 16356 27464
rect 14648 27344 14700 27396
rect 15476 27344 15528 27396
rect 17592 27489 17601 27523
rect 17601 27489 17635 27523
rect 17635 27489 17644 27523
rect 17592 27480 17644 27489
rect 17868 27480 17920 27532
rect 18972 27523 19024 27532
rect 18972 27489 18981 27523
rect 18981 27489 19015 27523
rect 19015 27489 19024 27523
rect 18972 27480 19024 27489
rect 19432 27548 19484 27600
rect 19984 27591 20036 27600
rect 19984 27557 19993 27591
rect 19993 27557 20027 27591
rect 20027 27557 20036 27591
rect 19984 27548 20036 27557
rect 20628 27548 20680 27600
rect 19524 27480 19576 27532
rect 21272 27616 21324 27668
rect 21916 27616 21968 27668
rect 22560 27616 22612 27668
rect 21640 27548 21692 27600
rect 21088 27523 21140 27532
rect 21088 27489 21094 27523
rect 21094 27489 21140 27523
rect 21088 27480 21140 27489
rect 21732 27480 21784 27532
rect 18052 27412 18104 27464
rect 21272 27455 21324 27464
rect 21272 27421 21281 27455
rect 21281 27421 21315 27455
rect 21315 27421 21324 27455
rect 21272 27412 21324 27421
rect 22008 27412 22060 27464
rect 22284 27412 22336 27464
rect 19156 27387 19208 27396
rect 19156 27353 19180 27387
rect 19180 27353 19208 27387
rect 19156 27344 19208 27353
rect 22744 27480 22796 27532
rect 23388 27412 23440 27464
rect 24124 27616 24176 27668
rect 24676 27616 24728 27668
rect 23664 27548 23716 27600
rect 24032 27591 24084 27600
rect 24032 27557 24041 27591
rect 24041 27557 24075 27591
rect 24075 27557 24084 27591
rect 24032 27548 24084 27557
rect 24492 27548 24544 27600
rect 25872 27616 25924 27668
rect 26792 27616 26844 27668
rect 27068 27616 27120 27668
rect 25320 27548 25372 27600
rect 27344 27591 27396 27600
rect 27344 27557 27353 27591
rect 27353 27557 27387 27591
rect 27387 27557 27396 27591
rect 27344 27548 27396 27557
rect 28908 27548 28960 27600
rect 23848 27480 23900 27532
rect 24676 27480 24728 27532
rect 27068 27480 27120 27532
rect 28080 27480 28132 27532
rect 28264 27480 28316 27532
rect 23664 27412 23716 27464
rect 24124 27412 24176 27464
rect 16856 27319 16908 27328
rect 16856 27285 16865 27319
rect 16865 27285 16899 27319
rect 16899 27285 16908 27319
rect 16856 27276 16908 27285
rect 19248 27319 19300 27328
rect 19248 27285 19257 27319
rect 19257 27285 19291 27319
rect 19291 27285 19300 27319
rect 19248 27276 19300 27285
rect 20904 27276 20956 27328
rect 21548 27319 21600 27328
rect 21548 27285 21557 27319
rect 21557 27285 21591 27319
rect 21591 27285 21600 27319
rect 21548 27276 21600 27285
rect 22284 27319 22336 27328
rect 22284 27285 22293 27319
rect 22293 27285 22327 27319
rect 22327 27285 22336 27319
rect 22284 27276 22336 27285
rect 22468 27276 22520 27328
rect 22744 27319 22796 27328
rect 22744 27285 22753 27319
rect 22753 27285 22787 27319
rect 22787 27285 22796 27319
rect 22744 27276 22796 27285
rect 23848 27319 23900 27328
rect 23848 27285 23857 27319
rect 23857 27285 23891 27319
rect 23891 27285 23900 27319
rect 23848 27276 23900 27285
rect 24860 27276 24912 27328
rect 25320 27276 25372 27328
rect 27804 27276 27856 27328
rect 4246 27174 4298 27226
rect 4310 27174 4362 27226
rect 4374 27174 4426 27226
rect 4438 27174 4490 27226
rect 34966 27174 35018 27226
rect 35030 27174 35082 27226
rect 35094 27174 35146 27226
rect 35158 27174 35210 27226
rect 6920 27072 6972 27124
rect 9588 27072 9640 27124
rect 14648 27115 14700 27124
rect 14648 27081 14657 27115
rect 14657 27081 14691 27115
rect 14691 27081 14700 27115
rect 14648 27072 14700 27081
rect 15660 27072 15712 27124
rect 1860 26979 1912 26988
rect 1860 26945 1869 26979
rect 1869 26945 1903 26979
rect 1903 26945 1912 26979
rect 1860 26936 1912 26945
rect 10416 26979 10468 26988
rect 10416 26945 10425 26979
rect 10425 26945 10459 26979
rect 10459 26945 10468 26979
rect 10416 26936 10468 26945
rect 10876 26979 10928 26988
rect 10876 26945 10885 26979
rect 10885 26945 10919 26979
rect 10919 26945 10928 26979
rect 10876 26936 10928 26945
rect 1676 26868 1728 26920
rect 4068 26800 4120 26852
rect 8668 26800 8720 26852
rect 9772 26800 9824 26852
rect 10140 26868 10192 26920
rect 10968 26911 11020 26920
rect 10968 26877 10977 26911
rect 10977 26877 11011 26911
rect 11011 26877 11020 26911
rect 10968 26868 11020 26877
rect 11704 27004 11756 27056
rect 12256 27047 12308 27056
rect 12256 27013 12265 27047
rect 12265 27013 12299 27047
rect 12299 27013 12308 27047
rect 12256 27004 12308 27013
rect 15108 27004 15160 27056
rect 15844 27072 15896 27124
rect 16212 27072 16264 27124
rect 16764 27072 16816 27124
rect 17408 27072 17460 27124
rect 18788 27115 18840 27124
rect 18788 27081 18797 27115
rect 18797 27081 18831 27115
rect 18831 27081 18840 27115
rect 18788 27072 18840 27081
rect 21088 27072 21140 27124
rect 17592 27004 17644 27056
rect 11888 26936 11940 26988
rect 14464 26936 14516 26988
rect 14924 26936 14976 26988
rect 16580 26979 16632 26988
rect 11244 26868 11296 26920
rect 10324 26800 10376 26852
rect 12808 26868 12860 26920
rect 13360 26868 13412 26920
rect 13728 26911 13780 26920
rect 13728 26877 13737 26911
rect 13737 26877 13771 26911
rect 13771 26877 13780 26911
rect 16580 26945 16589 26979
rect 16589 26945 16623 26979
rect 16623 26945 16632 26979
rect 16580 26936 16632 26945
rect 20260 26979 20312 26988
rect 20260 26945 20269 26979
rect 20269 26945 20303 26979
rect 20303 26945 20312 26979
rect 20260 26936 20312 26945
rect 23940 27047 23992 27056
rect 20628 26936 20680 26988
rect 20904 26936 20956 26988
rect 21088 26936 21140 26988
rect 13728 26868 13780 26877
rect 11612 26800 11664 26852
rect 15660 26911 15712 26920
rect 15660 26877 15669 26911
rect 15669 26877 15703 26911
rect 15703 26877 15712 26911
rect 15660 26868 15712 26877
rect 16396 26868 16448 26920
rect 16672 26911 16724 26920
rect 16672 26877 16681 26911
rect 16681 26877 16715 26911
rect 16715 26877 16724 26911
rect 16672 26868 16724 26877
rect 18788 26868 18840 26920
rect 19432 26911 19484 26920
rect 19432 26877 19441 26911
rect 19441 26877 19475 26911
rect 19475 26877 19484 26911
rect 19432 26868 19484 26877
rect 19984 26911 20036 26920
rect 7104 26775 7156 26784
rect 7104 26741 7113 26775
rect 7113 26741 7147 26775
rect 7147 26741 7156 26775
rect 7104 26732 7156 26741
rect 8484 26775 8536 26784
rect 8484 26741 8493 26775
rect 8493 26741 8527 26775
rect 8527 26741 8536 26775
rect 8484 26732 8536 26741
rect 9864 26775 9916 26784
rect 9864 26741 9873 26775
rect 9873 26741 9907 26775
rect 9907 26741 9916 26775
rect 9864 26732 9916 26741
rect 9956 26732 10008 26784
rect 10600 26732 10652 26784
rect 10968 26732 11020 26784
rect 13176 26732 13228 26784
rect 13820 26732 13872 26784
rect 14740 26732 14792 26784
rect 18880 26732 18932 26784
rect 19984 26877 19993 26911
rect 19993 26877 20027 26911
rect 20027 26877 20036 26911
rect 19984 26868 20036 26877
rect 20352 26868 20404 26920
rect 20628 26800 20680 26852
rect 20904 26800 20956 26852
rect 21456 26868 21508 26920
rect 22284 26843 22336 26852
rect 20812 26732 20864 26784
rect 21180 26732 21232 26784
rect 22284 26809 22293 26843
rect 22293 26809 22327 26843
rect 22327 26809 22336 26843
rect 22284 26800 22336 26809
rect 21732 26775 21784 26784
rect 21732 26741 21741 26775
rect 21741 26741 21775 26775
rect 21775 26741 21784 26775
rect 21732 26732 21784 26741
rect 22100 26732 22152 26784
rect 23388 26936 23440 26988
rect 23940 27013 23949 27047
rect 23949 27013 23983 27047
rect 23983 27013 23992 27047
rect 23940 27004 23992 27013
rect 25044 27072 25096 27124
rect 25872 27072 25924 27124
rect 26056 27115 26108 27124
rect 26056 27081 26065 27115
rect 26065 27081 26099 27115
rect 26099 27081 26108 27115
rect 26056 27072 26108 27081
rect 27068 27115 27120 27124
rect 27068 27081 27077 27115
rect 27077 27081 27111 27115
rect 27111 27081 27120 27115
rect 27068 27072 27120 27081
rect 28356 27072 28408 27124
rect 28724 27072 28776 27124
rect 25320 27004 25372 27056
rect 24308 26936 24360 26988
rect 23296 26868 23348 26920
rect 24676 26868 24728 26920
rect 25872 26868 25924 26920
rect 24032 26800 24084 26852
rect 26700 26868 26752 26920
rect 27068 26868 27120 26920
rect 28080 26911 28132 26920
rect 26792 26800 26844 26852
rect 28080 26877 28089 26911
rect 28089 26877 28123 26911
rect 28123 26877 28132 26911
rect 28080 26868 28132 26877
rect 23480 26732 23532 26784
rect 24308 26775 24360 26784
rect 24308 26741 24317 26775
rect 24317 26741 24351 26775
rect 24351 26741 24360 26775
rect 24308 26732 24360 26741
rect 24768 26775 24820 26784
rect 24768 26741 24777 26775
rect 24777 26741 24811 26775
rect 24811 26741 24820 26775
rect 24768 26732 24820 26741
rect 25872 26732 25924 26784
rect 26240 26732 26292 26784
rect 26700 26775 26752 26784
rect 26700 26741 26709 26775
rect 26709 26741 26743 26775
rect 26743 26741 26752 26775
rect 26700 26732 26752 26741
rect 27252 26732 27304 26784
rect 19606 26630 19658 26682
rect 19670 26630 19722 26682
rect 19734 26630 19786 26682
rect 19798 26630 19850 26682
rect 1860 26528 1912 26580
rect 7380 26528 7432 26580
rect 10140 26528 10192 26580
rect 11244 26528 11296 26580
rect 13452 26528 13504 26580
rect 14648 26571 14700 26580
rect 14648 26537 14657 26571
rect 14657 26537 14691 26571
rect 14691 26537 14700 26571
rect 14648 26528 14700 26537
rect 16120 26528 16172 26580
rect 16672 26528 16724 26580
rect 17224 26528 17276 26580
rect 18512 26528 18564 26580
rect 13268 26460 13320 26512
rect 1676 26392 1728 26444
rect 2044 26392 2096 26444
rect 2780 26392 2832 26444
rect 6000 26392 6052 26444
rect 6184 26392 6236 26444
rect 8668 26392 8720 26444
rect 9496 26435 9548 26444
rect 9496 26401 9505 26435
rect 9505 26401 9539 26435
rect 9539 26401 9548 26435
rect 9496 26392 9548 26401
rect 10876 26392 10928 26444
rect 12624 26392 12676 26444
rect 14740 26460 14792 26512
rect 15108 26503 15160 26512
rect 15108 26469 15117 26503
rect 15117 26469 15151 26503
rect 15151 26469 15160 26503
rect 15108 26460 15160 26469
rect 13820 26392 13872 26444
rect 14556 26392 14608 26444
rect 15016 26392 15068 26444
rect 15292 26392 15344 26444
rect 17316 26460 17368 26512
rect 18972 26460 19024 26512
rect 20444 26528 20496 26580
rect 21272 26528 21324 26580
rect 21732 26528 21784 26580
rect 21916 26528 21968 26580
rect 22560 26528 22612 26580
rect 23480 26528 23532 26580
rect 20812 26460 20864 26512
rect 21180 26460 21232 26512
rect 22008 26460 22060 26512
rect 22928 26460 22980 26512
rect 23940 26460 23992 26512
rect 16672 26435 16724 26444
rect 16672 26401 16681 26435
rect 16681 26401 16715 26435
rect 16715 26401 16724 26435
rect 16672 26392 16724 26401
rect 9680 26324 9732 26376
rect 10508 26367 10560 26376
rect 10508 26333 10517 26367
rect 10517 26333 10551 26367
rect 10551 26333 10560 26367
rect 10508 26324 10560 26333
rect 13360 26324 13412 26376
rect 10324 26299 10376 26308
rect 10324 26265 10333 26299
rect 10333 26265 10367 26299
rect 10367 26265 10376 26299
rect 10324 26256 10376 26265
rect 14004 26324 14056 26376
rect 16396 26324 16448 26376
rect 16856 26392 16908 26444
rect 17592 26435 17644 26444
rect 17592 26401 17601 26435
rect 17601 26401 17635 26435
rect 17635 26401 17644 26435
rect 17592 26392 17644 26401
rect 18512 26392 18564 26444
rect 17316 26324 17368 26376
rect 17776 26324 17828 26376
rect 18604 26324 18656 26376
rect 19248 26324 19300 26376
rect 19616 26367 19668 26376
rect 19616 26333 19625 26367
rect 19625 26333 19659 26367
rect 19659 26333 19668 26367
rect 19616 26324 19668 26333
rect 20352 26392 20404 26444
rect 21456 26392 21508 26444
rect 20628 26324 20680 26376
rect 21088 26367 21140 26376
rect 21088 26333 21094 26367
rect 21094 26333 21140 26367
rect 21088 26324 21140 26333
rect 14556 26256 14608 26308
rect 14740 26256 14792 26308
rect 15108 26256 15160 26308
rect 15844 26256 15896 26308
rect 17224 26256 17276 26308
rect 17868 26256 17920 26308
rect 8208 26188 8260 26240
rect 15568 26188 15620 26240
rect 16120 26231 16172 26240
rect 16120 26197 16129 26231
rect 16129 26197 16163 26231
rect 16163 26197 16172 26231
rect 16120 26188 16172 26197
rect 18236 26188 18288 26240
rect 20904 26256 20956 26308
rect 21180 26299 21232 26308
rect 19340 26188 19392 26240
rect 21180 26265 21189 26299
rect 21189 26265 21223 26299
rect 21223 26265 21232 26299
rect 21180 26256 21232 26265
rect 21916 26324 21968 26376
rect 22100 26392 22152 26444
rect 24216 26392 24268 26444
rect 24676 26460 24728 26512
rect 25136 26528 25188 26580
rect 26424 26528 26476 26580
rect 25688 26460 25740 26512
rect 24492 26392 24544 26444
rect 22836 26367 22888 26376
rect 22836 26333 22845 26367
rect 22845 26333 22879 26367
rect 22879 26333 22888 26367
rect 22836 26324 22888 26333
rect 23480 26324 23532 26376
rect 26976 26324 27028 26376
rect 28448 26528 28500 26580
rect 27528 26435 27580 26444
rect 27528 26401 27537 26435
rect 27537 26401 27571 26435
rect 27571 26401 27580 26435
rect 27528 26392 27580 26401
rect 27620 26324 27672 26376
rect 22100 26256 22152 26308
rect 22836 26188 22888 26240
rect 23296 26188 23348 26240
rect 24124 26256 24176 26308
rect 25044 26299 25096 26308
rect 25044 26265 25053 26299
rect 25053 26265 25087 26299
rect 25087 26265 25096 26299
rect 25044 26256 25096 26265
rect 25504 26299 25556 26308
rect 25504 26265 25513 26299
rect 25513 26265 25547 26299
rect 25547 26265 25556 26299
rect 25504 26256 25556 26265
rect 25872 26256 25924 26308
rect 26056 26188 26108 26240
rect 4246 26086 4298 26138
rect 4310 26086 4362 26138
rect 4374 26086 4426 26138
rect 4438 26086 4490 26138
rect 34966 26086 35018 26138
rect 35030 26086 35082 26138
rect 35094 26086 35146 26138
rect 35158 26086 35210 26138
rect 6000 25984 6052 26036
rect 8668 26027 8720 26036
rect 8668 25993 8677 26027
rect 8677 25993 8711 26027
rect 8711 25993 8720 26027
rect 8668 25984 8720 25993
rect 14004 25984 14056 26036
rect 15292 26027 15344 26036
rect 11520 25959 11572 25968
rect 11520 25925 11529 25959
rect 11529 25925 11563 25959
rect 11563 25925 11572 25959
rect 11520 25916 11572 25925
rect 12624 25916 12676 25968
rect 9220 25848 9272 25900
rect 9680 25780 9732 25832
rect 12624 25823 12676 25832
rect 12624 25789 12633 25823
rect 12633 25789 12667 25823
rect 12667 25789 12676 25823
rect 12624 25780 12676 25789
rect 14372 25916 14424 25968
rect 15292 25993 15301 26027
rect 15301 25993 15335 26027
rect 15335 25993 15344 26027
rect 15292 25984 15344 25993
rect 16672 26027 16724 26036
rect 16672 25993 16681 26027
rect 16681 25993 16715 26027
rect 16715 25993 16724 26027
rect 16672 25984 16724 25993
rect 17868 26027 17920 26036
rect 17868 25993 17877 26027
rect 17877 25993 17911 26027
rect 17911 25993 17920 26027
rect 17868 25984 17920 25993
rect 19064 25984 19116 26036
rect 21272 25984 21324 26036
rect 21456 26027 21508 26036
rect 21456 25993 21465 26027
rect 21465 25993 21499 26027
rect 21499 25993 21508 26027
rect 21456 25984 21508 25993
rect 22560 25984 22612 26036
rect 23480 25984 23532 26036
rect 25320 26027 25372 26036
rect 25320 25993 25329 26027
rect 25329 25993 25363 26027
rect 25363 25993 25372 26027
rect 25320 25984 25372 25993
rect 26976 25984 27028 26036
rect 27620 26027 27672 26036
rect 27620 25993 27629 26027
rect 27629 25993 27663 26027
rect 27663 25993 27672 26027
rect 27620 25984 27672 25993
rect 18512 25916 18564 25968
rect 19892 25916 19944 25968
rect 20628 25916 20680 25968
rect 21732 25916 21784 25968
rect 22928 25916 22980 25968
rect 14556 25848 14608 25900
rect 14648 25780 14700 25832
rect 6092 25687 6144 25696
rect 6092 25653 6101 25687
rect 6101 25653 6135 25687
rect 6135 25653 6144 25687
rect 6092 25644 6144 25653
rect 10600 25687 10652 25696
rect 10600 25653 10609 25687
rect 10609 25653 10643 25687
rect 10643 25653 10652 25687
rect 10600 25644 10652 25653
rect 11152 25687 11204 25696
rect 11152 25653 11161 25687
rect 11161 25653 11195 25687
rect 11195 25653 11204 25687
rect 11152 25644 11204 25653
rect 13728 25712 13780 25764
rect 14372 25712 14424 25764
rect 14556 25755 14608 25764
rect 14556 25721 14565 25755
rect 14565 25721 14599 25755
rect 14599 25721 14608 25755
rect 14556 25712 14608 25721
rect 15292 25848 15344 25900
rect 16120 25848 16172 25900
rect 15200 25780 15252 25832
rect 16212 25823 16264 25832
rect 16212 25789 16221 25823
rect 16221 25789 16255 25823
rect 16255 25789 16264 25823
rect 16212 25780 16264 25789
rect 16580 25780 16632 25832
rect 18236 25848 18288 25900
rect 19340 25848 19392 25900
rect 20076 25848 20128 25900
rect 21456 25848 21508 25900
rect 21640 25848 21692 25900
rect 23940 25848 23992 25900
rect 24952 25848 25004 25900
rect 18696 25823 18748 25832
rect 18696 25789 18705 25823
rect 18705 25789 18739 25823
rect 18739 25789 18748 25823
rect 18696 25780 18748 25789
rect 18788 25780 18840 25832
rect 19432 25780 19484 25832
rect 21364 25780 21416 25832
rect 21732 25780 21784 25832
rect 22468 25780 22520 25832
rect 24032 25780 24084 25832
rect 24860 25823 24912 25832
rect 24860 25789 24869 25823
rect 24869 25789 24903 25823
rect 24903 25789 24912 25823
rect 24860 25780 24912 25789
rect 20352 25712 20404 25764
rect 20812 25755 20864 25764
rect 20812 25721 20821 25755
rect 20821 25721 20855 25755
rect 20855 25721 20864 25755
rect 20812 25712 20864 25721
rect 26700 25891 26752 25900
rect 26700 25857 26709 25891
rect 26709 25857 26743 25891
rect 26743 25857 26752 25891
rect 26700 25848 26752 25857
rect 25872 25823 25924 25832
rect 25872 25789 25881 25823
rect 25881 25789 25915 25823
rect 25915 25789 25924 25823
rect 25872 25780 25924 25789
rect 26056 25823 26108 25832
rect 26056 25789 26065 25823
rect 26065 25789 26099 25823
rect 26099 25789 26108 25823
rect 26056 25780 26108 25789
rect 26424 25755 26476 25764
rect 13912 25644 13964 25696
rect 14740 25644 14792 25696
rect 17592 25644 17644 25696
rect 21640 25644 21692 25696
rect 22836 25687 22888 25696
rect 22836 25653 22845 25687
rect 22845 25653 22879 25687
rect 22879 25653 22888 25687
rect 22836 25644 22888 25653
rect 24124 25687 24176 25696
rect 24124 25653 24133 25687
rect 24133 25653 24167 25687
rect 24167 25653 24176 25687
rect 24124 25644 24176 25653
rect 26424 25721 26433 25755
rect 26433 25721 26467 25755
rect 26467 25721 26476 25755
rect 26424 25712 26476 25721
rect 27252 25644 27304 25696
rect 19606 25542 19658 25594
rect 19670 25542 19722 25594
rect 19734 25542 19786 25594
rect 19798 25542 19850 25594
rect 9220 25440 9272 25492
rect 9496 25483 9548 25492
rect 9496 25449 9505 25483
rect 9505 25449 9539 25483
rect 9539 25449 9548 25483
rect 9496 25440 9548 25449
rect 11336 25483 11388 25492
rect 11336 25449 11345 25483
rect 11345 25449 11379 25483
rect 11379 25449 11388 25483
rect 11336 25440 11388 25449
rect 12164 25483 12216 25492
rect 12164 25449 12173 25483
rect 12173 25449 12207 25483
rect 12207 25449 12216 25483
rect 12164 25440 12216 25449
rect 12348 25440 12400 25492
rect 13360 25440 13412 25492
rect 14740 25483 14792 25492
rect 14740 25449 14749 25483
rect 14749 25449 14783 25483
rect 14783 25449 14792 25483
rect 14740 25440 14792 25449
rect 15568 25483 15620 25492
rect 15568 25449 15577 25483
rect 15577 25449 15611 25483
rect 15611 25449 15620 25483
rect 15568 25440 15620 25449
rect 16488 25483 16540 25492
rect 16488 25449 16497 25483
rect 16497 25449 16531 25483
rect 16531 25449 16540 25483
rect 16488 25440 16540 25449
rect 16948 25440 17000 25492
rect 17684 25440 17736 25492
rect 20076 25483 20128 25492
rect 20076 25449 20085 25483
rect 20085 25449 20119 25483
rect 20119 25449 20128 25483
rect 20076 25440 20128 25449
rect 22744 25483 22796 25492
rect 22744 25449 22753 25483
rect 22753 25449 22787 25483
rect 22787 25449 22796 25483
rect 22744 25440 22796 25449
rect 25320 25483 25372 25492
rect 25320 25449 25329 25483
rect 25329 25449 25363 25483
rect 25363 25449 25372 25483
rect 25320 25440 25372 25449
rect 27344 25440 27396 25492
rect 10600 25372 10652 25424
rect 10232 25304 10284 25356
rect 18512 25372 18564 25424
rect 19432 25372 19484 25424
rect 19616 25372 19668 25424
rect 10784 25347 10836 25356
rect 10784 25313 10793 25347
rect 10793 25313 10827 25347
rect 10827 25313 10836 25347
rect 10784 25304 10836 25313
rect 11060 25304 11112 25356
rect 11888 25304 11940 25356
rect 14096 25304 14148 25356
rect 9680 25279 9732 25288
rect 9680 25245 9689 25279
rect 9689 25245 9723 25279
rect 9723 25245 9732 25279
rect 9680 25236 9732 25245
rect 13912 25236 13964 25288
rect 14464 25304 14516 25356
rect 15384 25347 15436 25356
rect 15384 25313 15393 25347
rect 15393 25313 15427 25347
rect 15427 25313 15436 25347
rect 15384 25304 15436 25313
rect 16672 25304 16724 25356
rect 16948 25347 17000 25356
rect 16948 25313 16957 25347
rect 16957 25313 16991 25347
rect 16991 25313 17000 25347
rect 16948 25304 17000 25313
rect 17040 25347 17092 25356
rect 17040 25313 17049 25347
rect 17049 25313 17083 25347
rect 17083 25313 17092 25347
rect 17224 25347 17276 25356
rect 17040 25304 17092 25313
rect 17224 25313 17233 25347
rect 17233 25313 17267 25347
rect 17267 25313 17276 25347
rect 17224 25304 17276 25313
rect 17500 25347 17552 25356
rect 17500 25313 17509 25347
rect 17509 25313 17543 25347
rect 17543 25313 17552 25347
rect 17500 25304 17552 25313
rect 17868 25347 17920 25356
rect 17868 25313 17877 25347
rect 17877 25313 17911 25347
rect 17911 25313 17920 25347
rect 17868 25304 17920 25313
rect 19248 25304 19300 25356
rect 19340 25304 19392 25356
rect 22836 25372 22888 25424
rect 26792 25372 26844 25424
rect 21088 25304 21140 25356
rect 21272 25304 21324 25356
rect 14372 25236 14424 25288
rect 22560 25304 22612 25356
rect 23756 25304 23808 25356
rect 23940 25304 23992 25356
rect 24032 25304 24084 25356
rect 25596 25304 25648 25356
rect 26608 25304 26660 25356
rect 22192 25236 22244 25288
rect 24768 25236 24820 25288
rect 26056 25279 26108 25288
rect 26056 25245 26065 25279
rect 26065 25245 26099 25279
rect 26099 25245 26108 25279
rect 26056 25236 26108 25245
rect 12348 25168 12400 25220
rect 13728 25168 13780 25220
rect 15568 25168 15620 25220
rect 17868 25168 17920 25220
rect 18052 25168 18104 25220
rect 19524 25211 19576 25220
rect 19524 25177 19533 25211
rect 19533 25177 19567 25211
rect 19567 25177 19576 25211
rect 19524 25168 19576 25177
rect 15108 25143 15160 25152
rect 15108 25109 15117 25143
rect 15117 25109 15151 25143
rect 15151 25109 15160 25143
rect 15108 25100 15160 25109
rect 15936 25143 15988 25152
rect 15936 25109 15945 25143
rect 15945 25109 15979 25143
rect 15979 25109 15988 25143
rect 15936 25100 15988 25109
rect 16488 25100 16540 25152
rect 18788 25100 18840 25152
rect 20444 25143 20496 25152
rect 20444 25109 20453 25143
rect 20453 25109 20487 25143
rect 20487 25109 20496 25143
rect 20444 25100 20496 25109
rect 21456 25143 21508 25152
rect 21456 25109 21465 25143
rect 21465 25109 21499 25143
rect 21499 25109 21508 25143
rect 21456 25100 21508 25109
rect 24860 25100 24912 25152
rect 4246 24998 4298 25050
rect 4310 24998 4362 25050
rect 4374 24998 4426 25050
rect 4438 24998 4490 25050
rect 34966 24998 35018 25050
rect 35030 24998 35082 25050
rect 35094 24998 35146 25050
rect 35158 24998 35210 25050
rect 11888 24939 11940 24948
rect 11888 24905 11897 24939
rect 11897 24905 11931 24939
rect 11931 24905 11940 24939
rect 11888 24896 11940 24905
rect 14188 24896 14240 24948
rect 15384 24939 15436 24948
rect 15384 24905 15393 24939
rect 15393 24905 15427 24939
rect 15427 24905 15436 24939
rect 15384 24896 15436 24905
rect 19616 24939 19668 24948
rect 19616 24905 19625 24939
rect 19625 24905 19659 24939
rect 19659 24905 19668 24939
rect 19616 24896 19668 24905
rect 20076 24896 20128 24948
rect 21180 24896 21232 24948
rect 23480 24939 23532 24948
rect 23480 24905 23489 24939
rect 23489 24905 23523 24939
rect 23523 24905 23532 24939
rect 23480 24896 23532 24905
rect 26608 24939 26660 24948
rect 26608 24905 26617 24939
rect 26617 24905 26651 24939
rect 26651 24905 26660 24939
rect 26608 24896 26660 24905
rect 10600 24828 10652 24880
rect 14096 24871 14148 24880
rect 2688 24760 2740 24812
rect 10048 24760 10100 24812
rect 14096 24837 14105 24871
rect 14105 24837 14139 24871
rect 14139 24837 14148 24871
rect 14096 24828 14148 24837
rect 15108 24828 15160 24880
rect 16948 24828 17000 24880
rect 17500 24828 17552 24880
rect 12440 24760 12492 24812
rect 14464 24803 14516 24812
rect 12624 24692 12676 24744
rect 13084 24692 13136 24744
rect 14464 24769 14473 24803
rect 14473 24769 14507 24803
rect 14507 24769 14516 24803
rect 14464 24760 14516 24769
rect 14924 24760 14976 24812
rect 16212 24760 16264 24812
rect 20076 24760 20128 24812
rect 21456 24828 21508 24880
rect 20444 24803 20496 24812
rect 20444 24769 20453 24803
rect 20453 24769 20487 24803
rect 20487 24769 20496 24803
rect 20444 24760 20496 24769
rect 13728 24735 13780 24744
rect 13728 24701 13737 24735
rect 13737 24701 13771 24735
rect 13771 24701 13780 24735
rect 13728 24692 13780 24701
rect 8668 24599 8720 24608
rect 8668 24565 8677 24599
rect 8677 24565 8711 24599
rect 8711 24565 8720 24599
rect 8668 24556 8720 24565
rect 10968 24556 11020 24608
rect 13820 24624 13872 24676
rect 15200 24692 15252 24744
rect 15476 24692 15528 24744
rect 16488 24692 16540 24744
rect 16764 24692 16816 24744
rect 17316 24692 17368 24744
rect 18696 24735 18748 24744
rect 18696 24701 18705 24735
rect 18705 24701 18739 24735
rect 18739 24701 18748 24735
rect 18696 24692 18748 24701
rect 19064 24735 19116 24744
rect 19064 24701 19073 24735
rect 19073 24701 19107 24735
rect 19107 24701 19116 24735
rect 19064 24692 19116 24701
rect 18052 24624 18104 24676
rect 19248 24692 19300 24744
rect 19984 24692 20036 24744
rect 22284 24760 22336 24812
rect 24676 24760 24728 24812
rect 24952 24803 25004 24812
rect 24952 24769 24961 24803
rect 24961 24769 24995 24803
rect 24995 24769 25004 24803
rect 24952 24760 25004 24769
rect 25780 24760 25832 24812
rect 20812 24735 20864 24744
rect 20812 24701 20821 24735
rect 20821 24701 20855 24735
rect 20855 24701 20864 24735
rect 20812 24692 20864 24701
rect 21088 24735 21140 24744
rect 21088 24701 21097 24735
rect 21097 24701 21131 24735
rect 21131 24701 21140 24735
rect 21088 24692 21140 24701
rect 21456 24692 21508 24744
rect 19800 24624 19852 24676
rect 21548 24624 21600 24676
rect 23756 24735 23808 24744
rect 23756 24701 23765 24735
rect 23765 24701 23799 24735
rect 23799 24701 23808 24735
rect 25044 24735 25096 24744
rect 23756 24692 23808 24701
rect 25044 24701 25053 24735
rect 25053 24701 25087 24735
rect 25087 24701 25096 24735
rect 25044 24692 25096 24701
rect 11980 24556 12032 24608
rect 12624 24556 12676 24608
rect 12808 24599 12860 24608
rect 12808 24565 12817 24599
rect 12817 24565 12851 24599
rect 12851 24565 12860 24599
rect 12808 24556 12860 24565
rect 14924 24556 14976 24608
rect 16396 24556 16448 24608
rect 17500 24599 17552 24608
rect 17500 24565 17509 24599
rect 17509 24565 17543 24599
rect 17543 24565 17552 24599
rect 17500 24556 17552 24565
rect 17776 24599 17828 24608
rect 17776 24565 17785 24599
rect 17785 24565 17819 24599
rect 17819 24565 17828 24599
rect 17776 24556 17828 24565
rect 19064 24556 19116 24608
rect 19984 24556 20036 24608
rect 20812 24556 20864 24608
rect 22008 24624 22060 24676
rect 24216 24667 24268 24676
rect 24216 24633 24225 24667
rect 24225 24633 24259 24667
rect 24259 24633 24268 24667
rect 24216 24624 24268 24633
rect 25228 24599 25280 24608
rect 25228 24565 25237 24599
rect 25237 24565 25271 24599
rect 25271 24565 25280 24599
rect 25228 24556 25280 24565
rect 19606 24454 19658 24506
rect 19670 24454 19722 24506
rect 19734 24454 19786 24506
rect 19798 24454 19850 24506
rect 7932 24395 7984 24404
rect 7932 24361 7941 24395
rect 7941 24361 7975 24395
rect 7975 24361 7984 24395
rect 7932 24352 7984 24361
rect 9220 24352 9272 24404
rect 10048 24352 10100 24404
rect 10232 24395 10284 24404
rect 10232 24361 10241 24395
rect 10241 24361 10275 24395
rect 10275 24361 10284 24395
rect 10232 24352 10284 24361
rect 10508 24352 10560 24404
rect 10968 24395 11020 24404
rect 10968 24361 10977 24395
rect 10977 24361 11011 24395
rect 11011 24361 11020 24395
rect 10968 24352 11020 24361
rect 11980 24395 12032 24404
rect 11980 24361 11989 24395
rect 11989 24361 12023 24395
rect 12023 24361 12032 24395
rect 11980 24352 12032 24361
rect 13912 24352 13964 24404
rect 14740 24395 14792 24404
rect 14740 24361 14749 24395
rect 14749 24361 14783 24395
rect 14783 24361 14792 24395
rect 14740 24352 14792 24361
rect 16948 24352 17000 24404
rect 17960 24352 18012 24404
rect 19340 24352 19392 24404
rect 19984 24352 20036 24404
rect 20628 24395 20680 24404
rect 20628 24361 20637 24395
rect 20637 24361 20671 24395
rect 20671 24361 20680 24395
rect 20628 24352 20680 24361
rect 13636 24327 13688 24336
rect 13636 24293 13645 24327
rect 13645 24293 13679 24327
rect 13679 24293 13688 24327
rect 13636 24284 13688 24293
rect 15292 24284 15344 24336
rect 17500 24284 17552 24336
rect 18788 24284 18840 24336
rect 8116 24259 8168 24268
rect 8116 24225 8125 24259
rect 8125 24225 8159 24259
rect 8159 24225 8168 24259
rect 8116 24216 8168 24225
rect 10876 24216 10928 24268
rect 12532 24216 12584 24268
rect 12808 24259 12860 24268
rect 12808 24225 12817 24259
rect 12817 24225 12851 24259
rect 12851 24225 12860 24259
rect 12808 24216 12860 24225
rect 12900 24216 12952 24268
rect 13912 24259 13964 24268
rect 13912 24225 13921 24259
rect 13921 24225 13955 24259
rect 13955 24225 13964 24259
rect 13912 24216 13964 24225
rect 15200 24216 15252 24268
rect 16396 24216 16448 24268
rect 16672 24216 16724 24268
rect 17592 24259 17644 24268
rect 17592 24225 17601 24259
rect 17601 24225 17635 24259
rect 17635 24225 17644 24259
rect 17592 24216 17644 24225
rect 17868 24216 17920 24268
rect 18972 24284 19024 24336
rect 21456 24352 21508 24404
rect 21548 24352 21600 24404
rect 22468 24352 22520 24404
rect 23112 24352 23164 24404
rect 23756 24395 23808 24404
rect 23756 24361 23765 24395
rect 23765 24361 23799 24395
rect 23799 24361 23808 24395
rect 23756 24352 23808 24361
rect 24676 24352 24728 24404
rect 24860 24352 24912 24404
rect 22008 24284 22060 24336
rect 25044 24284 25096 24336
rect 19984 24216 20036 24268
rect 20720 24216 20772 24268
rect 7656 24148 7708 24200
rect 8484 24148 8536 24200
rect 8760 24148 8812 24200
rect 9588 24148 9640 24200
rect 11152 24148 11204 24200
rect 14556 24148 14608 24200
rect 14832 24148 14884 24200
rect 15844 24191 15896 24200
rect 15844 24157 15853 24191
rect 15853 24157 15887 24191
rect 15887 24157 15896 24191
rect 15844 24148 15896 24157
rect 20904 24191 20956 24200
rect 10784 24080 10836 24132
rect 13728 24080 13780 24132
rect 16580 24080 16632 24132
rect 19340 24080 19392 24132
rect 20904 24157 20913 24191
rect 20913 24157 20947 24191
rect 20947 24157 20956 24191
rect 20904 24148 20956 24157
rect 21548 24216 21600 24268
rect 22192 24216 22244 24268
rect 22468 24259 22520 24268
rect 22468 24225 22477 24259
rect 22477 24225 22511 24259
rect 22511 24225 22520 24259
rect 22468 24216 22520 24225
rect 22560 24216 22612 24268
rect 23388 24216 23440 24268
rect 23480 24216 23532 24268
rect 24216 24216 24268 24268
rect 25228 24259 25280 24268
rect 25228 24225 25237 24259
rect 25237 24225 25271 24259
rect 25271 24225 25280 24259
rect 25228 24216 25280 24225
rect 21916 24148 21968 24200
rect 23572 24148 23624 24200
rect 23940 24080 23992 24132
rect 25596 24080 25648 24132
rect 11336 24055 11388 24064
rect 11336 24021 11345 24055
rect 11345 24021 11379 24055
rect 11379 24021 11388 24055
rect 11336 24012 11388 24021
rect 12992 24055 13044 24064
rect 12992 24021 13001 24055
rect 13001 24021 13035 24055
rect 13035 24021 13044 24055
rect 12992 24012 13044 24021
rect 14372 24012 14424 24064
rect 15108 24055 15160 24064
rect 15108 24021 15117 24055
rect 15117 24021 15151 24055
rect 15151 24021 15160 24055
rect 15108 24012 15160 24021
rect 17960 24055 18012 24064
rect 17960 24021 17969 24055
rect 17969 24021 18003 24055
rect 18003 24021 18012 24055
rect 17960 24012 18012 24021
rect 22468 24012 22520 24064
rect 25412 24055 25464 24064
rect 25412 24021 25421 24055
rect 25421 24021 25455 24055
rect 25455 24021 25464 24055
rect 25412 24012 25464 24021
rect 4246 23910 4298 23962
rect 4310 23910 4362 23962
rect 4374 23910 4426 23962
rect 4438 23910 4490 23962
rect 34966 23910 35018 23962
rect 35030 23910 35082 23962
rect 35094 23910 35146 23962
rect 35158 23910 35210 23962
rect 7012 23808 7064 23860
rect 8116 23808 8168 23860
rect 10876 23808 10928 23860
rect 12440 23808 12492 23860
rect 13820 23851 13872 23860
rect 12348 23740 12400 23792
rect 13820 23817 13829 23851
rect 13829 23817 13863 23851
rect 13863 23817 13872 23851
rect 13820 23808 13872 23817
rect 13912 23808 13964 23860
rect 15108 23808 15160 23860
rect 16764 23851 16816 23860
rect 16764 23817 16773 23851
rect 16773 23817 16807 23851
rect 16807 23817 16816 23851
rect 16764 23808 16816 23817
rect 17868 23851 17920 23860
rect 17868 23817 17877 23851
rect 17877 23817 17911 23851
rect 17911 23817 17920 23851
rect 17868 23808 17920 23817
rect 18328 23808 18380 23860
rect 21548 23808 21600 23860
rect 22560 23851 22612 23860
rect 22560 23817 22569 23851
rect 22569 23817 22603 23851
rect 22603 23817 22612 23851
rect 22560 23808 22612 23817
rect 23296 23808 23348 23860
rect 23848 23851 23900 23860
rect 23848 23817 23857 23851
rect 23857 23817 23891 23851
rect 23891 23817 23900 23851
rect 23848 23808 23900 23817
rect 24216 23851 24268 23860
rect 24216 23817 24225 23851
rect 24225 23817 24259 23851
rect 24259 23817 24268 23851
rect 24216 23808 24268 23817
rect 26240 23808 26292 23860
rect 14188 23740 14240 23792
rect 16672 23740 16724 23792
rect 17592 23740 17644 23792
rect 19524 23740 19576 23792
rect 21640 23740 21692 23792
rect 2044 23715 2096 23724
rect 2044 23681 2053 23715
rect 2053 23681 2087 23715
rect 2087 23681 2096 23715
rect 2044 23672 2096 23681
rect 9680 23672 9732 23724
rect 11336 23672 11388 23724
rect 13636 23672 13688 23724
rect 16212 23672 16264 23724
rect 17960 23672 18012 23724
rect 20720 23715 20772 23724
rect 1768 23468 1820 23520
rect 8668 23536 8720 23588
rect 12532 23604 12584 23656
rect 12808 23604 12860 23656
rect 14924 23647 14976 23656
rect 14924 23613 14933 23647
rect 14933 23613 14967 23647
rect 14967 23613 14976 23647
rect 14924 23604 14976 23613
rect 15568 23647 15620 23656
rect 15568 23613 15577 23647
rect 15577 23613 15611 23647
rect 15611 23613 15620 23647
rect 15568 23604 15620 23613
rect 9864 23536 9916 23588
rect 15108 23536 15160 23588
rect 20720 23681 20729 23715
rect 20729 23681 20763 23715
rect 20763 23681 20772 23715
rect 20720 23672 20772 23681
rect 16580 23647 16632 23656
rect 16580 23613 16589 23647
rect 16589 23613 16623 23647
rect 16623 23613 16632 23647
rect 18512 23647 18564 23656
rect 16580 23604 16632 23613
rect 18512 23613 18521 23647
rect 18521 23613 18555 23647
rect 18555 23613 18564 23647
rect 18512 23604 18564 23613
rect 19156 23647 19208 23656
rect 19156 23613 19165 23647
rect 19165 23613 19199 23647
rect 19199 23613 19208 23647
rect 19156 23604 19208 23613
rect 19432 23647 19484 23656
rect 19432 23613 19441 23647
rect 19441 23613 19475 23647
rect 19475 23613 19484 23647
rect 19432 23604 19484 23613
rect 20904 23604 20956 23656
rect 21456 23672 21508 23724
rect 21548 23647 21600 23656
rect 21548 23613 21557 23647
rect 21557 23613 21591 23647
rect 21591 23613 21600 23647
rect 21548 23604 21600 23613
rect 23664 23647 23716 23656
rect 18880 23536 18932 23588
rect 20996 23536 21048 23588
rect 23664 23613 23673 23647
rect 23673 23613 23707 23647
rect 23707 23613 23716 23647
rect 23664 23604 23716 23613
rect 23940 23604 23992 23656
rect 25044 23647 25096 23656
rect 25044 23613 25053 23647
rect 25053 23613 25087 23647
rect 25087 23613 25096 23647
rect 25044 23604 25096 23613
rect 21916 23536 21968 23588
rect 9680 23511 9732 23520
rect 9680 23477 9689 23511
rect 9689 23477 9723 23511
rect 9723 23477 9732 23511
rect 9680 23468 9732 23477
rect 11152 23511 11204 23520
rect 11152 23477 11161 23511
rect 11161 23477 11195 23511
rect 11195 23477 11204 23511
rect 11152 23468 11204 23477
rect 15660 23468 15712 23520
rect 16212 23468 16264 23520
rect 16396 23511 16448 23520
rect 16396 23477 16405 23511
rect 16405 23477 16439 23511
rect 16439 23477 16448 23511
rect 16396 23468 16448 23477
rect 19248 23468 19300 23520
rect 21548 23468 21600 23520
rect 22192 23468 22244 23520
rect 19606 23366 19658 23418
rect 19670 23366 19722 23418
rect 19734 23366 19786 23418
rect 19798 23366 19850 23418
rect 2044 23307 2096 23316
rect 2044 23273 2053 23307
rect 2053 23273 2087 23307
rect 2087 23273 2096 23307
rect 2044 23264 2096 23273
rect 11152 23264 11204 23316
rect 12808 23307 12860 23316
rect 12808 23273 12817 23307
rect 12817 23273 12851 23307
rect 12851 23273 12860 23307
rect 12808 23264 12860 23273
rect 14096 23264 14148 23316
rect 16304 23264 16356 23316
rect 16580 23307 16632 23316
rect 16580 23273 16589 23307
rect 16589 23273 16623 23307
rect 16623 23273 16632 23307
rect 16580 23264 16632 23273
rect 18512 23264 18564 23316
rect 10968 23128 11020 23180
rect 11612 23171 11664 23180
rect 11612 23137 11621 23171
rect 11621 23137 11655 23171
rect 11655 23137 11664 23171
rect 11612 23128 11664 23137
rect 13360 23128 13412 23180
rect 14832 23196 14884 23248
rect 14004 23128 14056 23180
rect 15568 23128 15620 23180
rect 18788 23239 18840 23248
rect 18788 23205 18797 23239
rect 18797 23205 18831 23239
rect 18831 23205 18840 23239
rect 18788 23196 18840 23205
rect 20812 23196 20864 23248
rect 21548 23196 21600 23248
rect 21732 23264 21784 23316
rect 25596 23307 25648 23316
rect 25596 23273 25605 23307
rect 25605 23273 25639 23307
rect 25639 23273 25648 23307
rect 25596 23264 25648 23273
rect 17224 23171 17276 23180
rect 17224 23137 17233 23171
rect 17233 23137 17267 23171
rect 17267 23137 17276 23171
rect 17224 23128 17276 23137
rect 17500 23128 17552 23180
rect 19432 23171 19484 23180
rect 19432 23137 19441 23171
rect 19441 23137 19475 23171
rect 19475 23137 19484 23171
rect 19432 23128 19484 23137
rect 19800 23171 19852 23180
rect 19800 23137 19809 23171
rect 19809 23137 19843 23171
rect 19843 23137 19852 23171
rect 19800 23128 19852 23137
rect 19892 23171 19944 23180
rect 19892 23137 19901 23171
rect 19901 23137 19935 23171
rect 19935 23137 19944 23171
rect 19892 23128 19944 23137
rect 20628 23128 20680 23180
rect 10600 23103 10652 23112
rect 10600 23069 10609 23103
rect 10609 23069 10643 23103
rect 10643 23069 10652 23103
rect 10600 23060 10652 23069
rect 13268 23103 13320 23112
rect 10784 22992 10836 23044
rect 13268 23069 13277 23103
rect 13277 23069 13311 23103
rect 13311 23069 13320 23103
rect 13268 23060 13320 23069
rect 13912 23103 13964 23112
rect 13912 23069 13921 23103
rect 13921 23069 13955 23103
rect 13955 23069 13964 23103
rect 13912 23060 13964 23069
rect 12624 22992 12676 23044
rect 13176 22992 13228 23044
rect 13728 22992 13780 23044
rect 15292 23060 15344 23112
rect 17868 23060 17920 23112
rect 19340 23103 19392 23112
rect 19340 23069 19349 23103
rect 19349 23069 19383 23103
rect 19383 23069 19392 23103
rect 19340 23060 19392 23069
rect 19984 23060 20036 23112
rect 15200 22992 15252 23044
rect 17040 23035 17092 23044
rect 17040 23001 17049 23035
rect 17049 23001 17083 23035
rect 17083 23001 17092 23035
rect 17040 22992 17092 23001
rect 1400 22924 1452 22976
rect 12532 22967 12584 22976
rect 12532 22933 12541 22967
rect 12541 22933 12575 22967
rect 12575 22933 12584 22967
rect 12532 22924 12584 22933
rect 14648 22967 14700 22976
rect 14648 22933 14657 22967
rect 14657 22933 14691 22967
rect 14691 22933 14700 22967
rect 14648 22924 14700 22933
rect 15476 22924 15528 22976
rect 18604 22967 18656 22976
rect 18604 22933 18613 22967
rect 18613 22933 18647 22967
rect 18647 22933 18656 22967
rect 18604 22924 18656 22933
rect 20904 22924 20956 22976
rect 21364 23128 21416 23180
rect 21916 23128 21968 23180
rect 22744 23128 22796 23180
rect 23388 23128 23440 23180
rect 22928 23060 22980 23112
rect 23572 23128 23624 23180
rect 24676 23171 24728 23180
rect 24676 23137 24685 23171
rect 24685 23137 24719 23171
rect 24719 23137 24728 23171
rect 24676 23128 24728 23137
rect 23848 23060 23900 23112
rect 22836 22992 22888 23044
rect 24492 23035 24544 23044
rect 24492 23001 24501 23035
rect 24501 23001 24535 23035
rect 24535 23001 24544 23035
rect 24492 22992 24544 23001
rect 21180 22924 21232 22976
rect 22192 22924 22244 22976
rect 25228 22967 25280 22976
rect 25228 22933 25237 22967
rect 25237 22933 25271 22967
rect 25271 22933 25280 22967
rect 25228 22924 25280 22933
rect 4246 22822 4298 22874
rect 4310 22822 4362 22874
rect 4374 22822 4426 22874
rect 4438 22822 4490 22874
rect 34966 22822 35018 22874
rect 35030 22822 35082 22874
rect 35094 22822 35146 22874
rect 35158 22822 35210 22874
rect 3148 22763 3200 22772
rect 3148 22729 3157 22763
rect 3157 22729 3191 22763
rect 3191 22729 3200 22763
rect 3148 22720 3200 22729
rect 11152 22720 11204 22772
rect 11796 22763 11848 22772
rect 11796 22729 11805 22763
rect 11805 22729 11839 22763
rect 11839 22729 11848 22763
rect 11796 22720 11848 22729
rect 12624 22763 12676 22772
rect 12624 22729 12633 22763
rect 12633 22729 12667 22763
rect 12667 22729 12676 22763
rect 12624 22720 12676 22729
rect 13360 22720 13412 22772
rect 15568 22763 15620 22772
rect 15568 22729 15577 22763
rect 15577 22729 15611 22763
rect 15611 22729 15620 22763
rect 15568 22720 15620 22729
rect 15752 22720 15804 22772
rect 10784 22652 10836 22704
rect 10968 22695 11020 22704
rect 10968 22661 10977 22695
rect 10977 22661 11011 22695
rect 11011 22661 11020 22695
rect 10968 22652 11020 22661
rect 11244 22652 11296 22704
rect 11612 22652 11664 22704
rect 15476 22652 15528 22704
rect 14004 22584 14056 22636
rect 17592 22720 17644 22772
rect 19800 22720 19852 22772
rect 20812 22720 20864 22772
rect 21364 22720 21416 22772
rect 22744 22763 22796 22772
rect 22744 22729 22753 22763
rect 22753 22729 22787 22763
rect 22787 22729 22796 22763
rect 22744 22720 22796 22729
rect 23848 22763 23900 22772
rect 23848 22729 23857 22763
rect 23857 22729 23891 22763
rect 23891 22729 23900 22763
rect 23848 22720 23900 22729
rect 24676 22720 24728 22772
rect 16120 22652 16172 22704
rect 16396 22652 16448 22704
rect 18420 22652 18472 22704
rect 19984 22652 20036 22704
rect 22008 22652 22060 22704
rect 23112 22652 23164 22704
rect 1400 22516 1452 22568
rect 1860 22559 1912 22568
rect 1860 22525 1869 22559
rect 1869 22525 1903 22559
rect 1903 22525 1912 22559
rect 1860 22516 1912 22525
rect 11796 22516 11848 22568
rect 12440 22559 12492 22568
rect 12440 22525 12449 22559
rect 12449 22525 12483 22559
rect 12483 22525 12492 22559
rect 13636 22559 13688 22568
rect 12440 22516 12492 22525
rect 13636 22525 13645 22559
rect 13645 22525 13679 22559
rect 13679 22525 13688 22559
rect 13636 22516 13688 22525
rect 13912 22559 13964 22568
rect 13912 22525 13921 22559
rect 13921 22525 13955 22559
rect 13955 22525 13964 22559
rect 13912 22516 13964 22525
rect 16304 22516 16356 22568
rect 18880 22627 18932 22636
rect 17868 22516 17920 22568
rect 18604 22516 18656 22568
rect 17684 22448 17736 22500
rect 18052 22448 18104 22500
rect 18328 22491 18380 22500
rect 18328 22457 18337 22491
rect 18337 22457 18371 22491
rect 18371 22457 18380 22491
rect 18328 22448 18380 22457
rect 18512 22491 18564 22500
rect 18512 22457 18521 22491
rect 18521 22457 18555 22491
rect 18555 22457 18564 22491
rect 18512 22448 18564 22457
rect 18880 22593 18889 22627
rect 18889 22593 18923 22627
rect 18923 22593 18932 22627
rect 18880 22584 18932 22593
rect 19064 22516 19116 22568
rect 20444 22627 20496 22636
rect 20444 22593 20453 22627
rect 20453 22593 20487 22627
rect 20487 22593 20496 22627
rect 20444 22584 20496 22593
rect 20904 22584 20956 22636
rect 25228 22584 25280 22636
rect 19156 22448 19208 22500
rect 20628 22516 20680 22568
rect 21732 22559 21784 22568
rect 21732 22525 21741 22559
rect 21741 22525 21775 22559
rect 21775 22525 21784 22559
rect 21732 22516 21784 22525
rect 23112 22559 23164 22568
rect 23112 22525 23121 22559
rect 23121 22525 23155 22559
rect 23155 22525 23164 22559
rect 23112 22516 23164 22525
rect 14372 22380 14424 22432
rect 16672 22380 16724 22432
rect 19984 22423 20036 22432
rect 19984 22389 19993 22423
rect 19993 22389 20027 22423
rect 20027 22389 20036 22423
rect 19984 22380 20036 22389
rect 19606 22278 19658 22330
rect 19670 22278 19722 22330
rect 19734 22278 19786 22330
rect 19798 22278 19850 22330
rect 11336 22176 11388 22228
rect 11888 22176 11940 22228
rect 13728 22176 13780 22228
rect 14832 22176 14884 22228
rect 17040 22176 17092 22228
rect 17684 22176 17736 22228
rect 18052 22176 18104 22228
rect 19248 22176 19300 22228
rect 20628 22176 20680 22228
rect 21732 22219 21784 22228
rect 21732 22185 21741 22219
rect 21741 22185 21775 22219
rect 21775 22185 21784 22219
rect 21732 22176 21784 22185
rect 5448 22108 5500 22160
rect 9864 22108 9916 22160
rect 10140 22040 10192 22092
rect 11336 22040 11388 22092
rect 13084 22040 13136 22092
rect 14004 22108 14056 22160
rect 15200 22108 15252 22160
rect 16856 22108 16908 22160
rect 17224 22108 17276 22160
rect 17316 22108 17368 22160
rect 14188 22083 14240 22092
rect 14188 22049 14197 22083
rect 14197 22049 14231 22083
rect 14231 22049 14240 22083
rect 14188 22040 14240 22049
rect 14740 22083 14792 22092
rect 14740 22049 14749 22083
rect 14749 22049 14783 22083
rect 14783 22049 14792 22083
rect 14740 22040 14792 22049
rect 16028 22083 16080 22092
rect 16028 22049 16037 22083
rect 16037 22049 16071 22083
rect 16071 22049 16080 22083
rect 16028 22040 16080 22049
rect 16304 22040 16356 22092
rect 17500 22083 17552 22092
rect 17500 22049 17509 22083
rect 17509 22049 17543 22083
rect 17543 22049 17552 22083
rect 17500 22040 17552 22049
rect 17868 22040 17920 22092
rect 19432 22108 19484 22160
rect 20444 22108 20496 22160
rect 21548 22108 21600 22160
rect 18880 22083 18932 22092
rect 18880 22049 18889 22083
rect 18889 22049 18923 22083
rect 18923 22049 18932 22083
rect 20996 22083 21048 22092
rect 18880 22040 18932 22049
rect 20996 22049 21005 22083
rect 21005 22049 21039 22083
rect 21039 22049 21048 22083
rect 20996 22040 21048 22049
rect 11612 22015 11664 22024
rect 11612 21981 11621 22015
rect 11621 21981 11655 22015
rect 11655 21981 11664 22015
rect 11612 21972 11664 21981
rect 12348 22015 12400 22024
rect 12348 21981 12357 22015
rect 12357 21981 12391 22015
rect 12391 21981 12400 22015
rect 12348 21972 12400 21981
rect 12532 22015 12584 22024
rect 12532 21981 12541 22015
rect 12541 21981 12575 22015
rect 12575 21981 12584 22015
rect 12532 21972 12584 21981
rect 15936 22015 15988 22024
rect 15936 21981 15945 22015
rect 15945 21981 15979 22015
rect 15979 21981 15988 22015
rect 15936 21972 15988 21981
rect 18052 21972 18104 22024
rect 18236 21972 18288 22024
rect 18788 22015 18840 22024
rect 18788 21981 18797 22015
rect 18797 21981 18831 22015
rect 18831 21981 18840 22015
rect 18788 21972 18840 21981
rect 21916 21972 21968 22024
rect 23112 22015 23164 22024
rect 23112 21981 23121 22015
rect 23121 21981 23155 22015
rect 23155 21981 23164 22015
rect 23112 21972 23164 21981
rect 23388 22015 23440 22024
rect 23388 21981 23397 22015
rect 23397 21981 23431 22015
rect 23431 21981 23440 22015
rect 23388 21972 23440 21981
rect 17960 21904 18012 21956
rect 1860 21836 1912 21888
rect 13912 21836 13964 21888
rect 15108 21836 15160 21888
rect 15568 21879 15620 21888
rect 15568 21845 15577 21879
rect 15577 21845 15611 21879
rect 15611 21845 15620 21879
rect 15568 21836 15620 21845
rect 17592 21836 17644 21888
rect 18696 21836 18748 21888
rect 20444 21879 20496 21888
rect 20444 21845 20453 21879
rect 20453 21845 20487 21879
rect 20487 21845 20496 21879
rect 20444 21836 20496 21845
rect 21088 21836 21140 21888
rect 22468 21879 22520 21888
rect 22468 21845 22477 21879
rect 22477 21845 22511 21879
rect 22511 21845 22520 21879
rect 22468 21836 22520 21845
rect 24492 21879 24544 21888
rect 24492 21845 24501 21879
rect 24501 21845 24535 21879
rect 24535 21845 24544 21879
rect 24492 21836 24544 21845
rect 4246 21734 4298 21786
rect 4310 21734 4362 21786
rect 4374 21734 4426 21786
rect 4438 21734 4490 21786
rect 34966 21734 35018 21786
rect 35030 21734 35082 21786
rect 35094 21734 35146 21786
rect 35158 21734 35210 21786
rect 11336 21675 11388 21684
rect 11336 21641 11345 21675
rect 11345 21641 11379 21675
rect 11379 21641 11388 21675
rect 11336 21632 11388 21641
rect 12256 21632 12308 21684
rect 13636 21675 13688 21684
rect 13636 21641 13645 21675
rect 13645 21641 13679 21675
rect 13679 21641 13688 21675
rect 13636 21632 13688 21641
rect 14188 21675 14240 21684
rect 14188 21641 14197 21675
rect 14197 21641 14231 21675
rect 14231 21641 14240 21675
rect 14188 21632 14240 21641
rect 15384 21632 15436 21684
rect 15752 21675 15804 21684
rect 15752 21641 15761 21675
rect 15761 21641 15795 21675
rect 15795 21641 15804 21675
rect 15752 21632 15804 21641
rect 16028 21632 16080 21684
rect 16304 21632 16356 21684
rect 17500 21675 17552 21684
rect 17500 21641 17509 21675
rect 17509 21641 17543 21675
rect 17543 21641 17552 21675
rect 17500 21632 17552 21641
rect 18880 21632 18932 21684
rect 20996 21632 21048 21684
rect 21916 21632 21968 21684
rect 23388 21632 23440 21684
rect 26424 21675 26476 21684
rect 26424 21641 26433 21675
rect 26433 21641 26467 21675
rect 26467 21641 26476 21675
rect 26424 21632 26476 21641
rect 11244 21564 11296 21616
rect 12532 21564 12584 21616
rect 12808 21564 12860 21616
rect 19892 21564 19944 21616
rect 14556 21496 14608 21548
rect 16396 21496 16448 21548
rect 17776 21496 17828 21548
rect 17960 21496 18012 21548
rect 19616 21539 19668 21548
rect 19616 21505 19625 21539
rect 19625 21505 19659 21539
rect 19659 21505 19668 21539
rect 19616 21496 19668 21505
rect 16672 21471 16724 21480
rect 16672 21437 16681 21471
rect 16681 21437 16715 21471
rect 16715 21437 16724 21471
rect 16672 21428 16724 21437
rect 18788 21471 18840 21480
rect 18788 21437 18797 21471
rect 18797 21437 18831 21471
rect 18831 21437 18840 21471
rect 18788 21428 18840 21437
rect 21272 21496 21324 21548
rect 20352 21471 20404 21480
rect 10968 21403 11020 21412
rect 10968 21369 10977 21403
rect 10977 21369 11011 21403
rect 11011 21369 11020 21403
rect 10968 21360 11020 21369
rect 19432 21292 19484 21344
rect 20352 21437 20361 21471
rect 20361 21437 20395 21471
rect 20395 21437 20404 21471
rect 20352 21428 20404 21437
rect 20444 21471 20496 21480
rect 20444 21437 20453 21471
rect 20453 21437 20487 21471
rect 20487 21437 20496 21471
rect 20444 21428 20496 21437
rect 22652 21360 22704 21412
rect 23112 21360 23164 21412
rect 25228 21428 25280 21480
rect 24952 21360 25004 21412
rect 22192 21335 22244 21344
rect 22192 21301 22201 21335
rect 22201 21301 22235 21335
rect 22235 21301 22244 21335
rect 22192 21292 22244 21301
rect 24676 21335 24728 21344
rect 24676 21301 24685 21335
rect 24685 21301 24719 21335
rect 24719 21301 24728 21335
rect 24676 21292 24728 21301
rect 25228 21292 25280 21344
rect 19606 21190 19658 21242
rect 19670 21190 19722 21242
rect 19734 21190 19786 21242
rect 19798 21190 19850 21242
rect 13084 21131 13136 21140
rect 13084 21097 13093 21131
rect 13093 21097 13127 21131
rect 13127 21097 13136 21131
rect 13084 21088 13136 21097
rect 16396 21131 16448 21140
rect 16396 21097 16405 21131
rect 16405 21097 16439 21131
rect 16439 21097 16448 21131
rect 16396 21088 16448 21097
rect 16856 21131 16908 21140
rect 16856 21097 16865 21131
rect 16865 21097 16899 21131
rect 16899 21097 16908 21131
rect 16856 21088 16908 21097
rect 18052 21131 18104 21140
rect 18052 21097 18061 21131
rect 18061 21097 18095 21131
rect 18095 21097 18104 21131
rect 18052 21088 18104 21097
rect 18604 21088 18656 21140
rect 19984 21088 20036 21140
rect 20628 21088 20680 21140
rect 21088 21131 21140 21140
rect 21088 21097 21097 21131
rect 21097 21097 21131 21131
rect 21131 21097 21140 21131
rect 21088 21088 21140 21097
rect 21364 21131 21416 21140
rect 21364 21097 21373 21131
rect 21373 21097 21407 21131
rect 21407 21097 21416 21131
rect 21364 21088 21416 21097
rect 12072 20952 12124 21004
rect 13636 20952 13688 21004
rect 17684 20995 17736 21004
rect 17684 20961 17693 20995
rect 17693 20961 17727 20995
rect 17727 20961 17736 20995
rect 17684 20952 17736 20961
rect 19064 21020 19116 21072
rect 19156 21020 19208 21072
rect 20444 21020 20496 21072
rect 11980 20927 12032 20936
rect 11980 20893 11989 20927
rect 11989 20893 12023 20927
rect 12023 20893 12032 20927
rect 11980 20884 12032 20893
rect 18328 20884 18380 20936
rect 19708 20952 19760 21004
rect 20352 20952 20404 21004
rect 21180 20952 21232 21004
rect 21364 20952 21416 21004
rect 20536 20884 20588 20936
rect 19340 20816 19392 20868
rect 20812 20816 20864 20868
rect 1860 20748 1912 20800
rect 2688 20748 2740 20800
rect 17960 20748 18012 20800
rect 19708 20748 19760 20800
rect 24952 20791 25004 20800
rect 24952 20757 24961 20791
rect 24961 20757 24995 20791
rect 24995 20757 25004 20791
rect 24952 20748 25004 20757
rect 4246 20646 4298 20698
rect 4310 20646 4362 20698
rect 4374 20646 4426 20698
rect 4438 20646 4490 20698
rect 34966 20646 35018 20698
rect 35030 20646 35082 20698
rect 35094 20646 35146 20698
rect 35158 20646 35210 20698
rect 12072 20587 12124 20596
rect 12072 20553 12081 20587
rect 12081 20553 12115 20587
rect 12115 20553 12124 20587
rect 12072 20544 12124 20553
rect 12256 20544 12308 20596
rect 13728 20544 13780 20596
rect 15568 20587 15620 20596
rect 15568 20553 15577 20587
rect 15577 20553 15611 20587
rect 15611 20553 15620 20587
rect 15568 20544 15620 20553
rect 17684 20544 17736 20596
rect 17868 20587 17920 20596
rect 17868 20553 17877 20587
rect 17877 20553 17911 20587
rect 17911 20553 17920 20587
rect 17868 20544 17920 20553
rect 19064 20587 19116 20596
rect 19064 20553 19073 20587
rect 19073 20553 19107 20587
rect 19107 20553 19116 20587
rect 19064 20544 19116 20553
rect 19340 20544 19392 20596
rect 13912 20519 13964 20528
rect 13912 20485 13921 20519
rect 13921 20485 13955 20519
rect 13955 20485 13964 20519
rect 13912 20476 13964 20485
rect 20720 20476 20772 20528
rect 11980 20340 12032 20392
rect 15660 20408 15712 20460
rect 16028 20408 16080 20460
rect 16120 20408 16172 20460
rect 17592 20408 17644 20460
rect 19432 20408 19484 20460
rect 20536 20408 20588 20460
rect 16948 20383 17000 20392
rect 16948 20349 16957 20383
rect 16957 20349 16991 20383
rect 16991 20349 17000 20383
rect 16948 20340 17000 20349
rect 17316 20340 17368 20392
rect 19984 20247 20036 20256
rect 19984 20213 19993 20247
rect 19993 20213 20027 20247
rect 20027 20213 20036 20247
rect 20260 20340 20312 20392
rect 20720 20340 20772 20392
rect 19984 20204 20036 20213
rect 19606 20102 19658 20154
rect 19670 20102 19722 20154
rect 19734 20102 19786 20154
rect 19798 20102 19850 20154
rect 12072 20000 12124 20052
rect 12440 20043 12492 20052
rect 12440 20009 12449 20043
rect 12449 20009 12483 20043
rect 12483 20009 12492 20043
rect 12440 20000 12492 20009
rect 14740 20000 14792 20052
rect 15476 20000 15528 20052
rect 19156 20043 19208 20052
rect 19156 20009 19165 20043
rect 19165 20009 19199 20043
rect 19199 20009 19208 20043
rect 19156 20000 19208 20009
rect 19432 20043 19484 20052
rect 19432 20009 19441 20043
rect 19441 20009 19475 20043
rect 19475 20009 19484 20043
rect 19432 20000 19484 20009
rect 20260 20043 20312 20052
rect 20260 20009 20269 20043
rect 20269 20009 20303 20043
rect 20303 20009 20312 20043
rect 20260 20000 20312 20009
rect 20536 20043 20588 20052
rect 20536 20009 20545 20043
rect 20545 20009 20579 20043
rect 20579 20009 20588 20043
rect 20536 20000 20588 20009
rect 21364 20043 21416 20052
rect 21364 20009 21373 20043
rect 21373 20009 21407 20043
rect 21407 20009 21416 20043
rect 21364 20000 21416 20009
rect 7840 19932 7892 19984
rect 17684 19932 17736 19984
rect 19984 19932 20036 19984
rect 5448 19864 5500 19916
rect 13636 19864 13688 19916
rect 16028 19907 16080 19916
rect 16028 19873 16037 19907
rect 16037 19873 16071 19907
rect 16071 19873 16080 19907
rect 16028 19864 16080 19873
rect 16304 19864 16356 19916
rect 17960 19864 18012 19916
rect 18144 19907 18196 19916
rect 18144 19873 18153 19907
rect 18153 19873 18187 19907
rect 18187 19873 18196 19907
rect 18144 19864 18196 19873
rect 18328 19907 18380 19916
rect 18328 19873 18337 19907
rect 18337 19873 18371 19907
rect 18371 19873 18380 19907
rect 18328 19864 18380 19873
rect 20996 19864 21048 19916
rect 22008 19864 22060 19916
rect 4712 19839 4764 19848
rect 4712 19805 4721 19839
rect 4721 19805 4755 19839
rect 4755 19805 4764 19839
rect 4712 19796 4764 19805
rect 4896 19796 4948 19848
rect 16212 19796 16264 19848
rect 17776 19796 17828 19848
rect 21088 19771 21140 19780
rect 21088 19737 21097 19771
rect 21097 19737 21131 19771
rect 21131 19737 21140 19771
rect 21088 19728 21140 19737
rect 14924 19703 14976 19712
rect 14924 19669 14933 19703
rect 14933 19669 14967 19703
rect 14967 19669 14976 19703
rect 14924 19660 14976 19669
rect 15936 19660 15988 19712
rect 16764 19660 16816 19712
rect 17316 19660 17368 19712
rect 4246 19558 4298 19610
rect 4310 19558 4362 19610
rect 4374 19558 4426 19610
rect 4438 19558 4490 19610
rect 34966 19558 35018 19610
rect 35030 19558 35082 19610
rect 35094 19558 35146 19610
rect 35158 19558 35210 19610
rect 16028 19499 16080 19508
rect 16028 19465 16037 19499
rect 16037 19465 16071 19499
rect 16071 19465 16080 19499
rect 16028 19456 16080 19465
rect 20076 19499 20128 19508
rect 20076 19465 20085 19499
rect 20085 19465 20119 19499
rect 20119 19465 20128 19499
rect 20076 19456 20128 19465
rect 20996 19499 21048 19508
rect 20996 19465 21005 19499
rect 21005 19465 21039 19499
rect 21039 19465 21048 19499
rect 20996 19456 21048 19465
rect 31484 19499 31536 19508
rect 31484 19465 31493 19499
rect 31493 19465 31527 19499
rect 31527 19465 31536 19499
rect 31484 19456 31536 19465
rect 12440 19363 12492 19372
rect 12440 19329 12449 19363
rect 12449 19329 12483 19363
rect 12483 19329 12492 19363
rect 12440 19320 12492 19329
rect 13636 19320 13688 19372
rect 14188 19320 14240 19372
rect 14924 19363 14976 19372
rect 14924 19329 14933 19363
rect 14933 19329 14967 19363
rect 14967 19329 14976 19363
rect 14924 19320 14976 19329
rect 14280 19252 14332 19304
rect 16580 19295 16632 19304
rect 14464 19227 14516 19236
rect 14464 19193 14473 19227
rect 14473 19193 14507 19227
rect 14507 19193 14516 19227
rect 14464 19184 14516 19193
rect 16580 19261 16589 19295
rect 16589 19261 16623 19295
rect 16623 19261 16632 19295
rect 16580 19252 16632 19261
rect 18144 19252 18196 19304
rect 18788 19295 18840 19304
rect 18788 19261 18797 19295
rect 18797 19261 18831 19295
rect 18831 19261 18840 19295
rect 18788 19252 18840 19261
rect 18972 19252 19024 19304
rect 19156 19295 19208 19304
rect 19156 19261 19165 19295
rect 19165 19261 19199 19295
rect 19199 19261 19208 19295
rect 19156 19252 19208 19261
rect 19432 19252 19484 19304
rect 30104 19295 30156 19304
rect 15476 19227 15528 19236
rect 15476 19193 15485 19227
rect 15485 19193 15519 19227
rect 15519 19193 15528 19227
rect 15476 19184 15528 19193
rect 18420 19184 18472 19236
rect 30104 19261 30113 19295
rect 30113 19261 30147 19295
rect 30147 19261 30156 19295
rect 30104 19252 30156 19261
rect 31668 19252 31720 19304
rect 4436 19159 4488 19168
rect 4436 19125 4445 19159
rect 4445 19125 4479 19159
rect 4479 19125 4488 19159
rect 4436 19116 4488 19125
rect 4712 19116 4764 19168
rect 4896 19159 4948 19168
rect 4896 19125 4905 19159
rect 4905 19125 4939 19159
rect 4939 19125 4948 19159
rect 4896 19116 4948 19125
rect 13820 19159 13872 19168
rect 13820 19125 13829 19159
rect 13829 19125 13863 19159
rect 13863 19125 13872 19159
rect 13820 19116 13872 19125
rect 16672 19116 16724 19168
rect 17684 19116 17736 19168
rect 17960 19116 18012 19168
rect 18972 19116 19024 19168
rect 19606 19014 19658 19066
rect 19670 19014 19722 19066
rect 19734 19014 19786 19066
rect 19798 19014 19850 19066
rect 12348 18844 12400 18896
rect 11336 18776 11388 18828
rect 12532 18819 12584 18828
rect 12532 18785 12541 18819
rect 12541 18785 12575 18819
rect 12575 18785 12584 18819
rect 12532 18776 12584 18785
rect 13912 18844 13964 18896
rect 15476 18912 15528 18964
rect 16580 18912 16632 18964
rect 17776 18955 17828 18964
rect 17776 18921 17785 18955
rect 17785 18921 17819 18955
rect 17819 18921 17828 18955
rect 17776 18912 17828 18921
rect 17960 18912 18012 18964
rect 19156 18912 19208 18964
rect 23848 18955 23900 18964
rect 23848 18921 23857 18955
rect 23857 18921 23891 18955
rect 23891 18921 23900 18955
rect 23848 18912 23900 18921
rect 15752 18844 15804 18896
rect 20260 18844 20312 18896
rect 13820 18776 13872 18828
rect 11888 18751 11940 18760
rect 11888 18717 11897 18751
rect 11897 18717 11931 18751
rect 11931 18717 11940 18751
rect 11888 18708 11940 18717
rect 12808 18751 12860 18760
rect 12072 18640 12124 18692
rect 12808 18717 12817 18751
rect 12817 18717 12851 18751
rect 12851 18717 12860 18751
rect 12808 18708 12860 18717
rect 13452 18751 13504 18760
rect 13452 18717 13461 18751
rect 13461 18717 13495 18751
rect 13495 18717 13504 18751
rect 14464 18776 14516 18828
rect 15936 18819 15988 18828
rect 15936 18785 15945 18819
rect 15945 18785 15979 18819
rect 15979 18785 15988 18819
rect 15936 18776 15988 18785
rect 16304 18819 16356 18828
rect 16304 18785 16313 18819
rect 16313 18785 16347 18819
rect 16347 18785 16356 18819
rect 16304 18776 16356 18785
rect 17316 18819 17368 18828
rect 17316 18785 17325 18819
rect 17325 18785 17359 18819
rect 17359 18785 17368 18819
rect 17316 18776 17368 18785
rect 18420 18776 18472 18828
rect 18788 18776 18840 18828
rect 19340 18776 19392 18828
rect 20444 18776 20496 18828
rect 22744 18819 22796 18828
rect 22744 18785 22753 18819
rect 22753 18785 22787 18819
rect 22787 18785 22796 18819
rect 22744 18776 22796 18785
rect 16396 18751 16448 18760
rect 13452 18708 13504 18717
rect 16396 18717 16405 18751
rect 16405 18717 16439 18751
rect 16439 18717 16448 18751
rect 16396 18708 16448 18717
rect 22468 18751 22520 18760
rect 22468 18717 22477 18751
rect 22477 18717 22511 18751
rect 22511 18717 22520 18751
rect 22468 18708 22520 18717
rect 14740 18640 14792 18692
rect 15752 18683 15804 18692
rect 15752 18649 15761 18683
rect 15761 18649 15795 18683
rect 15795 18649 15804 18683
rect 15752 18640 15804 18649
rect 12440 18572 12492 18624
rect 13360 18572 13412 18624
rect 17500 18615 17552 18624
rect 17500 18581 17509 18615
rect 17509 18581 17543 18615
rect 17543 18581 17552 18615
rect 17500 18572 17552 18581
rect 30104 18615 30156 18624
rect 30104 18581 30113 18615
rect 30113 18581 30147 18615
rect 30147 18581 30156 18615
rect 30104 18572 30156 18581
rect 4246 18470 4298 18522
rect 4310 18470 4362 18522
rect 4374 18470 4426 18522
rect 4438 18470 4490 18522
rect 34966 18470 35018 18522
rect 35030 18470 35082 18522
rect 35094 18470 35146 18522
rect 35158 18470 35210 18522
rect 12072 18368 12124 18420
rect 14464 18411 14516 18420
rect 14464 18377 14473 18411
rect 14473 18377 14507 18411
rect 14507 18377 14516 18411
rect 14464 18368 14516 18377
rect 14740 18411 14792 18420
rect 14740 18377 14749 18411
rect 14749 18377 14783 18411
rect 14783 18377 14792 18411
rect 14740 18368 14792 18377
rect 9864 18275 9916 18284
rect 9864 18241 9873 18275
rect 9873 18241 9907 18275
rect 9907 18241 9916 18275
rect 9864 18232 9916 18241
rect 12440 18275 12492 18284
rect 12440 18241 12449 18275
rect 12449 18241 12483 18275
rect 12483 18241 12492 18275
rect 12440 18232 12492 18241
rect 13452 18232 13504 18284
rect 9680 18071 9732 18080
rect 9680 18037 9689 18071
rect 9689 18037 9723 18071
rect 9723 18037 9732 18071
rect 12164 18164 12216 18216
rect 13820 18071 13872 18080
rect 9680 18028 9732 18037
rect 13820 18037 13829 18071
rect 13829 18037 13863 18071
rect 13863 18037 13872 18071
rect 13820 18028 13872 18037
rect 15476 18164 15528 18216
rect 15568 18207 15620 18216
rect 15568 18173 15577 18207
rect 15577 18173 15611 18207
rect 15611 18173 15620 18207
rect 15936 18368 15988 18420
rect 17316 18411 17368 18420
rect 17316 18377 17325 18411
rect 17325 18377 17359 18411
rect 17359 18377 17368 18411
rect 17316 18368 17368 18377
rect 18144 18368 18196 18420
rect 18972 18411 19024 18420
rect 16304 18343 16356 18352
rect 16304 18309 16313 18343
rect 16313 18309 16347 18343
rect 16347 18309 16356 18343
rect 16304 18300 16356 18309
rect 15568 18164 15620 18173
rect 18972 18377 18981 18411
rect 18981 18377 19015 18411
rect 19015 18377 19024 18411
rect 18972 18368 19024 18377
rect 22744 18368 22796 18420
rect 14924 18139 14976 18148
rect 14924 18105 14933 18139
rect 14933 18105 14967 18139
rect 14967 18105 14976 18139
rect 14924 18096 14976 18105
rect 16396 18096 16448 18148
rect 17040 18096 17092 18148
rect 17960 18096 18012 18148
rect 18788 18028 18840 18080
rect 22100 18028 22152 18080
rect 22468 18028 22520 18080
rect 19606 17926 19658 17978
rect 19670 17926 19722 17978
rect 19734 17926 19786 17978
rect 19798 17926 19850 17978
rect 9864 17867 9916 17876
rect 9864 17833 9873 17867
rect 9873 17833 9907 17867
rect 9907 17833 9916 17867
rect 9864 17824 9916 17833
rect 12348 17824 12400 17876
rect 14832 17824 14884 17876
rect 18420 17824 18472 17876
rect 19248 17824 19300 17876
rect 12808 17756 12860 17808
rect 17868 17756 17920 17808
rect 12624 17731 12676 17740
rect 12624 17697 12633 17731
rect 12633 17697 12667 17731
rect 12667 17697 12676 17731
rect 12624 17688 12676 17697
rect 11980 17663 12032 17672
rect 11980 17629 11989 17663
rect 11989 17629 12023 17663
rect 12023 17629 12032 17663
rect 11980 17620 12032 17629
rect 12992 17731 13044 17740
rect 12992 17697 13001 17731
rect 13001 17697 13035 17731
rect 13035 17697 13044 17731
rect 12992 17688 13044 17697
rect 13728 17688 13780 17740
rect 15384 17731 15436 17740
rect 15384 17697 15393 17731
rect 15393 17697 15427 17731
rect 15427 17697 15436 17731
rect 15384 17688 15436 17697
rect 17040 17731 17092 17740
rect 17040 17697 17049 17731
rect 17049 17697 17083 17731
rect 17083 17697 17092 17731
rect 17040 17688 17092 17697
rect 17500 17688 17552 17740
rect 17960 17688 18012 17740
rect 19156 17688 19208 17740
rect 20076 17688 20128 17740
rect 15292 17663 15344 17672
rect 12164 17552 12216 17604
rect 15292 17629 15301 17663
rect 15301 17629 15335 17663
rect 15335 17629 15344 17663
rect 15292 17620 15344 17629
rect 16948 17663 17000 17672
rect 16948 17629 16957 17663
rect 16957 17629 16991 17663
rect 16991 17629 17000 17663
rect 16948 17620 17000 17629
rect 13728 17552 13780 17604
rect 18604 17552 18656 17604
rect 9864 17484 9916 17536
rect 12900 17484 12952 17536
rect 15568 17527 15620 17536
rect 15568 17493 15577 17527
rect 15577 17493 15611 17527
rect 15611 17493 15620 17527
rect 15568 17484 15620 17493
rect 16488 17484 16540 17536
rect 18420 17484 18472 17536
rect 4246 17382 4298 17434
rect 4310 17382 4362 17434
rect 4374 17382 4426 17434
rect 4438 17382 4490 17434
rect 34966 17382 35018 17434
rect 35030 17382 35082 17434
rect 35094 17382 35146 17434
rect 35158 17382 35210 17434
rect 8392 17323 8444 17332
rect 8392 17289 8401 17323
rect 8401 17289 8435 17323
rect 8435 17289 8444 17323
rect 8392 17280 8444 17289
rect 12624 17280 12676 17332
rect 12808 17280 12860 17332
rect 15292 17280 15344 17332
rect 17500 17280 17552 17332
rect 18604 17323 18656 17332
rect 18604 17289 18613 17323
rect 18613 17289 18647 17323
rect 18647 17289 18656 17323
rect 18604 17280 18656 17289
rect 19156 17323 19208 17332
rect 19156 17289 19165 17323
rect 19165 17289 19199 17323
rect 19199 17289 19208 17323
rect 19156 17280 19208 17289
rect 12164 17212 12216 17264
rect 17868 17212 17920 17264
rect 12900 17187 12952 17196
rect 12900 17153 12909 17187
rect 12909 17153 12943 17187
rect 12943 17153 12952 17187
rect 12900 17144 12952 17153
rect 13544 17144 13596 17196
rect 15384 17144 15436 17196
rect 15844 17076 15896 17128
rect 16948 17144 17000 17196
rect 16396 17119 16448 17128
rect 16396 17085 16405 17119
rect 16405 17085 16439 17119
rect 16439 17085 16448 17119
rect 16396 17076 16448 17085
rect 16488 17119 16540 17128
rect 16488 17085 16497 17119
rect 16497 17085 16531 17119
rect 16531 17085 16540 17119
rect 16488 17076 16540 17085
rect 17500 17076 17552 17128
rect 17316 17008 17368 17060
rect 9496 16940 9548 16992
rect 19606 16838 19658 16890
rect 19670 16838 19722 16890
rect 19734 16838 19786 16890
rect 19798 16838 19850 16890
rect 1400 16736 1452 16788
rect 12992 16736 13044 16788
rect 15844 16779 15896 16788
rect 15844 16745 15853 16779
rect 15853 16745 15887 16779
rect 15887 16745 15896 16779
rect 15844 16736 15896 16745
rect 15568 16668 15620 16720
rect 25320 16711 25372 16720
rect 25320 16677 25329 16711
rect 25329 16677 25363 16711
rect 25363 16677 25372 16711
rect 25320 16668 25372 16677
rect 13544 16600 13596 16652
rect 13820 16643 13872 16652
rect 13820 16609 13829 16643
rect 13829 16609 13863 16643
rect 13863 16609 13872 16643
rect 13820 16600 13872 16609
rect 14096 16532 14148 16584
rect 13636 16507 13688 16516
rect 13636 16473 13645 16507
rect 13645 16473 13679 16507
rect 13679 16473 13688 16507
rect 13636 16464 13688 16473
rect 13728 16464 13780 16516
rect 15016 16600 15068 16652
rect 17500 16643 17552 16652
rect 17500 16609 17509 16643
rect 17509 16609 17543 16643
rect 17543 16609 17552 16643
rect 17500 16600 17552 16609
rect 17684 16643 17736 16652
rect 17684 16609 17693 16643
rect 17693 16609 17727 16643
rect 17727 16609 17736 16643
rect 17684 16600 17736 16609
rect 18328 16600 18380 16652
rect 24308 16600 24360 16652
rect 16396 16532 16448 16584
rect 16764 16575 16816 16584
rect 16764 16541 16773 16575
rect 16773 16541 16807 16575
rect 16807 16541 16816 16575
rect 16764 16532 16816 16541
rect 23848 16532 23900 16584
rect 17960 16439 18012 16448
rect 17960 16405 17969 16439
rect 17969 16405 18003 16439
rect 18003 16405 18012 16439
rect 17960 16396 18012 16405
rect 4246 16294 4298 16346
rect 4310 16294 4362 16346
rect 4374 16294 4426 16346
rect 4438 16294 4490 16346
rect 34966 16294 35018 16346
rect 35030 16294 35082 16346
rect 35094 16294 35146 16346
rect 35158 16294 35210 16346
rect 3240 16192 3292 16244
rect 13820 16235 13872 16244
rect 13820 16201 13829 16235
rect 13829 16201 13863 16235
rect 13863 16201 13872 16235
rect 13820 16192 13872 16201
rect 14096 16235 14148 16244
rect 14096 16201 14105 16235
rect 14105 16201 14139 16235
rect 14139 16201 14148 16235
rect 14096 16192 14148 16201
rect 17500 16235 17552 16244
rect 17500 16201 17509 16235
rect 17509 16201 17543 16235
rect 17543 16201 17552 16235
rect 17500 16192 17552 16201
rect 9496 16124 9548 16176
rect 10968 16124 11020 16176
rect 13728 16124 13780 16176
rect 17684 16124 17736 16176
rect 1400 16099 1452 16108
rect 1400 16065 1409 16099
rect 1409 16065 1443 16099
rect 1443 16065 1452 16099
rect 1400 16056 1452 16065
rect 1584 16056 1636 16108
rect 10232 16031 10284 16040
rect 10232 15997 10241 16031
rect 10241 15997 10275 16031
rect 10275 15997 10284 16031
rect 10232 15988 10284 15997
rect 15660 16031 15712 16040
rect 15660 15997 15669 16031
rect 15669 15997 15703 16031
rect 15703 15997 15712 16031
rect 15660 15988 15712 15997
rect 14832 15920 14884 15972
rect 16396 15963 16448 15972
rect 16396 15929 16405 15963
rect 16405 15929 16439 15963
rect 16439 15929 16448 15963
rect 16396 15920 16448 15929
rect 15384 15895 15436 15904
rect 15384 15861 15393 15895
rect 15393 15861 15427 15895
rect 15427 15861 15436 15895
rect 15384 15852 15436 15861
rect 23848 15895 23900 15904
rect 23848 15861 23857 15895
rect 23857 15861 23891 15895
rect 23891 15861 23900 15895
rect 23848 15852 23900 15861
rect 24308 15895 24360 15904
rect 24308 15861 24317 15895
rect 24317 15861 24351 15895
rect 24351 15861 24360 15895
rect 24308 15852 24360 15861
rect 24768 15852 24820 15904
rect 19606 15750 19658 15802
rect 19670 15750 19722 15802
rect 19734 15750 19786 15802
rect 19798 15750 19850 15802
rect 17960 15648 18012 15700
rect 18052 15623 18104 15632
rect 18052 15589 18061 15623
rect 18061 15589 18095 15623
rect 18095 15589 18104 15623
rect 18052 15580 18104 15589
rect 21180 15555 21232 15564
rect 21180 15521 21189 15555
rect 21189 15521 21223 15555
rect 21223 15521 21232 15555
rect 21180 15512 21232 15521
rect 21272 15444 21324 15496
rect 22008 15444 22060 15496
rect 1584 15351 1636 15360
rect 1584 15317 1593 15351
rect 1593 15317 1627 15351
rect 1627 15317 1636 15351
rect 1584 15308 1636 15317
rect 15844 15308 15896 15360
rect 22468 15351 22520 15360
rect 22468 15317 22477 15351
rect 22477 15317 22511 15351
rect 22511 15317 22520 15351
rect 22468 15308 22520 15317
rect 4246 15206 4298 15258
rect 4310 15206 4362 15258
rect 4374 15206 4426 15258
rect 4438 15206 4490 15258
rect 34966 15206 35018 15258
rect 35030 15206 35082 15258
rect 35094 15206 35146 15258
rect 35158 15206 35210 15258
rect 15200 15104 15252 15156
rect 16856 15104 16908 15156
rect 18328 15147 18380 15156
rect 18328 15113 18337 15147
rect 18337 15113 18371 15147
rect 18371 15113 18380 15147
rect 18328 15104 18380 15113
rect 21180 15104 21232 15156
rect 16028 15036 16080 15088
rect 13360 14968 13412 15020
rect 13820 15011 13872 15020
rect 13820 14977 13829 15011
rect 13829 14977 13863 15011
rect 13863 14977 13872 15011
rect 13820 14968 13872 14977
rect 15292 14968 15344 15020
rect 18604 15036 18656 15088
rect 17960 14968 18012 15020
rect 15200 14875 15252 14884
rect 15200 14841 15209 14875
rect 15209 14841 15243 14875
rect 15243 14841 15252 14875
rect 15200 14832 15252 14841
rect 15844 14900 15896 14952
rect 16856 14943 16908 14952
rect 16856 14909 16865 14943
rect 16865 14909 16899 14943
rect 16899 14909 16908 14943
rect 16856 14900 16908 14909
rect 18052 14900 18104 14952
rect 18972 14832 19024 14884
rect 21272 14807 21324 14816
rect 21272 14773 21281 14807
rect 21281 14773 21315 14807
rect 21315 14773 21324 14807
rect 21272 14764 21324 14773
rect 19606 14662 19658 14714
rect 19670 14662 19722 14714
rect 19734 14662 19786 14714
rect 19798 14662 19850 14714
rect 13360 14560 13412 14612
rect 18972 14603 19024 14612
rect 18972 14569 18981 14603
rect 18981 14569 19015 14603
rect 19015 14569 19024 14603
rect 18972 14560 19024 14569
rect 15844 14535 15896 14544
rect 15844 14501 15853 14535
rect 15853 14501 15887 14535
rect 15887 14501 15896 14535
rect 15844 14492 15896 14501
rect 11060 14424 11112 14476
rect 11520 14424 11572 14476
rect 15200 14424 15252 14476
rect 17960 14424 18012 14476
rect 23296 14467 23348 14476
rect 23296 14433 23305 14467
rect 23305 14433 23339 14467
rect 23339 14433 23348 14467
rect 23296 14424 23348 14433
rect 15292 14399 15344 14408
rect 15292 14365 15301 14399
rect 15301 14365 15335 14399
rect 15335 14365 15344 14399
rect 15292 14356 15344 14365
rect 17500 14356 17552 14408
rect 18328 14356 18380 14408
rect 22100 14220 22152 14272
rect 23112 14263 23164 14272
rect 23112 14229 23121 14263
rect 23121 14229 23155 14263
rect 23155 14229 23164 14263
rect 23112 14220 23164 14229
rect 4246 14118 4298 14170
rect 4310 14118 4362 14170
rect 4374 14118 4426 14170
rect 4438 14118 4490 14170
rect 34966 14118 35018 14170
rect 35030 14118 35082 14170
rect 35094 14118 35146 14170
rect 35158 14118 35210 14170
rect 11520 14059 11572 14068
rect 11520 14025 11529 14059
rect 11529 14025 11563 14059
rect 11563 14025 11572 14059
rect 11520 14016 11572 14025
rect 15200 14016 15252 14068
rect 17960 14016 18012 14068
rect 18328 14059 18380 14068
rect 18328 14025 18337 14059
rect 18337 14025 18371 14059
rect 18371 14025 18380 14059
rect 18328 14016 18380 14025
rect 23296 14016 23348 14068
rect 15292 13991 15344 14000
rect 15292 13957 15301 13991
rect 15301 13957 15335 13991
rect 15335 13957 15344 13991
rect 15292 13948 15344 13957
rect 24952 13991 25004 14000
rect 24952 13957 24961 13991
rect 24961 13957 24995 13991
rect 24995 13957 25004 13991
rect 24952 13948 25004 13957
rect 25136 13855 25188 13864
rect 25136 13821 25145 13855
rect 25145 13821 25179 13855
rect 25179 13821 25188 13855
rect 25136 13812 25188 13821
rect 19606 13574 19658 13626
rect 19670 13574 19722 13626
rect 19734 13574 19786 13626
rect 19798 13574 19850 13626
rect 13360 13472 13412 13524
rect 21272 13472 21324 13524
rect 17868 13404 17920 13456
rect 16764 13379 16816 13388
rect 16764 13345 16773 13379
rect 16773 13345 16807 13379
rect 16807 13345 16816 13379
rect 16764 13336 16816 13345
rect 16948 13379 17000 13388
rect 16948 13345 16957 13379
rect 16957 13345 16991 13379
rect 16991 13345 17000 13379
rect 16948 13336 17000 13345
rect 17316 13379 17368 13388
rect 17316 13345 17325 13379
rect 17325 13345 17359 13379
rect 17359 13345 17368 13379
rect 17316 13336 17368 13345
rect 21916 13336 21968 13388
rect 16488 13311 16540 13320
rect 16488 13277 16497 13311
rect 16497 13277 16531 13311
rect 16531 13277 16540 13311
rect 16488 13268 16540 13277
rect 16580 13268 16632 13320
rect 4246 13030 4298 13082
rect 4310 13030 4362 13082
rect 4374 13030 4426 13082
rect 4438 13030 4490 13082
rect 34966 13030 35018 13082
rect 35030 13030 35082 13082
rect 35094 13030 35146 13082
rect 35158 13030 35210 13082
rect 15016 12928 15068 12980
rect 16580 12928 16632 12980
rect 16948 12928 17000 12980
rect 17132 12928 17184 12980
rect 21916 12971 21968 12980
rect 21916 12937 21925 12971
rect 21925 12937 21959 12971
rect 21959 12937 21968 12971
rect 21916 12928 21968 12937
rect 15936 12860 15988 12912
rect 17316 12860 17368 12912
rect 13912 12835 13964 12844
rect 13912 12801 13921 12835
rect 13921 12801 13955 12835
rect 13955 12801 13964 12835
rect 13912 12792 13964 12801
rect 14924 12792 14976 12844
rect 16764 12835 16816 12844
rect 16764 12801 16773 12835
rect 16773 12801 16807 12835
rect 16807 12801 16816 12835
rect 16764 12792 16816 12801
rect 12440 12724 12492 12776
rect 13360 12724 13412 12776
rect 14740 12724 14792 12776
rect 15108 12588 15160 12640
rect 30288 12588 30340 12640
rect 30472 12588 30524 12640
rect 19606 12486 19658 12538
rect 19670 12486 19722 12538
rect 19734 12486 19786 12538
rect 19798 12486 19850 12538
rect 17132 12384 17184 12436
rect 34704 12384 34756 12436
rect 35348 12384 35400 12436
rect 13176 12359 13228 12368
rect 13176 12325 13185 12359
rect 13185 12325 13219 12359
rect 13219 12325 13228 12359
rect 13176 12316 13228 12325
rect 13728 12248 13780 12300
rect 14004 12316 14056 12368
rect 15108 12316 15160 12368
rect 18420 12316 18472 12368
rect 13912 12248 13964 12300
rect 12716 12180 12768 12232
rect 13360 12180 13412 12232
rect 15016 12248 15068 12300
rect 17500 12248 17552 12300
rect 19248 12291 19300 12300
rect 19248 12257 19257 12291
rect 19257 12257 19291 12291
rect 19291 12257 19300 12291
rect 19248 12248 19300 12257
rect 16396 12223 16448 12232
rect 16396 12189 16405 12223
rect 16405 12189 16439 12223
rect 16439 12189 16448 12223
rect 16396 12180 16448 12189
rect 18052 12180 18104 12232
rect 18328 12180 18380 12232
rect 18604 12112 18656 12164
rect 15292 12044 15344 12096
rect 15752 12044 15804 12096
rect 17868 12044 17920 12096
rect 18420 12087 18472 12096
rect 18420 12053 18429 12087
rect 18429 12053 18463 12087
rect 18463 12053 18472 12087
rect 18420 12044 18472 12053
rect 18880 12087 18932 12096
rect 18880 12053 18889 12087
rect 18889 12053 18923 12087
rect 18923 12053 18932 12087
rect 18880 12044 18932 12053
rect 4246 11942 4298 11994
rect 4310 11942 4362 11994
rect 4374 11942 4426 11994
rect 4438 11942 4490 11994
rect 34966 11942 35018 11994
rect 35030 11942 35082 11994
rect 35094 11942 35146 11994
rect 35158 11942 35210 11994
rect 13360 11840 13412 11892
rect 14004 11883 14056 11892
rect 14004 11849 14013 11883
rect 14013 11849 14047 11883
rect 14047 11849 14056 11883
rect 14004 11840 14056 11849
rect 14740 11840 14792 11892
rect 13912 11772 13964 11824
rect 15936 11840 15988 11892
rect 16396 11840 16448 11892
rect 17500 11883 17552 11892
rect 17500 11849 17509 11883
rect 17509 11849 17543 11883
rect 17543 11849 17552 11883
rect 17500 11840 17552 11849
rect 18328 11883 18380 11892
rect 18328 11849 18337 11883
rect 18337 11849 18371 11883
rect 18371 11849 18380 11883
rect 18328 11840 18380 11849
rect 21548 11840 21600 11892
rect 15292 11636 15344 11688
rect 19432 11679 19484 11688
rect 19432 11645 19441 11679
rect 19441 11645 19475 11679
rect 19475 11645 19484 11679
rect 19432 11636 19484 11645
rect 19984 11636 20036 11688
rect 19248 11568 19300 11620
rect 13728 11500 13780 11552
rect 16212 11500 16264 11552
rect 18604 11543 18656 11552
rect 18604 11509 18613 11543
rect 18613 11509 18647 11543
rect 18647 11509 18656 11543
rect 18604 11500 18656 11509
rect 19606 11398 19658 11450
rect 19670 11398 19722 11450
rect 19734 11398 19786 11450
rect 19798 11398 19850 11450
rect 15292 11228 15344 11280
rect 19248 11271 19300 11280
rect 16212 11203 16264 11212
rect 16212 11169 16221 11203
rect 16221 11169 16255 11203
rect 16255 11169 16264 11203
rect 16212 11160 16264 11169
rect 19248 11237 19257 11271
rect 19257 11237 19291 11271
rect 19291 11237 19300 11271
rect 19248 11228 19300 11237
rect 13728 11092 13780 11144
rect 16396 11092 16448 11144
rect 16488 11135 16540 11144
rect 16488 11101 16497 11135
rect 16497 11101 16531 11135
rect 16531 11101 16540 11135
rect 18604 11160 18656 11212
rect 16488 11092 16540 11101
rect 17500 11092 17552 11144
rect 17868 11135 17920 11144
rect 17868 11101 17877 11135
rect 17877 11101 17911 11135
rect 17911 11101 17920 11135
rect 17868 11092 17920 11101
rect 15844 11067 15896 11076
rect 15844 11033 15853 11067
rect 15853 11033 15887 11067
rect 15887 11033 15896 11067
rect 15844 11024 15896 11033
rect 18604 11024 18656 11076
rect 19432 11024 19484 11076
rect 4246 10854 4298 10906
rect 4310 10854 4362 10906
rect 4374 10854 4426 10906
rect 4438 10854 4490 10906
rect 34966 10854 35018 10906
rect 35030 10854 35082 10906
rect 35094 10854 35146 10906
rect 35158 10854 35210 10906
rect 15292 10795 15344 10804
rect 15292 10761 15301 10795
rect 15301 10761 15335 10795
rect 15335 10761 15344 10795
rect 15292 10752 15344 10761
rect 16212 10752 16264 10804
rect 17868 10752 17920 10804
rect 16396 10684 16448 10736
rect 17500 10684 17552 10736
rect 18236 10727 18288 10736
rect 18236 10693 18245 10727
rect 18245 10693 18279 10727
rect 18279 10693 18288 10727
rect 18236 10684 18288 10693
rect 18604 10684 18656 10736
rect 16488 10616 16540 10668
rect 19606 10310 19658 10362
rect 19670 10310 19722 10362
rect 19734 10310 19786 10362
rect 19798 10310 19850 10362
rect 9404 10140 9456 10192
rect 1584 10072 1636 10124
rect 2044 10072 2096 10124
rect 7104 10115 7156 10124
rect 7104 10081 7113 10115
rect 7113 10081 7147 10115
rect 7147 10081 7156 10115
rect 7104 10072 7156 10081
rect 7196 10072 7248 10124
rect 1400 10004 1452 10056
rect 3148 10047 3200 10056
rect 3148 10013 3157 10047
rect 3157 10013 3191 10047
rect 3191 10013 3200 10047
rect 3148 10004 3200 10013
rect 4246 9766 4298 9818
rect 4310 9766 4362 9818
rect 4374 9766 4426 9818
rect 4438 9766 4490 9818
rect 34966 9766 35018 9818
rect 35030 9766 35082 9818
rect 35094 9766 35146 9818
rect 35158 9766 35210 9818
rect 2044 9707 2096 9716
rect 2044 9673 2053 9707
rect 2053 9673 2087 9707
rect 2087 9673 2096 9707
rect 2044 9664 2096 9673
rect 7104 9664 7156 9716
rect 2872 9596 2924 9648
rect 3332 9596 3384 9648
rect 1584 9367 1636 9376
rect 1584 9333 1593 9367
rect 1593 9333 1627 9367
rect 1627 9333 1636 9367
rect 1584 9324 1636 9333
rect 7196 9367 7248 9376
rect 7196 9333 7205 9367
rect 7205 9333 7239 9367
rect 7239 9333 7248 9367
rect 7196 9324 7248 9333
rect 19606 9222 19658 9274
rect 19670 9222 19722 9274
rect 19734 9222 19786 9274
rect 19798 9222 19850 9274
rect 4246 8678 4298 8730
rect 4310 8678 4362 8730
rect 4374 8678 4426 8730
rect 4438 8678 4490 8730
rect 34966 8678 35018 8730
rect 35030 8678 35082 8730
rect 35094 8678 35146 8730
rect 35158 8678 35210 8730
rect 19606 8134 19658 8186
rect 19670 8134 19722 8186
rect 19734 8134 19786 8186
rect 19798 8134 19850 8186
rect 37464 7692 37516 7744
rect 39580 7692 39632 7744
rect 4246 7590 4298 7642
rect 4310 7590 4362 7642
rect 4374 7590 4426 7642
rect 4438 7590 4490 7642
rect 34966 7590 35018 7642
rect 35030 7590 35082 7642
rect 35094 7590 35146 7642
rect 35158 7590 35210 7642
rect 4620 7488 4672 7540
rect 5080 7488 5132 7540
rect 37556 7488 37608 7540
rect 39120 7488 39172 7540
rect 12348 7284 12400 7336
rect 13452 7284 13504 7336
rect 19606 7046 19658 7098
rect 19670 7046 19722 7098
rect 19734 7046 19786 7098
rect 19798 7046 19850 7098
rect 4246 6502 4298 6554
rect 4310 6502 4362 6554
rect 4374 6502 4426 6554
rect 4438 6502 4490 6554
rect 34966 6502 35018 6554
rect 35030 6502 35082 6554
rect 35094 6502 35146 6554
rect 35158 6502 35210 6554
rect 36268 6307 36320 6316
rect 36268 6273 36277 6307
rect 36277 6273 36311 6307
rect 36311 6273 36320 6307
rect 36268 6264 36320 6273
rect 35992 6239 36044 6248
rect 35992 6205 36001 6239
rect 36001 6205 36035 6239
rect 36035 6205 36044 6239
rect 35992 6196 36044 6205
rect 37372 6103 37424 6112
rect 37372 6069 37381 6103
rect 37381 6069 37415 6103
rect 37415 6069 37424 6103
rect 37372 6060 37424 6069
rect 19606 5958 19658 6010
rect 19670 5958 19722 6010
rect 19734 5958 19786 6010
rect 19798 5958 19850 6010
rect 35992 5695 36044 5704
rect 35992 5661 36001 5695
rect 36001 5661 36035 5695
rect 36035 5661 36044 5695
rect 35992 5652 36044 5661
rect 4246 5414 4298 5466
rect 4310 5414 4362 5466
rect 4374 5414 4426 5466
rect 4438 5414 4490 5466
rect 34966 5414 35018 5466
rect 35030 5414 35082 5466
rect 35094 5414 35146 5466
rect 35158 5414 35210 5466
rect 19606 4870 19658 4922
rect 19670 4870 19722 4922
rect 19734 4870 19786 4922
rect 19798 4870 19850 4922
rect 14004 4811 14056 4820
rect 14004 4777 14013 4811
rect 14013 4777 14047 4811
rect 14047 4777 14056 4811
rect 14004 4768 14056 4777
rect 21732 4768 21784 4820
rect 22008 4768 22060 4820
rect 29000 4768 29052 4820
rect 29368 4768 29420 4820
rect 33140 4768 33192 4820
rect 33508 4768 33560 4820
rect 12440 4675 12492 4684
rect 12440 4641 12449 4675
rect 12449 4641 12483 4675
rect 12483 4641 12492 4675
rect 12440 4632 12492 4641
rect 12716 4607 12768 4616
rect 12716 4573 12725 4607
rect 12725 4573 12759 4607
rect 12759 4573 12768 4607
rect 12716 4564 12768 4573
rect 4246 4326 4298 4378
rect 4310 4326 4362 4378
rect 4374 4326 4426 4378
rect 4438 4326 4490 4378
rect 34966 4326 35018 4378
rect 35030 4326 35082 4378
rect 35094 4326 35146 4378
rect 35158 4326 35210 4378
rect 12716 4267 12768 4276
rect 12716 4233 12725 4267
rect 12725 4233 12759 4267
rect 12759 4233 12768 4267
rect 12716 4224 12768 4233
rect 12440 4156 12492 4208
rect 6920 4088 6972 4140
rect 8208 4088 8260 4140
rect 8392 4088 8444 4140
rect 9220 4088 9272 4140
rect 10140 4088 10192 4140
rect 10692 4088 10744 4140
rect 17960 4088 18012 4140
rect 19156 4088 19208 4140
rect 21824 4088 21876 4140
rect 19432 3952 19484 4004
rect 22744 4020 22796 4072
rect 11980 3884 12032 3936
rect 12716 3884 12768 3936
rect 19606 3782 19658 3834
rect 19670 3782 19722 3834
rect 19734 3782 19786 3834
rect 19798 3782 19850 3834
rect 14280 3723 14332 3732
rect 14280 3689 14289 3723
rect 14289 3689 14323 3723
rect 14323 3689 14332 3723
rect 14280 3680 14332 3689
rect 12440 3544 12492 3596
rect 12808 3544 12860 3596
rect 20 3476 72 3528
rect 1308 3476 1360 3528
rect 19432 3340 19484 3392
rect 20812 3340 20864 3392
rect 4246 3238 4298 3290
rect 4310 3238 4362 3290
rect 4374 3238 4426 3290
rect 4438 3238 4490 3290
rect 34966 3238 35018 3290
rect 35030 3238 35082 3290
rect 35094 3238 35146 3290
rect 35158 3238 35210 3290
rect 12440 3136 12492 3188
rect 14832 3136 14884 3188
rect 22376 3136 22428 3188
rect 20720 3068 20772 3120
rect 13820 3043 13872 3052
rect 13820 3009 13829 3043
rect 13829 3009 13863 3043
rect 13863 3009 13872 3043
rect 13820 3000 13872 3009
rect 12532 2932 12584 2984
rect 20812 2932 20864 2984
rect 11060 2864 11112 2916
rect 12440 2864 12492 2916
rect 12808 2839 12860 2848
rect 12808 2805 12817 2839
rect 12817 2805 12851 2839
rect 12851 2805 12860 2839
rect 12808 2796 12860 2805
rect 19606 2694 19658 2746
rect 19670 2694 19722 2746
rect 19734 2694 19786 2746
rect 19798 2694 19850 2746
rect 12440 2635 12492 2644
rect 12440 2601 12449 2635
rect 12449 2601 12483 2635
rect 12483 2601 12492 2635
rect 14188 2635 14240 2644
rect 12440 2592 12492 2601
rect 14188 2601 14197 2635
rect 14197 2601 14231 2635
rect 14231 2601 14240 2635
rect 14188 2592 14240 2601
rect 20812 2635 20864 2644
rect 20812 2601 20821 2635
rect 20821 2601 20855 2635
rect 20855 2601 20864 2635
rect 20812 2592 20864 2601
rect 28448 2635 28500 2644
rect 28448 2601 28457 2635
rect 28457 2601 28491 2635
rect 28491 2601 28500 2635
rect 28448 2592 28500 2601
rect 18236 2456 18288 2508
rect 12532 2388 12584 2440
rect 18972 2388 19024 2440
rect 27620 2456 27672 2508
rect 23756 2363 23808 2372
rect 23756 2329 23765 2363
rect 23765 2329 23799 2363
rect 23799 2329 23808 2363
rect 23756 2320 23808 2329
rect 19800 2252 19852 2304
rect 26148 2388 26200 2440
rect 27160 2431 27212 2440
rect 27160 2397 27169 2431
rect 27169 2397 27203 2431
rect 27203 2397 27212 2431
rect 27160 2388 27212 2397
rect 28540 2388 28592 2440
rect 27160 2252 27212 2304
rect 4246 2150 4298 2202
rect 4310 2150 4362 2202
rect 4374 2150 4426 2202
rect 4438 2150 4490 2202
rect 34966 2150 35018 2202
rect 35030 2150 35082 2202
rect 35094 2150 35146 2202
rect 35158 2150 35210 2202
rect 23480 1368 23532 1420
rect 24584 1368 24636 1420
rect 480 1232 532 1284
rect 4804 1232 4856 1284
rect 3240 892 3292 944
rect 3332 892 3384 944
<< metal2 >>
rect 478 79200 534 80000
rect 938 79200 994 80000
rect 1858 79200 1914 80000
rect 2778 79200 2834 80000
rect 3698 79200 3754 80000
rect 3974 79656 4030 79665
rect 3974 79591 4030 79600
rect 112 75880 164 75886
rect 492 75857 520 79200
rect 952 75886 980 79200
rect 940 75880 992 75886
rect 112 75822 164 75828
rect 478 75848 534 75857
rect 124 69873 152 75822
rect 940 75822 992 75828
rect 1674 75848 1730 75857
rect 478 75783 534 75792
rect 1674 75783 1730 75792
rect 110 69864 166 69873
rect 110 69799 166 69808
rect 1582 66736 1638 66745
rect 1582 66671 1638 66680
rect 1596 65210 1624 66671
rect 1584 65204 1636 65210
rect 1584 65146 1636 65152
rect 1584 65068 1636 65074
rect 1584 65010 1636 65016
rect 1596 64326 1624 65010
rect 1584 64320 1636 64326
rect 1584 64262 1636 64268
rect 1596 63918 1624 64262
rect 1584 63912 1636 63918
rect 1584 63854 1636 63860
rect 1596 59226 1624 63854
rect 1584 59220 1636 59226
rect 1584 59162 1636 59168
rect 1596 58546 1624 59162
rect 1584 58540 1636 58546
rect 1584 58482 1636 58488
rect 1400 46912 1452 46918
rect 1400 46854 1452 46860
rect 1412 46510 1440 46854
rect 1688 46578 1716 75783
rect 1872 75449 1900 79200
rect 2410 76936 2466 76945
rect 2410 76871 2466 76880
rect 1858 75440 1914 75449
rect 1858 75375 1914 75384
rect 1768 65408 1820 65414
rect 1768 65350 1820 65356
rect 1780 65074 1808 65350
rect 1768 65068 1820 65074
rect 1768 65010 1820 65016
rect 1858 64016 1914 64025
rect 1858 63951 1860 63960
rect 1912 63951 1914 63960
rect 1860 63922 1912 63928
rect 1872 63578 1900 63922
rect 1860 63572 1912 63578
rect 1860 63514 1912 63520
rect 1858 59936 1914 59945
rect 1858 59871 1914 59880
rect 1872 58546 1900 59871
rect 1860 58540 1912 58546
rect 1860 58482 1912 58488
rect 1872 58138 1900 58482
rect 1860 58132 1912 58138
rect 1860 58074 1912 58080
rect 1676 46572 1728 46578
rect 1676 46514 1728 46520
rect 1400 46504 1452 46510
rect 1400 46446 1452 46452
rect 1306 46064 1362 46073
rect 1306 45999 1362 46008
rect 1320 3534 1348 45999
rect 1412 44878 1440 46446
rect 1688 46170 1716 46514
rect 1766 46336 1822 46345
rect 1766 46271 1822 46280
rect 1676 46164 1728 46170
rect 1676 46106 1728 46112
rect 1780 44946 1808 46271
rect 1768 44940 1820 44946
rect 1768 44882 1820 44888
rect 1400 44872 1452 44878
rect 1400 44814 1452 44820
rect 1780 44538 1808 44882
rect 1952 44872 2004 44878
rect 2004 44820 2084 44826
rect 1952 44814 2084 44820
rect 1964 44798 2084 44814
rect 1768 44532 1820 44538
rect 1768 44474 1820 44480
rect 2056 44334 2084 44798
rect 2044 44328 2096 44334
rect 2042 44296 2044 44305
rect 2096 44296 2098 44305
rect 2042 44231 2098 44240
rect 2424 40662 2452 76871
rect 2792 74662 2820 79200
rect 3330 75576 3386 75585
rect 3330 75511 3386 75520
rect 2780 74656 2832 74662
rect 2780 74598 2832 74604
rect 3238 69456 3294 69465
rect 3238 69391 3294 69400
rect 2870 65376 2926 65385
rect 2870 65311 2926 65320
rect 2688 63912 2740 63918
rect 2688 63854 2740 63860
rect 2700 63374 2728 63854
rect 2688 63368 2740 63374
rect 2688 63310 2740 63316
rect 2412 40656 2464 40662
rect 1950 40624 2006 40633
rect 2412 40598 2464 40604
rect 1950 40559 2006 40568
rect 1964 40390 1992 40559
rect 2228 40520 2280 40526
rect 2228 40462 2280 40468
rect 1952 40384 2004 40390
rect 1952 40326 2004 40332
rect 1964 40050 1992 40326
rect 1952 40044 2004 40050
rect 1952 39986 2004 39992
rect 1676 39976 1728 39982
rect 1596 39924 1676 39930
rect 1596 39918 1728 39924
rect 1596 39902 1716 39918
rect 1596 39574 1624 39902
rect 1584 39568 1636 39574
rect 1582 39536 1584 39545
rect 1636 39536 1638 39545
rect 1582 39471 1638 39480
rect 1676 38956 1728 38962
rect 1676 38898 1728 38904
rect 1688 38554 1716 38898
rect 1964 38894 1992 39986
rect 2240 39302 2268 40462
rect 2424 39642 2452 40598
rect 2412 39636 2464 39642
rect 2412 39578 2464 39584
rect 2228 39296 2280 39302
rect 2228 39238 2280 39244
rect 1952 38888 2004 38894
rect 1952 38830 2004 38836
rect 1964 38554 1992 38830
rect 1676 38548 1728 38554
rect 1676 38490 1728 38496
rect 1952 38548 2004 38554
rect 1952 38490 2004 38496
rect 1964 35290 1992 38490
rect 1676 35284 1728 35290
rect 1676 35226 1728 35232
rect 1952 35284 2004 35290
rect 1952 35226 2004 35232
rect 1688 34610 1716 35226
rect 1676 34604 1728 34610
rect 1676 34546 1728 34552
rect 1688 32570 1716 34546
rect 1952 34536 2004 34542
rect 1952 34478 2004 34484
rect 1964 33862 1992 34478
rect 1952 33856 2004 33862
rect 1952 33798 2004 33804
rect 1676 32564 1728 32570
rect 1676 32506 1728 32512
rect 1688 29850 1716 32506
rect 1676 29844 1728 29850
rect 1728 29804 1808 29832
rect 1676 29786 1728 29792
rect 1676 29640 1728 29646
rect 1676 29582 1728 29588
rect 1688 28966 1716 29582
rect 1780 29306 1808 29804
rect 1858 29336 1914 29345
rect 1768 29300 1820 29306
rect 1858 29271 1914 29280
rect 1768 29242 1820 29248
rect 1676 28960 1728 28966
rect 1676 28902 1728 28908
rect 1688 28218 1716 28902
rect 1676 28212 1728 28218
rect 1676 28154 1728 28160
rect 1584 28008 1636 28014
rect 1584 27950 1636 27956
rect 1596 27334 1624 27950
rect 1584 27328 1636 27334
rect 1584 27270 1636 27276
rect 1596 26625 1624 27270
rect 1872 26994 1900 29271
rect 1860 26988 1912 26994
rect 1860 26930 1912 26936
rect 1676 26920 1728 26926
rect 1676 26862 1728 26868
rect 1582 26616 1638 26625
rect 1582 26551 1638 26560
rect 1688 26450 1716 26862
rect 1872 26586 1900 26930
rect 1860 26580 1912 26586
rect 1860 26522 1912 26528
rect 1676 26444 1728 26450
rect 1676 26386 1728 26392
rect 1768 23520 1820 23526
rect 1768 23462 1820 23468
rect 1400 22976 1452 22982
rect 1400 22918 1452 22924
rect 1412 22574 1440 22918
rect 1400 22568 1452 22574
rect 1400 22510 1452 22516
rect 1412 16969 1440 22510
rect 1780 19145 1808 23462
rect 1860 22568 1912 22574
rect 1860 22510 1912 22516
rect 1872 21894 1900 22510
rect 1860 21888 1912 21894
rect 1860 21830 1912 21836
rect 1872 20806 1900 21830
rect 1860 20800 1912 20806
rect 1860 20742 1912 20748
rect 1766 19136 1822 19145
rect 1766 19071 1822 19080
rect 1398 16960 1454 16969
rect 1398 16895 1454 16904
rect 1412 16794 1440 16895
rect 1400 16788 1452 16794
rect 1400 16730 1452 16736
rect 1412 16114 1440 16730
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 1584 16108 1636 16114
rect 1584 16050 1636 16056
rect 1412 10062 1440 16050
rect 1596 15366 1624 16050
rect 1584 15360 1636 15366
rect 1582 15328 1584 15337
rect 1636 15328 1638 15337
rect 1582 15263 1638 15272
rect 1964 13841 1992 33798
rect 2240 28218 2268 39238
rect 2424 38962 2452 39578
rect 2412 38956 2464 38962
rect 2412 38898 2464 38904
rect 2780 38752 2832 38758
rect 2780 38694 2832 38700
rect 2792 38185 2820 38694
rect 2778 38176 2834 38185
rect 2778 38111 2834 38120
rect 2884 29850 2912 65311
rect 2964 58336 3016 58342
rect 2964 58278 3016 58284
rect 2976 36553 3004 58278
rect 3056 46436 3108 46442
rect 3056 46378 3108 46384
rect 3068 46209 3096 46378
rect 3054 46200 3110 46209
rect 3054 46135 3110 46144
rect 3056 44736 3108 44742
rect 3056 44678 3108 44684
rect 3068 43353 3096 44678
rect 3054 43344 3110 43353
rect 3054 43279 3110 43288
rect 3054 36816 3110 36825
rect 3054 36751 3110 36760
rect 2962 36544 3018 36553
rect 2962 36479 3018 36488
rect 3068 34746 3096 36751
rect 3056 34740 3108 34746
rect 3056 34682 3108 34688
rect 2872 29844 2924 29850
rect 2872 29786 2924 29792
rect 2780 29300 2832 29306
rect 2780 29242 2832 29248
rect 2228 28212 2280 28218
rect 2228 28154 2280 28160
rect 2044 26444 2096 26450
rect 2044 26386 2096 26392
rect 2056 23730 2084 26386
rect 2044 23724 2096 23730
rect 2044 23666 2096 23672
rect 2056 23322 2084 23666
rect 2044 23316 2096 23322
rect 2044 23258 2096 23264
rect 2240 16561 2268 28154
rect 2792 26450 2820 29242
rect 2780 26444 2832 26450
rect 2780 26386 2832 26392
rect 2688 24812 2740 24818
rect 2688 24754 2740 24760
rect 2700 23361 2728 24754
rect 2686 23352 2742 23361
rect 2686 23287 2742 23296
rect 3146 23352 3202 23361
rect 3146 23287 3202 23296
rect 3160 22778 3188 23287
rect 3148 22772 3200 22778
rect 3148 22714 3200 22720
rect 2688 20800 2740 20806
rect 2688 20742 2740 20748
rect 2226 16552 2282 16561
rect 2226 16487 2282 16496
rect 2700 15314 2728 20742
rect 2870 19136 2926 19145
rect 2870 19071 2926 19080
rect 2700 15286 2820 15314
rect 1950 13832 2006 13841
rect 1950 13767 2006 13776
rect 2792 13705 2820 15286
rect 2778 13696 2834 13705
rect 2778 13631 2834 13640
rect 2778 12336 2834 12345
rect 2778 12271 2834 12280
rect 2792 11801 2820 12271
rect 2778 11792 2834 11801
rect 2778 11727 2834 11736
rect 2686 10568 2742 10577
rect 2686 10503 2742 10512
rect 2042 10160 2098 10169
rect 1584 10124 1636 10130
rect 2042 10095 2044 10104
rect 1584 10066 1636 10072
rect 2096 10095 2098 10104
rect 2044 10066 2096 10072
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1596 9382 1624 10066
rect 2056 9722 2084 10066
rect 2044 9716 2096 9722
rect 2044 9658 2096 9664
rect 1584 9376 1636 9382
rect 1584 9318 1636 9324
rect 1596 8945 1624 9318
rect 1582 8936 1638 8945
rect 1582 8871 1638 8880
rect 1398 7848 1454 7857
rect 1398 7783 1454 7792
rect 20 3528 72 3534
rect 20 3470 72 3476
rect 1308 3528 1360 3534
rect 1308 3470 1360 3476
rect 32 800 60 3470
rect 480 1284 532 1290
rect 480 1226 532 1232
rect 492 800 520 1226
rect 1412 800 1440 7783
rect 2700 3346 2728 10503
rect 2884 9654 2912 19071
rect 3252 16250 3280 69391
rect 3344 68241 3372 75511
rect 3712 74746 3740 79200
rect 3988 77722 4016 79591
rect 4618 79200 4674 80000
rect 5538 79200 5594 80000
rect 6458 79200 6514 80000
rect 7378 79200 7434 80000
rect 8298 79200 8354 80000
rect 8758 79200 8814 80000
rect 9678 79200 9734 80000
rect 10598 79200 10654 80000
rect 11518 79200 11574 80000
rect 12438 79200 12494 80000
rect 13358 79200 13414 80000
rect 14278 79200 14334 80000
rect 15198 79200 15254 80000
rect 16118 79200 16174 80000
rect 16578 79200 16634 80000
rect 17498 79200 17554 80000
rect 18418 79200 18474 80000
rect 19338 79200 19394 80000
rect 20258 79200 20314 80000
rect 21178 79200 21234 80000
rect 22098 79200 22154 80000
rect 23018 79200 23074 80000
rect 23938 79200 23994 80000
rect 24398 79200 24454 80000
rect 25318 79200 25374 80000
rect 26238 79200 26294 80000
rect 27158 79200 27214 80000
rect 28078 79200 28134 80000
rect 28998 79200 29054 80000
rect 29918 79200 29974 80000
rect 30838 79200 30894 80000
rect 31758 79200 31814 80000
rect 32218 79200 32274 80000
rect 33138 79200 33194 80000
rect 34058 79200 34114 80000
rect 34978 79200 35034 80000
rect 35438 79656 35494 79665
rect 35438 79591 35494 79600
rect 4066 78296 4122 78305
rect 4066 78231 4122 78240
rect 3976 77716 4028 77722
rect 3976 77658 4028 77664
rect 4080 77586 4108 78231
rect 4068 77580 4120 77586
rect 4068 77522 4120 77528
rect 4220 77276 4516 77296
rect 4276 77274 4300 77276
rect 4356 77274 4380 77276
rect 4436 77274 4460 77276
rect 4298 77222 4300 77274
rect 4362 77222 4374 77274
rect 4436 77222 4438 77274
rect 4276 77220 4300 77222
rect 4356 77220 4380 77222
rect 4436 77220 4460 77222
rect 4220 77200 4516 77220
rect 4220 76188 4516 76208
rect 4276 76186 4300 76188
rect 4356 76186 4380 76188
rect 4436 76186 4460 76188
rect 4298 76134 4300 76186
rect 4362 76134 4374 76186
rect 4436 76134 4438 76186
rect 4276 76132 4300 76134
rect 4356 76132 4380 76134
rect 4436 76132 4460 76134
rect 4220 76112 4516 76132
rect 4220 75100 4516 75120
rect 4276 75098 4300 75100
rect 4356 75098 4380 75100
rect 4436 75098 4460 75100
rect 4298 75046 4300 75098
rect 4362 75046 4374 75098
rect 4436 75046 4438 75098
rect 4276 75044 4300 75046
rect 4356 75044 4380 75046
rect 4436 75044 4460 75046
rect 4220 75024 4516 75044
rect 4632 74769 4660 79200
rect 5552 79098 5580 79200
rect 5552 79070 5672 79098
rect 4618 74760 4674 74769
rect 3712 74718 4016 74746
rect 3884 74656 3936 74662
rect 3884 74598 3936 74604
rect 3790 74216 3846 74225
rect 3790 74151 3846 74160
rect 3804 72593 3832 74151
rect 3790 72584 3846 72593
rect 3790 72519 3846 72528
rect 3330 68232 3386 68241
rect 3330 68167 3386 68176
rect 3422 68096 3478 68105
rect 3422 68031 3478 68040
rect 3436 60625 3464 68031
rect 3896 63986 3924 74598
rect 3988 67153 4016 74718
rect 4618 74695 4674 74704
rect 4220 74012 4516 74032
rect 4276 74010 4300 74012
rect 4356 74010 4380 74012
rect 4436 74010 4460 74012
rect 4298 73958 4300 74010
rect 4362 73958 4374 74010
rect 4436 73958 4438 74010
rect 4276 73956 4300 73958
rect 4356 73956 4380 73958
rect 4436 73956 4460 73958
rect 4220 73936 4516 73956
rect 4220 72924 4516 72944
rect 4276 72922 4300 72924
rect 4356 72922 4380 72924
rect 4436 72922 4460 72924
rect 4298 72870 4300 72922
rect 4362 72870 4374 72922
rect 4436 72870 4438 72922
rect 4276 72868 4300 72870
rect 4356 72868 4380 72870
rect 4436 72868 4460 72870
rect 4066 72856 4122 72865
rect 4220 72848 4516 72868
rect 4066 72791 4122 72800
rect 4080 72049 4108 72791
rect 4066 72040 4122 72049
rect 4066 71975 4122 71984
rect 4220 71836 4516 71856
rect 4276 71834 4300 71836
rect 4356 71834 4380 71836
rect 4436 71834 4460 71836
rect 4298 71782 4300 71834
rect 4362 71782 4374 71834
rect 4436 71782 4438 71834
rect 4276 71780 4300 71782
rect 4356 71780 4380 71782
rect 4436 71780 4460 71782
rect 4220 71760 4516 71780
rect 4802 71632 4858 71641
rect 4802 71567 4858 71576
rect 4816 70825 4844 71567
rect 4802 70816 4858 70825
rect 4220 70748 4516 70768
rect 4802 70751 4858 70760
rect 4276 70746 4300 70748
rect 4356 70746 4380 70748
rect 4436 70746 4460 70748
rect 4298 70694 4300 70746
rect 4362 70694 4374 70746
rect 4436 70694 4438 70746
rect 4276 70692 4300 70694
rect 4356 70692 4380 70694
rect 4436 70692 4460 70694
rect 4220 70672 4516 70692
rect 4894 70136 4950 70145
rect 4894 70071 4950 70080
rect 4220 69660 4516 69680
rect 4276 69658 4300 69660
rect 4356 69658 4380 69660
rect 4436 69658 4460 69660
rect 4298 69606 4300 69658
rect 4362 69606 4374 69658
rect 4436 69606 4438 69658
rect 4276 69604 4300 69606
rect 4356 69604 4380 69606
rect 4436 69604 4460 69606
rect 4220 69584 4516 69604
rect 4220 68572 4516 68592
rect 4276 68570 4300 68572
rect 4356 68570 4380 68572
rect 4436 68570 4460 68572
rect 4298 68518 4300 68570
rect 4362 68518 4374 68570
rect 4436 68518 4438 68570
rect 4276 68516 4300 68518
rect 4356 68516 4380 68518
rect 4436 68516 4460 68518
rect 4220 68496 4516 68516
rect 4220 67484 4516 67504
rect 4276 67482 4300 67484
rect 4356 67482 4380 67484
rect 4436 67482 4460 67484
rect 4298 67430 4300 67482
rect 4362 67430 4374 67482
rect 4436 67430 4438 67482
rect 4276 67428 4300 67430
rect 4356 67428 4380 67430
rect 4436 67428 4460 67430
rect 4220 67408 4516 67428
rect 3974 67144 4030 67153
rect 3974 67079 4030 67088
rect 4220 66396 4516 66416
rect 4276 66394 4300 66396
rect 4356 66394 4380 66396
rect 4436 66394 4460 66396
rect 4298 66342 4300 66394
rect 4362 66342 4374 66394
rect 4436 66342 4438 66394
rect 4276 66340 4300 66342
rect 4356 66340 4380 66342
rect 4436 66340 4460 66342
rect 4220 66320 4516 66340
rect 4220 65308 4516 65328
rect 4276 65306 4300 65308
rect 4356 65306 4380 65308
rect 4436 65306 4460 65308
rect 4298 65254 4300 65306
rect 4362 65254 4374 65306
rect 4436 65254 4438 65306
rect 4276 65252 4300 65254
rect 4356 65252 4380 65254
rect 4436 65252 4460 65254
rect 4220 65232 4516 65252
rect 4620 64932 4672 64938
rect 4620 64874 4672 64880
rect 4220 64220 4516 64240
rect 4276 64218 4300 64220
rect 4356 64218 4380 64220
rect 4436 64218 4460 64220
rect 4298 64166 4300 64218
rect 4362 64166 4374 64218
rect 4436 64166 4438 64218
rect 4276 64164 4300 64166
rect 4356 64164 4380 64166
rect 4436 64164 4460 64166
rect 4220 64144 4516 64164
rect 4158 64016 4214 64025
rect 3884 63980 3936 63986
rect 4158 63951 4214 63960
rect 3884 63922 3936 63928
rect 4172 63918 4200 63951
rect 4160 63912 4212 63918
rect 4160 63854 4212 63860
rect 4252 63844 4304 63850
rect 4252 63786 4304 63792
rect 4264 63578 4292 63786
rect 4252 63572 4304 63578
rect 4252 63514 4304 63520
rect 4632 63442 4660 64874
rect 4620 63436 4672 63442
rect 4620 63378 4672 63384
rect 4220 63132 4516 63152
rect 4276 63130 4300 63132
rect 4356 63130 4380 63132
rect 4436 63130 4460 63132
rect 4298 63078 4300 63130
rect 4362 63078 4374 63130
rect 4436 63078 4438 63130
rect 4276 63076 4300 63078
rect 4356 63076 4380 63078
rect 4436 63076 4460 63078
rect 4220 63056 4516 63076
rect 4632 63034 4660 63378
rect 4620 63028 4672 63034
rect 4620 62970 4672 62976
rect 4220 62044 4516 62064
rect 4276 62042 4300 62044
rect 4356 62042 4380 62044
rect 4436 62042 4460 62044
rect 4298 61990 4300 62042
rect 4362 61990 4374 62042
rect 4436 61990 4438 62042
rect 4276 61988 4300 61990
rect 4356 61988 4380 61990
rect 4436 61988 4460 61990
rect 4220 61968 4516 61988
rect 4220 60956 4516 60976
rect 4276 60954 4300 60956
rect 4356 60954 4380 60956
rect 4436 60954 4460 60956
rect 4298 60902 4300 60954
rect 4362 60902 4374 60954
rect 4436 60902 4438 60954
rect 4276 60900 4300 60902
rect 4356 60900 4380 60902
rect 4436 60900 4460 60902
rect 4220 60880 4516 60900
rect 3422 60616 3478 60625
rect 3422 60551 3478 60560
rect 4908 59945 4936 70071
rect 5644 69601 5672 79070
rect 6472 75177 6500 79200
rect 6458 75168 6514 75177
rect 6458 75103 6514 75112
rect 7392 74905 7420 79200
rect 8312 79098 8340 79200
rect 8312 79070 8432 79098
rect 7378 74896 7434 74905
rect 7378 74831 7434 74840
rect 6182 74760 6238 74769
rect 6182 74695 6238 74704
rect 5630 69592 5686 69601
rect 5630 69527 5686 69536
rect 5080 63912 5132 63918
rect 5080 63854 5132 63860
rect 5092 63782 5120 63854
rect 5080 63776 5132 63782
rect 5080 63718 5132 63724
rect 4894 59936 4950 59945
rect 4220 59868 4516 59888
rect 4894 59871 4950 59880
rect 4276 59866 4300 59868
rect 4356 59866 4380 59868
rect 4436 59866 4460 59868
rect 4298 59814 4300 59866
rect 4362 59814 4374 59866
rect 4436 59814 4438 59866
rect 4276 59812 4300 59814
rect 4356 59812 4380 59814
rect 4436 59812 4460 59814
rect 4220 59792 4516 59812
rect 4220 58780 4516 58800
rect 4276 58778 4300 58780
rect 4356 58778 4380 58780
rect 4436 58778 4460 58780
rect 4298 58726 4300 58778
rect 4362 58726 4374 58778
rect 4436 58726 4438 58778
rect 4276 58724 4300 58726
rect 4356 58724 4380 58726
rect 4436 58724 4460 58726
rect 4220 58704 4516 58724
rect 4220 57692 4516 57712
rect 4276 57690 4300 57692
rect 4356 57690 4380 57692
rect 4436 57690 4460 57692
rect 4298 57638 4300 57690
rect 4362 57638 4374 57690
rect 4436 57638 4438 57690
rect 4276 57636 4300 57638
rect 4356 57636 4380 57638
rect 4436 57636 4460 57638
rect 4220 57616 4516 57636
rect 4220 56604 4516 56624
rect 4276 56602 4300 56604
rect 4356 56602 4380 56604
rect 4436 56602 4460 56604
rect 4298 56550 4300 56602
rect 4362 56550 4374 56602
rect 4436 56550 4438 56602
rect 4276 56548 4300 56550
rect 4356 56548 4380 56550
rect 4436 56548 4460 56550
rect 4220 56528 4516 56548
rect 3882 56400 3938 56409
rect 3882 56335 3938 56344
rect 3330 55176 3386 55185
rect 3330 55111 3386 55120
rect 3344 53145 3372 55111
rect 3698 53816 3754 53825
rect 3698 53751 3754 53760
rect 3330 53136 3386 53145
rect 3330 53071 3386 53080
rect 3330 52456 3386 52465
rect 3330 52391 3386 52400
rect 3344 49609 3372 52391
rect 3330 49600 3386 49609
rect 3330 49535 3386 49544
rect 3514 48648 3570 48657
rect 3514 48583 3570 48592
rect 3528 47025 3556 48583
rect 3712 47025 3740 53751
rect 3896 48385 3924 56335
rect 4220 55516 4516 55536
rect 4276 55514 4300 55516
rect 4356 55514 4380 55516
rect 4436 55514 4460 55516
rect 4298 55462 4300 55514
rect 4362 55462 4374 55514
rect 4436 55462 4438 55514
rect 4276 55460 4300 55462
rect 4356 55460 4380 55462
rect 4436 55460 4460 55462
rect 4220 55440 4516 55460
rect 4220 54428 4516 54448
rect 4276 54426 4300 54428
rect 4356 54426 4380 54428
rect 4436 54426 4460 54428
rect 4298 54374 4300 54426
rect 4362 54374 4374 54426
rect 4436 54374 4438 54426
rect 4276 54372 4300 54374
rect 4356 54372 4380 54374
rect 4436 54372 4460 54374
rect 4220 54352 4516 54372
rect 4220 53340 4516 53360
rect 4276 53338 4300 53340
rect 4356 53338 4380 53340
rect 4436 53338 4460 53340
rect 4298 53286 4300 53338
rect 4362 53286 4374 53338
rect 4436 53286 4438 53338
rect 4276 53284 4300 53286
rect 4356 53284 4380 53286
rect 4436 53284 4460 53286
rect 4220 53264 4516 53284
rect 4220 52252 4516 52272
rect 4276 52250 4300 52252
rect 4356 52250 4380 52252
rect 4436 52250 4460 52252
rect 4298 52198 4300 52250
rect 4362 52198 4374 52250
rect 4436 52198 4438 52250
rect 4276 52196 4300 52198
rect 4356 52196 4380 52198
rect 4436 52196 4460 52198
rect 4220 52176 4516 52196
rect 4220 51164 4516 51184
rect 4276 51162 4300 51164
rect 4356 51162 4380 51164
rect 4436 51162 4460 51164
rect 4298 51110 4300 51162
rect 4362 51110 4374 51162
rect 4436 51110 4438 51162
rect 4276 51108 4300 51110
rect 4356 51108 4380 51110
rect 4436 51108 4460 51110
rect 4220 51088 4516 51108
rect 4220 50076 4516 50096
rect 4276 50074 4300 50076
rect 4356 50074 4380 50076
rect 4436 50074 4460 50076
rect 4298 50022 4300 50074
rect 4362 50022 4374 50074
rect 4436 50022 4438 50074
rect 4276 50020 4300 50022
rect 4356 50020 4380 50022
rect 4436 50020 4460 50022
rect 4220 50000 4516 50020
rect 5092 49745 5120 63718
rect 5172 63368 5224 63374
rect 5172 63310 5224 63316
rect 5184 62694 5212 63310
rect 5172 62688 5224 62694
rect 5172 62630 5224 62636
rect 5184 62121 5212 62630
rect 5170 62112 5226 62121
rect 5170 62047 5226 62056
rect 6196 54505 6224 74695
rect 7378 69864 7434 69873
rect 7378 69799 7434 69808
rect 6920 63232 6972 63238
rect 6920 63174 6972 63180
rect 6182 54496 6238 54505
rect 6182 54431 6238 54440
rect 4066 49736 4122 49745
rect 4066 49671 4122 49680
rect 5078 49736 5134 49745
rect 5078 49671 5134 49680
rect 4080 48793 4108 49671
rect 4220 48988 4516 49008
rect 4276 48986 4300 48988
rect 4356 48986 4380 48988
rect 4436 48986 4460 48988
rect 4298 48934 4300 48986
rect 4362 48934 4374 48986
rect 4436 48934 4438 48986
rect 4276 48932 4300 48934
rect 4356 48932 4380 48934
rect 4436 48932 4460 48934
rect 4220 48912 4516 48932
rect 4066 48784 4122 48793
rect 4066 48719 4122 48728
rect 3882 48376 3938 48385
rect 3882 48311 3938 48320
rect 4220 47900 4516 47920
rect 4276 47898 4300 47900
rect 4356 47898 4380 47900
rect 4436 47898 4460 47900
rect 4298 47846 4300 47898
rect 4362 47846 4374 47898
rect 4436 47846 4438 47898
rect 4276 47844 4300 47846
rect 4356 47844 4380 47846
rect 4436 47844 4460 47846
rect 4220 47824 4516 47844
rect 3514 47016 3570 47025
rect 3514 46951 3570 46960
rect 3698 47016 3754 47025
rect 3698 46951 3754 46960
rect 6274 47016 6330 47025
rect 6274 46951 6330 46960
rect 4220 46812 4516 46832
rect 4276 46810 4300 46812
rect 4356 46810 4380 46812
rect 4436 46810 4460 46812
rect 4298 46758 4300 46810
rect 4362 46758 4374 46810
rect 4436 46758 4438 46810
rect 4276 46756 4300 46758
rect 4356 46756 4380 46758
rect 4436 46756 4460 46758
rect 4220 46736 4516 46756
rect 4220 45724 4516 45744
rect 4276 45722 4300 45724
rect 4356 45722 4380 45724
rect 4436 45722 4460 45724
rect 4298 45670 4300 45722
rect 4362 45670 4374 45722
rect 4436 45670 4438 45722
rect 4276 45668 4300 45670
rect 4356 45668 4380 45670
rect 4436 45668 4460 45670
rect 4220 45648 4516 45668
rect 4220 44636 4516 44656
rect 4276 44634 4300 44636
rect 4356 44634 4380 44636
rect 4436 44634 4460 44636
rect 4298 44582 4300 44634
rect 4362 44582 4374 44634
rect 4436 44582 4438 44634
rect 4276 44580 4300 44582
rect 4356 44580 4380 44582
rect 4436 44580 4460 44582
rect 4220 44560 4516 44580
rect 4220 43548 4516 43568
rect 4276 43546 4300 43548
rect 4356 43546 4380 43548
rect 4436 43546 4460 43548
rect 4298 43494 4300 43546
rect 4362 43494 4374 43546
rect 4436 43494 4438 43546
rect 4276 43492 4300 43494
rect 4356 43492 4380 43494
rect 4436 43492 4460 43494
rect 4220 43472 4516 43492
rect 4220 42460 4516 42480
rect 4276 42458 4300 42460
rect 4356 42458 4380 42460
rect 4436 42458 4460 42460
rect 4298 42406 4300 42458
rect 4362 42406 4374 42458
rect 4436 42406 4438 42458
rect 4276 42404 4300 42406
rect 4356 42404 4380 42406
rect 4436 42404 4460 42406
rect 4220 42384 4516 42404
rect 5722 41848 5778 41857
rect 5722 41783 5778 41792
rect 5736 41750 5764 41783
rect 5724 41744 5776 41750
rect 5724 41686 5776 41692
rect 4160 41676 4212 41682
rect 4160 41618 4212 41624
rect 3976 41608 4028 41614
rect 4172 41562 4200 41618
rect 3976 41550 4028 41556
rect 3988 41002 4016 41550
rect 4080 41534 4200 41562
rect 3976 40996 4028 41002
rect 3976 40938 4028 40944
rect 3882 40896 3938 40905
rect 3882 40831 3938 40840
rect 3790 40760 3846 40769
rect 3790 40695 3846 40704
rect 3514 37904 3570 37913
rect 3514 37839 3570 37848
rect 3330 32056 3386 32065
rect 3330 31991 3386 32000
rect 3344 30297 3372 31991
rect 3330 30288 3386 30297
rect 3330 30223 3386 30232
rect 3528 25265 3556 37839
rect 3698 37360 3754 37369
rect 3698 37295 3754 37304
rect 3712 27985 3740 37295
rect 3804 35465 3832 40695
rect 3896 39409 3924 40831
rect 3988 40633 4016 40938
rect 4080 40934 4108 41534
rect 4220 41372 4516 41392
rect 4276 41370 4300 41372
rect 4356 41370 4380 41372
rect 4436 41370 4460 41372
rect 4298 41318 4300 41370
rect 4362 41318 4374 41370
rect 4436 41318 4438 41370
rect 4276 41316 4300 41318
rect 4356 41316 4380 41318
rect 4436 41316 4460 41318
rect 4220 41296 4516 41316
rect 4068 40928 4120 40934
rect 4068 40870 4120 40876
rect 4080 40662 4108 40870
rect 4068 40656 4120 40662
rect 3974 40624 4030 40633
rect 4068 40598 4120 40604
rect 3974 40559 4030 40568
rect 4220 40284 4516 40304
rect 4276 40282 4300 40284
rect 4356 40282 4380 40284
rect 4436 40282 4460 40284
rect 4298 40230 4300 40282
rect 4362 40230 4374 40282
rect 4436 40230 4438 40282
rect 4276 40228 4300 40230
rect 4356 40228 4380 40230
rect 4436 40228 4460 40230
rect 4220 40208 4516 40228
rect 4068 39908 4120 39914
rect 4068 39850 4120 39856
rect 4080 39681 4108 39850
rect 4066 39672 4122 39681
rect 4066 39607 4122 39616
rect 3882 39400 3938 39409
rect 3882 39335 3938 39344
rect 4220 39196 4516 39216
rect 4276 39194 4300 39196
rect 4356 39194 4380 39196
rect 4436 39194 4460 39196
rect 4298 39142 4300 39194
rect 4362 39142 4374 39194
rect 4436 39142 4438 39194
rect 4276 39140 4300 39142
rect 4356 39140 4380 39142
rect 4436 39140 4460 39142
rect 4220 39120 4516 39140
rect 4220 38108 4516 38128
rect 4276 38106 4300 38108
rect 4356 38106 4380 38108
rect 4436 38106 4460 38108
rect 4298 38054 4300 38106
rect 4362 38054 4374 38106
rect 4436 38054 4438 38106
rect 4276 38052 4300 38054
rect 4356 38052 4380 38054
rect 4436 38052 4460 38054
rect 4220 38032 4516 38052
rect 4220 37020 4516 37040
rect 4276 37018 4300 37020
rect 4356 37018 4380 37020
rect 4436 37018 4460 37020
rect 4298 36966 4300 37018
rect 4362 36966 4374 37018
rect 4436 36966 4438 37018
rect 4276 36964 4300 36966
rect 4356 36964 4380 36966
rect 4436 36964 4460 36966
rect 4220 36944 4516 36964
rect 3882 36136 3938 36145
rect 3882 36071 3938 36080
rect 3790 35456 3846 35465
rect 3790 35391 3846 35400
rect 3896 34785 3924 36071
rect 4220 35932 4516 35952
rect 4276 35930 4300 35932
rect 4356 35930 4380 35932
rect 4436 35930 4460 35932
rect 4298 35878 4300 35930
rect 4362 35878 4374 35930
rect 4436 35878 4438 35930
rect 4276 35876 4300 35878
rect 4356 35876 4380 35878
rect 4436 35876 4460 35878
rect 4220 35856 4516 35876
rect 4220 34844 4516 34864
rect 4276 34842 4300 34844
rect 4356 34842 4380 34844
rect 4436 34842 4460 34844
rect 4298 34790 4300 34842
rect 4362 34790 4374 34842
rect 4436 34790 4438 34842
rect 4276 34788 4300 34790
rect 4356 34788 4380 34790
rect 4436 34788 4460 34790
rect 3882 34776 3938 34785
rect 4220 34768 4516 34788
rect 3882 34711 3938 34720
rect 4220 33756 4516 33776
rect 4276 33754 4300 33756
rect 4356 33754 4380 33756
rect 4436 33754 4460 33756
rect 4298 33702 4300 33754
rect 4362 33702 4374 33754
rect 4436 33702 4438 33754
rect 4276 33700 4300 33702
rect 4356 33700 4380 33702
rect 4436 33700 4460 33702
rect 4220 33680 4516 33700
rect 5448 33652 5500 33658
rect 5448 33594 5500 33600
rect 4220 32668 4516 32688
rect 4276 32666 4300 32668
rect 4356 32666 4380 32668
rect 4436 32666 4460 32668
rect 4298 32614 4300 32666
rect 4362 32614 4374 32666
rect 4436 32614 4438 32666
rect 4276 32612 4300 32614
rect 4356 32612 4380 32614
rect 4436 32612 4460 32614
rect 4220 32592 4516 32612
rect 5460 32570 5488 33594
rect 5448 32564 5500 32570
rect 5448 32506 5500 32512
rect 5460 32366 5488 32506
rect 5448 32360 5500 32366
rect 5448 32302 5500 32308
rect 4220 31580 4516 31600
rect 4276 31578 4300 31580
rect 4356 31578 4380 31580
rect 4436 31578 4460 31580
rect 4298 31526 4300 31578
rect 4362 31526 4374 31578
rect 4436 31526 4438 31578
rect 4276 31524 4300 31526
rect 4356 31524 4380 31526
rect 4436 31524 4460 31526
rect 4220 31504 4516 31524
rect 4066 30696 4122 30705
rect 4066 30631 4122 30640
rect 4080 28937 4108 30631
rect 4220 30492 4516 30512
rect 4276 30490 4300 30492
rect 4356 30490 4380 30492
rect 4436 30490 4460 30492
rect 4298 30438 4300 30490
rect 4362 30438 4374 30490
rect 4436 30438 4438 30490
rect 4276 30436 4300 30438
rect 4356 30436 4380 30438
rect 4436 30436 4460 30438
rect 4220 30416 4516 30436
rect 4220 29404 4516 29424
rect 4276 29402 4300 29404
rect 4356 29402 4380 29404
rect 4436 29402 4460 29404
rect 4298 29350 4300 29402
rect 4362 29350 4374 29402
rect 4436 29350 4438 29402
rect 4276 29348 4300 29350
rect 4356 29348 4380 29350
rect 4436 29348 4460 29350
rect 4220 29328 4516 29348
rect 4066 28928 4122 28937
rect 4066 28863 4122 28872
rect 4220 28316 4516 28336
rect 4276 28314 4300 28316
rect 4356 28314 4380 28316
rect 4436 28314 4460 28316
rect 4298 28262 4300 28314
rect 4362 28262 4374 28314
rect 4436 28262 4438 28314
rect 4276 28260 4300 28262
rect 4356 28260 4380 28262
rect 4436 28260 4460 28262
rect 4220 28240 4516 28260
rect 3698 27976 3754 27985
rect 3698 27911 3754 27920
rect 6000 27532 6052 27538
rect 6000 27474 6052 27480
rect 4220 27228 4516 27248
rect 4276 27226 4300 27228
rect 4356 27226 4380 27228
rect 4436 27226 4460 27228
rect 4298 27174 4300 27226
rect 4362 27174 4374 27226
rect 4436 27174 4438 27226
rect 4276 27172 4300 27174
rect 4356 27172 4380 27174
rect 4436 27172 4460 27174
rect 4220 27152 4516 27172
rect 4068 26852 4120 26858
rect 4068 26794 4120 26800
rect 4080 26353 4108 26794
rect 6012 26450 6040 27474
rect 6000 26444 6052 26450
rect 6184 26444 6236 26450
rect 6000 26386 6052 26392
rect 6104 26404 6184 26432
rect 4066 26344 4122 26353
rect 4066 26279 4122 26288
rect 4220 26140 4516 26160
rect 4276 26138 4300 26140
rect 4356 26138 4380 26140
rect 4436 26138 4460 26140
rect 4298 26086 4300 26138
rect 4362 26086 4374 26138
rect 4436 26086 4438 26138
rect 4276 26084 4300 26086
rect 4356 26084 4380 26086
rect 4436 26084 4460 26086
rect 4220 26064 4516 26084
rect 6012 26042 6040 26386
rect 6000 26036 6052 26042
rect 6000 25978 6052 25984
rect 6104 25702 6132 26404
rect 6184 26386 6236 26392
rect 6092 25696 6144 25702
rect 6092 25638 6144 25644
rect 3514 25256 3570 25265
rect 3514 25191 3570 25200
rect 4066 25256 4122 25265
rect 4066 25191 4122 25200
rect 4080 23905 4108 25191
rect 4220 25052 4516 25072
rect 4276 25050 4300 25052
rect 4356 25050 4380 25052
rect 4436 25050 4460 25052
rect 4298 24998 4300 25050
rect 4362 24998 4374 25050
rect 4436 24998 4438 25050
rect 4276 24996 4300 24998
rect 4356 24996 4380 24998
rect 4436 24996 4460 24998
rect 4220 24976 4516 24996
rect 4220 23964 4516 23984
rect 4276 23962 4300 23964
rect 4356 23962 4380 23964
rect 4436 23962 4460 23964
rect 4298 23910 4300 23962
rect 4362 23910 4374 23962
rect 4436 23910 4438 23962
rect 4276 23908 4300 23910
rect 4356 23908 4380 23910
rect 4436 23908 4460 23910
rect 4066 23896 4122 23905
rect 4220 23888 4516 23908
rect 4066 23831 4122 23840
rect 4220 22876 4516 22896
rect 4276 22874 4300 22876
rect 4356 22874 4380 22876
rect 4436 22874 4460 22876
rect 4298 22822 4300 22874
rect 4362 22822 4374 22874
rect 4436 22822 4438 22874
rect 4276 22820 4300 22822
rect 4356 22820 4380 22822
rect 4436 22820 4460 22822
rect 4220 22800 4516 22820
rect 5448 22160 5500 22166
rect 5448 22102 5500 22108
rect 4220 21788 4516 21808
rect 4276 21786 4300 21788
rect 4356 21786 4380 21788
rect 4436 21786 4460 21788
rect 4298 21734 4300 21786
rect 4362 21734 4374 21786
rect 4436 21734 4438 21786
rect 4276 21732 4300 21734
rect 4356 21732 4380 21734
rect 4436 21732 4460 21734
rect 4220 21712 4516 21732
rect 4220 20700 4516 20720
rect 4276 20698 4300 20700
rect 4356 20698 4380 20700
rect 4436 20698 4460 20700
rect 4298 20646 4300 20698
rect 4362 20646 4374 20698
rect 4436 20646 4438 20698
rect 4276 20644 4300 20646
rect 4356 20644 4380 20646
rect 4436 20644 4460 20646
rect 4220 20624 4516 20644
rect 5460 19922 5488 22102
rect 5448 19916 5500 19922
rect 5448 19858 5500 19864
rect 4712 19848 4764 19854
rect 4712 19790 4764 19796
rect 4896 19848 4948 19854
rect 4896 19790 4948 19796
rect 4220 19612 4516 19632
rect 4276 19610 4300 19612
rect 4356 19610 4380 19612
rect 4436 19610 4460 19612
rect 4298 19558 4300 19610
rect 4362 19558 4374 19610
rect 4436 19558 4438 19610
rect 4276 19556 4300 19558
rect 4356 19556 4380 19558
rect 4436 19556 4460 19558
rect 4220 19536 4516 19556
rect 4618 19408 4674 19417
rect 4618 19343 4674 19352
rect 4436 19168 4488 19174
rect 4434 19136 4436 19145
rect 4488 19136 4490 19145
rect 4434 19071 4490 19080
rect 4220 18524 4516 18544
rect 4276 18522 4300 18524
rect 4356 18522 4380 18524
rect 4436 18522 4460 18524
rect 4298 18470 4300 18522
rect 4362 18470 4374 18522
rect 4436 18470 4438 18522
rect 4276 18468 4300 18470
rect 4356 18468 4380 18470
rect 4436 18468 4460 18470
rect 4220 18448 4516 18468
rect 3882 18048 3938 18057
rect 3882 17983 3938 17992
rect 3240 16244 3292 16250
rect 3240 16186 3292 16192
rect 3422 15056 3478 15065
rect 3422 14991 3478 15000
rect 3330 13424 3386 13433
rect 3330 13359 3386 13368
rect 3344 11665 3372 13359
rect 3330 11656 3386 11665
rect 3330 11591 3386 11600
rect 3148 10056 3200 10062
rect 3146 10024 3148 10033
rect 3200 10024 3202 10033
rect 3146 9959 3202 9968
rect 2872 9648 2924 9654
rect 2872 9590 2924 9596
rect 3332 9648 3384 9654
rect 3332 9590 3384 9596
rect 2332 3318 2728 3346
rect 2332 800 2360 3318
rect 3344 950 3372 9590
rect 3436 4865 3464 14991
rect 3698 12336 3754 12345
rect 3698 12271 3754 12280
rect 3514 5128 3570 5137
rect 3514 5063 3570 5072
rect 3422 4856 3478 4865
rect 3422 4791 3478 4800
rect 3528 2802 3556 5063
rect 3712 3505 3740 12271
rect 3896 10305 3924 17983
rect 4220 17436 4516 17456
rect 4276 17434 4300 17436
rect 4356 17434 4380 17436
rect 4436 17434 4460 17436
rect 4298 17382 4300 17434
rect 4362 17382 4374 17434
rect 4436 17382 4438 17434
rect 4276 17380 4300 17382
rect 4356 17380 4380 17382
rect 4436 17380 4460 17382
rect 4220 17360 4516 17380
rect 4220 16348 4516 16368
rect 4276 16346 4300 16348
rect 4356 16346 4380 16348
rect 4436 16346 4460 16348
rect 4298 16294 4300 16346
rect 4362 16294 4374 16346
rect 4436 16294 4438 16346
rect 4276 16292 4300 16294
rect 4356 16292 4380 16294
rect 4436 16292 4460 16294
rect 4220 16272 4516 16292
rect 4220 15260 4516 15280
rect 4276 15258 4300 15260
rect 4356 15258 4380 15260
rect 4436 15258 4460 15260
rect 4298 15206 4300 15258
rect 4362 15206 4374 15258
rect 4436 15206 4438 15258
rect 4276 15204 4300 15206
rect 4356 15204 4380 15206
rect 4436 15204 4460 15206
rect 4220 15184 4516 15204
rect 4220 14172 4516 14192
rect 4276 14170 4300 14172
rect 4356 14170 4380 14172
rect 4436 14170 4460 14172
rect 4298 14118 4300 14170
rect 4362 14118 4374 14170
rect 4436 14118 4438 14170
rect 4276 14116 4300 14118
rect 4356 14116 4380 14118
rect 4436 14116 4460 14118
rect 4220 14096 4516 14116
rect 4220 13084 4516 13104
rect 4276 13082 4300 13084
rect 4356 13082 4380 13084
rect 4436 13082 4460 13084
rect 4298 13030 4300 13082
rect 4362 13030 4374 13082
rect 4436 13030 4438 13082
rect 4276 13028 4300 13030
rect 4356 13028 4380 13030
rect 4436 13028 4460 13030
rect 4220 13008 4516 13028
rect 4220 11996 4516 12016
rect 4276 11994 4300 11996
rect 4356 11994 4380 11996
rect 4436 11994 4460 11996
rect 4298 11942 4300 11994
rect 4362 11942 4374 11994
rect 4436 11942 4438 11994
rect 4276 11940 4300 11942
rect 4356 11940 4380 11942
rect 4436 11940 4460 11942
rect 4220 11920 4516 11940
rect 4220 10908 4516 10928
rect 4276 10906 4300 10908
rect 4356 10906 4380 10908
rect 4436 10906 4460 10908
rect 4298 10854 4300 10906
rect 4362 10854 4374 10906
rect 4436 10854 4438 10906
rect 4276 10852 4300 10854
rect 4356 10852 4380 10854
rect 4436 10852 4460 10854
rect 4220 10832 4516 10852
rect 3882 10296 3938 10305
rect 3882 10231 3938 10240
rect 4220 9820 4516 9840
rect 4276 9818 4300 9820
rect 4356 9818 4380 9820
rect 4436 9818 4460 9820
rect 4298 9766 4300 9818
rect 4362 9766 4374 9818
rect 4436 9766 4438 9818
rect 4276 9764 4300 9766
rect 4356 9764 4380 9766
rect 4436 9764 4460 9766
rect 4220 9744 4516 9764
rect 4220 8732 4516 8752
rect 4276 8730 4300 8732
rect 4356 8730 4380 8732
rect 4436 8730 4460 8732
rect 4298 8678 4300 8730
rect 4362 8678 4374 8730
rect 4436 8678 4438 8730
rect 4276 8676 4300 8678
rect 4356 8676 4380 8678
rect 4436 8676 4460 8678
rect 4220 8656 4516 8676
rect 4220 7644 4516 7664
rect 4276 7642 4300 7644
rect 4356 7642 4380 7644
rect 4436 7642 4460 7644
rect 4298 7590 4300 7642
rect 4362 7590 4374 7642
rect 4436 7590 4438 7642
rect 4276 7588 4300 7590
rect 4356 7588 4380 7590
rect 4436 7588 4460 7590
rect 4220 7568 4516 7588
rect 4632 7546 4660 19343
rect 4724 19174 4752 19790
rect 4908 19174 4936 19790
rect 6104 19417 6132 25638
rect 6288 21865 6316 46951
rect 6734 33824 6790 33833
rect 6734 33759 6790 33768
rect 6748 29850 6776 33759
rect 6932 32026 6960 63174
rect 7392 62257 7420 69799
rect 8404 67697 8432 79070
rect 8772 74769 8800 79200
rect 9402 74896 9458 74905
rect 9402 74831 9458 74840
rect 8758 74760 8814 74769
rect 8758 74695 8814 74704
rect 8942 72856 8998 72865
rect 8942 72791 8998 72800
rect 8390 67688 8446 67697
rect 8390 67623 8446 67632
rect 7378 62248 7434 62257
rect 7378 62183 7434 62192
rect 8758 49736 8814 49745
rect 8758 49671 8814 49680
rect 8772 45558 8800 49671
rect 8850 46200 8906 46209
rect 8850 46135 8852 46144
rect 8904 46135 8906 46144
rect 8852 46106 8904 46112
rect 8760 45552 8812 45558
rect 8760 45494 8812 45500
rect 8576 45348 8628 45354
rect 8576 45290 8628 45296
rect 8114 44976 8170 44985
rect 8114 44911 8170 44920
rect 8128 44538 8156 44911
rect 8116 44532 8168 44538
rect 8116 44474 8168 44480
rect 8300 44328 8352 44334
rect 8298 44296 8300 44305
rect 8352 44296 8354 44305
rect 8298 44231 8354 44240
rect 8312 43994 8340 44231
rect 8300 43988 8352 43994
rect 8300 43930 8352 43936
rect 8588 38706 8616 45290
rect 8772 45082 8800 45494
rect 8760 45076 8812 45082
rect 8760 45018 8812 45024
rect 8850 42392 8906 42401
rect 8850 42327 8906 42336
rect 8496 38678 8616 38706
rect 8496 34513 8524 38678
rect 8666 36544 8722 36553
rect 8666 36479 8722 36488
rect 8482 34504 8538 34513
rect 8482 34439 8538 34448
rect 8484 34400 8536 34406
rect 8484 34342 8536 34348
rect 7564 34060 7616 34066
rect 7564 34002 7616 34008
rect 7576 33658 7604 34002
rect 8496 33862 8524 34342
rect 8574 33960 8630 33969
rect 8574 33895 8630 33904
rect 8116 33856 8168 33862
rect 8484 33856 8536 33862
rect 8116 33798 8168 33804
rect 8482 33824 8484 33833
rect 8536 33824 8538 33833
rect 7564 33652 7616 33658
rect 7564 33594 7616 33600
rect 7932 33380 7984 33386
rect 7932 33322 7984 33328
rect 7746 32736 7802 32745
rect 7746 32671 7802 32680
rect 7760 32570 7788 32671
rect 7748 32564 7800 32570
rect 7748 32506 7800 32512
rect 7564 32224 7616 32230
rect 7564 32166 7616 32172
rect 6920 32020 6972 32026
rect 6920 31962 6972 31968
rect 7288 31952 7340 31958
rect 7576 31929 7604 32166
rect 7840 32020 7892 32026
rect 7840 31962 7892 31968
rect 7288 31894 7340 31900
rect 7562 31920 7618 31929
rect 7010 31240 7066 31249
rect 7010 31175 7066 31184
rect 7024 31142 7052 31175
rect 7012 31136 7064 31142
rect 7012 31078 7064 31084
rect 7024 30938 7052 31078
rect 7012 30932 7064 30938
rect 7012 30874 7064 30880
rect 6736 29844 6788 29850
rect 6736 29786 6788 29792
rect 7196 29708 7248 29714
rect 7196 29650 7248 29656
rect 6644 29640 6696 29646
rect 6644 29582 6696 29588
rect 6656 29306 6684 29582
rect 7208 29306 7236 29650
rect 6644 29300 6696 29306
rect 6644 29242 6696 29248
rect 7012 29300 7064 29306
rect 7012 29242 7064 29248
rect 7196 29300 7248 29306
rect 7196 29242 7248 29248
rect 6656 29102 6684 29242
rect 6644 29096 6696 29102
rect 6644 29038 6696 29044
rect 6920 29096 6972 29102
rect 6920 29038 6972 29044
rect 6932 28422 6960 29038
rect 6920 28416 6972 28422
rect 6920 28358 6972 28364
rect 6932 27554 6960 28358
rect 6840 27538 6960 27554
rect 6828 27532 6960 27538
rect 6880 27526 6960 27532
rect 6828 27474 6880 27480
rect 6932 27130 6960 27526
rect 6920 27124 6972 27130
rect 6920 27066 6972 27072
rect 7024 23866 7052 29242
rect 7300 29238 7328 31894
rect 7562 31855 7618 31864
rect 7576 31686 7604 31855
rect 7656 31816 7708 31822
rect 7654 31784 7656 31793
rect 7708 31784 7710 31793
rect 7654 31719 7710 31728
rect 7564 31680 7616 31686
rect 7564 31622 7616 31628
rect 7576 31346 7604 31622
rect 7852 31346 7880 31962
rect 7564 31340 7616 31346
rect 7564 31282 7616 31288
rect 7840 31340 7892 31346
rect 7840 31282 7892 31288
rect 7472 31136 7524 31142
rect 7470 31104 7472 31113
rect 7524 31104 7526 31113
rect 7470 31039 7526 31048
rect 7748 30932 7800 30938
rect 7748 30874 7800 30880
rect 7760 30841 7788 30874
rect 7746 30832 7802 30841
rect 7564 30796 7616 30802
rect 7746 30767 7802 30776
rect 7564 30738 7616 30744
rect 7576 30394 7604 30738
rect 7564 30388 7616 30394
rect 7564 30330 7616 30336
rect 7472 30048 7524 30054
rect 7576 30025 7604 30330
rect 7654 30288 7710 30297
rect 7654 30223 7656 30232
rect 7708 30223 7710 30232
rect 7656 30194 7708 30200
rect 7472 29990 7524 29996
rect 7562 30016 7618 30025
rect 7288 29232 7340 29238
rect 7288 29174 7340 29180
rect 7484 29170 7512 29990
rect 7562 29951 7618 29960
rect 7472 29164 7524 29170
rect 7472 29106 7524 29112
rect 7840 29096 7892 29102
rect 7840 29038 7892 29044
rect 7380 29028 7432 29034
rect 7380 28970 7432 28976
rect 7288 28416 7340 28422
rect 7288 28358 7340 28364
rect 7300 27946 7328 28358
rect 7288 27940 7340 27946
rect 7288 27882 7340 27888
rect 7104 27464 7156 27470
rect 7104 27406 7156 27412
rect 7392 27452 7420 28970
rect 7656 28960 7708 28966
rect 7562 28928 7618 28937
rect 7656 28902 7708 28908
rect 7562 28863 7618 28872
rect 7576 28694 7604 28863
rect 7564 28688 7616 28694
rect 7564 28630 7616 28636
rect 7472 27464 7524 27470
rect 7392 27424 7472 27452
rect 7116 26790 7144 27406
rect 7104 26784 7156 26790
rect 7102 26752 7104 26761
rect 7156 26752 7158 26761
rect 7102 26687 7158 26696
rect 7392 26586 7420 27424
rect 7472 27406 7524 27412
rect 7380 26580 7432 26586
rect 7380 26522 7432 26528
rect 7668 24206 7696 28902
rect 7852 28558 7880 29038
rect 7840 28552 7892 28558
rect 7840 28494 7892 28500
rect 7944 24410 7972 33322
rect 8128 33114 8156 33798
rect 8482 33759 8538 33768
rect 8484 33312 8536 33318
rect 8588 33300 8616 33895
rect 8536 33272 8616 33300
rect 8484 33254 8536 33260
rect 8116 33108 8168 33114
rect 8116 33050 8168 33056
rect 8128 32881 8156 33050
rect 8114 32872 8170 32881
rect 8114 32807 8170 32816
rect 8116 32224 8168 32230
rect 8116 32166 8168 32172
rect 8024 31816 8076 31822
rect 8024 31758 8076 31764
rect 8036 31113 8064 31758
rect 8022 31104 8078 31113
rect 8022 31039 8078 31048
rect 8128 30954 8156 32166
rect 8496 31482 8524 33254
rect 8576 32972 8628 32978
rect 8576 32914 8628 32920
rect 8588 32745 8616 32914
rect 8574 32736 8630 32745
rect 8574 32671 8630 32680
rect 8576 31884 8628 31890
rect 8576 31826 8628 31832
rect 8484 31476 8536 31482
rect 8484 31418 8536 31424
rect 8036 30926 8156 30954
rect 8588 30938 8616 31826
rect 8576 30932 8628 30938
rect 8036 29186 8064 30926
rect 8576 30874 8628 30880
rect 8116 30728 8168 30734
rect 8116 30670 8168 30676
rect 8128 30258 8156 30670
rect 8208 30660 8260 30666
rect 8208 30602 8260 30608
rect 8220 30258 8248 30602
rect 8300 30592 8352 30598
rect 8300 30534 8352 30540
rect 8484 30592 8536 30598
rect 8484 30534 8536 30540
rect 8116 30252 8168 30258
rect 8116 30194 8168 30200
rect 8208 30252 8260 30258
rect 8208 30194 8260 30200
rect 8128 29714 8156 30194
rect 8116 29708 8168 29714
rect 8116 29650 8168 29656
rect 8220 29345 8248 30194
rect 8312 30190 8340 30534
rect 8496 30190 8524 30534
rect 8300 30184 8352 30190
rect 8300 30126 8352 30132
rect 8484 30184 8536 30190
rect 8484 30126 8536 30132
rect 8312 29458 8340 30126
rect 8496 29782 8524 30126
rect 8484 29776 8536 29782
rect 8484 29718 8536 29724
rect 8312 29430 8524 29458
rect 8206 29336 8262 29345
rect 8496 29306 8524 29430
rect 8206 29271 8262 29280
rect 8484 29300 8536 29306
rect 8484 29242 8536 29248
rect 8206 29200 8262 29209
rect 8036 29158 8156 29186
rect 8024 29096 8076 29102
rect 8024 29038 8076 29044
rect 8036 28762 8064 29038
rect 8128 28937 8156 29158
rect 8206 29135 8262 29144
rect 8390 29200 8446 29209
rect 8390 29135 8446 29144
rect 8114 28928 8170 28937
rect 8114 28863 8170 28872
rect 8114 28792 8170 28801
rect 8024 28756 8076 28762
rect 8114 28727 8170 28736
rect 8220 28744 8248 29135
rect 8300 29028 8352 29034
rect 8300 28970 8352 28976
rect 8312 28937 8340 28970
rect 8404 28966 8432 29135
rect 8680 29050 8708 36479
rect 8758 33144 8814 33153
rect 8758 33079 8760 33088
rect 8812 33079 8814 33088
rect 8760 33050 8812 33056
rect 8758 32736 8814 32745
rect 8758 32671 8814 32680
rect 8772 31754 8800 32671
rect 8760 31748 8812 31754
rect 8760 31690 8812 31696
rect 8760 31476 8812 31482
rect 8760 31418 8812 31424
rect 8772 29170 8800 31418
rect 8760 29164 8812 29170
rect 8760 29106 8812 29112
rect 8484 29028 8536 29034
rect 8484 28970 8536 28976
rect 8576 29028 8628 29034
rect 8680 29022 8800 29050
rect 8576 28970 8628 28976
rect 8392 28960 8444 28966
rect 8298 28928 8354 28937
rect 8496 28937 8524 28970
rect 8392 28902 8444 28908
rect 8482 28928 8538 28937
rect 8298 28863 8354 28872
rect 8482 28863 8538 28872
rect 8484 28756 8536 28762
rect 8024 28698 8076 28704
rect 8024 28620 8076 28626
rect 8128 28608 8156 28727
rect 8220 28716 8340 28744
rect 8076 28580 8156 28608
rect 8206 28656 8262 28665
rect 8206 28591 8262 28600
rect 8024 28562 8076 28568
rect 8036 27878 8064 28562
rect 8024 27872 8076 27878
rect 8022 27840 8024 27849
rect 8076 27840 8078 27849
rect 8022 27775 8078 27784
rect 8220 26246 8248 28591
rect 8312 27674 8340 28716
rect 8484 28698 8536 28704
rect 8392 28552 8444 28558
rect 8392 28494 8444 28500
rect 8404 27946 8432 28494
rect 8496 28082 8524 28698
rect 8588 28150 8616 28970
rect 8668 28960 8720 28966
rect 8668 28902 8720 28908
rect 8680 28626 8708 28902
rect 8668 28620 8720 28626
rect 8668 28562 8720 28568
rect 8680 28218 8708 28562
rect 8668 28212 8720 28218
rect 8668 28154 8720 28160
rect 8576 28144 8628 28150
rect 8576 28086 8628 28092
rect 8484 28076 8536 28082
rect 8484 28018 8536 28024
rect 8392 27940 8444 27946
rect 8392 27882 8444 27888
rect 8300 27668 8352 27674
rect 8300 27610 8352 27616
rect 8404 27334 8432 27882
rect 8300 27328 8352 27334
rect 8300 27270 8352 27276
rect 8392 27328 8444 27334
rect 8392 27270 8444 27276
rect 8208 26240 8260 26246
rect 8208 26182 8260 26188
rect 7932 24404 7984 24410
rect 7932 24346 7984 24352
rect 7656 24200 7708 24206
rect 7656 24142 7708 24148
rect 7012 23860 7064 23866
rect 7012 23802 7064 23808
rect 7838 23760 7894 23769
rect 7838 23695 7894 23704
rect 6274 21856 6330 21865
rect 6274 21791 6330 21800
rect 7852 19990 7880 23695
rect 7840 19984 7892 19990
rect 7840 19926 7892 19932
rect 6090 19408 6146 19417
rect 6090 19343 6146 19352
rect 4712 19168 4764 19174
rect 4712 19110 4764 19116
rect 4896 19168 4948 19174
rect 4896 19110 4948 19116
rect 4908 17785 4936 19110
rect 4894 17776 4950 17785
rect 4894 17711 4950 17720
rect 4908 16969 4936 17711
rect 4894 16960 4950 16969
rect 4894 16895 4950 16904
rect 7944 16289 7972 24346
rect 8116 24268 8168 24274
rect 8116 24210 8168 24216
rect 8128 24041 8156 24210
rect 8114 24032 8170 24041
rect 8114 23967 8170 23976
rect 8128 23866 8156 23967
rect 8116 23860 8168 23866
rect 8116 23802 8168 23808
rect 7930 16280 7986 16289
rect 7930 16215 7986 16224
rect 8312 15178 8340 27270
rect 8668 26852 8720 26858
rect 8668 26794 8720 26800
rect 8484 26784 8536 26790
rect 8484 26726 8536 26732
rect 8496 26489 8524 26726
rect 8482 26480 8538 26489
rect 8680 26450 8708 26794
rect 8482 26415 8538 26424
rect 8668 26444 8720 26450
rect 8668 26386 8720 26392
rect 8680 26042 8708 26386
rect 8668 26036 8720 26042
rect 8668 25978 8720 25984
rect 8668 24608 8720 24614
rect 8668 24550 8720 24556
rect 8484 24200 8536 24206
rect 8484 24142 8536 24148
rect 8390 17776 8446 17785
rect 8390 17711 8446 17720
rect 8404 17338 8432 17711
rect 8392 17332 8444 17338
rect 8392 17274 8444 17280
rect 8220 15150 8340 15178
rect 4710 13832 4766 13841
rect 4710 13767 4766 13776
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 4066 6896 4122 6905
rect 4066 6831 4122 6840
rect 4080 6225 4108 6831
rect 4220 6556 4516 6576
rect 4276 6554 4300 6556
rect 4356 6554 4380 6556
rect 4436 6554 4460 6556
rect 4298 6502 4300 6554
rect 4362 6502 4374 6554
rect 4436 6502 4438 6554
rect 4276 6500 4300 6502
rect 4356 6500 4380 6502
rect 4436 6500 4460 6502
rect 4220 6480 4516 6500
rect 4066 6216 4122 6225
rect 4066 6151 4122 6160
rect 4220 5468 4516 5488
rect 4276 5466 4300 5468
rect 4356 5466 4380 5468
rect 4436 5466 4460 5468
rect 4298 5414 4300 5466
rect 4362 5414 4374 5466
rect 4436 5414 4438 5466
rect 4276 5412 4300 5414
rect 4356 5412 4380 5414
rect 4436 5412 4460 5414
rect 4220 5392 4516 5412
rect 4220 4380 4516 4400
rect 4276 4378 4300 4380
rect 4356 4378 4380 4380
rect 4436 4378 4460 4380
rect 4298 4326 4300 4378
rect 4362 4326 4374 4378
rect 4436 4326 4438 4378
rect 4276 4324 4300 4326
rect 4356 4324 4380 4326
rect 4436 4324 4460 4326
rect 4220 4304 4516 4324
rect 3698 3496 3754 3505
rect 3698 3431 3754 3440
rect 4220 3292 4516 3312
rect 4276 3290 4300 3292
rect 4356 3290 4380 3292
rect 4436 3290 4460 3292
rect 4298 3238 4300 3290
rect 4362 3238 4374 3290
rect 4436 3238 4438 3290
rect 4276 3236 4300 3238
rect 4356 3236 4380 3238
rect 4436 3236 4460 3238
rect 4220 3216 4516 3236
rect 3436 2774 3556 2802
rect 3240 944 3292 950
rect 3240 886 3292 892
rect 3332 944 3384 950
rect 3332 886 3384 892
rect 3252 800 3280 886
rect 18 0 74 800
rect 478 0 534 800
rect 1398 0 1454 800
rect 2318 0 2374 800
rect 3238 0 3294 800
rect 3436 785 3464 2774
rect 4220 2204 4516 2224
rect 4276 2202 4300 2204
rect 4356 2202 4380 2204
rect 4436 2202 4460 2204
rect 4298 2150 4300 2202
rect 4362 2150 4374 2202
rect 4436 2150 4438 2202
rect 4276 2148 4300 2150
rect 4356 2148 4380 2150
rect 4436 2148 4460 2150
rect 4220 2128 4516 2148
rect 4724 1986 4752 13767
rect 7102 10160 7158 10169
rect 7102 10095 7104 10104
rect 7156 10095 7158 10104
rect 7196 10124 7248 10130
rect 7104 10066 7156 10072
rect 7196 10066 7248 10072
rect 7116 9722 7144 10066
rect 7104 9716 7156 9722
rect 7104 9658 7156 9664
rect 7208 9382 7236 10066
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7208 8401 7236 9318
rect 7194 8392 7250 8401
rect 7194 8327 7250 8336
rect 5998 7576 6054 7585
rect 5080 7540 5132 7546
rect 5998 7511 6054 7520
rect 5080 7482 5132 7488
rect 4802 6216 4858 6225
rect 4802 6151 4858 6160
rect 4172 1958 4752 1986
rect 4172 800 4200 1958
rect 4816 1290 4844 6151
rect 4804 1284 4856 1290
rect 4804 1226 4856 1232
rect 5092 800 5120 7482
rect 6012 800 6040 7511
rect 7838 6352 7894 6361
rect 7838 6287 7894 6296
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 6932 800 6960 4082
rect 7852 800 7880 6287
rect 8220 4146 8248 15150
rect 8496 12458 8524 24142
rect 8680 23594 8708 24550
rect 8772 24206 8800 29022
rect 8760 24200 8812 24206
rect 8760 24142 8812 24148
rect 8668 23588 8720 23594
rect 8668 23530 8720 23536
rect 8864 22001 8892 42327
rect 8956 41857 8984 72791
rect 9416 60790 9444 74831
rect 9692 74798 9720 79200
rect 10612 75313 10640 79200
rect 10598 75304 10654 75313
rect 10598 75239 10654 75248
rect 9680 74792 9732 74798
rect 10876 74792 10928 74798
rect 9680 74734 9732 74740
rect 10414 74760 10470 74769
rect 10876 74734 10928 74740
rect 10414 74695 10470 74704
rect 9404 60784 9456 60790
rect 9404 60726 9456 60732
rect 9496 60648 9548 60654
rect 9218 60616 9274 60625
rect 9496 60590 9548 60596
rect 9218 60551 9274 60560
rect 9128 57928 9180 57934
rect 9128 57870 9180 57876
rect 9140 48346 9168 57870
rect 9128 48340 9180 48346
rect 9128 48282 9180 48288
rect 9128 45416 9180 45422
rect 9128 45358 9180 45364
rect 9140 43761 9168 45358
rect 9126 43752 9182 43761
rect 9126 43687 9182 43696
rect 8942 41848 8998 41857
rect 8942 41783 8998 41792
rect 9034 36952 9090 36961
rect 9034 36887 9090 36896
rect 8942 35184 8998 35193
rect 8942 35119 8998 35128
rect 8956 34746 8984 35119
rect 8944 34740 8996 34746
rect 8944 34682 8996 34688
rect 9048 33046 9076 36887
rect 9232 34746 9260 60551
rect 9508 57934 9536 60590
rect 9496 57928 9548 57934
rect 9496 57870 9548 57876
rect 9954 53136 10010 53145
rect 9954 53071 10010 53080
rect 9968 52562 9996 53071
rect 9956 52556 10008 52562
rect 9956 52498 10008 52504
rect 9968 52154 9996 52498
rect 9956 52148 10008 52154
rect 9956 52090 10008 52096
rect 9404 48340 9456 48346
rect 9404 48282 9456 48288
rect 9416 43602 9444 48282
rect 9680 46164 9732 46170
rect 9680 46106 9732 46112
rect 9692 45422 9720 46106
rect 9864 45484 9916 45490
rect 9864 45426 9916 45432
rect 9680 45416 9732 45422
rect 9876 45393 9904 45426
rect 9680 45358 9732 45364
rect 9862 45384 9918 45393
rect 9862 45319 9918 45328
rect 9416 43574 9536 43602
rect 9402 39400 9458 39409
rect 9402 39335 9458 39344
rect 9416 39098 9444 39335
rect 9404 39092 9456 39098
rect 9404 39034 9456 39040
rect 9404 38888 9456 38894
rect 9404 38830 9456 38836
rect 9416 37330 9444 38830
rect 9404 37324 9456 37330
rect 9404 37266 9456 37272
rect 9310 36408 9366 36417
rect 9310 36343 9366 36352
rect 9220 34740 9272 34746
rect 9220 34682 9272 34688
rect 9220 34536 9272 34542
rect 9220 34478 9272 34484
rect 9232 33862 9260 34478
rect 9220 33856 9272 33862
rect 9220 33798 9272 33804
rect 9036 33040 9088 33046
rect 9036 32982 9088 32988
rect 9048 32366 9076 32982
rect 9232 32910 9260 33798
rect 9220 32904 9272 32910
rect 9220 32846 9272 32852
rect 9218 32600 9274 32609
rect 9218 32535 9220 32544
rect 9272 32535 9274 32544
rect 9220 32506 9272 32512
rect 9324 32434 9352 36343
rect 9416 34950 9444 37266
rect 9404 34944 9456 34950
rect 9404 34886 9456 34892
rect 9416 34542 9444 34886
rect 9404 34536 9456 34542
rect 9404 34478 9456 34484
rect 9402 33824 9458 33833
rect 9402 33759 9458 33768
rect 9416 33658 9444 33759
rect 9404 33652 9456 33658
rect 9404 33594 9456 33600
rect 9508 33538 9536 43574
rect 10324 41608 10376 41614
rect 10324 41550 10376 41556
rect 10336 40934 10364 41550
rect 10324 40928 10376 40934
rect 10324 40870 10376 40876
rect 9680 40112 9732 40118
rect 9680 40054 9732 40060
rect 9692 38894 9720 40054
rect 10230 39944 10286 39953
rect 10230 39879 10286 39888
rect 9680 38888 9732 38894
rect 9680 38830 9732 38836
rect 10140 36576 10192 36582
rect 10140 36518 10192 36524
rect 10152 35494 10180 36518
rect 10140 35488 10192 35494
rect 10140 35430 10192 35436
rect 10152 34921 10180 35430
rect 10138 34912 10194 34921
rect 10138 34847 10194 34856
rect 10046 34776 10102 34785
rect 10046 34711 10102 34720
rect 9588 33856 9640 33862
rect 9588 33798 9640 33804
rect 9956 33856 10008 33862
rect 9956 33798 10008 33804
rect 9600 33561 9628 33798
rect 9416 33510 9536 33538
rect 9586 33552 9642 33561
rect 9312 32428 9364 32434
rect 9312 32370 9364 32376
rect 9036 32360 9088 32366
rect 9036 32302 9088 32308
rect 9048 32026 9076 32302
rect 9036 32020 9088 32026
rect 9036 31962 9088 31968
rect 8944 31816 8996 31822
rect 8944 31758 8996 31764
rect 8956 28762 8984 31758
rect 9036 31136 9088 31142
rect 9036 31078 9088 31084
rect 8944 28756 8996 28762
rect 8944 28698 8996 28704
rect 8942 28656 8998 28665
rect 8942 28591 8944 28600
rect 8996 28591 8998 28600
rect 8944 28562 8996 28568
rect 8956 28014 8984 28562
rect 8944 28008 8996 28014
rect 8942 27976 8944 27985
rect 8996 27976 8998 27985
rect 8942 27911 8998 27920
rect 8956 27885 8984 27911
rect 8944 27328 8996 27334
rect 8944 27270 8996 27276
rect 8956 23769 8984 27270
rect 8942 23760 8998 23769
rect 8942 23695 8998 23704
rect 8850 21992 8906 22001
rect 8850 21927 8906 21936
rect 9048 19961 9076 31078
rect 9128 30796 9180 30802
rect 9128 30738 9180 30744
rect 9140 30666 9168 30738
rect 9128 30660 9180 30666
rect 9128 30602 9180 30608
rect 9140 30394 9168 30602
rect 9312 30592 9364 30598
rect 9312 30534 9364 30540
rect 9128 30388 9180 30394
rect 9128 30330 9180 30336
rect 9220 30116 9272 30122
rect 9220 30058 9272 30064
rect 9126 29744 9182 29753
rect 9126 29679 9128 29688
rect 9180 29679 9182 29688
rect 9128 29650 9180 29656
rect 9140 28694 9168 29650
rect 9232 29306 9260 30058
rect 9324 29306 9352 30534
rect 9220 29300 9272 29306
rect 9220 29242 9272 29248
rect 9312 29300 9364 29306
rect 9312 29242 9364 29248
rect 9220 29096 9272 29102
rect 9220 29038 9272 29044
rect 9128 28688 9180 28694
rect 9128 28630 9180 28636
rect 9126 28248 9182 28257
rect 9126 28183 9182 28192
rect 9140 28082 9168 28183
rect 9128 28076 9180 28082
rect 9128 28018 9180 28024
rect 9128 27464 9180 27470
rect 9128 27406 9180 27412
rect 9140 27033 9168 27406
rect 9126 27024 9182 27033
rect 9126 26959 9182 26968
rect 9232 25906 9260 29038
rect 9220 25900 9272 25906
rect 9220 25842 9272 25848
rect 9232 25498 9260 25842
rect 9324 25537 9352 29242
rect 9310 25528 9366 25537
rect 9220 25492 9272 25498
rect 9310 25463 9366 25472
rect 9220 25434 9272 25440
rect 9232 24410 9260 25434
rect 9220 24404 9272 24410
rect 9220 24346 9272 24352
rect 9034 19952 9090 19961
rect 9034 19887 9090 19896
rect 8404 12430 8524 12458
rect 8298 9072 8354 9081
rect 8298 9007 8354 9016
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8312 800 8340 9007
rect 8404 4146 8432 12430
rect 9416 10198 9444 33510
rect 9586 33487 9642 33496
rect 9588 33448 9640 33454
rect 9588 33390 9640 33396
rect 9600 33114 9628 33390
rect 9968 33318 9996 33798
rect 10060 33658 10088 34711
rect 10048 33652 10100 33658
rect 10048 33594 10100 33600
rect 10060 33386 10088 33594
rect 10048 33380 10100 33386
rect 10048 33322 10100 33328
rect 9956 33312 10008 33318
rect 10152 33266 10180 34847
rect 9956 33254 10008 33260
rect 9588 33108 9640 33114
rect 9588 33050 9640 33056
rect 9862 33008 9918 33017
rect 9862 32943 9918 32952
rect 9876 32910 9904 32943
rect 9680 32904 9732 32910
rect 9864 32904 9916 32910
rect 9732 32852 9812 32858
rect 9680 32846 9812 32852
rect 9864 32846 9916 32852
rect 9692 32830 9812 32846
rect 9586 32600 9642 32609
rect 9586 32535 9642 32544
rect 9600 32042 9628 32535
rect 9680 32360 9732 32366
rect 9680 32302 9732 32308
rect 9692 32201 9720 32302
rect 9678 32192 9734 32201
rect 9678 32127 9734 32136
rect 9600 32014 9720 32042
rect 9496 31748 9548 31754
rect 9496 31690 9548 31696
rect 9508 31521 9536 31690
rect 9494 31512 9550 31521
rect 9494 31447 9550 31456
rect 9588 31136 9640 31142
rect 9588 31078 9640 31084
rect 9600 30938 9628 31078
rect 9588 30932 9640 30938
rect 9588 30874 9640 30880
rect 9494 30696 9550 30705
rect 9494 30631 9550 30640
rect 9508 29850 9536 30631
rect 9600 30569 9628 30874
rect 9586 30560 9642 30569
rect 9586 30495 9642 30504
rect 9692 30394 9720 32014
rect 9784 31906 9812 32830
rect 9876 32570 9904 32846
rect 9864 32564 9916 32570
rect 9864 32506 9916 32512
rect 9862 31920 9918 31929
rect 9784 31878 9862 31906
rect 9862 31855 9918 31864
rect 9876 31822 9904 31855
rect 9772 31816 9824 31822
rect 9772 31758 9824 31764
rect 9864 31816 9916 31822
rect 9864 31758 9916 31764
rect 9680 30388 9732 30394
rect 9680 30330 9732 30336
rect 9588 30320 9640 30326
rect 9588 30262 9640 30268
rect 9496 29844 9548 29850
rect 9496 29786 9548 29792
rect 9600 29345 9628 30262
rect 9680 30048 9732 30054
rect 9680 29990 9732 29996
rect 9586 29336 9642 29345
rect 9586 29271 9642 29280
rect 9600 29238 9628 29271
rect 9588 29232 9640 29238
rect 9588 29174 9640 29180
rect 9692 28801 9720 29990
rect 9784 29714 9812 31758
rect 9772 29708 9824 29714
rect 9772 29650 9824 29656
rect 9784 29306 9812 29650
rect 9772 29300 9824 29306
rect 9772 29242 9824 29248
rect 9678 28792 9734 28801
rect 9678 28727 9734 28736
rect 9784 28626 9812 29242
rect 9772 28620 9824 28626
rect 9772 28562 9824 28568
rect 9494 28384 9550 28393
rect 9494 28319 9550 28328
rect 9508 28218 9536 28319
rect 9496 28212 9548 28218
rect 9496 28154 9548 28160
rect 9588 28076 9640 28082
rect 9588 28018 9640 28024
rect 9600 27130 9628 28018
rect 9876 27962 9904 31758
rect 9968 31142 9996 33254
rect 10060 33238 10180 33266
rect 9956 31136 10008 31142
rect 9956 31078 10008 31084
rect 9956 30388 10008 30394
rect 9956 30330 10008 30336
rect 9968 29481 9996 30330
rect 9954 29472 10010 29481
rect 9954 29407 10010 29416
rect 9692 27934 9904 27962
rect 9588 27124 9640 27130
rect 9588 27066 9640 27072
rect 9496 26444 9548 26450
rect 9496 26386 9548 26392
rect 9508 25498 9536 26386
rect 9692 26382 9720 27934
rect 9864 27872 9916 27878
rect 9864 27814 9916 27820
rect 9876 27713 9904 27814
rect 9862 27704 9918 27713
rect 9862 27639 9918 27648
rect 9784 26858 9996 26874
rect 9772 26852 9996 26858
rect 9824 26846 9996 26852
rect 9772 26794 9824 26800
rect 9968 26790 9996 26846
rect 9864 26784 9916 26790
rect 9864 26726 9916 26732
rect 9956 26784 10008 26790
rect 9956 26726 10008 26732
rect 9680 26376 9732 26382
rect 9876 26353 9904 26726
rect 9680 26318 9732 26324
rect 9862 26344 9918 26353
rect 9692 25838 9720 26318
rect 9862 26279 9918 26288
rect 9680 25832 9732 25838
rect 9680 25774 9732 25780
rect 9496 25492 9548 25498
rect 9496 25434 9548 25440
rect 9680 25288 9732 25294
rect 9678 25256 9680 25265
rect 9732 25256 9734 25265
rect 9678 25191 9734 25200
rect 10060 24818 10088 33238
rect 10140 32292 10192 32298
rect 10140 32234 10192 32240
rect 10152 32026 10180 32234
rect 10140 32020 10192 32026
rect 10140 31962 10192 31968
rect 10244 31958 10272 39879
rect 10232 31952 10284 31958
rect 10232 31894 10284 31900
rect 10232 31136 10284 31142
rect 10232 31078 10284 31084
rect 10244 30666 10272 31078
rect 10232 30660 10284 30666
rect 10232 30602 10284 30608
rect 10244 29306 10272 30602
rect 10324 30048 10376 30054
rect 10324 29990 10376 29996
rect 10232 29300 10284 29306
rect 10232 29242 10284 29248
rect 10336 29102 10364 29990
rect 10324 29096 10376 29102
rect 10324 29038 10376 29044
rect 10322 28520 10378 28529
rect 10322 28455 10378 28464
rect 10336 28218 10364 28455
rect 10324 28212 10376 28218
rect 10324 28154 10376 28160
rect 10230 27840 10286 27849
rect 10230 27775 10286 27784
rect 10140 27464 10192 27470
rect 10138 27432 10140 27441
rect 10192 27432 10194 27441
rect 10138 27367 10194 27376
rect 10140 26920 10192 26926
rect 10140 26862 10192 26868
rect 10152 26586 10180 26862
rect 10140 26580 10192 26586
rect 10140 26522 10192 26528
rect 10048 24812 10100 24818
rect 10048 24754 10100 24760
rect 10048 24404 10100 24410
rect 10048 24346 10100 24352
rect 9588 24200 9640 24206
rect 9588 24142 9640 24148
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9508 16182 9536 16934
rect 9496 16176 9548 16182
rect 9496 16118 9548 16124
rect 9404 10192 9456 10198
rect 9404 10134 9456 10140
rect 9600 4321 9628 24142
rect 9680 23724 9732 23730
rect 9680 23666 9732 23672
rect 9692 23526 9720 23666
rect 9864 23588 9916 23594
rect 9864 23530 9916 23536
rect 9680 23520 9732 23526
rect 9680 23462 9732 23468
rect 9692 23361 9720 23462
rect 9678 23352 9734 23361
rect 9678 23287 9734 23296
rect 9876 22166 9904 23530
rect 10060 22273 10088 24346
rect 10046 22264 10102 22273
rect 10046 22199 10102 22208
rect 9864 22160 9916 22166
rect 9864 22102 9916 22108
rect 9876 18290 9904 22102
rect 10152 22098 10180 26522
rect 10244 25362 10272 27775
rect 10428 26994 10456 74695
rect 10690 69728 10746 69737
rect 10690 69663 10746 69672
rect 10506 59936 10562 59945
rect 10506 59871 10562 59880
rect 10520 41614 10548 59871
rect 10508 41608 10560 41614
rect 10508 41550 10560 41556
rect 10520 41274 10548 41550
rect 10508 41268 10560 41274
rect 10508 41210 10560 41216
rect 10600 36576 10652 36582
rect 10600 36518 10652 36524
rect 10612 34202 10640 36518
rect 10600 34196 10652 34202
rect 10600 34138 10652 34144
rect 10612 34105 10640 34138
rect 10598 34096 10654 34105
rect 10598 34031 10654 34040
rect 10506 33688 10562 33697
rect 10506 33623 10562 33632
rect 10520 33454 10548 33623
rect 10508 33448 10560 33454
rect 10508 33390 10560 33396
rect 10600 32020 10652 32026
rect 10600 31962 10652 31968
rect 10612 31657 10640 31962
rect 10598 31648 10654 31657
rect 10598 31583 10654 31592
rect 10508 31204 10560 31210
rect 10508 31146 10560 31152
rect 10520 29306 10548 31146
rect 10600 30252 10652 30258
rect 10600 30194 10652 30200
rect 10508 29300 10560 29306
rect 10508 29242 10560 29248
rect 10612 29170 10640 30194
rect 10600 29164 10652 29170
rect 10600 29106 10652 29112
rect 10598 28928 10654 28937
rect 10598 28863 10654 28872
rect 10612 28762 10640 28863
rect 10600 28756 10652 28762
rect 10600 28698 10652 28704
rect 10506 28656 10562 28665
rect 10506 28591 10562 28600
rect 10520 28218 10548 28591
rect 10508 28212 10560 28218
rect 10508 28154 10560 28160
rect 10508 27600 10560 27606
rect 10506 27568 10508 27577
rect 10560 27568 10562 27577
rect 10506 27503 10562 27512
rect 10600 27532 10652 27538
rect 10600 27474 10652 27480
rect 10416 26988 10468 26994
rect 10416 26930 10468 26936
rect 10324 26852 10376 26858
rect 10324 26794 10376 26800
rect 10336 26314 10364 26794
rect 10612 26790 10640 27474
rect 10600 26784 10652 26790
rect 10600 26726 10652 26732
rect 10508 26376 10560 26382
rect 10508 26318 10560 26324
rect 10324 26308 10376 26314
rect 10324 26250 10376 26256
rect 10232 25356 10284 25362
rect 10232 25298 10284 25304
rect 10244 24410 10272 25298
rect 10520 24410 10548 26318
rect 10600 25696 10652 25702
rect 10600 25638 10652 25644
rect 10612 25430 10640 25638
rect 10600 25424 10652 25430
rect 10600 25366 10652 25372
rect 10612 24886 10640 25366
rect 10600 24880 10652 24886
rect 10600 24822 10652 24828
rect 10232 24404 10284 24410
rect 10232 24346 10284 24352
rect 10508 24404 10560 24410
rect 10508 24346 10560 24352
rect 10600 23112 10652 23118
rect 10600 23054 10652 23060
rect 10140 22092 10192 22098
rect 10140 22034 10192 22040
rect 9864 18284 9916 18290
rect 9864 18226 9916 18232
rect 9680 18080 9732 18086
rect 9680 18022 9732 18028
rect 9692 17921 9720 18022
rect 9678 17912 9734 17921
rect 9876 17882 9904 18226
rect 9678 17847 9734 17856
rect 9864 17876 9916 17882
rect 9864 17818 9916 17824
rect 9876 17542 9904 17818
rect 9864 17536 9916 17542
rect 9864 17478 9916 17484
rect 10230 16280 10286 16289
rect 10230 16215 10286 16224
rect 10244 16046 10272 16215
rect 10232 16040 10284 16046
rect 10232 15982 10284 15988
rect 10612 15065 10640 23054
rect 10598 15056 10654 15065
rect 10598 14991 10654 15000
rect 9586 4312 9642 4321
rect 9586 4247 9642 4256
rect 10704 4146 10732 69663
rect 10888 67289 10916 74734
rect 11532 70553 11560 79200
rect 12346 75440 12402 75449
rect 12346 75375 12402 75384
rect 11518 70544 11574 70553
rect 11518 70479 11574 70488
rect 12360 68377 12388 75375
rect 12346 68368 12402 68377
rect 12346 68303 12402 68312
rect 11242 67688 11298 67697
rect 11242 67623 11298 67632
rect 10874 67280 10930 67289
rect 10874 67215 10930 67224
rect 10782 62112 10838 62121
rect 10782 62047 10838 62056
rect 10796 61062 10824 62047
rect 10966 61568 11022 61577
rect 10966 61503 11022 61512
rect 10980 61266 11008 61503
rect 10968 61260 11020 61266
rect 10968 61202 11020 61208
rect 10784 61056 10836 61062
rect 10784 60998 10836 61004
rect 10796 57633 10824 60998
rect 10980 60858 11008 61202
rect 10968 60852 11020 60858
rect 10968 60794 11020 60800
rect 10782 57624 10838 57633
rect 10782 57559 10838 57568
rect 10796 52562 10824 57559
rect 10784 52556 10836 52562
rect 10784 52498 10836 52504
rect 10796 52154 10824 52498
rect 10784 52148 10836 52154
rect 10784 52090 10836 52096
rect 10968 48204 11020 48210
rect 10968 48146 11020 48152
rect 10980 47802 11008 48146
rect 10968 47796 11020 47802
rect 10968 47738 11020 47744
rect 10968 44260 11020 44266
rect 11020 44220 11192 44248
rect 10968 44202 11020 44208
rect 11164 43790 11192 44220
rect 11152 43784 11204 43790
rect 11152 43726 11204 43732
rect 11164 43450 11192 43726
rect 11152 43444 11204 43450
rect 11152 43386 11204 43392
rect 11152 38752 11204 38758
rect 11152 38694 11204 38700
rect 11060 38208 11112 38214
rect 11060 38150 11112 38156
rect 11072 37330 11100 38150
rect 11060 37324 11112 37330
rect 11060 37266 11112 37272
rect 11072 36922 11100 37266
rect 11060 36916 11112 36922
rect 11060 36858 11112 36864
rect 10966 36680 11022 36689
rect 10966 36615 11022 36624
rect 10980 36378 11008 36615
rect 10968 36372 11020 36378
rect 10968 36314 11020 36320
rect 11060 36236 11112 36242
rect 11060 36178 11112 36184
rect 10782 35864 10838 35873
rect 11072 35834 11100 36178
rect 10782 35799 10784 35808
rect 10836 35799 10838 35808
rect 11060 35828 11112 35834
rect 10784 35770 10836 35776
rect 11060 35770 11112 35776
rect 10966 35728 11022 35737
rect 10966 35663 10968 35672
rect 11020 35663 11022 35672
rect 11060 35692 11112 35698
rect 10968 35634 11020 35640
rect 11060 35634 11112 35640
rect 10876 34468 10928 34474
rect 10876 34410 10928 34416
rect 10784 33448 10836 33454
rect 10784 33390 10836 33396
rect 10796 32178 10824 33390
rect 10888 32609 10916 34410
rect 10968 34196 11020 34202
rect 10968 34138 11020 34144
rect 10980 33969 11008 34138
rect 11072 34134 11100 35634
rect 11164 35193 11192 38694
rect 11150 35184 11206 35193
rect 11150 35119 11206 35128
rect 11060 34128 11112 34134
rect 11060 34070 11112 34076
rect 10966 33960 11022 33969
rect 10966 33895 11022 33904
rect 11072 33454 11100 34070
rect 11152 34060 11204 34066
rect 11152 34002 11204 34008
rect 11060 33448 11112 33454
rect 11060 33390 11112 33396
rect 11164 33300 11192 34002
rect 11072 33272 11192 33300
rect 11072 33114 11100 33272
rect 11060 33108 11112 33114
rect 11060 33050 11112 33056
rect 10968 32972 11020 32978
rect 10968 32914 11020 32920
rect 10874 32600 10930 32609
rect 10874 32535 10930 32544
rect 10980 32473 11008 32914
rect 11072 32881 11100 33050
rect 11150 33008 11206 33017
rect 11150 32943 11206 32952
rect 11058 32872 11114 32881
rect 11058 32807 11114 32816
rect 10966 32464 11022 32473
rect 10966 32399 10968 32408
rect 11020 32399 11022 32408
rect 10968 32370 11020 32376
rect 11060 32360 11112 32366
rect 10874 32328 10930 32337
rect 11060 32302 11112 32308
rect 10874 32263 10876 32272
rect 10928 32263 10930 32272
rect 10876 32234 10928 32240
rect 10796 32150 10916 32178
rect 10784 31816 10836 31822
rect 10784 31758 10836 31764
rect 10796 31249 10824 31758
rect 10888 31414 10916 32150
rect 10968 31816 11020 31822
rect 10968 31758 11020 31764
rect 10876 31408 10928 31414
rect 10876 31350 10928 31356
rect 10980 31346 11008 31758
rect 11072 31498 11100 32302
rect 11164 31890 11192 32943
rect 11152 31884 11204 31890
rect 11152 31826 11204 31832
rect 11164 31686 11192 31826
rect 11152 31680 11204 31686
rect 11152 31622 11204 31628
rect 11072 31470 11192 31498
rect 10968 31340 11020 31346
rect 10968 31282 11020 31288
rect 11060 31340 11112 31346
rect 11060 31282 11112 31288
rect 10782 31240 10838 31249
rect 10782 31175 10838 31184
rect 10968 31136 11020 31142
rect 10966 31104 10968 31113
rect 11020 31104 11022 31113
rect 10966 31039 11022 31048
rect 10784 30932 10836 30938
rect 10784 30874 10836 30880
rect 10796 30122 10824 30874
rect 10876 30796 10928 30802
rect 10876 30738 10928 30744
rect 10888 30161 10916 30738
rect 10980 30598 11008 31039
rect 10968 30592 11020 30598
rect 10968 30534 11020 30540
rect 10980 30433 11008 30534
rect 10966 30424 11022 30433
rect 10966 30359 11022 30368
rect 10874 30152 10930 30161
rect 10784 30116 10836 30122
rect 10874 30087 10930 30096
rect 10784 30058 10836 30064
rect 10888 29850 10916 30087
rect 10968 30048 11020 30054
rect 10968 29990 11020 29996
rect 10980 29889 11008 29990
rect 10966 29880 11022 29889
rect 10876 29844 10928 29850
rect 11072 29850 11100 31282
rect 10966 29815 11022 29824
rect 11060 29844 11112 29850
rect 10876 29786 10928 29792
rect 11060 29786 11112 29792
rect 11060 29708 11112 29714
rect 11060 29650 11112 29656
rect 10966 29608 11022 29617
rect 10966 29543 10968 29552
rect 11020 29543 11022 29552
rect 10968 29514 11020 29520
rect 10876 29504 10928 29510
rect 10876 29446 10928 29452
rect 10888 29209 10916 29446
rect 10874 29200 10930 29209
rect 10874 29135 10930 29144
rect 10876 29096 10928 29102
rect 10874 29064 10876 29073
rect 10928 29064 10930 29073
rect 11072 29034 11100 29650
rect 10874 28999 10930 29008
rect 11060 29028 11112 29034
rect 11060 28970 11112 28976
rect 11164 28914 11192 31470
rect 11256 30938 11284 67623
rect 12256 55820 12308 55826
rect 12256 55762 12308 55768
rect 12268 55457 12296 55762
rect 12452 55706 12480 79200
rect 13372 75857 13400 79200
rect 13358 75848 13414 75857
rect 13358 75783 13414 75792
rect 14292 73953 14320 79200
rect 15212 74798 15240 79200
rect 16132 77042 16160 79200
rect 16592 79098 16620 79200
rect 16592 79070 17080 79098
rect 16120 77036 16172 77042
rect 16120 76978 16172 76984
rect 15476 76968 15528 76974
rect 15476 76910 15528 76916
rect 15488 76430 15516 76910
rect 15476 76424 15528 76430
rect 15476 76366 15528 76372
rect 16394 75848 16450 75857
rect 16394 75783 16450 75792
rect 15200 74792 15252 74798
rect 15200 74734 15252 74740
rect 14278 73944 14334 73953
rect 14278 73879 14334 73888
rect 15382 73808 15438 73817
rect 15382 73743 15438 73752
rect 14094 71904 14150 71913
rect 14094 71839 14150 71848
rect 12622 67824 12678 67833
rect 12622 67759 12678 67768
rect 12360 55678 12480 55706
rect 12254 55448 12310 55457
rect 12254 55383 12256 55392
rect 12308 55383 12310 55392
rect 12256 55354 12308 55360
rect 12360 55282 12388 55678
rect 12440 55616 12492 55622
rect 12440 55558 12492 55564
rect 12348 55276 12400 55282
rect 12348 55218 12400 55224
rect 12452 54126 12480 55558
rect 12532 55276 12584 55282
rect 12532 55218 12584 55224
rect 12440 54120 12492 54126
rect 12440 54062 12492 54068
rect 11888 52488 11940 52494
rect 11888 52430 11940 52436
rect 11900 50561 11928 52430
rect 11886 50552 11942 50561
rect 11886 50487 11942 50496
rect 11610 49600 11666 49609
rect 11610 49535 11666 49544
rect 11624 48278 11652 49535
rect 11612 48272 11664 48278
rect 11612 48214 11664 48220
rect 12256 48204 12308 48210
rect 12256 48146 12308 48152
rect 12164 48136 12216 48142
rect 12164 48078 12216 48084
rect 11428 48000 11480 48006
rect 11428 47942 11480 47948
rect 11440 47122 11468 47942
rect 12176 47734 12204 48078
rect 12164 47728 12216 47734
rect 12164 47670 12216 47676
rect 12268 47258 12296 48146
rect 12256 47252 12308 47258
rect 12256 47194 12308 47200
rect 11428 47116 11480 47122
rect 11428 47058 11480 47064
rect 11440 46374 11468 47058
rect 11704 47048 11756 47054
rect 11704 46990 11756 46996
rect 11716 46714 11744 46990
rect 11704 46708 11756 46714
rect 11704 46650 11756 46656
rect 11716 46510 11744 46650
rect 11704 46504 11756 46510
rect 11704 46446 11756 46452
rect 12440 46504 12492 46510
rect 12440 46446 12492 46452
rect 11428 46368 11480 46374
rect 11426 46336 11428 46345
rect 12348 46368 12400 46374
rect 11480 46336 11482 46345
rect 12348 46310 12400 46316
rect 11426 46271 11482 46280
rect 12256 44328 12308 44334
rect 12256 44270 12308 44276
rect 11796 44192 11848 44198
rect 11796 44134 11848 44140
rect 11336 43852 11388 43858
rect 11336 43794 11388 43800
rect 11348 43450 11376 43794
rect 11336 43444 11388 43450
rect 11336 43386 11388 43392
rect 11612 41472 11664 41478
rect 11612 41414 11664 41420
rect 11336 40928 11388 40934
rect 11336 40870 11388 40876
rect 11348 40526 11376 40870
rect 11624 40610 11652 41414
rect 11532 40582 11652 40610
rect 11336 40520 11388 40526
rect 11336 40462 11388 40468
rect 11348 40118 11376 40462
rect 11336 40112 11388 40118
rect 11336 40054 11388 40060
rect 11336 38344 11388 38350
rect 11336 38286 11388 38292
rect 11348 37369 11376 38286
rect 11334 37360 11390 37369
rect 11334 37295 11390 37304
rect 11428 36848 11480 36854
rect 11428 36790 11480 36796
rect 11334 36272 11390 36281
rect 11440 36242 11468 36790
rect 11334 36207 11390 36216
rect 11428 36236 11480 36242
rect 11348 35290 11376 36207
rect 11428 36178 11480 36184
rect 11428 36032 11480 36038
rect 11428 35974 11480 35980
rect 11440 35834 11468 35974
rect 11428 35828 11480 35834
rect 11428 35770 11480 35776
rect 11336 35284 11388 35290
rect 11336 35226 11388 35232
rect 11348 32858 11376 35226
rect 11532 33946 11560 40582
rect 11612 40520 11664 40526
rect 11612 40462 11664 40468
rect 11624 39846 11652 40462
rect 11612 39840 11664 39846
rect 11612 39782 11664 39788
rect 11808 38570 11836 44134
rect 12268 43790 12296 44270
rect 12256 43784 12308 43790
rect 12256 43726 12308 43732
rect 12164 42288 12216 42294
rect 12164 42230 12216 42236
rect 11716 38542 11836 38570
rect 11716 35816 11744 38542
rect 12176 38486 12204 42230
rect 12268 40905 12296 43726
rect 12254 40896 12310 40905
rect 12254 40831 12310 40840
rect 12164 38480 12216 38486
rect 12164 38422 12216 38428
rect 11796 38412 11848 38418
rect 11796 38354 11848 38360
rect 11980 38412 12032 38418
rect 11980 38354 12032 38360
rect 12256 38412 12308 38418
rect 12256 38354 12308 38360
rect 11808 37942 11836 38354
rect 11796 37936 11848 37942
rect 11796 37878 11848 37884
rect 11992 37738 12020 38354
rect 12268 38214 12296 38354
rect 12256 38208 12308 38214
rect 12256 38150 12308 38156
rect 11980 37732 12032 37738
rect 11980 37674 12032 37680
rect 11992 37466 12020 37674
rect 11980 37460 12032 37466
rect 11980 37402 12032 37408
rect 11888 37256 11940 37262
rect 11888 37198 11940 37204
rect 11796 37188 11848 37194
rect 11796 37130 11848 37136
rect 11808 36786 11836 37130
rect 11796 36780 11848 36786
rect 11796 36722 11848 36728
rect 11900 36378 11928 37198
rect 12268 36378 12296 38150
rect 11888 36372 11940 36378
rect 11888 36314 11940 36320
rect 12256 36372 12308 36378
rect 12256 36314 12308 36320
rect 12164 36236 12216 36242
rect 12164 36178 12216 36184
rect 11980 36032 12032 36038
rect 11980 35974 12032 35980
rect 11716 35788 11836 35816
rect 11702 35592 11758 35601
rect 11702 35527 11758 35536
rect 11716 35290 11744 35527
rect 11704 35284 11756 35290
rect 11704 35226 11756 35232
rect 11612 35080 11664 35086
rect 11612 35022 11664 35028
rect 11624 34746 11652 35022
rect 11612 34740 11664 34746
rect 11612 34682 11664 34688
rect 11440 33918 11560 33946
rect 11440 33017 11468 33918
rect 11518 33824 11574 33833
rect 11518 33759 11574 33768
rect 11532 33522 11560 33759
rect 11624 33538 11652 34682
rect 11520 33516 11572 33522
rect 11624 33510 11744 33538
rect 11520 33458 11572 33464
rect 11612 33448 11664 33454
rect 11612 33390 11664 33396
rect 11426 33008 11482 33017
rect 11426 32943 11482 32952
rect 11520 32904 11572 32910
rect 11348 32830 11468 32858
rect 11520 32846 11572 32852
rect 11336 32768 11388 32774
rect 11336 32710 11388 32716
rect 11348 31793 11376 32710
rect 11334 31784 11390 31793
rect 11334 31719 11390 31728
rect 11244 30932 11296 30938
rect 11244 30874 11296 30880
rect 11242 30832 11298 30841
rect 11242 30767 11298 30776
rect 11256 30394 11284 30767
rect 11244 30388 11296 30394
rect 11244 30330 11296 30336
rect 11348 30326 11376 31719
rect 11336 30320 11388 30326
rect 11336 30262 11388 30268
rect 11336 30116 11388 30122
rect 11336 30058 11388 30064
rect 11244 30048 11296 30054
rect 11244 29990 11296 29996
rect 11256 29850 11284 29990
rect 11244 29844 11296 29850
rect 11244 29786 11296 29792
rect 11244 29708 11296 29714
rect 11244 29650 11296 29656
rect 10980 28886 11192 28914
rect 10980 28665 11008 28886
rect 10966 28656 11022 28665
rect 10784 28620 10836 28626
rect 10966 28591 11022 28600
rect 10784 28562 10836 28568
rect 10796 28218 10824 28562
rect 11060 28416 11112 28422
rect 11060 28358 11112 28364
rect 10784 28212 10836 28218
rect 10784 28154 10836 28160
rect 10968 28076 11020 28082
rect 10968 28018 11020 28024
rect 10782 27976 10838 27985
rect 10782 27911 10838 27920
rect 10796 27674 10824 27911
rect 10784 27668 10836 27674
rect 10784 27610 10836 27616
rect 10796 25362 10824 27610
rect 10876 26988 10928 26994
rect 10876 26930 10928 26936
rect 10888 26897 10916 26930
rect 10980 26926 11008 28018
rect 10968 26920 11020 26926
rect 10874 26888 10930 26897
rect 10968 26862 11020 26868
rect 10874 26823 10930 26832
rect 10888 26450 10916 26823
rect 10968 26784 11020 26790
rect 11072 26772 11100 28358
rect 11256 27010 11284 29650
rect 11348 29345 11376 30058
rect 11334 29336 11390 29345
rect 11334 29271 11390 29280
rect 11440 27878 11468 32830
rect 11532 32434 11560 32846
rect 11520 32428 11572 32434
rect 11520 32370 11572 32376
rect 11624 32201 11652 33390
rect 11716 32881 11744 33510
rect 11702 32872 11758 32881
rect 11702 32807 11758 32816
rect 11704 32768 11756 32774
rect 11704 32710 11756 32716
rect 11716 32609 11744 32710
rect 11702 32600 11758 32609
rect 11702 32535 11758 32544
rect 11808 32450 11836 35788
rect 11888 35148 11940 35154
rect 11888 35090 11940 35096
rect 11900 35057 11928 35090
rect 11886 35048 11942 35057
rect 11886 34983 11942 34992
rect 11992 34610 12020 35974
rect 12176 35834 12204 36178
rect 12254 36000 12310 36009
rect 12254 35935 12310 35944
rect 12164 35828 12216 35834
rect 12164 35770 12216 35776
rect 12268 35222 12296 35935
rect 12256 35216 12308 35222
rect 12256 35158 12308 35164
rect 12256 34944 12308 34950
rect 12256 34886 12308 34892
rect 11980 34604 12032 34610
rect 11980 34546 12032 34552
rect 12072 34400 12124 34406
rect 12072 34342 12124 34348
rect 11888 33992 11940 33998
rect 11886 33960 11888 33969
rect 11940 33960 11942 33969
rect 11886 33895 11942 33904
rect 11886 33416 11942 33425
rect 11886 33351 11942 33360
rect 11900 32570 11928 33351
rect 12084 33318 12112 34342
rect 12268 34134 12296 34886
rect 12256 34128 12308 34134
rect 12256 34070 12308 34076
rect 11980 33312 12032 33318
rect 11980 33254 12032 33260
rect 12072 33312 12124 33318
rect 12072 33254 12124 33260
rect 11992 32586 12020 33254
rect 12162 33008 12218 33017
rect 12162 32943 12164 32952
rect 12216 32943 12218 32952
rect 12164 32914 12216 32920
rect 12072 32768 12124 32774
rect 12070 32736 12072 32745
rect 12124 32736 12126 32745
rect 12070 32671 12126 32680
rect 11888 32564 11940 32570
rect 11992 32558 12112 32586
rect 12176 32570 12204 32914
rect 12256 32768 12308 32774
rect 12256 32710 12308 32716
rect 11888 32506 11940 32512
rect 11716 32422 11836 32450
rect 11610 32192 11666 32201
rect 11610 32127 11666 32136
rect 11520 31680 11572 31686
rect 11520 31622 11572 31628
rect 11532 31346 11560 31622
rect 11520 31340 11572 31346
rect 11520 31282 11572 31288
rect 11520 30932 11572 30938
rect 11520 30874 11572 30880
rect 11336 27872 11388 27878
rect 11336 27814 11388 27820
rect 11428 27872 11480 27878
rect 11428 27814 11480 27820
rect 11020 26744 11100 26772
rect 10968 26726 11020 26732
rect 10876 26444 10928 26450
rect 10876 26386 10928 26392
rect 11072 25362 11100 26744
rect 11164 26982 11284 27010
rect 11164 25702 11192 26982
rect 11244 26920 11296 26926
rect 11244 26862 11296 26868
rect 11256 26586 11284 26862
rect 11348 26625 11376 27814
rect 11334 26616 11390 26625
rect 11244 26580 11296 26586
rect 11334 26551 11390 26560
rect 11244 26522 11296 26528
rect 11242 26480 11298 26489
rect 11242 26415 11298 26424
rect 11152 25696 11204 25702
rect 11152 25638 11204 25644
rect 10784 25356 10836 25362
rect 10784 25298 10836 25304
rect 11060 25356 11112 25362
rect 11060 25298 11112 25304
rect 10796 24138 10824 25298
rect 10968 24608 11020 24614
rect 10968 24550 11020 24556
rect 10980 24410 11008 24550
rect 10968 24404 11020 24410
rect 10968 24346 11020 24352
rect 10876 24268 10928 24274
rect 10876 24210 10928 24216
rect 10784 24132 10836 24138
rect 10784 24074 10836 24080
rect 10888 23866 10916 24210
rect 10876 23860 10928 23866
rect 10876 23802 10928 23808
rect 10980 23186 11008 24346
rect 11164 24206 11192 25638
rect 11152 24200 11204 24206
rect 11152 24142 11204 24148
rect 11256 23610 11284 26415
rect 11334 25528 11390 25537
rect 11334 25463 11336 25472
rect 11388 25463 11390 25472
rect 11336 25434 11388 25440
rect 11336 24064 11388 24070
rect 11336 24006 11388 24012
rect 11348 23730 11376 24006
rect 11336 23724 11388 23730
rect 11336 23666 11388 23672
rect 11256 23582 11376 23610
rect 11152 23520 11204 23526
rect 11152 23462 11204 23468
rect 11164 23322 11192 23462
rect 11152 23316 11204 23322
rect 11152 23258 11204 23264
rect 10968 23180 11020 23186
rect 10968 23122 11020 23128
rect 10784 23044 10836 23050
rect 10784 22986 10836 22992
rect 10796 22710 10824 22986
rect 10980 22710 11008 23122
rect 11164 22778 11192 23258
rect 11152 22772 11204 22778
rect 11152 22714 11204 22720
rect 10784 22704 10836 22710
rect 10784 22646 10836 22652
rect 10968 22704 11020 22710
rect 10968 22646 11020 22652
rect 11244 22704 11296 22710
rect 11244 22646 11296 22652
rect 11256 21622 11284 22646
rect 11348 22234 11376 23582
rect 11336 22228 11388 22234
rect 11336 22170 11388 22176
rect 11336 22092 11388 22098
rect 11336 22034 11388 22040
rect 11348 21690 11376 22034
rect 11336 21684 11388 21690
rect 11336 21626 11388 21632
rect 11244 21616 11296 21622
rect 11244 21558 11296 21564
rect 10966 21448 11022 21457
rect 10966 21383 10968 21392
rect 11020 21383 11022 21392
rect 10968 21354 11020 21360
rect 11348 18834 11376 21626
rect 11336 18828 11388 18834
rect 11336 18770 11388 18776
rect 11440 18193 11468 27814
rect 11532 26489 11560 30874
rect 11624 28150 11652 32127
rect 11716 30938 11744 32422
rect 11900 32366 11928 32506
rect 11888 32360 11940 32366
rect 11888 32302 11940 32308
rect 11886 32192 11942 32201
rect 11886 32127 11942 32136
rect 11796 31680 11848 31686
rect 11796 31622 11848 31628
rect 11704 30932 11756 30938
rect 11704 30874 11756 30880
rect 11808 30802 11836 31622
rect 11900 31482 11928 32127
rect 11888 31476 11940 31482
rect 11888 31418 11940 31424
rect 11980 31272 12032 31278
rect 11978 31240 11980 31249
rect 12032 31240 12034 31249
rect 11888 31204 11940 31210
rect 11978 31175 12034 31184
rect 11888 31146 11940 31152
rect 11900 30841 11928 31146
rect 11886 30832 11942 30841
rect 11796 30796 11848 30802
rect 11992 30802 12020 31175
rect 11886 30767 11942 30776
rect 11980 30796 12032 30802
rect 11796 30738 11848 30744
rect 11980 30738 12032 30744
rect 11704 30728 11756 30734
rect 11808 30705 11836 30738
rect 11704 30670 11756 30676
rect 11794 30696 11850 30705
rect 11716 29646 11744 30670
rect 11794 30631 11850 30640
rect 12084 30394 12112 32558
rect 12164 32564 12216 32570
rect 12164 32506 12216 32512
rect 12268 32065 12296 32710
rect 12254 32056 12310 32065
rect 12254 31991 12310 32000
rect 12256 31748 12308 31754
rect 12256 31690 12308 31696
rect 12268 31521 12296 31690
rect 12254 31512 12310 31521
rect 12254 31447 12310 31456
rect 12162 31240 12218 31249
rect 12162 31175 12218 31184
rect 12072 30388 12124 30394
rect 12072 30330 12124 30336
rect 11980 30116 12032 30122
rect 11980 30058 12032 30064
rect 11886 30016 11942 30025
rect 11886 29951 11942 29960
rect 11900 29866 11928 29951
rect 11808 29850 11928 29866
rect 11808 29844 11940 29850
rect 11808 29838 11888 29844
rect 11704 29640 11756 29646
rect 11704 29582 11756 29588
rect 11716 29510 11744 29582
rect 11704 29504 11756 29510
rect 11704 29446 11756 29452
rect 11612 28144 11664 28150
rect 11612 28086 11664 28092
rect 11716 27656 11744 29446
rect 11808 28762 11836 29838
rect 11888 29786 11940 29792
rect 11888 29572 11940 29578
rect 11888 29514 11940 29520
rect 11900 29345 11928 29514
rect 11886 29336 11942 29345
rect 11886 29271 11888 29280
rect 11940 29271 11942 29280
rect 11888 29242 11940 29248
rect 11900 29211 11928 29242
rect 11796 28756 11848 28762
rect 11796 28698 11848 28704
rect 11716 27628 11836 27656
rect 11704 27532 11756 27538
rect 11704 27474 11756 27480
rect 11716 27062 11744 27474
rect 11704 27056 11756 27062
rect 11704 26998 11756 27004
rect 11612 26852 11664 26858
rect 11612 26794 11664 26800
rect 11518 26480 11574 26489
rect 11518 26415 11574 26424
rect 11520 25968 11572 25974
rect 11518 25936 11520 25945
rect 11572 25936 11574 25945
rect 11518 25871 11574 25880
rect 11624 23186 11652 26794
rect 11808 24324 11836 27628
rect 11888 27328 11940 27334
rect 11888 27270 11940 27276
rect 11900 26994 11928 27270
rect 11888 26988 11940 26994
rect 11888 26930 11940 26936
rect 11992 25401 12020 30058
rect 12072 29844 12124 29850
rect 12072 29786 12124 29792
rect 12084 29753 12112 29786
rect 12070 29744 12126 29753
rect 12070 29679 12126 29688
rect 12176 29696 12204 31175
rect 12256 31136 12308 31142
rect 12254 31104 12256 31113
rect 12308 31104 12310 31113
rect 12254 31039 12310 31048
rect 12176 29668 12296 29696
rect 12268 29306 12296 29668
rect 12256 29300 12308 29306
rect 12256 29242 12308 29248
rect 12164 29232 12216 29238
rect 12164 29174 12216 29180
rect 12176 28014 12204 29174
rect 12268 29102 12296 29242
rect 12256 29096 12308 29102
rect 12256 29038 12308 29044
rect 12360 28762 12388 46310
rect 12452 46170 12480 46446
rect 12440 46164 12492 46170
rect 12440 46106 12492 46112
rect 12544 44402 12572 55218
rect 12636 47666 12664 67759
rect 14108 67658 14136 71839
rect 15198 70816 15254 70825
rect 15198 70751 15254 70760
rect 15212 69873 15240 70751
rect 15198 69864 15254 69873
rect 15198 69799 15254 69808
rect 14004 67652 14056 67658
rect 14004 67594 14056 67600
rect 14096 67652 14148 67658
rect 14096 67594 14148 67600
rect 13820 63436 13872 63442
rect 13820 63378 13872 63384
rect 13832 62694 13860 63378
rect 14016 63306 14044 67594
rect 14094 65512 14150 65521
rect 14094 65447 14150 65456
rect 14004 63300 14056 63306
rect 14004 63242 14056 63248
rect 13820 62688 13872 62694
rect 13820 62630 13872 62636
rect 13176 61600 13228 61606
rect 13174 61568 13176 61577
rect 13832 61577 13860 62630
rect 13912 61600 13964 61606
rect 13228 61568 13230 61577
rect 13174 61503 13230 61512
rect 13818 61568 13874 61577
rect 13912 61542 13964 61548
rect 13818 61503 13874 61512
rect 13358 58032 13414 58041
rect 13358 57967 13414 57976
rect 13266 56672 13322 56681
rect 13266 56607 13322 56616
rect 13280 56506 13308 56607
rect 13268 56500 13320 56506
rect 13268 56442 13320 56448
rect 13280 56302 13308 56442
rect 13268 56296 13320 56302
rect 13268 56238 13320 56244
rect 12716 55888 12768 55894
rect 12716 55830 12768 55836
rect 12728 55418 12756 55830
rect 13176 55820 13228 55826
rect 13176 55762 13228 55768
rect 12716 55412 12768 55418
rect 12716 55354 12768 55360
rect 13188 55282 13216 55762
rect 13176 55276 13228 55282
rect 13176 55218 13228 55224
rect 13372 54738 13400 57967
rect 13924 57934 13952 61542
rect 13728 57928 13780 57934
rect 13728 57870 13780 57876
rect 13912 57928 13964 57934
rect 13912 57870 13964 57876
rect 13740 56658 13768 57870
rect 14016 56710 14044 63242
rect 13648 56630 13768 56658
rect 14004 56704 14056 56710
rect 14004 56646 14056 56652
rect 13544 56160 13596 56166
rect 13544 56102 13596 56108
rect 13452 55616 13504 55622
rect 13452 55558 13504 55564
rect 13464 55185 13492 55558
rect 13450 55176 13506 55185
rect 13450 55111 13506 55120
rect 13176 54732 13228 54738
rect 13176 54674 13228 54680
rect 13360 54732 13412 54738
rect 13360 54674 13412 54680
rect 13188 54330 13216 54674
rect 13360 54528 13412 54534
rect 13266 54496 13322 54505
rect 13556 54505 13584 56102
rect 13648 55842 13676 56630
rect 14016 56302 14044 56646
rect 14004 56296 14056 56302
rect 14004 56238 14056 56244
rect 13648 55814 13860 55842
rect 13636 55752 13688 55758
rect 13636 55694 13688 55700
rect 13648 54874 13676 55694
rect 13636 54868 13688 54874
rect 13636 54810 13688 54816
rect 13360 54470 13412 54476
rect 13542 54496 13598 54505
rect 13266 54431 13322 54440
rect 13176 54324 13228 54330
rect 13176 54266 13228 54272
rect 13280 49366 13308 54431
rect 13372 54097 13400 54470
rect 13542 54431 13598 54440
rect 13358 54088 13414 54097
rect 13358 54023 13414 54032
rect 13832 53242 13860 55814
rect 13912 55616 13964 55622
rect 13912 55558 13964 55564
rect 13924 55418 13952 55558
rect 13912 55412 13964 55418
rect 13912 55354 13964 55360
rect 14016 54194 14044 56238
rect 14004 54188 14056 54194
rect 14004 54130 14056 54136
rect 13820 53236 13872 53242
rect 13820 53178 13872 53184
rect 13820 49768 13872 49774
rect 13820 49710 13872 49716
rect 13268 49360 13320 49366
rect 13268 49302 13320 49308
rect 13728 49292 13780 49298
rect 13728 49234 13780 49240
rect 13544 49224 13596 49230
rect 13544 49166 13596 49172
rect 13268 49156 13320 49162
rect 13268 49098 13320 49104
rect 13280 48686 13308 49098
rect 13556 48686 13584 49166
rect 13268 48680 13320 48686
rect 13268 48622 13320 48628
rect 13544 48680 13596 48686
rect 13544 48622 13596 48628
rect 12808 48204 12860 48210
rect 12808 48146 12860 48152
rect 12820 47802 12848 48146
rect 12808 47796 12860 47802
rect 12808 47738 12860 47744
rect 13176 47796 13228 47802
rect 13176 47738 13228 47744
rect 12624 47660 12676 47666
rect 12624 47602 12676 47608
rect 12992 47592 13044 47598
rect 12992 47534 13044 47540
rect 13004 47190 13032 47534
rect 12992 47184 13044 47190
rect 12992 47126 13044 47132
rect 12806 46880 12862 46889
rect 12806 46815 12862 46824
rect 12716 46572 12768 46578
rect 12716 46514 12768 46520
rect 12728 46374 12756 46514
rect 12716 46368 12768 46374
rect 12716 46310 12768 46316
rect 12820 46034 12848 46815
rect 12808 46028 12860 46034
rect 12808 45970 12860 45976
rect 12820 45286 12848 45970
rect 12808 45280 12860 45286
rect 12808 45222 12860 45228
rect 12532 44396 12584 44402
rect 12532 44338 12584 44344
rect 12532 44260 12584 44266
rect 12532 44202 12584 44208
rect 12544 43994 12572 44202
rect 12820 44198 12848 45222
rect 13084 44804 13136 44810
rect 13084 44746 13136 44752
rect 12900 44736 12952 44742
rect 12900 44678 12952 44684
rect 12912 44402 12940 44678
rect 12900 44396 12952 44402
rect 12900 44338 12952 44344
rect 13096 44334 13124 44746
rect 13084 44328 13136 44334
rect 13004 44288 13084 44316
rect 12808 44192 12860 44198
rect 12808 44134 12860 44140
rect 12532 43988 12584 43994
rect 12532 43930 12584 43936
rect 12624 43104 12676 43110
rect 12624 43046 12676 43052
rect 12440 41812 12492 41818
rect 12440 41754 12492 41760
rect 12452 39846 12480 41754
rect 12636 41614 12664 43046
rect 12900 42764 12952 42770
rect 12900 42706 12952 42712
rect 12714 42664 12770 42673
rect 12714 42599 12716 42608
rect 12768 42599 12770 42608
rect 12716 42570 12768 42576
rect 12716 42356 12768 42362
rect 12716 42298 12768 42304
rect 12624 41608 12676 41614
rect 12624 41550 12676 41556
rect 12622 40352 12678 40361
rect 12622 40287 12678 40296
rect 12440 39840 12492 39846
rect 12440 39782 12492 39788
rect 12452 34202 12480 39782
rect 12636 38418 12664 40287
rect 12624 38412 12676 38418
rect 12624 38354 12676 38360
rect 12532 38208 12584 38214
rect 12532 38150 12584 38156
rect 12544 37874 12572 38150
rect 12636 38010 12664 38354
rect 12624 38004 12676 38010
rect 12624 37946 12676 37952
rect 12532 37868 12584 37874
rect 12532 37810 12584 37816
rect 12544 35680 12572 37810
rect 12636 36802 12664 37946
rect 12728 36922 12756 42298
rect 12912 42022 12940 42706
rect 13004 42362 13032 44288
rect 13084 44270 13136 44276
rect 13084 43852 13136 43858
rect 13084 43794 13136 43800
rect 13096 43314 13124 43794
rect 13084 43308 13136 43314
rect 13084 43250 13136 43256
rect 13084 42764 13136 42770
rect 13084 42706 13136 42712
rect 12992 42356 13044 42362
rect 12992 42298 13044 42304
rect 12992 42220 13044 42226
rect 12992 42162 13044 42168
rect 12900 42016 12952 42022
rect 12900 41958 12952 41964
rect 12912 41750 12940 41958
rect 12900 41744 12952 41750
rect 12900 41686 12952 41692
rect 12900 41608 12952 41614
rect 12900 41550 12952 41556
rect 12808 37664 12860 37670
rect 12808 37606 12860 37612
rect 12820 37126 12848 37606
rect 12808 37120 12860 37126
rect 12808 37062 12860 37068
rect 12716 36916 12768 36922
rect 12716 36858 12768 36864
rect 12636 36774 12756 36802
rect 12820 36786 12848 37062
rect 12624 36712 12676 36718
rect 12624 36654 12676 36660
rect 12636 35834 12664 36654
rect 12624 35828 12676 35834
rect 12624 35770 12676 35776
rect 12544 35652 12664 35680
rect 12532 35556 12584 35562
rect 12532 35498 12584 35504
rect 12544 35290 12572 35498
rect 12532 35284 12584 35290
rect 12532 35226 12584 35232
rect 12636 34474 12664 35652
rect 12624 34468 12676 34474
rect 12624 34410 12676 34416
rect 12440 34196 12492 34202
rect 12440 34138 12492 34144
rect 12532 33992 12584 33998
rect 12532 33934 12584 33940
rect 12544 33561 12572 33934
rect 12636 33862 12664 34410
rect 12624 33856 12676 33862
rect 12624 33798 12676 33804
rect 12530 33552 12586 33561
rect 12530 33487 12532 33496
rect 12584 33487 12586 33496
rect 12532 33458 12584 33464
rect 12544 33427 12572 33458
rect 12440 33380 12492 33386
rect 12636 33368 12664 33798
rect 12728 33538 12756 36774
rect 12808 36780 12860 36786
rect 12808 36722 12860 36728
rect 12820 36242 12848 36722
rect 12808 36236 12860 36242
rect 12808 36178 12860 36184
rect 12806 34640 12862 34649
rect 12806 34575 12808 34584
rect 12860 34575 12862 34584
rect 12808 34546 12860 34552
rect 12808 33992 12860 33998
rect 12808 33934 12860 33940
rect 12820 33697 12848 33934
rect 12806 33688 12862 33697
rect 12806 33623 12862 33632
rect 12728 33510 12848 33538
rect 12440 33322 12492 33328
rect 12544 33340 12664 33368
rect 12452 32298 12480 33322
rect 12440 32292 12492 32298
rect 12440 32234 12492 32240
rect 12544 31754 12572 33340
rect 12714 32872 12770 32881
rect 12624 32836 12676 32842
rect 12714 32807 12716 32816
rect 12624 32778 12676 32784
rect 12768 32807 12770 32816
rect 12716 32778 12768 32784
rect 12636 32366 12664 32778
rect 12624 32360 12676 32366
rect 12624 32302 12676 32308
rect 12728 31958 12756 32778
rect 12820 32774 12848 33510
rect 12808 32768 12860 32774
rect 12808 32710 12860 32716
rect 12716 31952 12768 31958
rect 12716 31894 12768 31900
rect 12912 31906 12940 41550
rect 13004 40338 13032 42162
rect 13096 41818 13124 42706
rect 13084 41812 13136 41818
rect 13084 41754 13136 41760
rect 13084 41608 13136 41614
rect 13084 41550 13136 41556
rect 13096 41002 13124 41550
rect 13084 40996 13136 41002
rect 13084 40938 13136 40944
rect 13188 40361 13216 47738
rect 13280 47682 13308 48622
rect 13556 48346 13584 48622
rect 13544 48340 13596 48346
rect 13544 48282 13596 48288
rect 13740 48074 13768 49234
rect 13728 48068 13780 48074
rect 13728 48010 13780 48016
rect 13832 47802 13860 49710
rect 14004 49292 14056 49298
rect 14004 49234 14056 49240
rect 14016 48890 14044 49234
rect 14004 48884 14056 48890
rect 14004 48826 14056 48832
rect 14004 48136 14056 48142
rect 14004 48078 14056 48084
rect 13820 47796 13872 47802
rect 13820 47738 13872 47744
rect 13280 47654 13400 47682
rect 13268 47592 13320 47598
rect 13268 47534 13320 47540
rect 13280 45830 13308 47534
rect 13372 46170 13400 47654
rect 13452 47592 13504 47598
rect 13452 47534 13504 47540
rect 13464 47258 13492 47534
rect 14016 47462 14044 48078
rect 14004 47456 14056 47462
rect 14004 47398 14056 47404
rect 13452 47252 13504 47258
rect 13452 47194 13504 47200
rect 13464 46578 13492 47194
rect 13912 47116 13964 47122
rect 13912 47058 13964 47064
rect 13924 46714 13952 47058
rect 14016 47054 14044 47398
rect 14004 47048 14056 47054
rect 14004 46990 14056 46996
rect 13912 46708 13964 46714
rect 13912 46650 13964 46656
rect 13452 46572 13504 46578
rect 13452 46514 13504 46520
rect 13634 46336 13690 46345
rect 13634 46271 13690 46280
rect 13360 46164 13412 46170
rect 13360 46106 13412 46112
rect 13268 45824 13320 45830
rect 13268 45766 13320 45772
rect 13280 43874 13308 45766
rect 13372 45490 13400 46106
rect 13360 45484 13412 45490
rect 13360 45426 13412 45432
rect 13372 45082 13400 45426
rect 13452 45416 13504 45422
rect 13452 45358 13504 45364
rect 13360 45076 13412 45082
rect 13360 45018 13412 45024
rect 13372 43994 13400 45018
rect 13464 44810 13492 45358
rect 13452 44804 13504 44810
rect 13452 44746 13504 44752
rect 13360 43988 13412 43994
rect 13360 43930 13412 43936
rect 13280 43846 13400 43874
rect 13372 42770 13400 43846
rect 13360 42764 13412 42770
rect 13360 42706 13412 42712
rect 13372 42294 13400 42706
rect 13360 42288 13412 42294
rect 13360 42230 13412 42236
rect 13452 41676 13504 41682
rect 13452 41618 13504 41624
rect 13464 40934 13492 41618
rect 13452 40928 13504 40934
rect 13452 40870 13504 40876
rect 13464 40662 13492 40870
rect 13452 40656 13504 40662
rect 13452 40598 13504 40604
rect 13174 40352 13230 40361
rect 13004 40310 13124 40338
rect 13096 39982 13124 40310
rect 13174 40287 13230 40296
rect 13084 39976 13136 39982
rect 13082 39944 13084 39953
rect 13136 39944 13138 39953
rect 13082 39879 13138 39888
rect 13452 39840 13504 39846
rect 13452 39782 13504 39788
rect 13084 38752 13136 38758
rect 13084 38694 13136 38700
rect 12990 36816 13046 36825
rect 12990 36751 13046 36760
rect 13004 36242 13032 36751
rect 12992 36236 13044 36242
rect 12992 36178 13044 36184
rect 13004 35222 13032 36178
rect 12992 35216 13044 35222
rect 12992 35158 13044 35164
rect 12992 34536 13044 34542
rect 12992 34478 13044 34484
rect 13004 32978 13032 34478
rect 13096 33046 13124 38694
rect 13360 38344 13412 38350
rect 13360 38286 13412 38292
rect 13268 37664 13320 37670
rect 13268 37606 13320 37612
rect 13176 36916 13228 36922
rect 13176 36858 13228 36864
rect 13084 33040 13136 33046
rect 13084 32982 13136 32988
rect 12992 32972 13044 32978
rect 12992 32914 13044 32920
rect 13004 32026 13032 32914
rect 13082 32872 13138 32881
rect 13082 32807 13138 32816
rect 13096 32502 13124 32807
rect 13084 32496 13136 32502
rect 13084 32438 13136 32444
rect 13084 32224 13136 32230
rect 13084 32166 13136 32172
rect 12992 32020 13044 32026
rect 12992 31962 13044 31968
rect 12912 31878 13032 31906
rect 12440 31748 12492 31754
rect 12440 31690 12492 31696
rect 12532 31748 12584 31754
rect 12532 31690 12584 31696
rect 12808 31748 12860 31754
rect 12808 31690 12860 31696
rect 12452 31482 12480 31690
rect 12440 31476 12492 31482
rect 12440 31418 12492 31424
rect 12820 31124 12848 31690
rect 12898 31648 12954 31657
rect 12898 31583 12954 31592
rect 12912 31278 12940 31583
rect 12900 31272 12952 31278
rect 12900 31214 12952 31220
rect 12820 31096 12940 31124
rect 12530 30968 12586 30977
rect 12440 30932 12492 30938
rect 12530 30903 12586 30912
rect 12440 30874 12492 30880
rect 12452 29617 12480 30874
rect 12544 30870 12572 30903
rect 12532 30864 12584 30870
rect 12532 30806 12584 30812
rect 12438 29608 12494 29617
rect 12438 29543 12494 29552
rect 12440 29504 12492 29510
rect 12440 29446 12492 29452
rect 12452 29306 12480 29446
rect 12440 29300 12492 29306
rect 12440 29242 12492 29248
rect 12440 28960 12492 28966
rect 12440 28902 12492 28908
rect 12348 28756 12400 28762
rect 12348 28698 12400 28704
rect 12256 28688 12308 28694
rect 12256 28630 12308 28636
rect 12164 28008 12216 28014
rect 12164 27950 12216 27956
rect 12268 27470 12296 28630
rect 12452 28218 12480 28902
rect 12440 28212 12492 28218
rect 12440 28154 12492 28160
rect 12440 27872 12492 27878
rect 12440 27814 12492 27820
rect 12452 27674 12480 27814
rect 12440 27668 12492 27674
rect 12440 27610 12492 27616
rect 12256 27464 12308 27470
rect 12256 27406 12308 27412
rect 12268 27062 12296 27406
rect 12256 27056 12308 27062
rect 12544 27044 12572 30806
rect 12624 30796 12676 30802
rect 12624 30738 12676 30744
rect 12636 30394 12664 30738
rect 12912 30734 12940 31096
rect 12900 30728 12952 30734
rect 12714 30696 12770 30705
rect 12898 30696 12900 30705
rect 12952 30696 12954 30705
rect 12714 30631 12770 30640
rect 12808 30660 12860 30666
rect 12624 30388 12676 30394
rect 12624 30330 12676 30336
rect 12728 30326 12756 30631
rect 12898 30631 12954 30640
rect 12808 30602 12860 30608
rect 12716 30320 12768 30326
rect 12622 30288 12678 30297
rect 12716 30262 12768 30268
rect 12622 30223 12678 30232
rect 12636 29782 12664 30223
rect 12820 30172 12848 30602
rect 12728 30144 12848 30172
rect 12900 30184 12952 30190
rect 12624 29776 12676 29782
rect 12624 29718 12676 29724
rect 12622 29472 12678 29481
rect 12622 29407 12678 29416
rect 12636 27538 12664 29407
rect 12624 27532 12676 27538
rect 12624 27474 12676 27480
rect 12256 26998 12308 27004
rect 12360 27016 12572 27044
rect 12162 25800 12218 25809
rect 12162 25735 12218 25744
rect 12176 25498 12204 25735
rect 12164 25492 12216 25498
rect 12164 25434 12216 25440
rect 11978 25392 12034 25401
rect 11888 25356 11940 25362
rect 11978 25327 12034 25336
rect 11888 25298 11940 25304
rect 11900 24954 11928 25298
rect 11888 24948 11940 24954
rect 11888 24890 11940 24896
rect 11980 24608 12032 24614
rect 11980 24550 12032 24556
rect 11992 24410 12020 24550
rect 11980 24404 12032 24410
rect 11980 24346 12032 24352
rect 11808 24296 11928 24324
rect 11794 23352 11850 23361
rect 11794 23287 11850 23296
rect 11612 23180 11664 23186
rect 11612 23122 11664 23128
rect 11624 22710 11652 23122
rect 11808 22778 11836 23287
rect 11796 22772 11848 22778
rect 11796 22714 11848 22720
rect 11612 22704 11664 22710
rect 11612 22646 11664 22652
rect 11808 22574 11836 22714
rect 11796 22568 11848 22574
rect 11796 22510 11848 22516
rect 11900 22386 11928 24296
rect 12162 22808 12218 22817
rect 12162 22743 12218 22752
rect 11716 22358 11928 22386
rect 11612 22024 11664 22030
rect 11612 21966 11664 21972
rect 11624 21865 11652 21966
rect 11610 21856 11666 21865
rect 11610 21791 11666 21800
rect 11426 18184 11482 18193
rect 11426 18119 11482 18128
rect 10968 16176 11020 16182
rect 10968 16118 11020 16124
rect 10980 15994 11008 16118
rect 10980 15966 11100 15994
rect 11072 14482 11100 15966
rect 11716 14521 11744 22358
rect 11888 22228 11940 22234
rect 11888 22170 11940 22176
rect 11900 20369 11928 22170
rect 12072 21004 12124 21010
rect 12072 20946 12124 20952
rect 11980 20936 12032 20942
rect 11980 20878 12032 20884
rect 11992 20398 12020 20878
rect 12084 20602 12112 20946
rect 12072 20596 12124 20602
rect 12072 20538 12124 20544
rect 11980 20392 12032 20398
rect 11886 20360 11942 20369
rect 11980 20334 12032 20340
rect 11886 20295 11942 20304
rect 12084 20058 12112 20538
rect 12072 20052 12124 20058
rect 12072 19994 12124 20000
rect 11888 18760 11940 18766
rect 11888 18702 11940 18708
rect 11900 18057 11928 18702
rect 12072 18692 12124 18698
rect 12072 18634 12124 18640
rect 12084 18426 12112 18634
rect 12072 18420 12124 18426
rect 12072 18362 12124 18368
rect 12176 18222 12204 22743
rect 12268 22012 12296 26998
rect 12360 25498 12388 27016
rect 12728 26840 12756 30144
rect 12900 30126 12952 30132
rect 12912 29578 12940 30126
rect 12900 29572 12952 29578
rect 12900 29514 12952 29520
rect 12808 29504 12860 29510
rect 12808 29446 12860 29452
rect 12820 28694 12848 29446
rect 13004 29034 13032 31878
rect 13096 30666 13124 32166
rect 13084 30660 13136 30666
rect 13084 30602 13136 30608
rect 13082 30560 13138 30569
rect 13082 30495 13138 30504
rect 13096 30190 13124 30495
rect 13084 30184 13136 30190
rect 13084 30126 13136 30132
rect 13084 30048 13136 30054
rect 13084 29990 13136 29996
rect 12992 29028 13044 29034
rect 12992 28970 13044 28976
rect 12900 28756 12952 28762
rect 12900 28698 12952 28704
rect 12808 28688 12860 28694
rect 12808 28630 12860 28636
rect 12808 28552 12860 28558
rect 12806 28520 12808 28529
rect 12860 28520 12862 28529
rect 12806 28455 12862 28464
rect 12820 26926 12848 28455
rect 12912 27878 12940 28698
rect 12992 28620 13044 28626
rect 12992 28562 13044 28568
rect 12900 27872 12952 27878
rect 12900 27814 12952 27820
rect 13004 27606 13032 28562
rect 12992 27600 13044 27606
rect 12990 27568 12992 27577
rect 13044 27568 13046 27577
rect 12990 27503 13046 27512
rect 12808 26920 12860 26926
rect 12808 26862 12860 26868
rect 12544 26812 12756 26840
rect 12348 25492 12400 25498
rect 12348 25434 12400 25440
rect 12348 25220 12400 25226
rect 12348 25162 12400 25168
rect 12360 24698 12388 25162
rect 12440 24812 12492 24818
rect 12440 24754 12492 24760
rect 12452 24698 12480 24754
rect 12360 24670 12480 24698
rect 12544 24392 12572 26812
rect 13096 26772 13124 29990
rect 13188 28082 13216 36858
rect 13280 35766 13308 37606
rect 13372 37262 13400 38286
rect 13360 37256 13412 37262
rect 13360 37198 13412 37204
rect 13360 36712 13412 36718
rect 13360 36654 13412 36660
rect 13372 35834 13400 36654
rect 13360 35828 13412 35834
rect 13360 35770 13412 35776
rect 13268 35760 13320 35766
rect 13268 35702 13320 35708
rect 13268 35624 13320 35630
rect 13268 35566 13320 35572
rect 13280 33454 13308 35566
rect 13360 35012 13412 35018
rect 13360 34954 13412 34960
rect 13372 34746 13400 34954
rect 13360 34740 13412 34746
rect 13360 34682 13412 34688
rect 13360 34060 13412 34066
rect 13360 34002 13412 34008
rect 13268 33448 13320 33454
rect 13268 33390 13320 33396
rect 13372 32858 13400 34002
rect 13280 32830 13400 32858
rect 13280 32026 13308 32830
rect 13360 32768 13412 32774
rect 13360 32710 13412 32716
rect 13268 32020 13320 32026
rect 13268 31962 13320 31968
rect 13266 31648 13322 31657
rect 13266 31583 13322 31592
rect 13280 31482 13308 31583
rect 13268 31476 13320 31482
rect 13268 31418 13320 31424
rect 13280 31278 13308 31418
rect 13268 31272 13320 31278
rect 13268 31214 13320 31220
rect 13268 31136 13320 31142
rect 13268 31078 13320 31084
rect 13280 30258 13308 31078
rect 13268 30252 13320 30258
rect 13268 30194 13320 30200
rect 13280 29850 13308 30194
rect 13372 30054 13400 32710
rect 13464 32230 13492 39782
rect 13542 38312 13598 38321
rect 13542 38247 13598 38256
rect 13556 37806 13584 38247
rect 13648 38010 13676 46271
rect 13924 46170 13952 46650
rect 14016 46374 14044 46990
rect 14004 46368 14056 46374
rect 14004 46310 14056 46316
rect 13912 46164 13964 46170
rect 13912 46106 13964 46112
rect 14016 45966 14044 46310
rect 14004 45960 14056 45966
rect 14004 45902 14056 45908
rect 14016 45286 14044 45902
rect 14004 45280 14056 45286
rect 14004 45222 14056 45228
rect 13728 44940 13780 44946
rect 13728 44882 13780 44888
rect 13740 44538 13768 44882
rect 14016 44742 14044 45222
rect 14108 44946 14136 65447
rect 14554 63880 14610 63889
rect 14554 63815 14610 63824
rect 14278 57624 14334 57633
rect 14278 57559 14280 57568
rect 14332 57559 14334 57568
rect 14280 57530 14332 57536
rect 14280 56908 14332 56914
rect 14280 56850 14332 56856
rect 14186 56400 14242 56409
rect 14186 56335 14188 56344
rect 14240 56335 14242 56344
rect 14188 56306 14240 56312
rect 14292 56234 14320 56850
rect 14370 56808 14426 56817
rect 14370 56743 14426 56752
rect 14280 56228 14332 56234
rect 14280 56170 14332 56176
rect 14384 55962 14412 56743
rect 14464 56704 14516 56710
rect 14464 56646 14516 56652
rect 14372 55956 14424 55962
rect 14372 55898 14424 55904
rect 14278 55312 14334 55321
rect 14476 55282 14504 56646
rect 14278 55247 14334 55256
rect 14464 55276 14516 55282
rect 14188 55208 14240 55214
rect 14188 55150 14240 55156
rect 14200 54738 14228 55150
rect 14188 54732 14240 54738
rect 14188 54674 14240 54680
rect 14200 54330 14228 54674
rect 14188 54324 14240 54330
rect 14188 54266 14240 54272
rect 14292 53650 14320 55247
rect 14464 55218 14516 55224
rect 14370 54632 14426 54641
rect 14370 54567 14372 54576
rect 14424 54567 14426 54576
rect 14372 54538 14424 54544
rect 14464 54188 14516 54194
rect 14464 54130 14516 54136
rect 14372 54120 14424 54126
rect 14372 54062 14424 54068
rect 14384 53650 14412 54062
rect 14476 53786 14504 54130
rect 14464 53780 14516 53786
rect 14464 53722 14516 53728
rect 14280 53644 14332 53650
rect 14280 53586 14332 53592
rect 14372 53644 14424 53650
rect 14372 53586 14424 53592
rect 14292 53174 14320 53586
rect 14280 53168 14332 53174
rect 14280 53110 14332 53116
rect 14280 48204 14332 48210
rect 14280 48146 14332 48152
rect 14292 47802 14320 48146
rect 14280 47796 14332 47802
rect 14280 47738 14332 47744
rect 14568 46578 14596 63815
rect 15108 57996 15160 58002
rect 15108 57938 15160 57944
rect 15120 57594 15148 57938
rect 15108 57588 15160 57594
rect 15108 57530 15160 57536
rect 15014 57352 15070 57361
rect 15014 57287 15016 57296
rect 15068 57287 15070 57296
rect 15016 57258 15068 57264
rect 15016 56704 15068 56710
rect 15016 56646 15068 56652
rect 14646 55992 14702 56001
rect 14646 55927 14702 55936
rect 14660 55418 14688 55927
rect 15028 55894 15056 56646
rect 15016 55888 15068 55894
rect 15016 55830 15068 55836
rect 14832 55820 14884 55826
rect 14832 55762 14884 55768
rect 14648 55412 14700 55418
rect 14648 55354 14700 55360
rect 14660 53786 14688 55354
rect 14844 55146 14872 55762
rect 15016 55616 15068 55622
rect 15016 55558 15068 55564
rect 15028 55350 15056 55558
rect 15016 55344 15068 55350
rect 15016 55286 15068 55292
rect 14832 55140 14884 55146
rect 14832 55082 14884 55088
rect 14844 54806 14872 55082
rect 14832 54800 14884 54806
rect 14832 54742 14884 54748
rect 15028 54534 15056 55286
rect 15120 55214 15148 57530
rect 15108 55208 15160 55214
rect 15108 55150 15160 55156
rect 15292 55208 15344 55214
rect 15292 55150 15344 55156
rect 15200 55072 15252 55078
rect 15200 55014 15252 55020
rect 15016 54528 15068 54534
rect 15016 54470 15068 54476
rect 14832 54052 14884 54058
rect 14832 53994 14884 54000
rect 14740 53984 14792 53990
rect 14738 53952 14740 53961
rect 14792 53952 14794 53961
rect 14844 53938 14872 53994
rect 14922 53952 14978 53961
rect 14844 53910 14922 53938
rect 14738 53887 14794 53896
rect 14922 53887 14978 53896
rect 15106 53816 15162 53825
rect 14648 53780 14700 53786
rect 15106 53751 15162 53760
rect 14648 53722 14700 53728
rect 14660 53174 14688 53722
rect 15120 53718 15148 53751
rect 15108 53712 15160 53718
rect 15028 53660 15108 53666
rect 15028 53654 15160 53660
rect 15028 53638 15148 53654
rect 14924 53508 14976 53514
rect 14924 53450 14976 53456
rect 14740 53440 14792 53446
rect 14740 53382 14792 53388
rect 14648 53168 14700 53174
rect 14648 53110 14700 53116
rect 14752 52737 14780 53382
rect 14738 52728 14794 52737
rect 14738 52663 14740 52672
rect 14792 52663 14794 52672
rect 14740 52634 14792 52640
rect 14752 52603 14780 52634
rect 14936 51542 14964 53450
rect 14924 51536 14976 51542
rect 14924 51478 14976 51484
rect 14740 51264 14792 51270
rect 14738 51232 14740 51241
rect 14792 51232 14794 51241
rect 14738 51167 14794 51176
rect 15028 51066 15056 53638
rect 15212 53417 15240 55014
rect 15304 54670 15332 55150
rect 15292 54664 15344 54670
rect 15292 54606 15344 54612
rect 15198 53408 15254 53417
rect 15198 53343 15254 53352
rect 15212 52494 15240 53343
rect 15292 53032 15344 53038
rect 15292 52974 15344 52980
rect 15304 52601 15332 52974
rect 15290 52592 15346 52601
rect 15290 52527 15346 52536
rect 15200 52488 15252 52494
rect 15200 52430 15252 52436
rect 15106 52184 15162 52193
rect 15212 52154 15240 52430
rect 15106 52119 15162 52128
rect 15200 52148 15252 52154
rect 15120 51610 15148 52119
rect 15200 52090 15252 52096
rect 15108 51604 15160 51610
rect 15108 51546 15160 51552
rect 15016 51060 15068 51066
rect 15016 51002 15068 51008
rect 15108 50856 15160 50862
rect 15108 50798 15160 50804
rect 14830 50552 14886 50561
rect 14830 50487 14886 50496
rect 14844 50182 14872 50487
rect 14832 50176 14884 50182
rect 14832 50118 14884 50124
rect 14844 49094 14872 50118
rect 15016 49360 15068 49366
rect 15016 49302 15068 49308
rect 14832 49088 14884 49094
rect 14832 49030 14884 49036
rect 14648 48544 14700 48550
rect 14648 48486 14700 48492
rect 14660 48210 14688 48486
rect 14648 48204 14700 48210
rect 14648 48146 14700 48152
rect 14648 48000 14700 48006
rect 14648 47942 14700 47948
rect 14660 47598 14688 47942
rect 14648 47592 14700 47598
rect 14648 47534 14700 47540
rect 14556 46572 14608 46578
rect 14556 46514 14608 46520
rect 14462 45520 14518 45529
rect 14462 45455 14518 45464
rect 14096 44940 14148 44946
rect 14096 44882 14148 44888
rect 14004 44736 14056 44742
rect 14004 44678 14056 44684
rect 13728 44532 13780 44538
rect 13728 44474 13780 44480
rect 14108 44470 14136 44882
rect 14476 44810 14504 45455
rect 14464 44804 14516 44810
rect 14464 44746 14516 44752
rect 13820 44464 13872 44470
rect 13820 44406 13872 44412
rect 14096 44464 14148 44470
rect 14096 44406 14148 44412
rect 13832 44180 13860 44406
rect 13740 44152 13860 44180
rect 13740 42226 13768 44152
rect 14096 43240 14148 43246
rect 14096 43182 14148 43188
rect 14108 42906 14136 43182
rect 14096 42900 14148 42906
rect 14096 42842 14148 42848
rect 14096 42764 14148 42770
rect 14096 42706 14148 42712
rect 13728 42220 13780 42226
rect 13728 42162 13780 42168
rect 13820 40996 13872 41002
rect 13820 40938 13872 40944
rect 13832 40594 13860 40938
rect 13820 40588 13872 40594
rect 13820 40530 13872 40536
rect 13832 39846 13860 40530
rect 14004 40384 14056 40390
rect 14002 40352 14004 40361
rect 14056 40352 14058 40361
rect 14002 40287 14058 40296
rect 14108 40202 14136 42706
rect 14372 42288 14424 42294
rect 14372 42230 14424 42236
rect 14188 42152 14240 42158
rect 14188 42094 14240 42100
rect 14200 41818 14228 42094
rect 14384 41857 14412 42230
rect 14370 41848 14426 41857
rect 14188 41812 14240 41818
rect 14370 41783 14426 41792
rect 14188 41754 14240 41760
rect 14016 40174 14136 40202
rect 13820 39840 13872 39846
rect 13820 39782 13872 39788
rect 13912 38888 13964 38894
rect 13912 38830 13964 38836
rect 13924 38554 13952 38830
rect 13728 38548 13780 38554
rect 13728 38490 13780 38496
rect 13912 38548 13964 38554
rect 13912 38490 13964 38496
rect 13636 38004 13688 38010
rect 13636 37946 13688 37952
rect 13544 37800 13596 37806
rect 13544 37742 13596 37748
rect 13556 37466 13584 37742
rect 13544 37460 13596 37466
rect 13740 37448 13768 38490
rect 13912 38344 13964 38350
rect 13912 38286 13964 38292
rect 13924 38010 13952 38286
rect 13912 38004 13964 38010
rect 13912 37946 13964 37952
rect 13544 37402 13596 37408
rect 13648 37420 13768 37448
rect 13648 36768 13676 37420
rect 13726 37360 13782 37369
rect 13726 37295 13728 37304
rect 13780 37295 13782 37304
rect 13728 37266 13780 37272
rect 14016 36961 14044 40174
rect 14188 39432 14240 39438
rect 14188 39374 14240 39380
rect 14096 38412 14148 38418
rect 14096 38354 14148 38360
rect 14108 37097 14136 38354
rect 14094 37088 14150 37097
rect 14094 37023 14150 37032
rect 14002 36952 14058 36961
rect 14002 36887 14058 36896
rect 13648 36740 13768 36768
rect 13636 36644 13688 36650
rect 13636 36586 13688 36592
rect 13542 36544 13598 36553
rect 13542 36479 13598 36488
rect 13556 35222 13584 36479
rect 13544 35216 13596 35222
rect 13544 35158 13596 35164
rect 13542 34096 13598 34105
rect 13542 34031 13598 34040
rect 13556 33697 13584 34031
rect 13542 33688 13598 33697
rect 13542 33623 13598 33632
rect 13556 33386 13584 33623
rect 13544 33380 13596 33386
rect 13544 33322 13596 33328
rect 13556 33046 13584 33322
rect 13544 33040 13596 33046
rect 13544 32982 13596 32988
rect 13544 32428 13596 32434
rect 13544 32370 13596 32376
rect 13452 32224 13504 32230
rect 13452 32166 13504 32172
rect 13556 31822 13584 32370
rect 13544 31816 13596 31822
rect 13544 31758 13596 31764
rect 13452 31680 13504 31686
rect 13452 31622 13504 31628
rect 13464 31278 13492 31622
rect 13556 31414 13584 31758
rect 13544 31408 13596 31414
rect 13544 31350 13596 31356
rect 13452 31272 13504 31278
rect 13452 31214 13504 31220
rect 13464 30598 13492 31214
rect 13452 30592 13504 30598
rect 13452 30534 13504 30540
rect 13542 30560 13598 30569
rect 13360 30048 13412 30054
rect 13360 29990 13412 29996
rect 13268 29844 13320 29850
rect 13268 29786 13320 29792
rect 13280 29510 13308 29786
rect 13360 29640 13412 29646
rect 13360 29582 13412 29588
rect 13268 29504 13320 29510
rect 13268 29446 13320 29452
rect 13266 29200 13322 29209
rect 13372 29170 13400 29582
rect 13266 29135 13322 29144
rect 13360 29164 13412 29170
rect 13176 28076 13228 28082
rect 13176 28018 13228 28024
rect 12728 26744 13124 26772
rect 13176 26784 13228 26790
rect 12624 26444 12676 26450
rect 12624 26386 12676 26392
rect 12636 25974 12664 26386
rect 12624 25968 12676 25974
rect 12624 25910 12676 25916
rect 12624 25832 12676 25838
rect 12624 25774 12676 25780
rect 12636 25673 12664 25774
rect 12622 25664 12678 25673
rect 12622 25599 12678 25608
rect 12624 24744 12676 24750
rect 12624 24686 12676 24692
rect 12636 24614 12664 24686
rect 12624 24608 12676 24614
rect 12624 24550 12676 24556
rect 12452 24364 12572 24392
rect 12452 23866 12480 24364
rect 12532 24268 12584 24274
rect 12532 24210 12584 24216
rect 12440 23860 12492 23866
rect 12440 23802 12492 23808
rect 12348 23792 12400 23798
rect 12346 23760 12348 23769
rect 12400 23760 12402 23769
rect 12346 23695 12402 23704
rect 12544 23662 12572 24210
rect 12532 23656 12584 23662
rect 12532 23598 12584 23604
rect 12544 22982 12572 23598
rect 12624 23044 12676 23050
rect 12624 22986 12676 22992
rect 12532 22976 12584 22982
rect 12530 22944 12532 22953
rect 12584 22944 12586 22953
rect 12530 22879 12586 22888
rect 12636 22778 12664 22986
rect 12624 22772 12676 22778
rect 12624 22714 12676 22720
rect 12440 22568 12492 22574
rect 12440 22510 12492 22516
rect 12452 22409 12480 22510
rect 12438 22400 12494 22409
rect 12438 22335 12494 22344
rect 12348 22024 12400 22030
rect 12268 21984 12348 22012
rect 12268 21690 12296 21984
rect 12348 21966 12400 21972
rect 12532 22024 12584 22030
rect 12532 21966 12584 21972
rect 12256 21684 12308 21690
rect 12256 21626 12308 21632
rect 12268 20602 12296 21626
rect 12544 21622 12572 21966
rect 12532 21616 12584 21622
rect 12532 21558 12584 21564
rect 12256 20596 12308 20602
rect 12256 20538 12308 20544
rect 12440 20052 12492 20058
rect 12440 19994 12492 20000
rect 12452 19378 12480 19994
rect 12440 19372 12492 19378
rect 12440 19314 12492 19320
rect 12348 18896 12400 18902
rect 12348 18838 12400 18844
rect 12164 18216 12216 18222
rect 12164 18158 12216 18164
rect 11886 18048 11942 18057
rect 11886 17983 11942 17992
rect 12360 17882 12388 18838
rect 12452 18630 12480 19314
rect 12532 18828 12584 18834
rect 12532 18770 12584 18776
rect 12544 18680 12572 18770
rect 12544 18652 12664 18680
rect 12440 18624 12492 18630
rect 12440 18566 12492 18572
rect 12452 18290 12480 18566
rect 12440 18284 12492 18290
rect 12440 18226 12492 18232
rect 12348 17876 12400 17882
rect 12348 17818 12400 17824
rect 12636 17746 12664 18652
rect 12624 17740 12676 17746
rect 12624 17682 12676 17688
rect 11980 17672 12032 17678
rect 11980 17614 12032 17620
rect 11992 16153 12020 17614
rect 12164 17604 12216 17610
rect 12164 17546 12216 17552
rect 12176 17270 12204 17546
rect 12636 17338 12664 17682
rect 12624 17332 12676 17338
rect 12624 17274 12676 17280
rect 12164 17264 12216 17270
rect 12164 17206 12216 17212
rect 11978 16144 12034 16153
rect 11978 16079 12034 16088
rect 11702 14512 11758 14521
rect 11060 14476 11112 14482
rect 11060 14418 11112 14424
rect 11520 14476 11572 14482
rect 11702 14447 11758 14456
rect 11520 14418 11572 14424
rect 11532 14074 11560 14418
rect 11520 14068 11572 14074
rect 11520 14010 11572 14016
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12348 7336 12400 7342
rect 12346 7304 12348 7313
rect 12400 7304 12402 7313
rect 12346 7239 12402 7248
rect 12452 4690 12480 12718
rect 12728 12238 12756 26744
rect 13176 26726 13228 26732
rect 13188 26602 13216 26726
rect 13004 26574 13216 26602
rect 12898 26344 12954 26353
rect 12898 26279 12954 26288
rect 12806 24848 12862 24857
rect 12806 24783 12862 24792
rect 12820 24614 12848 24783
rect 12808 24608 12860 24614
rect 12808 24550 12860 24556
rect 12912 24274 12940 26279
rect 12808 24268 12860 24274
rect 12808 24210 12860 24216
rect 12900 24268 12952 24274
rect 12900 24210 12952 24216
rect 12820 23662 12848 24210
rect 13004 24070 13032 26574
rect 13280 26518 13308 29135
rect 13360 29106 13412 29112
rect 13372 28937 13400 29106
rect 13358 28928 13414 28937
rect 13358 28863 13414 28872
rect 13464 28762 13492 30534
rect 13542 30495 13598 30504
rect 13556 28966 13584 30495
rect 13544 28960 13596 28966
rect 13544 28902 13596 28908
rect 13452 28756 13504 28762
rect 13452 28698 13504 28704
rect 13452 28552 13504 28558
rect 13452 28494 13504 28500
rect 13464 28257 13492 28494
rect 13450 28248 13506 28257
rect 13450 28183 13506 28192
rect 13544 28076 13596 28082
rect 13544 28018 13596 28024
rect 13452 27872 13504 27878
rect 13450 27840 13452 27849
rect 13504 27840 13506 27849
rect 13450 27775 13506 27784
rect 13360 27668 13412 27674
rect 13360 27610 13412 27616
rect 13372 26926 13400 27610
rect 13556 27470 13584 28018
rect 13544 27464 13596 27470
rect 13464 27424 13544 27452
rect 13360 26920 13412 26926
rect 13360 26862 13412 26868
rect 13268 26512 13320 26518
rect 13082 26480 13138 26489
rect 13268 26454 13320 26460
rect 13082 26415 13138 26424
rect 13096 24750 13124 26415
rect 13372 26382 13400 26862
rect 13464 26586 13492 27424
rect 13544 27406 13596 27412
rect 13544 27328 13596 27334
rect 13544 27270 13596 27276
rect 13556 27033 13584 27270
rect 13542 27024 13598 27033
rect 13542 26959 13598 26968
rect 13648 26874 13676 36586
rect 13740 35290 13768 36740
rect 14016 36632 14044 36887
rect 13924 36604 14044 36632
rect 13924 35766 13952 36604
rect 14200 36553 14228 39374
rect 14280 39296 14332 39302
rect 14280 39238 14332 39244
rect 14292 38894 14320 39238
rect 14280 38888 14332 38894
rect 14280 38830 14332 38836
rect 14292 37874 14320 38830
rect 14370 38448 14426 38457
rect 14370 38383 14372 38392
rect 14424 38383 14426 38392
rect 14372 38354 14424 38360
rect 14280 37868 14332 37874
rect 14280 37810 14332 37816
rect 14280 37324 14332 37330
rect 14280 37266 14332 37272
rect 14186 36544 14242 36553
rect 14186 36479 14242 36488
rect 14096 35828 14148 35834
rect 14096 35770 14148 35776
rect 13912 35760 13964 35766
rect 13912 35702 13964 35708
rect 14108 35698 14136 35770
rect 14096 35692 14148 35698
rect 14096 35634 14148 35640
rect 13912 35556 13964 35562
rect 13912 35498 13964 35504
rect 13728 35284 13780 35290
rect 13728 35226 13780 35232
rect 13820 35148 13872 35154
rect 13820 35090 13872 35096
rect 13728 34944 13780 34950
rect 13728 34886 13780 34892
rect 13740 34406 13768 34886
rect 13728 34400 13780 34406
rect 13728 34342 13780 34348
rect 13832 33522 13860 35090
rect 13924 34649 13952 35498
rect 14108 34746 14136 35634
rect 14188 35148 14240 35154
rect 14188 35090 14240 35096
rect 14096 34740 14148 34746
rect 14096 34682 14148 34688
rect 13910 34640 13966 34649
rect 13910 34575 13966 34584
rect 14096 34468 14148 34474
rect 14096 34410 14148 34416
rect 13912 33992 13964 33998
rect 13912 33934 13964 33940
rect 13820 33516 13872 33522
rect 13820 33458 13872 33464
rect 13924 33318 13952 33934
rect 14108 33862 14136 34410
rect 14200 34066 14228 35090
rect 14292 34626 14320 37266
rect 14372 37188 14424 37194
rect 14372 37130 14424 37136
rect 14384 35630 14412 37130
rect 14476 36922 14504 44746
rect 14556 42016 14608 42022
rect 14556 41958 14608 41964
rect 14464 36916 14516 36922
rect 14464 36858 14516 36864
rect 14464 36644 14516 36650
rect 14464 36586 14516 36592
rect 14476 35630 14504 36586
rect 14372 35624 14424 35630
rect 14370 35592 14372 35601
rect 14464 35624 14516 35630
rect 14424 35592 14426 35601
rect 14464 35566 14516 35572
rect 14370 35527 14426 35536
rect 14476 35222 14504 35566
rect 14464 35216 14516 35222
rect 14464 35158 14516 35164
rect 14464 34944 14516 34950
rect 14464 34886 14516 34892
rect 14292 34598 14412 34626
rect 14188 34060 14240 34066
rect 14188 34002 14240 34008
rect 14096 33856 14148 33862
rect 14096 33798 14148 33804
rect 14280 33856 14332 33862
rect 14280 33798 14332 33804
rect 14108 33318 14136 33798
rect 14188 33652 14240 33658
rect 14188 33594 14240 33600
rect 13912 33312 13964 33318
rect 13912 33254 13964 33260
rect 14096 33312 14148 33318
rect 14096 33254 14148 33260
rect 13924 33153 13952 33254
rect 13910 33144 13966 33153
rect 13910 33079 13966 33088
rect 13912 33040 13964 33046
rect 13912 32982 13964 32988
rect 13820 32768 13872 32774
rect 13820 32710 13872 32716
rect 13832 32366 13860 32710
rect 13820 32360 13872 32366
rect 13820 32302 13872 32308
rect 13820 32224 13872 32230
rect 13820 32166 13872 32172
rect 13832 32065 13860 32166
rect 13818 32056 13874 32065
rect 13924 32042 13952 32982
rect 13924 32014 14044 32042
rect 13818 31991 13874 32000
rect 13832 31958 13860 31991
rect 13820 31952 13872 31958
rect 13820 31894 13872 31900
rect 13832 31482 13860 31894
rect 13912 31884 13964 31890
rect 13912 31826 13964 31832
rect 13820 31476 13872 31482
rect 13820 31418 13872 31424
rect 13924 31226 13952 31826
rect 13740 31198 13952 31226
rect 13740 30938 13768 31198
rect 13728 30932 13780 30938
rect 13728 30874 13780 30880
rect 13740 30818 13768 30874
rect 13740 30790 13952 30818
rect 13728 30728 13780 30734
rect 13728 30670 13780 30676
rect 13740 30326 13768 30670
rect 13728 30320 13780 30326
rect 13728 30262 13780 30268
rect 13820 30252 13872 30258
rect 13820 30194 13872 30200
rect 13728 30116 13780 30122
rect 13728 30058 13780 30064
rect 13740 29866 13768 30058
rect 13832 30054 13860 30194
rect 13924 30122 13952 30790
rect 13912 30116 13964 30122
rect 13912 30058 13964 30064
rect 13820 30048 13872 30054
rect 13820 29990 13872 29996
rect 13740 29838 13952 29866
rect 13728 29708 13780 29714
rect 13728 29650 13780 29656
rect 13740 29238 13768 29650
rect 13728 29232 13780 29238
rect 13728 29174 13780 29180
rect 13818 29200 13874 29209
rect 13740 28914 13768 29174
rect 13818 29135 13874 29144
rect 13832 29102 13860 29135
rect 13820 29096 13872 29102
rect 13820 29038 13872 29044
rect 13924 29034 13952 29838
rect 14016 29646 14044 32014
rect 14200 30954 14228 33594
rect 14292 33538 14320 33798
rect 14384 33697 14412 34598
rect 14476 34542 14504 34886
rect 14464 34536 14516 34542
rect 14464 34478 14516 34484
rect 14370 33688 14426 33697
rect 14370 33623 14426 33632
rect 14292 33522 14412 33538
rect 14292 33516 14424 33522
rect 14292 33510 14372 33516
rect 14292 33425 14320 33510
rect 14372 33458 14424 33464
rect 14278 33416 14334 33425
rect 14278 33351 14334 33360
rect 14372 33312 14424 33318
rect 14372 33254 14424 33260
rect 14384 32502 14412 33254
rect 14476 32774 14504 34478
rect 14464 32768 14516 32774
rect 14464 32710 14516 32716
rect 14372 32496 14424 32502
rect 14372 32438 14424 32444
rect 14384 32366 14412 32438
rect 14372 32360 14424 32366
rect 14372 32302 14424 32308
rect 14464 32020 14516 32026
rect 14464 31962 14516 31968
rect 14370 31920 14426 31929
rect 14370 31855 14372 31864
rect 14424 31855 14426 31864
rect 14372 31826 14424 31832
rect 14278 31648 14334 31657
rect 14278 31583 14334 31592
rect 14108 30926 14228 30954
rect 14108 29714 14136 30926
rect 14188 30864 14240 30870
rect 14188 30806 14240 30812
rect 14200 30394 14228 30806
rect 14188 30388 14240 30394
rect 14188 30330 14240 30336
rect 14200 30190 14228 30330
rect 14188 30184 14240 30190
rect 14188 30126 14240 30132
rect 14096 29708 14148 29714
rect 14096 29650 14148 29656
rect 14004 29640 14056 29646
rect 14004 29582 14056 29588
rect 14186 29608 14242 29617
rect 13912 29028 13964 29034
rect 13912 28970 13964 28976
rect 13910 28928 13966 28937
rect 13740 28886 13860 28914
rect 13728 28484 13780 28490
rect 13728 28426 13780 28432
rect 13740 28014 13768 28426
rect 13728 28008 13780 28014
rect 13728 27950 13780 27956
rect 13832 27538 13860 28886
rect 13910 28863 13966 28872
rect 13924 28422 13952 28863
rect 14016 28762 14044 29582
rect 14096 29572 14148 29578
rect 14186 29543 14242 29552
rect 14096 29514 14148 29520
rect 14108 29209 14136 29514
rect 14094 29200 14150 29209
rect 14200 29170 14228 29543
rect 14094 29135 14150 29144
rect 14188 29164 14240 29170
rect 14188 29106 14240 29112
rect 14096 29096 14148 29102
rect 14096 29038 14148 29044
rect 14004 28756 14056 28762
rect 14004 28698 14056 28704
rect 14016 28490 14044 28698
rect 14004 28484 14056 28490
rect 14004 28426 14056 28432
rect 13912 28416 13964 28422
rect 13912 28358 13964 28364
rect 13728 27532 13780 27538
rect 13728 27474 13780 27480
rect 13820 27532 13872 27538
rect 13820 27474 13872 27480
rect 13740 26926 13768 27474
rect 13556 26846 13676 26874
rect 13728 26920 13780 26926
rect 13728 26862 13780 26868
rect 13452 26580 13504 26586
rect 13452 26522 13504 26528
rect 13360 26376 13412 26382
rect 13174 26344 13230 26353
rect 13360 26318 13412 26324
rect 13174 26279 13230 26288
rect 13084 24744 13136 24750
rect 13084 24686 13136 24692
rect 13096 24177 13124 24686
rect 13082 24168 13138 24177
rect 13082 24103 13138 24112
rect 12992 24064 13044 24070
rect 12992 24006 13044 24012
rect 12808 23656 12860 23662
rect 12808 23598 12860 23604
rect 12820 23322 12848 23598
rect 12808 23316 12860 23322
rect 12808 23258 12860 23264
rect 12808 21616 12860 21622
rect 12808 21558 12860 21564
rect 12820 18766 12848 21558
rect 13004 19417 13032 24006
rect 13188 23050 13216 26279
rect 13372 25498 13400 26318
rect 13360 25492 13412 25498
rect 13360 25434 13412 25440
rect 13360 23180 13412 23186
rect 13360 23122 13412 23128
rect 13268 23112 13320 23118
rect 13268 23054 13320 23060
rect 13176 23044 13228 23050
rect 13176 22986 13228 22992
rect 13188 22681 13216 22986
rect 13174 22672 13230 22681
rect 13174 22607 13230 22616
rect 13084 22092 13136 22098
rect 13084 22034 13136 22040
rect 13096 21457 13124 22034
rect 13082 21448 13138 21457
rect 13082 21383 13138 21392
rect 13096 21146 13124 21383
rect 13084 21140 13136 21146
rect 13084 21082 13136 21088
rect 12990 19408 13046 19417
rect 12990 19343 13046 19352
rect 12808 18760 12860 18766
rect 12808 18702 12860 18708
rect 12820 17814 12848 18702
rect 12808 17808 12860 17814
rect 12808 17750 12860 17756
rect 12820 17338 12848 17750
rect 12992 17740 13044 17746
rect 12992 17682 13044 17688
rect 12900 17536 12952 17542
rect 12900 17478 12952 17484
rect 12808 17332 12860 17338
rect 12808 17274 12860 17280
rect 12912 17202 12940 17478
rect 12900 17196 12952 17202
rect 12900 17138 12952 17144
rect 13004 16794 13032 17682
rect 12992 16788 13044 16794
rect 12992 16730 13044 16736
rect 13176 12368 13228 12374
rect 13174 12336 13176 12345
rect 13228 12336 13230 12345
rect 13174 12271 13230 12280
rect 12716 12232 12768 12238
rect 12716 12174 12768 12180
rect 13280 8537 13308 23054
rect 13372 22778 13400 23122
rect 13360 22772 13412 22778
rect 13360 22714 13412 22720
rect 13452 18760 13504 18766
rect 13452 18702 13504 18708
rect 13360 18624 13412 18630
rect 13360 18566 13412 18572
rect 13372 15026 13400 18566
rect 13464 18290 13492 18702
rect 13452 18284 13504 18290
rect 13452 18226 13504 18232
rect 13556 17202 13584 26846
rect 13832 26790 13860 27474
rect 13820 26784 13872 26790
rect 13820 26726 13872 26732
rect 13820 26444 13872 26450
rect 13820 26386 13872 26392
rect 13832 25786 13860 26386
rect 13740 25770 13860 25786
rect 13728 25764 13860 25770
rect 13780 25758 13860 25764
rect 13728 25706 13780 25712
rect 13728 25220 13780 25226
rect 13832 25208 13860 25758
rect 13924 25702 13952 28358
rect 14016 28082 14044 28426
rect 14004 28076 14056 28082
rect 14004 28018 14056 28024
rect 14004 27940 14056 27946
rect 14004 27882 14056 27888
rect 14016 27441 14044 27882
rect 14108 27674 14136 29038
rect 14188 29028 14240 29034
rect 14188 28970 14240 28976
rect 14200 28257 14228 28970
rect 14186 28248 14242 28257
rect 14186 28183 14242 28192
rect 14188 28144 14240 28150
rect 14188 28086 14240 28092
rect 14200 27878 14228 28086
rect 14188 27872 14240 27878
rect 14188 27814 14240 27820
rect 14096 27668 14148 27674
rect 14096 27610 14148 27616
rect 14002 27432 14058 27441
rect 14002 27367 14058 27376
rect 14094 27296 14150 27305
rect 14094 27231 14150 27240
rect 14004 26376 14056 26382
rect 14004 26318 14056 26324
rect 14016 26217 14044 26318
rect 14002 26208 14058 26217
rect 14002 26143 14058 26152
rect 14016 26042 14044 26143
rect 14004 26036 14056 26042
rect 14004 25978 14056 25984
rect 14108 25922 14136 27231
rect 14016 25894 14136 25922
rect 13912 25696 13964 25702
rect 13912 25638 13964 25644
rect 13912 25288 13964 25294
rect 13912 25230 13964 25236
rect 13780 25180 13860 25208
rect 13728 25162 13780 25168
rect 13728 24744 13780 24750
rect 13728 24686 13780 24692
rect 13634 24576 13690 24585
rect 13634 24511 13690 24520
rect 13648 24342 13676 24511
rect 13636 24336 13688 24342
rect 13636 24278 13688 24284
rect 13740 24138 13768 24686
rect 13820 24676 13872 24682
rect 13820 24618 13872 24624
rect 13728 24132 13780 24138
rect 13728 24074 13780 24080
rect 13636 23724 13688 23730
rect 13636 23666 13688 23672
rect 13648 22574 13676 23666
rect 13740 23050 13768 24074
rect 13832 23866 13860 24618
rect 13924 24449 13952 25230
rect 13910 24440 13966 24449
rect 13910 24375 13912 24384
rect 13964 24375 13966 24384
rect 13912 24346 13964 24352
rect 13924 24315 13952 24346
rect 13912 24268 13964 24274
rect 13912 24210 13964 24216
rect 13924 23866 13952 24210
rect 13820 23860 13872 23866
rect 13820 23802 13872 23808
rect 13912 23860 13964 23866
rect 13912 23802 13964 23808
rect 14016 23361 14044 25894
rect 14096 25356 14148 25362
rect 14096 25298 14148 25304
rect 14108 24886 14136 25298
rect 14200 24954 14228 27814
rect 14188 24948 14240 24954
rect 14188 24890 14240 24896
rect 14096 24880 14148 24886
rect 14096 24822 14148 24828
rect 14094 24440 14150 24449
rect 14094 24375 14150 24384
rect 14002 23352 14058 23361
rect 14108 23322 14136 24375
rect 14188 23792 14240 23798
rect 14188 23734 14240 23740
rect 14002 23287 14058 23296
rect 14096 23316 14148 23322
rect 14096 23258 14148 23264
rect 14004 23180 14056 23186
rect 14004 23122 14056 23128
rect 13912 23112 13964 23118
rect 13912 23054 13964 23060
rect 13728 23044 13780 23050
rect 13728 22986 13780 22992
rect 13636 22568 13688 22574
rect 13636 22510 13688 22516
rect 13648 21690 13676 22510
rect 13740 22234 13768 22986
rect 13924 22574 13952 23054
rect 14016 22642 14044 23122
rect 14004 22636 14056 22642
rect 14004 22578 14056 22584
rect 13912 22568 13964 22574
rect 13912 22510 13964 22516
rect 13728 22228 13780 22234
rect 13728 22170 13780 22176
rect 13924 21894 13952 22510
rect 14016 22166 14044 22578
rect 14004 22160 14056 22166
rect 14004 22102 14056 22108
rect 14200 22098 14228 23734
rect 14188 22092 14240 22098
rect 14188 22034 14240 22040
rect 13912 21888 13964 21894
rect 13912 21830 13964 21836
rect 14200 21690 14228 22034
rect 13636 21684 13688 21690
rect 13636 21626 13688 21632
rect 14188 21684 14240 21690
rect 14188 21626 14240 21632
rect 13648 21010 13676 21626
rect 13636 21004 13688 21010
rect 13636 20946 13688 20952
rect 14292 20641 14320 31583
rect 14476 31346 14504 31962
rect 14464 31340 14516 31346
rect 14464 31282 14516 31288
rect 14372 31272 14424 31278
rect 14372 31214 14424 31220
rect 14384 29238 14412 31214
rect 14464 30796 14516 30802
rect 14464 30738 14516 30744
rect 14372 29232 14424 29238
rect 14372 29174 14424 29180
rect 14372 29096 14424 29102
rect 14372 29038 14424 29044
rect 14384 28694 14412 29038
rect 14372 28688 14424 28694
rect 14372 28630 14424 28636
rect 14384 27928 14412 28630
rect 14476 28626 14504 30738
rect 14464 28620 14516 28626
rect 14464 28562 14516 28568
rect 14464 27940 14516 27946
rect 14384 27900 14464 27928
rect 14464 27882 14516 27888
rect 14370 27840 14426 27849
rect 14370 27775 14426 27784
rect 14384 25974 14412 27775
rect 14464 27464 14516 27470
rect 14462 27432 14464 27441
rect 14516 27432 14518 27441
rect 14462 27367 14518 27376
rect 14464 26988 14516 26994
rect 14464 26930 14516 26936
rect 14372 25968 14424 25974
rect 14372 25910 14424 25916
rect 14372 25764 14424 25770
rect 14372 25706 14424 25712
rect 14384 25294 14412 25706
rect 14476 25362 14504 26930
rect 14568 26450 14596 41958
rect 14660 36786 14688 47534
rect 14740 46028 14792 46034
rect 14740 45970 14792 45976
rect 14752 45626 14780 45970
rect 14740 45620 14792 45626
rect 14740 45562 14792 45568
rect 14752 45082 14780 45562
rect 14740 45076 14792 45082
rect 14740 45018 14792 45024
rect 14740 42900 14792 42906
rect 14740 42842 14792 42848
rect 14752 42158 14780 42842
rect 14844 42770 14872 49030
rect 15028 47444 15056 49302
rect 15120 48929 15148 50798
rect 15292 50312 15344 50318
rect 15292 50254 15344 50260
rect 15200 50176 15252 50182
rect 15200 50118 15252 50124
rect 15212 49910 15240 50118
rect 15200 49904 15252 49910
rect 15200 49846 15252 49852
rect 15304 49298 15332 50254
rect 15396 49842 15424 73743
rect 16408 72865 16436 75783
rect 16488 74792 16540 74798
rect 16488 74734 16540 74740
rect 16394 72856 16450 72865
rect 16394 72791 16450 72800
rect 15842 72040 15898 72049
rect 15842 71975 15898 71984
rect 15566 71632 15622 71641
rect 15566 71567 15622 71576
rect 15476 56908 15528 56914
rect 15476 56850 15528 56856
rect 15488 55758 15516 56850
rect 15476 55752 15528 55758
rect 15474 55720 15476 55729
rect 15528 55720 15530 55729
rect 15474 55655 15530 55664
rect 15476 55412 15528 55418
rect 15476 55354 15528 55360
rect 15488 54874 15516 55354
rect 15476 54868 15528 54874
rect 15476 54810 15528 54816
rect 15474 53680 15530 53689
rect 15474 53615 15530 53624
rect 15488 52902 15516 53615
rect 15476 52896 15528 52902
rect 15476 52838 15528 52844
rect 15488 52630 15516 52838
rect 15476 52624 15528 52630
rect 15476 52566 15528 52572
rect 15488 51610 15516 52566
rect 15476 51604 15528 51610
rect 15476 51546 15528 51552
rect 15384 49836 15436 49842
rect 15384 49778 15436 49784
rect 15292 49292 15344 49298
rect 15292 49234 15344 49240
rect 15476 49292 15528 49298
rect 15476 49234 15528 49240
rect 15106 48920 15162 48929
rect 15304 48890 15332 49234
rect 15488 49178 15516 49234
rect 15396 49150 15516 49178
rect 15106 48855 15162 48864
rect 15292 48884 15344 48890
rect 15292 48826 15344 48832
rect 15304 48362 15332 48826
rect 15396 48822 15424 49150
rect 15384 48816 15436 48822
rect 15382 48784 15384 48793
rect 15436 48784 15438 48793
rect 15382 48719 15438 48728
rect 15120 48334 15332 48362
rect 15476 48340 15528 48346
rect 15120 48278 15148 48334
rect 15476 48282 15528 48288
rect 15108 48272 15160 48278
rect 15108 48214 15160 48220
rect 15120 47666 15148 48214
rect 15108 47660 15160 47666
rect 15108 47602 15160 47608
rect 15292 47592 15344 47598
rect 15212 47540 15292 47546
rect 15212 47534 15344 47540
rect 15212 47518 15332 47534
rect 15212 47444 15240 47518
rect 15028 47416 15240 47444
rect 14924 46912 14976 46918
rect 14924 46854 14976 46860
rect 14936 46492 14964 46854
rect 15016 46504 15068 46510
rect 14936 46464 15016 46492
rect 14936 46102 14964 46464
rect 15016 46446 15068 46452
rect 15120 46356 15148 47416
rect 15028 46328 15148 46356
rect 14924 46096 14976 46102
rect 14924 46038 14976 46044
rect 14832 42764 14884 42770
rect 14832 42706 14884 42712
rect 15028 42158 15056 46328
rect 15108 44736 15160 44742
rect 15160 44684 15332 44690
rect 15108 44678 15332 44684
rect 15120 44662 15332 44678
rect 15304 43790 15332 44662
rect 15384 43852 15436 43858
rect 15384 43794 15436 43800
rect 15292 43784 15344 43790
rect 15292 43726 15344 43732
rect 15108 43648 15160 43654
rect 15108 43590 15160 43596
rect 15120 42226 15148 43590
rect 15304 43450 15332 43726
rect 15292 43444 15344 43450
rect 15292 43386 15344 43392
rect 15396 43314 15424 43794
rect 15488 43466 15516 48282
rect 15580 48074 15608 71567
rect 15750 70952 15806 70961
rect 15750 70887 15806 70896
rect 15660 58132 15712 58138
rect 15660 58074 15712 58080
rect 15672 55690 15700 58074
rect 15764 56506 15792 70887
rect 15856 64161 15884 71975
rect 15934 70544 15990 70553
rect 15934 70479 15990 70488
rect 15842 64152 15898 64161
rect 15842 64087 15898 64096
rect 15948 63481 15976 70479
rect 15934 63472 15990 63481
rect 15934 63407 15990 63416
rect 16500 59401 16528 74734
rect 16486 59392 16542 59401
rect 16486 59327 16542 59336
rect 16580 59084 16632 59090
rect 16580 59026 16632 59032
rect 16592 58342 16620 59026
rect 16764 58880 16816 58886
rect 16764 58822 16816 58828
rect 16580 58336 16632 58342
rect 16580 58278 16632 58284
rect 16488 57792 16540 57798
rect 16488 57734 16540 57740
rect 16500 56914 16528 57734
rect 16592 57390 16620 58278
rect 16672 57792 16724 57798
rect 16672 57734 16724 57740
rect 16580 57384 16632 57390
rect 16580 57326 16632 57332
rect 16488 56908 16540 56914
rect 16488 56850 16540 56856
rect 16500 56710 16528 56850
rect 16488 56704 16540 56710
rect 16488 56646 16540 56652
rect 15752 56500 15804 56506
rect 15752 56442 15804 56448
rect 15660 55684 15712 55690
rect 15660 55626 15712 55632
rect 16028 55684 16080 55690
rect 16028 55626 16080 55632
rect 15936 55208 15988 55214
rect 15936 55150 15988 55156
rect 15660 54868 15712 54874
rect 15660 54810 15712 54816
rect 15672 53718 15700 54810
rect 15844 54528 15896 54534
rect 15844 54470 15896 54476
rect 15856 54262 15884 54470
rect 15844 54256 15896 54262
rect 15844 54198 15896 54204
rect 15948 53718 15976 55150
rect 16040 54602 16068 55626
rect 16500 55622 16528 56646
rect 16684 56273 16712 57734
rect 16670 56264 16726 56273
rect 16670 56199 16726 56208
rect 16488 55616 16540 55622
rect 16302 55584 16358 55593
rect 16488 55558 16540 55564
rect 16302 55519 16358 55528
rect 16120 55140 16172 55146
rect 16120 55082 16172 55088
rect 16028 54596 16080 54602
rect 16028 54538 16080 54544
rect 16132 54233 16160 55082
rect 16118 54224 16174 54233
rect 16118 54159 16174 54168
rect 16316 53718 16344 55519
rect 16776 55418 16804 58822
rect 16948 58472 17000 58478
rect 16948 58414 17000 58420
rect 16854 55856 16910 55865
rect 16854 55791 16856 55800
rect 16908 55791 16910 55800
rect 16856 55762 16908 55768
rect 16960 55758 16988 58414
rect 16948 55752 17000 55758
rect 16948 55694 17000 55700
rect 16960 55418 16988 55694
rect 16764 55412 16816 55418
rect 16764 55354 16816 55360
rect 16948 55412 17000 55418
rect 16948 55354 17000 55360
rect 16578 55176 16634 55185
rect 16578 55111 16634 55120
rect 16592 55078 16620 55111
rect 16580 55072 16632 55078
rect 16580 55014 16632 55020
rect 16592 54874 16620 55014
rect 16580 54868 16632 54874
rect 16580 54810 16632 54816
rect 16856 54664 16908 54670
rect 16856 54606 16908 54612
rect 16580 54596 16632 54602
rect 16580 54538 16632 54544
rect 16488 54528 16540 54534
rect 16488 54470 16540 54476
rect 16396 53780 16448 53786
rect 16396 53722 16448 53728
rect 15660 53712 15712 53718
rect 15660 53654 15712 53660
rect 15936 53712 15988 53718
rect 15936 53654 15988 53660
rect 16304 53712 16356 53718
rect 16304 53654 16356 53660
rect 15672 53446 15700 53654
rect 15660 53440 15712 53446
rect 15660 53382 15712 53388
rect 15672 53106 15700 53382
rect 15844 53236 15896 53242
rect 15844 53178 15896 53184
rect 15660 53100 15712 53106
rect 15660 53042 15712 53048
rect 15856 52884 15884 53178
rect 15948 53038 15976 53654
rect 16408 53038 16436 53722
rect 15936 53032 15988 53038
rect 16396 53032 16448 53038
rect 15936 52974 15988 52980
rect 16210 53000 16266 53009
rect 16396 52974 16448 52980
rect 16210 52935 16266 52944
rect 15856 52856 15976 52884
rect 15660 52556 15712 52562
rect 15660 52498 15712 52504
rect 15752 52556 15804 52562
rect 15752 52498 15804 52504
rect 15672 52154 15700 52498
rect 15660 52148 15712 52154
rect 15660 52090 15712 52096
rect 15672 51105 15700 52090
rect 15764 51814 15792 52498
rect 15752 51808 15804 51814
rect 15752 51750 15804 51756
rect 15658 51096 15714 51105
rect 15658 51031 15714 51040
rect 15660 50380 15712 50386
rect 15660 50322 15712 50328
rect 15672 49910 15700 50322
rect 15660 49904 15712 49910
rect 15660 49846 15712 49852
rect 15660 49768 15712 49774
rect 15660 49710 15712 49716
rect 15568 48068 15620 48074
rect 15568 48010 15620 48016
rect 15672 46889 15700 49710
rect 15844 48204 15896 48210
rect 15844 48146 15896 48152
rect 15752 47456 15804 47462
rect 15752 47398 15804 47404
rect 15764 47122 15792 47398
rect 15856 47190 15884 48146
rect 15844 47184 15896 47190
rect 15844 47126 15896 47132
rect 15752 47116 15804 47122
rect 15752 47058 15804 47064
rect 15658 46880 15714 46889
rect 15658 46815 15714 46824
rect 15568 46504 15620 46510
rect 15568 46446 15620 46452
rect 15660 46504 15712 46510
rect 15660 46446 15712 46452
rect 15580 45529 15608 46446
rect 15672 45830 15700 46446
rect 15764 46170 15792 47058
rect 15752 46164 15804 46170
rect 15752 46106 15804 46112
rect 15660 45824 15712 45830
rect 15660 45766 15712 45772
rect 15566 45520 15622 45529
rect 15566 45455 15622 45464
rect 15948 44538 15976 52856
rect 16224 52630 16252 52935
rect 16212 52624 16264 52630
rect 16212 52566 16264 52572
rect 16118 52048 16174 52057
rect 16118 51983 16120 51992
rect 16172 51983 16174 51992
rect 16120 51954 16172 51960
rect 16500 51921 16528 54470
rect 16592 53718 16620 54538
rect 16868 54369 16896 54606
rect 16854 54360 16910 54369
rect 16854 54295 16856 54304
rect 16908 54295 16910 54304
rect 16856 54266 16908 54272
rect 16960 54210 16988 55354
rect 16776 54182 16988 54210
rect 16580 53712 16632 53718
rect 16580 53654 16632 53660
rect 16592 53242 16620 53654
rect 16776 53650 16804 54182
rect 16854 54088 16910 54097
rect 16854 54023 16910 54032
rect 16868 53650 16896 54023
rect 16948 53712 17000 53718
rect 16948 53654 17000 53660
rect 16764 53644 16816 53650
rect 16764 53586 16816 53592
rect 16856 53644 16908 53650
rect 16856 53586 16908 53592
rect 16580 53236 16632 53242
rect 16580 53178 16632 53184
rect 16592 52698 16620 53178
rect 16776 53106 16804 53586
rect 16868 53242 16896 53586
rect 16856 53236 16908 53242
rect 16856 53178 16908 53184
rect 16764 53100 16816 53106
rect 16764 53042 16816 53048
rect 16580 52692 16632 52698
rect 16580 52634 16632 52640
rect 16776 52562 16804 53042
rect 16960 52737 16988 53654
rect 16946 52728 17002 52737
rect 16946 52663 17002 52672
rect 16960 52630 16988 52663
rect 16948 52624 17000 52630
rect 16948 52566 17000 52572
rect 16764 52556 16816 52562
rect 16764 52498 16816 52504
rect 16578 52456 16634 52465
rect 16578 52391 16634 52400
rect 16486 51912 16542 51921
rect 16486 51847 16542 51856
rect 16028 51468 16080 51474
rect 16028 51410 16080 51416
rect 16040 51066 16068 51410
rect 16592 51406 16620 52391
rect 16948 52352 17000 52358
rect 16948 52294 17000 52300
rect 16670 52184 16726 52193
rect 16670 52119 16726 52128
rect 16684 52018 16712 52119
rect 16672 52012 16724 52018
rect 16672 51954 16724 51960
rect 16960 51950 16988 52294
rect 16948 51944 17000 51950
rect 16948 51886 17000 51892
rect 16580 51400 16632 51406
rect 16580 51342 16632 51348
rect 16212 51264 16264 51270
rect 16212 51206 16264 51212
rect 16028 51060 16080 51066
rect 16028 51002 16080 51008
rect 16224 50998 16252 51206
rect 16212 50992 16264 50998
rect 16212 50934 16264 50940
rect 16592 50930 16620 51342
rect 16580 50924 16632 50930
rect 16580 50866 16632 50872
rect 16672 50856 16724 50862
rect 16672 50798 16724 50804
rect 16304 50176 16356 50182
rect 16304 50118 16356 50124
rect 16316 49774 16344 50118
rect 16304 49768 16356 49774
rect 16304 49710 16356 49716
rect 16684 49337 16712 50798
rect 16670 49328 16726 49337
rect 16670 49263 16726 49272
rect 16120 48204 16172 48210
rect 16120 48146 16172 48152
rect 16132 47598 16160 48146
rect 16672 48136 16724 48142
rect 16672 48078 16724 48084
rect 16684 47802 16712 48078
rect 16672 47796 16724 47802
rect 16672 47738 16724 47744
rect 16120 47592 16172 47598
rect 16120 47534 16172 47540
rect 16856 47592 16908 47598
rect 16856 47534 16908 47540
rect 16868 46889 16896 47534
rect 16948 47048 17000 47054
rect 16948 46990 17000 46996
rect 16854 46880 16910 46889
rect 16854 46815 16910 46824
rect 16960 46442 16988 46990
rect 17052 46481 17080 79070
rect 17512 77217 17540 79200
rect 18052 77376 18104 77382
rect 18052 77318 18104 77324
rect 17498 77208 17554 77217
rect 17498 77143 17554 77152
rect 18064 76974 18092 77318
rect 18432 77042 18460 79200
rect 18420 77036 18472 77042
rect 18420 76978 18472 76984
rect 17592 76968 17644 76974
rect 17592 76910 17644 76916
rect 18052 76968 18104 76974
rect 18052 76910 18104 76916
rect 19352 76922 19380 79200
rect 19580 77820 19876 77840
rect 19636 77818 19660 77820
rect 19716 77818 19740 77820
rect 19796 77818 19820 77820
rect 19658 77766 19660 77818
rect 19722 77766 19734 77818
rect 19796 77766 19798 77818
rect 19636 77764 19660 77766
rect 19716 77764 19740 77766
rect 19796 77764 19820 77766
rect 19580 77744 19876 77764
rect 17604 76430 17632 76910
rect 17684 76900 17736 76906
rect 19352 76894 19472 76922
rect 17684 76842 17736 76848
rect 17592 76424 17644 76430
rect 17592 76366 17644 76372
rect 17604 75954 17632 76366
rect 17500 75948 17552 75954
rect 17420 75908 17500 75936
rect 17420 75834 17448 75908
rect 17500 75890 17552 75896
rect 17592 75948 17644 75954
rect 17592 75890 17644 75896
rect 17420 75806 17540 75834
rect 17512 66298 17540 75806
rect 17224 66292 17276 66298
rect 17224 66234 17276 66240
rect 17500 66292 17552 66298
rect 17500 66234 17552 66240
rect 17236 66162 17264 66234
rect 17224 66156 17276 66162
rect 17224 66098 17276 66104
rect 17592 66156 17644 66162
rect 17592 66098 17644 66104
rect 17408 59084 17460 59090
rect 17408 59026 17460 59032
rect 17224 59016 17276 59022
rect 17224 58958 17276 58964
rect 17236 58682 17264 58958
rect 17420 58886 17448 59026
rect 17408 58880 17460 58886
rect 17408 58822 17460 58828
rect 17224 58676 17276 58682
rect 17224 58618 17276 58624
rect 17420 57798 17448 58822
rect 17132 57792 17184 57798
rect 17130 57760 17132 57769
rect 17408 57792 17460 57798
rect 17184 57760 17186 57769
rect 17408 57734 17460 57740
rect 17130 57695 17186 57704
rect 17420 57322 17448 57734
rect 17408 57316 17460 57322
rect 17408 57258 17460 57264
rect 17604 57066 17632 66098
rect 17328 57038 17632 57066
rect 17224 56160 17276 56166
rect 17224 56102 17276 56108
rect 17236 55758 17264 56102
rect 17224 55752 17276 55758
rect 17222 55720 17224 55729
rect 17276 55720 17278 55729
rect 17222 55655 17278 55664
rect 17236 55457 17264 55655
rect 17222 55448 17278 55457
rect 17222 55383 17278 55392
rect 17236 54738 17264 55383
rect 17224 54732 17276 54738
rect 17224 54674 17276 54680
rect 17236 54194 17264 54674
rect 17224 54188 17276 54194
rect 17224 54130 17276 54136
rect 17328 53156 17356 57038
rect 17500 56772 17552 56778
rect 17500 56714 17552 56720
rect 17512 56506 17540 56714
rect 17500 56500 17552 56506
rect 17500 56442 17552 56448
rect 17512 55962 17540 56442
rect 17592 56160 17644 56166
rect 17592 56102 17644 56108
rect 17500 55956 17552 55962
rect 17500 55898 17552 55904
rect 17500 55072 17552 55078
rect 17500 55014 17552 55020
rect 17512 54777 17540 55014
rect 17604 54874 17632 56102
rect 17592 54868 17644 54874
rect 17592 54810 17644 54816
rect 17498 54768 17554 54777
rect 17498 54703 17554 54712
rect 17500 54596 17552 54602
rect 17500 54538 17552 54544
rect 17512 53825 17540 54538
rect 17592 54324 17644 54330
rect 17592 54266 17644 54272
rect 17498 53816 17554 53825
rect 17604 53786 17632 54266
rect 17498 53751 17554 53760
rect 17592 53780 17644 53786
rect 17512 53650 17540 53751
rect 17592 53722 17644 53728
rect 17500 53644 17552 53650
rect 17500 53586 17552 53592
rect 17408 53236 17460 53242
rect 17408 53178 17460 53184
rect 17144 53128 17356 53156
rect 17038 46472 17094 46481
rect 16948 46436 17000 46442
rect 17038 46407 17094 46416
rect 16948 46378 17000 46384
rect 15936 44532 15988 44538
rect 15936 44474 15988 44480
rect 15948 44334 15976 44474
rect 16580 44464 16632 44470
rect 16580 44406 16632 44412
rect 15936 44328 15988 44334
rect 15936 44270 15988 44276
rect 16592 43858 16620 44406
rect 16580 43852 16632 43858
rect 16580 43794 16632 43800
rect 17144 43636 17172 53128
rect 17420 51474 17448 53178
rect 17592 52488 17644 52494
rect 17592 52430 17644 52436
rect 17408 51468 17460 51474
rect 17408 51410 17460 51416
rect 17222 50960 17278 50969
rect 17222 50895 17224 50904
rect 17276 50895 17278 50904
rect 17224 50866 17276 50872
rect 17316 50788 17368 50794
rect 17316 50730 17368 50736
rect 17222 50008 17278 50017
rect 17328 49978 17356 50730
rect 17420 50318 17448 51410
rect 17500 51400 17552 51406
rect 17500 51342 17552 51348
rect 17512 50794 17540 51342
rect 17604 51241 17632 52430
rect 17590 51232 17646 51241
rect 17590 51167 17646 51176
rect 17604 50833 17632 51167
rect 17590 50824 17646 50833
rect 17500 50788 17552 50794
rect 17590 50759 17646 50768
rect 17500 50730 17552 50736
rect 17408 50312 17460 50318
rect 17406 50280 17408 50289
rect 17460 50280 17462 50289
rect 17406 50215 17462 50224
rect 17222 49943 17224 49952
rect 17276 49943 17278 49952
rect 17316 49972 17368 49978
rect 17224 49914 17276 49920
rect 17316 49914 17368 49920
rect 17408 49292 17460 49298
rect 17408 49234 17460 49240
rect 17420 48929 17448 49234
rect 17406 48920 17462 48929
rect 17406 48855 17408 48864
rect 17460 48855 17462 48864
rect 17408 48826 17460 48832
rect 17224 48544 17276 48550
rect 17224 48486 17276 48492
rect 17236 48346 17264 48486
rect 17224 48340 17276 48346
rect 17224 48282 17276 48288
rect 17316 47116 17368 47122
rect 17316 47058 17368 47064
rect 17328 46374 17356 47058
rect 17500 46436 17552 46442
rect 17500 46378 17552 46384
rect 17316 46368 17368 46374
rect 17316 46310 17368 46316
rect 17328 43994 17356 46310
rect 17316 43988 17368 43994
rect 17316 43930 17368 43936
rect 17052 43608 17172 43636
rect 15488 43438 15608 43466
rect 15384 43308 15436 43314
rect 15384 43250 15436 43256
rect 15108 42220 15160 42226
rect 15108 42162 15160 42168
rect 14740 42152 14792 42158
rect 14740 42094 14792 42100
rect 15016 42152 15068 42158
rect 15016 42094 15068 42100
rect 15580 41290 15608 43438
rect 15580 41262 15884 41290
rect 15200 40384 15252 40390
rect 15200 40326 15252 40332
rect 14830 39808 14886 39817
rect 14830 39743 14886 39752
rect 14740 38208 14792 38214
rect 14740 38150 14792 38156
rect 14752 37398 14780 38150
rect 14844 37913 14872 39743
rect 15212 39522 15240 40326
rect 15476 39840 15528 39846
rect 15476 39782 15528 39788
rect 14936 39494 15424 39522
rect 14936 38894 14964 39494
rect 15108 39364 15160 39370
rect 15108 39306 15160 39312
rect 15016 39296 15068 39302
rect 15016 39238 15068 39244
rect 14924 38888 14976 38894
rect 14924 38830 14976 38836
rect 15028 37913 15056 39238
rect 15120 38894 15148 39306
rect 15108 38888 15160 38894
rect 15108 38830 15160 38836
rect 15120 38593 15148 38830
rect 15106 38584 15162 38593
rect 15106 38519 15162 38528
rect 15108 38208 15160 38214
rect 15108 38150 15160 38156
rect 15292 38208 15344 38214
rect 15292 38150 15344 38156
rect 14830 37904 14886 37913
rect 14830 37839 14886 37848
rect 15014 37904 15070 37913
rect 15014 37839 15070 37848
rect 15120 37505 15148 38150
rect 15106 37496 15162 37505
rect 15106 37431 15162 37440
rect 14740 37392 14792 37398
rect 14740 37334 14792 37340
rect 14832 37256 14884 37262
rect 14832 37198 14884 37204
rect 14740 37120 14792 37126
rect 14738 37088 14740 37097
rect 14792 37088 14794 37097
rect 14738 37023 14794 37032
rect 14740 36916 14792 36922
rect 14740 36858 14792 36864
rect 14648 36780 14700 36786
rect 14648 36722 14700 36728
rect 14646 35456 14702 35465
rect 14646 35391 14702 35400
rect 14660 35193 14688 35391
rect 14646 35184 14702 35193
rect 14646 35119 14702 35128
rect 14660 35086 14688 35119
rect 14648 35080 14700 35086
rect 14648 35022 14700 35028
rect 14648 33448 14700 33454
rect 14646 33416 14648 33425
rect 14700 33416 14702 33425
rect 14646 33351 14702 33360
rect 14648 32360 14700 32366
rect 14648 32302 14700 32308
rect 14660 32026 14688 32302
rect 14648 32020 14700 32026
rect 14648 31962 14700 31968
rect 14648 31884 14700 31890
rect 14648 31826 14700 31832
rect 14660 30258 14688 31826
rect 14648 30252 14700 30258
rect 14648 30194 14700 30200
rect 14648 30048 14700 30054
rect 14648 29990 14700 29996
rect 14660 29034 14688 29990
rect 14648 29028 14700 29034
rect 14648 28970 14700 28976
rect 14648 28552 14700 28558
rect 14648 28494 14700 28500
rect 14660 28014 14688 28494
rect 14752 28218 14780 36858
rect 14844 36378 14872 37198
rect 15108 36848 15160 36854
rect 15108 36790 15160 36796
rect 14924 36712 14976 36718
rect 14922 36680 14924 36689
rect 14976 36680 14978 36689
rect 14922 36615 14978 36624
rect 15016 36644 15068 36650
rect 15016 36586 15068 36592
rect 15028 36530 15056 36586
rect 14936 36502 15056 36530
rect 14832 36372 14884 36378
rect 14832 36314 14884 36320
rect 14936 36174 14964 36502
rect 14924 36168 14976 36174
rect 14924 36110 14976 36116
rect 14936 36038 14964 36110
rect 14924 36032 14976 36038
rect 14924 35974 14976 35980
rect 14936 35630 14964 35974
rect 14924 35624 14976 35630
rect 14924 35566 14976 35572
rect 14936 34950 14964 35566
rect 14924 34944 14976 34950
rect 14924 34886 14976 34892
rect 14936 34785 14964 34886
rect 14922 34776 14978 34785
rect 14832 34740 14884 34746
rect 15120 34728 15148 36790
rect 15200 36712 15252 36718
rect 15200 36654 15252 36660
rect 15212 36553 15240 36654
rect 15198 36544 15254 36553
rect 15198 36479 15254 36488
rect 15198 36408 15254 36417
rect 15198 36343 15254 36352
rect 15212 35562 15240 36343
rect 15304 36281 15332 38150
rect 15396 37330 15424 39494
rect 15488 37777 15516 39782
rect 15568 39500 15620 39506
rect 15568 39442 15620 39448
rect 15580 39098 15608 39442
rect 15568 39092 15620 39098
rect 15568 39034 15620 39040
rect 15474 37768 15530 37777
rect 15474 37703 15530 37712
rect 15752 37392 15804 37398
rect 15752 37334 15804 37340
rect 15384 37324 15436 37330
rect 15384 37266 15436 37272
rect 15396 36922 15424 37266
rect 15660 37120 15712 37126
rect 15660 37062 15712 37068
rect 15384 36916 15436 36922
rect 15384 36858 15436 36864
rect 15672 36718 15700 37062
rect 15660 36712 15712 36718
rect 15660 36654 15712 36660
rect 15384 36372 15436 36378
rect 15384 36314 15436 36320
rect 15290 36272 15346 36281
rect 15290 36207 15346 36216
rect 15304 35698 15332 36207
rect 15292 35692 15344 35698
rect 15292 35634 15344 35640
rect 15200 35556 15252 35562
rect 15200 35498 15252 35504
rect 15198 35184 15254 35193
rect 15198 35119 15254 35128
rect 14922 34711 14978 34720
rect 14832 34682 14884 34688
rect 15028 34700 15148 34728
rect 14844 34649 14872 34682
rect 14924 34672 14976 34678
rect 14830 34640 14886 34649
rect 14924 34614 14976 34620
rect 14830 34575 14886 34584
rect 14844 34542 14872 34575
rect 14832 34536 14884 34542
rect 14832 34478 14884 34484
rect 14830 33960 14886 33969
rect 14830 33895 14886 33904
rect 14844 33697 14872 33895
rect 14830 33688 14886 33697
rect 14830 33623 14886 33632
rect 14844 33454 14872 33623
rect 14832 33448 14884 33454
rect 14832 33390 14884 33396
rect 14832 32360 14884 32366
rect 14832 32302 14884 32308
rect 14844 32065 14872 32302
rect 14830 32056 14886 32065
rect 14830 31991 14886 32000
rect 14936 31890 14964 34614
rect 15028 33658 15056 34700
rect 15212 34626 15240 35119
rect 15120 34598 15240 34626
rect 15016 33652 15068 33658
rect 15016 33594 15068 33600
rect 15016 33448 15068 33454
rect 15016 33390 15068 33396
rect 15028 32774 15056 33390
rect 15016 32768 15068 32774
rect 15016 32710 15068 32716
rect 14924 31884 14976 31890
rect 14924 31826 14976 31832
rect 14922 31784 14978 31793
rect 14922 31719 14978 31728
rect 14936 30870 14964 31719
rect 15028 31278 15056 32710
rect 15120 31793 15148 34598
rect 15200 34536 15252 34542
rect 15200 34478 15252 34484
rect 15212 33522 15240 34478
rect 15200 33516 15252 33522
rect 15200 33458 15252 33464
rect 15200 33312 15252 33318
rect 15200 33254 15252 33260
rect 15106 31784 15162 31793
rect 15106 31719 15162 31728
rect 15106 31512 15162 31521
rect 15106 31447 15162 31456
rect 15016 31272 15068 31278
rect 15016 31214 15068 31220
rect 14924 30864 14976 30870
rect 14830 30832 14886 30841
rect 14924 30806 14976 30812
rect 14830 30767 14832 30776
rect 14884 30767 14886 30776
rect 14832 30738 14884 30744
rect 14922 30696 14978 30705
rect 14922 30631 14978 30640
rect 14832 30320 14884 30326
rect 14832 30262 14884 30268
rect 14844 29850 14872 30262
rect 14832 29844 14884 29850
rect 14832 29786 14884 29792
rect 14830 29608 14886 29617
rect 14830 29543 14886 29552
rect 14740 28212 14792 28218
rect 14740 28154 14792 28160
rect 14844 28098 14872 29543
rect 14752 28070 14872 28098
rect 14648 28008 14700 28014
rect 14648 27950 14700 27956
rect 14752 27538 14780 28070
rect 14832 28008 14884 28014
rect 14832 27950 14884 27956
rect 14740 27532 14792 27538
rect 14740 27474 14792 27480
rect 14648 27396 14700 27402
rect 14648 27338 14700 27344
rect 14660 27130 14688 27338
rect 14648 27124 14700 27130
rect 14648 27066 14700 27072
rect 14740 26784 14792 26790
rect 14740 26726 14792 26732
rect 14646 26616 14702 26625
rect 14646 26551 14648 26560
rect 14700 26551 14702 26560
rect 14648 26522 14700 26528
rect 14556 26444 14608 26450
rect 14556 26386 14608 26392
rect 14556 26308 14608 26314
rect 14556 26250 14608 26256
rect 14568 25906 14596 26250
rect 14556 25900 14608 25906
rect 14556 25842 14608 25848
rect 14660 25838 14688 26522
rect 14752 26518 14780 26726
rect 14740 26512 14792 26518
rect 14740 26454 14792 26460
rect 14752 26314 14780 26454
rect 14740 26308 14792 26314
rect 14740 26250 14792 26256
rect 14648 25832 14700 25838
rect 14648 25774 14700 25780
rect 14556 25764 14608 25770
rect 14556 25706 14608 25712
rect 14464 25356 14516 25362
rect 14464 25298 14516 25304
rect 14372 25288 14424 25294
rect 14372 25230 14424 25236
rect 14462 25256 14518 25265
rect 14384 24070 14412 25230
rect 14462 25191 14518 25200
rect 14476 24818 14504 25191
rect 14568 24993 14596 25706
rect 14740 25696 14792 25702
rect 14740 25638 14792 25644
rect 14752 25498 14780 25638
rect 14740 25492 14792 25498
rect 14740 25434 14792 25440
rect 14646 25120 14702 25129
rect 14646 25055 14702 25064
rect 14554 24984 14610 24993
rect 14554 24919 14610 24928
rect 14660 24834 14688 25055
rect 14464 24812 14516 24818
rect 14464 24754 14516 24760
rect 14568 24806 14688 24834
rect 14568 24290 14596 24806
rect 14738 24712 14794 24721
rect 14738 24647 14794 24656
rect 14752 24410 14780 24647
rect 14740 24404 14792 24410
rect 14740 24346 14792 24352
rect 14568 24262 14780 24290
rect 14556 24200 14608 24206
rect 14556 24142 14608 24148
rect 14372 24064 14424 24070
rect 14372 24006 14424 24012
rect 14384 22438 14412 24006
rect 14568 23769 14596 24142
rect 14554 23760 14610 23769
rect 14554 23695 14610 23704
rect 14372 22432 14424 22438
rect 14372 22374 14424 22380
rect 14568 21554 14596 23695
rect 14752 23474 14780 24262
rect 14844 24206 14872 27950
rect 14936 27606 14964 30631
rect 15028 30190 15056 31214
rect 15120 30734 15148 31447
rect 15212 30938 15240 33254
rect 15396 32994 15424 36314
rect 15568 33856 15620 33862
rect 15568 33798 15620 33804
rect 15476 33380 15528 33386
rect 15476 33322 15528 33328
rect 15488 33114 15516 33322
rect 15476 33108 15528 33114
rect 15476 33050 15528 33056
rect 15396 32966 15516 32994
rect 15384 32904 15436 32910
rect 15384 32846 15436 32852
rect 15290 32736 15346 32745
rect 15290 32671 15346 32680
rect 15304 32502 15332 32671
rect 15396 32570 15424 32846
rect 15384 32564 15436 32570
rect 15384 32506 15436 32512
rect 15292 32496 15344 32502
rect 15292 32438 15344 32444
rect 15396 32314 15424 32506
rect 15304 32286 15424 32314
rect 15304 31414 15332 32286
rect 15488 32212 15516 32966
rect 15396 32184 15516 32212
rect 15292 31408 15344 31414
rect 15292 31350 15344 31356
rect 15292 31204 15344 31210
rect 15292 31146 15344 31152
rect 15200 30932 15252 30938
rect 15200 30874 15252 30880
rect 15108 30728 15160 30734
rect 15108 30670 15160 30676
rect 15304 30546 15332 31146
rect 15120 30518 15332 30546
rect 15016 30184 15068 30190
rect 15016 30126 15068 30132
rect 15016 30048 15068 30054
rect 15016 29990 15068 29996
rect 15028 29782 15056 29990
rect 15016 29776 15068 29782
rect 15016 29718 15068 29724
rect 15120 29617 15148 30518
rect 15292 30116 15344 30122
rect 15292 30058 15344 30064
rect 15200 29708 15252 29714
rect 15200 29650 15252 29656
rect 15106 29608 15162 29617
rect 15106 29543 15162 29552
rect 15106 29336 15162 29345
rect 15106 29271 15162 29280
rect 15016 29164 15068 29170
rect 15016 29106 15068 29112
rect 14924 27600 14976 27606
rect 14924 27542 14976 27548
rect 14936 26994 14964 27542
rect 14924 26988 14976 26994
rect 14924 26930 14976 26936
rect 15028 26840 15056 29106
rect 15120 29102 15148 29271
rect 15108 29096 15160 29102
rect 15108 29038 15160 29044
rect 15108 28756 15160 28762
rect 15212 28744 15240 29650
rect 15304 29306 15332 30058
rect 15292 29300 15344 29306
rect 15292 29242 15344 29248
rect 15396 28948 15424 32184
rect 15474 31376 15530 31385
rect 15474 31311 15476 31320
rect 15528 31311 15530 31320
rect 15476 31282 15528 31288
rect 15580 30326 15608 33798
rect 15672 33658 15700 36654
rect 15764 36242 15792 37334
rect 15856 36310 15884 41262
rect 15936 40588 15988 40594
rect 15936 40530 15988 40536
rect 15948 39982 15976 40530
rect 16486 40080 16542 40089
rect 16486 40015 16542 40024
rect 16500 39982 16528 40015
rect 15936 39976 15988 39982
rect 15936 39918 15988 39924
rect 16488 39976 16540 39982
rect 16488 39918 16540 39924
rect 15936 39840 15988 39846
rect 15936 39782 15988 39788
rect 15948 38554 15976 39782
rect 16580 39500 16632 39506
rect 16580 39442 16632 39448
rect 16028 39432 16080 39438
rect 16028 39374 16080 39380
rect 16120 39432 16172 39438
rect 16120 39374 16172 39380
rect 15936 38548 15988 38554
rect 15936 38490 15988 38496
rect 15948 37874 15976 38490
rect 16040 38418 16068 39374
rect 16132 38894 16160 39374
rect 16212 39364 16264 39370
rect 16212 39306 16264 39312
rect 16120 38888 16172 38894
rect 16120 38830 16172 38836
rect 16224 38758 16252 39306
rect 16592 39302 16620 39442
rect 16304 39296 16356 39302
rect 16580 39296 16632 39302
rect 16304 39238 16356 39244
rect 16408 39256 16580 39284
rect 16316 38894 16344 39238
rect 16304 38888 16356 38894
rect 16304 38830 16356 38836
rect 16212 38752 16264 38758
rect 16212 38694 16264 38700
rect 16028 38412 16080 38418
rect 16028 38354 16080 38360
rect 16120 38412 16172 38418
rect 16120 38354 16172 38360
rect 16040 38010 16068 38354
rect 16028 38004 16080 38010
rect 16028 37946 16080 37952
rect 15936 37868 15988 37874
rect 15936 37810 15988 37816
rect 15936 37732 15988 37738
rect 15936 37674 15988 37680
rect 15948 36689 15976 37674
rect 16132 37330 16160 38354
rect 16120 37324 16172 37330
rect 16120 37266 16172 37272
rect 16028 36916 16080 36922
rect 16028 36858 16080 36864
rect 15934 36680 15990 36689
rect 15934 36615 15990 36624
rect 15844 36304 15896 36310
rect 15844 36246 15896 36252
rect 15752 36236 15804 36242
rect 15752 36178 15804 36184
rect 15936 36236 15988 36242
rect 15936 36178 15988 36184
rect 15948 35873 15976 36178
rect 15934 35864 15990 35873
rect 16040 35834 16068 36858
rect 15934 35799 15990 35808
rect 16028 35828 16080 35834
rect 16028 35770 16080 35776
rect 15844 35760 15896 35766
rect 15844 35702 15896 35708
rect 15856 33969 15884 35702
rect 16040 35154 16068 35770
rect 15936 35148 15988 35154
rect 15936 35090 15988 35096
rect 16028 35148 16080 35154
rect 16028 35090 16080 35096
rect 15948 34610 15976 35090
rect 16040 35018 16068 35090
rect 16028 35012 16080 35018
rect 16028 34954 16080 34960
rect 16040 34746 16068 34954
rect 16028 34740 16080 34746
rect 16028 34682 16080 34688
rect 15936 34604 15988 34610
rect 15936 34546 15988 34552
rect 15934 34096 15990 34105
rect 15934 34031 15990 34040
rect 15842 33960 15898 33969
rect 15842 33895 15898 33904
rect 15660 33652 15712 33658
rect 15660 33594 15712 33600
rect 15672 33386 15700 33594
rect 15660 33380 15712 33386
rect 15660 33322 15712 33328
rect 15660 32972 15712 32978
rect 15660 32914 15712 32920
rect 15568 30320 15620 30326
rect 15568 30262 15620 30268
rect 15672 30122 15700 32914
rect 15752 32768 15804 32774
rect 15752 32710 15804 32716
rect 15764 32026 15792 32710
rect 15856 32434 15884 33895
rect 15948 33862 15976 34031
rect 15936 33856 15988 33862
rect 15936 33798 15988 33804
rect 15844 32428 15896 32434
rect 15844 32370 15896 32376
rect 15842 32328 15898 32337
rect 15842 32263 15844 32272
rect 15896 32263 15898 32272
rect 15844 32234 15896 32240
rect 15752 32020 15804 32026
rect 15752 31962 15804 31968
rect 15856 31958 15884 32234
rect 15844 31952 15896 31958
rect 15844 31894 15896 31900
rect 15752 31884 15804 31890
rect 15752 31826 15804 31832
rect 15764 30841 15792 31826
rect 15842 31784 15898 31793
rect 15842 31719 15898 31728
rect 15856 31482 15884 31719
rect 15844 31476 15896 31482
rect 15844 31418 15896 31424
rect 15844 31204 15896 31210
rect 15844 31146 15896 31152
rect 15750 30832 15806 30841
rect 15750 30767 15806 30776
rect 15856 30682 15884 31146
rect 15764 30654 15884 30682
rect 15764 30598 15792 30654
rect 15752 30592 15804 30598
rect 15752 30534 15804 30540
rect 15660 30116 15712 30122
rect 15660 30058 15712 30064
rect 15476 30048 15528 30054
rect 15476 29990 15528 29996
rect 15488 29889 15516 29990
rect 15474 29880 15530 29889
rect 15672 29850 15700 30058
rect 15474 29815 15476 29824
rect 15528 29815 15530 29824
rect 15660 29844 15712 29850
rect 15476 29786 15528 29792
rect 15660 29786 15712 29792
rect 15488 29306 15516 29786
rect 15764 29730 15792 30534
rect 15842 30016 15898 30025
rect 15842 29951 15898 29960
rect 15580 29702 15792 29730
rect 15476 29300 15528 29306
rect 15476 29242 15528 29248
rect 15580 29073 15608 29702
rect 15660 29640 15712 29646
rect 15660 29582 15712 29588
rect 15672 29238 15700 29582
rect 15752 29504 15804 29510
rect 15752 29446 15804 29452
rect 15764 29306 15792 29446
rect 15752 29300 15804 29306
rect 15752 29242 15804 29248
rect 15660 29232 15712 29238
rect 15660 29174 15712 29180
rect 15566 29064 15622 29073
rect 15566 28999 15622 29008
rect 15396 28920 15516 28948
rect 15160 28716 15240 28744
rect 15108 28698 15160 28704
rect 15120 28665 15148 28698
rect 15106 28656 15162 28665
rect 15106 28591 15162 28600
rect 15200 28620 15252 28626
rect 15200 28562 15252 28568
rect 15212 28506 15240 28562
rect 15488 28506 15516 28920
rect 15120 28478 15240 28506
rect 15396 28478 15516 28506
rect 15120 28218 15148 28478
rect 15108 28212 15160 28218
rect 15108 28154 15160 28160
rect 15108 28076 15160 28082
rect 15160 28036 15240 28064
rect 15108 28018 15160 28024
rect 15108 27600 15160 27606
rect 15108 27542 15160 27548
rect 15120 27062 15148 27542
rect 15108 27056 15160 27062
rect 15108 26998 15160 27004
rect 14936 26812 15056 26840
rect 14936 24818 14964 26812
rect 15120 26518 15148 26998
rect 15108 26512 15160 26518
rect 15108 26454 15160 26460
rect 15016 26444 15068 26450
rect 15016 26386 15068 26392
rect 14924 24812 14976 24818
rect 14924 24754 14976 24760
rect 14924 24608 14976 24614
rect 14924 24550 14976 24556
rect 14832 24200 14884 24206
rect 14832 24142 14884 24148
rect 14936 23662 14964 24550
rect 14924 23656 14976 23662
rect 14924 23598 14976 23604
rect 14752 23446 14964 23474
rect 14832 23248 14884 23254
rect 14832 23190 14884 23196
rect 14648 22976 14700 22982
rect 14648 22918 14700 22924
rect 14660 22817 14688 22918
rect 14844 22817 14872 23190
rect 14646 22808 14702 22817
rect 14646 22743 14702 22752
rect 14830 22808 14886 22817
rect 14830 22743 14886 22752
rect 14738 22400 14794 22409
rect 14738 22335 14794 22344
rect 14752 22098 14780 22335
rect 14844 22234 14872 22743
rect 14832 22228 14884 22234
rect 14832 22170 14884 22176
rect 14740 22092 14792 22098
rect 14740 22034 14792 22040
rect 14556 21548 14608 21554
rect 14556 21490 14608 21496
rect 14278 20632 14334 20641
rect 13728 20596 13780 20602
rect 14278 20567 14334 20576
rect 13728 20538 13780 20544
rect 13636 19916 13688 19922
rect 13636 19858 13688 19864
rect 13648 19553 13676 19858
rect 13634 19544 13690 19553
rect 13634 19479 13690 19488
rect 13648 19378 13676 19479
rect 13636 19372 13688 19378
rect 13636 19314 13688 19320
rect 13740 18873 13768 20538
rect 13912 20528 13964 20534
rect 13910 20496 13912 20505
rect 13964 20496 13966 20505
rect 13910 20431 13966 20440
rect 14188 19372 14240 19378
rect 14188 19314 14240 19320
rect 13820 19168 13872 19174
rect 13820 19110 13872 19116
rect 13726 18864 13782 18873
rect 13832 18834 13860 19110
rect 13912 18896 13964 18902
rect 13912 18838 13964 18844
rect 13726 18799 13782 18808
rect 13820 18828 13872 18834
rect 13820 18770 13872 18776
rect 13820 18080 13872 18086
rect 13820 18022 13872 18028
rect 13832 17762 13860 18022
rect 13740 17746 13860 17762
rect 13728 17740 13860 17746
rect 13780 17734 13860 17740
rect 13728 17682 13780 17688
rect 13728 17604 13780 17610
rect 13924 17592 13952 18838
rect 13780 17564 13952 17592
rect 13728 17546 13780 17552
rect 13544 17196 13596 17202
rect 13544 17138 13596 17144
rect 13556 16658 13584 17138
rect 13544 16652 13596 16658
rect 13544 16594 13596 16600
rect 13820 16652 13872 16658
rect 13820 16594 13872 16600
rect 13636 16516 13688 16522
rect 13636 16458 13688 16464
rect 13728 16516 13780 16522
rect 13728 16458 13780 16464
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 13372 14618 13400 14962
rect 13360 14612 13412 14618
rect 13360 14554 13412 14560
rect 13372 13530 13400 14554
rect 13360 13524 13412 13530
rect 13360 13466 13412 13472
rect 13372 12782 13400 13466
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 13360 12232 13412 12238
rect 13360 12174 13412 12180
rect 13372 11898 13400 12174
rect 13360 11892 13412 11898
rect 13360 11834 13412 11840
rect 13266 8528 13322 8537
rect 13266 8463 13322 8472
rect 13452 7336 13504 7342
rect 13450 7304 13452 7313
rect 13504 7304 13506 7313
rect 13450 7239 13506 7248
rect 13648 5545 13676 16458
rect 13740 16182 13768 16458
rect 13832 16250 13860 16594
rect 14096 16584 14148 16590
rect 14096 16526 14148 16532
rect 14108 16250 14136 16526
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 14096 16244 14148 16250
rect 14096 16186 14148 16192
rect 13728 16176 13780 16182
rect 13728 16118 13780 16124
rect 13818 15056 13874 15065
rect 13818 14991 13820 15000
rect 13872 14991 13874 15000
rect 13820 14962 13872 14968
rect 13912 12844 13964 12850
rect 13912 12786 13964 12792
rect 13924 12306 13952 12786
rect 14004 12368 14056 12374
rect 14004 12310 14056 12316
rect 13728 12300 13780 12306
rect 13728 12242 13780 12248
rect 13912 12300 13964 12306
rect 13912 12242 13964 12248
rect 13740 11558 13768 12242
rect 13924 11830 13952 12242
rect 14016 11898 14044 12310
rect 14004 11892 14056 11898
rect 14004 11834 14056 11840
rect 13912 11824 13964 11830
rect 13912 11766 13964 11772
rect 13728 11552 13780 11558
rect 13728 11494 13780 11500
rect 13740 11150 13768 11494
rect 13728 11144 13780 11150
rect 13728 11086 13780 11092
rect 13634 5536 13690 5545
rect 13634 5471 13690 5480
rect 14002 4856 14058 4865
rect 14002 4791 14004 4800
rect 14056 4791 14058 4800
rect 14004 4762 14056 4768
rect 12440 4684 12492 4690
rect 12440 4626 12492 4632
rect 12452 4214 12480 4626
rect 12716 4616 12768 4622
rect 12716 4558 12768 4564
rect 12728 4282 12756 4558
rect 12716 4276 12768 4282
rect 12716 4218 12768 4224
rect 12440 4208 12492 4214
rect 12440 4150 12492 4156
rect 8392 4140 8444 4146
rect 8392 4082 8444 4088
rect 9220 4140 9272 4146
rect 9220 4082 9272 4088
rect 10140 4140 10192 4146
rect 10140 4082 10192 4088
rect 10692 4140 10744 4146
rect 10692 4082 10744 4088
rect 9232 800 9260 4082
rect 10152 800 10180 4082
rect 11980 3936 12032 3942
rect 11980 3878 12032 3884
rect 11060 2916 11112 2922
rect 11060 2858 11112 2864
rect 11072 800 11100 2858
rect 11992 800 12020 3878
rect 12452 3602 12480 4150
rect 12728 3942 12756 4218
rect 12716 3936 12768 3942
rect 12716 3878 12768 3884
rect 12440 3596 12492 3602
rect 12440 3538 12492 3544
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 12452 3194 12480 3538
rect 12440 3188 12492 3194
rect 12440 3130 12492 3136
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 12440 2916 12492 2922
rect 12440 2858 12492 2864
rect 12452 2650 12480 2858
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12544 2446 12572 2926
rect 12820 2854 12848 3538
rect 13820 3052 13872 3058
rect 13820 2994 13872 3000
rect 12808 2848 12860 2854
rect 12808 2790 12860 2796
rect 12532 2440 12584 2446
rect 12532 2382 12584 2388
rect 12820 898 12848 2790
rect 12820 870 12940 898
rect 12912 800 12940 870
rect 13832 800 13860 2994
rect 14200 2650 14228 19314
rect 14292 19310 14320 20567
rect 14740 20052 14792 20058
rect 14740 19994 14792 20000
rect 14462 19544 14518 19553
rect 14462 19479 14518 19488
rect 14280 19304 14332 19310
rect 14280 19246 14332 19252
rect 14476 19242 14504 19479
rect 14464 19236 14516 19242
rect 14464 19178 14516 19184
rect 14464 18828 14516 18834
rect 14464 18770 14516 18776
rect 14476 18465 14504 18770
rect 14752 18698 14780 19994
rect 14936 19718 14964 23446
rect 14924 19712 14976 19718
rect 14924 19654 14976 19660
rect 14936 19378 14964 19654
rect 14924 19372 14976 19378
rect 14924 19314 14976 19320
rect 14740 18692 14792 18698
rect 14740 18634 14792 18640
rect 14462 18456 14518 18465
rect 14752 18426 14780 18634
rect 14462 18391 14464 18400
rect 14516 18391 14518 18400
rect 14740 18420 14792 18426
rect 14464 18362 14516 18368
rect 14740 18362 14792 18368
rect 14924 18148 14976 18154
rect 14924 18090 14976 18096
rect 14830 18048 14886 18057
rect 14830 17983 14886 17992
rect 14844 17882 14872 17983
rect 14832 17876 14884 17882
rect 14832 17818 14884 17824
rect 14832 15972 14884 15978
rect 14832 15914 14884 15920
rect 14740 12776 14792 12782
rect 14740 12718 14792 12724
rect 14752 11898 14780 12718
rect 14740 11892 14792 11898
rect 14740 11834 14792 11840
rect 14738 5536 14794 5545
rect 14738 5471 14794 5480
rect 14278 4040 14334 4049
rect 14278 3975 14334 3984
rect 14292 3738 14320 3975
rect 14280 3732 14332 3738
rect 14280 3674 14332 3680
rect 14188 2644 14240 2650
rect 14188 2586 14240 2592
rect 14752 800 14780 5471
rect 14844 3194 14872 15914
rect 14936 12850 14964 18090
rect 15028 16658 15056 26386
rect 15108 26308 15160 26314
rect 15108 26250 15160 26256
rect 15120 25650 15148 26250
rect 15212 25838 15240 28036
rect 15292 26444 15344 26450
rect 15292 26386 15344 26392
rect 15304 26042 15332 26386
rect 15292 26036 15344 26042
rect 15292 25978 15344 25984
rect 15292 25900 15344 25906
rect 15292 25842 15344 25848
rect 15200 25832 15252 25838
rect 15200 25774 15252 25780
rect 15120 25622 15240 25650
rect 15108 25152 15160 25158
rect 15108 25094 15160 25100
rect 15120 24886 15148 25094
rect 15108 24880 15160 24886
rect 15106 24848 15108 24857
rect 15160 24848 15162 24857
rect 15106 24783 15162 24792
rect 15120 24757 15148 24783
rect 15212 24750 15240 25622
rect 15200 24744 15252 24750
rect 15200 24686 15252 24692
rect 15304 24342 15332 25842
rect 15396 25650 15424 28478
rect 15476 28416 15528 28422
rect 15476 28358 15528 28364
rect 15488 27402 15516 28358
rect 15476 27396 15528 27402
rect 15476 27338 15528 27344
rect 15580 27112 15608 28999
rect 15672 28393 15700 29174
rect 15752 29164 15804 29170
rect 15752 29106 15804 29112
rect 15658 28384 15714 28393
rect 15658 28319 15714 28328
rect 15672 27130 15700 28319
rect 15488 27084 15608 27112
rect 15660 27124 15712 27130
rect 15488 25752 15516 27084
rect 15660 27066 15712 27072
rect 15764 27010 15792 29106
rect 15856 27538 15884 29951
rect 15948 29170 15976 33798
rect 16028 32836 16080 32842
rect 16028 32778 16080 32784
rect 16040 32609 16068 32778
rect 16026 32600 16082 32609
rect 16026 32535 16028 32544
rect 16080 32535 16082 32544
rect 16028 32506 16080 32512
rect 16132 32026 16160 37266
rect 16224 37194 16252 38694
rect 16212 37188 16264 37194
rect 16212 37130 16264 37136
rect 16224 36825 16252 37130
rect 16210 36816 16266 36825
rect 16210 36751 16266 36760
rect 16304 36168 16356 36174
rect 16304 36110 16356 36116
rect 16316 35737 16344 36110
rect 16302 35728 16358 35737
rect 16408 35714 16436 39256
rect 16580 39238 16632 39244
rect 16764 39092 16816 39098
rect 16764 39034 16816 39040
rect 16488 38888 16540 38894
rect 16488 38830 16540 38836
rect 16580 38888 16632 38894
rect 16580 38830 16632 38836
rect 16670 38856 16726 38865
rect 16500 38321 16528 38830
rect 16486 38312 16542 38321
rect 16486 38247 16542 38256
rect 16592 37992 16620 38830
rect 16670 38791 16726 38800
rect 16500 37964 16620 37992
rect 16500 37618 16528 37964
rect 16578 37904 16634 37913
rect 16578 37839 16634 37848
rect 16592 37806 16620 37839
rect 16580 37800 16632 37806
rect 16580 37742 16632 37748
rect 16500 37590 16620 37618
rect 16486 36000 16542 36009
rect 16486 35935 16542 35944
rect 16500 35834 16528 35935
rect 16488 35828 16540 35834
rect 16488 35770 16540 35776
rect 16408 35686 16528 35714
rect 16302 35663 16358 35672
rect 16210 35048 16266 35057
rect 16210 34983 16266 34992
rect 16224 34542 16252 34983
rect 16316 34785 16344 35663
rect 16396 35080 16448 35086
rect 16396 35022 16448 35028
rect 16408 34921 16436 35022
rect 16394 34912 16450 34921
rect 16394 34847 16450 34856
rect 16302 34776 16358 34785
rect 16302 34711 16358 34720
rect 16396 34672 16448 34678
rect 16394 34640 16396 34649
rect 16448 34640 16450 34649
rect 16394 34575 16450 34584
rect 16212 34536 16264 34542
rect 16212 34478 16264 34484
rect 16304 34468 16356 34474
rect 16304 34410 16356 34416
rect 16212 34060 16264 34066
rect 16212 34002 16264 34008
rect 16224 33318 16252 34002
rect 16316 33425 16344 34410
rect 16302 33416 16358 33425
rect 16302 33351 16358 33360
rect 16212 33312 16264 33318
rect 16212 33254 16264 33260
rect 16396 33312 16448 33318
rect 16396 33254 16448 33260
rect 16408 32978 16436 33254
rect 16396 32972 16448 32978
rect 16396 32914 16448 32920
rect 16304 32768 16356 32774
rect 16304 32710 16356 32716
rect 16212 32496 16264 32502
rect 16212 32438 16264 32444
rect 16028 32020 16080 32026
rect 16028 31962 16080 31968
rect 16120 32020 16172 32026
rect 16120 31962 16172 31968
rect 16040 31793 16068 31962
rect 16120 31884 16172 31890
rect 16120 31826 16172 31832
rect 16026 31784 16082 31793
rect 16026 31719 16082 31728
rect 16026 31648 16082 31657
rect 16026 31583 16082 31592
rect 15936 29164 15988 29170
rect 15936 29106 15988 29112
rect 15936 28960 15988 28966
rect 15936 28902 15988 28908
rect 15948 28558 15976 28902
rect 15936 28552 15988 28558
rect 15936 28494 15988 28500
rect 15948 27985 15976 28494
rect 15934 27976 15990 27985
rect 15934 27911 15990 27920
rect 15936 27872 15988 27878
rect 15936 27814 15988 27820
rect 15844 27532 15896 27538
rect 15844 27474 15896 27480
rect 15856 27130 15884 27474
rect 15844 27124 15896 27130
rect 15844 27066 15896 27072
rect 15580 26982 15792 27010
rect 15580 26246 15608 26982
rect 15660 26920 15712 26926
rect 15660 26862 15712 26868
rect 15568 26240 15620 26246
rect 15568 26182 15620 26188
rect 15488 25724 15608 25752
rect 15396 25622 15516 25650
rect 15384 25356 15436 25362
rect 15384 25298 15436 25304
rect 15396 24954 15424 25298
rect 15384 24948 15436 24954
rect 15384 24890 15436 24896
rect 15488 24834 15516 25622
rect 15580 25498 15608 25724
rect 15672 25537 15700 26862
rect 15658 25528 15714 25537
rect 15568 25492 15620 25498
rect 15658 25463 15714 25472
rect 15568 25434 15620 25440
rect 15580 25226 15608 25434
rect 15568 25220 15620 25226
rect 15568 25162 15620 25168
rect 15488 24806 15608 24834
rect 15476 24744 15528 24750
rect 15476 24686 15528 24692
rect 15292 24336 15344 24342
rect 15292 24278 15344 24284
rect 15200 24268 15252 24274
rect 15200 24210 15252 24216
rect 15108 24064 15160 24070
rect 15106 24032 15108 24041
rect 15160 24032 15162 24041
rect 15106 23967 15162 23976
rect 15106 23896 15162 23905
rect 15106 23831 15108 23840
rect 15160 23831 15162 23840
rect 15108 23802 15160 23808
rect 15108 23588 15160 23594
rect 15108 23530 15160 23536
rect 15120 21894 15148 23530
rect 15212 23050 15240 24210
rect 15290 23352 15346 23361
rect 15290 23287 15346 23296
rect 15304 23118 15332 23287
rect 15292 23112 15344 23118
rect 15292 23054 15344 23060
rect 15200 23044 15252 23050
rect 15200 22986 15252 22992
rect 15304 22930 15332 23054
rect 15488 22982 15516 24686
rect 15580 23662 15608 24806
rect 15568 23656 15620 23662
rect 15568 23598 15620 23604
rect 15580 23304 15608 23598
rect 15672 23526 15700 25463
rect 15660 23520 15712 23526
rect 15660 23462 15712 23468
rect 15580 23276 15700 23304
rect 15568 23180 15620 23186
rect 15568 23122 15620 23128
rect 15212 22902 15332 22930
rect 15476 22976 15528 22982
rect 15476 22918 15528 22924
rect 15212 22166 15240 22902
rect 15580 22778 15608 23122
rect 15568 22772 15620 22778
rect 15568 22714 15620 22720
rect 15476 22704 15528 22710
rect 15476 22646 15528 22652
rect 15200 22160 15252 22166
rect 15198 22128 15200 22137
rect 15252 22128 15254 22137
rect 15198 22063 15254 22072
rect 15108 21888 15160 21894
rect 15108 21830 15160 21836
rect 15384 21684 15436 21690
rect 15384 21626 15436 21632
rect 15396 17746 15424 21626
rect 15488 20058 15516 22646
rect 15568 21888 15620 21894
rect 15566 21856 15568 21865
rect 15620 21856 15622 21865
rect 15566 21791 15622 21800
rect 15566 20632 15622 20641
rect 15566 20567 15568 20576
rect 15620 20567 15622 20576
rect 15568 20538 15620 20544
rect 15672 20466 15700 23276
rect 15764 22778 15792 26982
rect 15856 26314 15884 27066
rect 15844 26308 15896 26314
rect 15844 26250 15896 26256
rect 15948 25158 15976 27814
rect 15936 25152 15988 25158
rect 15936 25094 15988 25100
rect 15842 24440 15898 24449
rect 15842 24375 15898 24384
rect 15856 24206 15884 24375
rect 15844 24200 15896 24206
rect 15844 24142 15896 24148
rect 15752 22772 15804 22778
rect 15752 22714 15804 22720
rect 15934 22672 15990 22681
rect 15934 22607 15990 22616
rect 15948 22030 15976 22607
rect 16040 22098 16068 31583
rect 16132 28082 16160 31826
rect 16224 30938 16252 32438
rect 16316 32434 16344 32710
rect 16304 32428 16356 32434
rect 16304 32370 16356 32376
rect 16396 31952 16448 31958
rect 16396 31894 16448 31900
rect 16304 31408 16356 31414
rect 16304 31350 16356 31356
rect 16212 30932 16264 30938
rect 16212 30874 16264 30880
rect 16316 30870 16344 31350
rect 16408 31113 16436 31894
rect 16394 31104 16450 31113
rect 16394 31039 16450 31048
rect 16304 30864 16356 30870
rect 16304 30806 16356 30812
rect 16212 30796 16264 30802
rect 16212 30738 16264 30744
rect 16224 30598 16252 30738
rect 16212 30592 16264 30598
rect 16212 30534 16264 30540
rect 16224 30054 16252 30534
rect 16316 30394 16344 30806
rect 16304 30388 16356 30394
rect 16304 30330 16356 30336
rect 16408 30258 16436 31039
rect 16396 30252 16448 30258
rect 16396 30194 16448 30200
rect 16212 30048 16264 30054
rect 16212 29990 16264 29996
rect 16396 29844 16448 29850
rect 16396 29786 16448 29792
rect 16304 29776 16356 29782
rect 16304 29718 16356 29724
rect 16212 29028 16264 29034
rect 16212 28970 16264 28976
rect 16120 28076 16172 28082
rect 16120 28018 16172 28024
rect 16120 27532 16172 27538
rect 16120 27474 16172 27480
rect 16132 26586 16160 27474
rect 16224 27470 16252 28970
rect 16316 28762 16344 29718
rect 16304 28756 16356 28762
rect 16304 28698 16356 28704
rect 16316 28082 16344 28698
rect 16304 28076 16356 28082
rect 16304 28018 16356 28024
rect 16212 27464 16264 27470
rect 16212 27406 16264 27412
rect 16304 27464 16356 27470
rect 16304 27406 16356 27412
rect 16224 27130 16252 27406
rect 16212 27124 16264 27130
rect 16212 27066 16264 27072
rect 16120 26580 16172 26586
rect 16120 26522 16172 26528
rect 16132 26330 16160 26522
rect 16132 26302 16252 26330
rect 16120 26240 16172 26246
rect 16120 26182 16172 26188
rect 16132 25906 16160 26182
rect 16224 25922 16252 26302
rect 16316 26081 16344 27406
rect 16408 26926 16436 29786
rect 16396 26920 16448 26926
rect 16396 26862 16448 26868
rect 16396 26376 16448 26382
rect 16396 26318 16448 26324
rect 16302 26072 16358 26081
rect 16302 26007 16358 26016
rect 16120 25900 16172 25906
rect 16224 25894 16344 25922
rect 16120 25842 16172 25848
rect 16212 25832 16264 25838
rect 16210 25800 16212 25809
rect 16264 25800 16266 25809
rect 16210 25735 16266 25744
rect 16212 24812 16264 24818
rect 16212 24754 16264 24760
rect 16224 23730 16252 24754
rect 16212 23724 16264 23730
rect 16212 23666 16264 23672
rect 16212 23520 16264 23526
rect 16212 23462 16264 23468
rect 16120 22704 16172 22710
rect 16120 22646 16172 22652
rect 16028 22092 16080 22098
rect 16028 22034 16080 22040
rect 15936 22024 15988 22030
rect 15936 21966 15988 21972
rect 16040 21690 16068 22034
rect 15752 21684 15804 21690
rect 15752 21626 15804 21632
rect 16028 21684 16080 21690
rect 16028 21626 16080 21632
rect 15660 20460 15712 20466
rect 15660 20402 15712 20408
rect 15658 20360 15714 20369
rect 15658 20295 15714 20304
rect 15476 20052 15528 20058
rect 15476 19994 15528 20000
rect 15476 19236 15528 19242
rect 15476 19178 15528 19184
rect 15488 18970 15516 19178
rect 15476 18964 15528 18970
rect 15476 18906 15528 18912
rect 15488 18222 15516 18906
rect 15476 18216 15528 18222
rect 15476 18158 15528 18164
rect 15568 18216 15620 18222
rect 15568 18158 15620 18164
rect 15580 18057 15608 18158
rect 15566 18048 15622 18057
rect 15566 17983 15622 17992
rect 15384 17740 15436 17746
rect 15384 17682 15436 17688
rect 15292 17672 15344 17678
rect 15292 17614 15344 17620
rect 15304 17338 15332 17614
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 15396 17202 15424 17682
rect 15568 17536 15620 17542
rect 15568 17478 15620 17484
rect 15384 17196 15436 17202
rect 15384 17138 15436 17144
rect 15580 16726 15608 17478
rect 15568 16720 15620 16726
rect 15568 16662 15620 16668
rect 15016 16652 15068 16658
rect 15016 16594 15068 16600
rect 15028 15314 15056 16594
rect 15672 16046 15700 20295
rect 15764 18902 15792 21626
rect 16132 20466 16160 22646
rect 16028 20460 16080 20466
rect 16028 20402 16080 20408
rect 16120 20460 16172 20466
rect 16120 20402 16172 20408
rect 16040 19922 16068 20402
rect 16028 19916 16080 19922
rect 16028 19858 16080 19864
rect 15936 19712 15988 19718
rect 15936 19654 15988 19660
rect 15752 18896 15804 18902
rect 15804 18856 15884 18884
rect 15752 18838 15804 18844
rect 15752 18692 15804 18698
rect 15752 18634 15804 18640
rect 15660 16040 15712 16046
rect 15660 15982 15712 15988
rect 15384 15904 15436 15910
rect 15384 15846 15436 15852
rect 15396 15745 15424 15846
rect 15382 15736 15438 15745
rect 15382 15671 15438 15680
rect 15028 15286 15240 15314
rect 15212 15162 15240 15286
rect 15200 15156 15252 15162
rect 15200 15098 15252 15104
rect 15292 15020 15344 15026
rect 15292 14962 15344 14968
rect 15200 14884 15252 14890
rect 15200 14826 15252 14832
rect 15212 14482 15240 14826
rect 15304 14521 15332 14962
rect 15290 14512 15346 14521
rect 15200 14476 15252 14482
rect 15290 14447 15346 14456
rect 15200 14418 15252 14424
rect 15212 14074 15240 14418
rect 15304 14414 15332 14447
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 15200 14068 15252 14074
rect 15200 14010 15252 14016
rect 15304 14006 15332 14350
rect 15292 14000 15344 14006
rect 15292 13942 15344 13948
rect 15016 12980 15068 12986
rect 15016 12922 15068 12928
rect 14924 12844 14976 12850
rect 14924 12786 14976 12792
rect 15028 12306 15056 12922
rect 15108 12640 15160 12646
rect 15108 12582 15160 12588
rect 15120 12374 15148 12582
rect 15108 12368 15160 12374
rect 15108 12310 15160 12316
rect 15016 12300 15068 12306
rect 15016 12242 15068 12248
rect 15764 12102 15792 18634
rect 15856 17134 15884 18856
rect 15948 18834 15976 19654
rect 16040 19514 16068 19858
rect 16224 19854 16252 23462
rect 16316 23322 16344 25894
rect 16408 24614 16436 26318
rect 16500 25498 16528 35686
rect 16592 35601 16620 37590
rect 16684 36378 16712 38791
rect 16776 38457 16804 39034
rect 16854 38584 16910 38593
rect 16854 38519 16910 38528
rect 16762 38448 16818 38457
rect 16762 38383 16818 38392
rect 16868 38282 16896 38519
rect 16856 38276 16908 38282
rect 16856 38218 16908 38224
rect 16948 37800 17000 37806
rect 16946 37768 16948 37777
rect 17000 37768 17002 37777
rect 16946 37703 17002 37712
rect 16856 37664 16908 37670
rect 16856 37606 16908 37612
rect 16868 37262 16896 37606
rect 16946 37496 17002 37505
rect 16946 37431 17002 37440
rect 16960 37330 16988 37431
rect 16948 37324 17000 37330
rect 16948 37266 17000 37272
rect 16856 37256 16908 37262
rect 16854 37224 16856 37233
rect 16908 37224 16910 37233
rect 16854 37159 16910 37168
rect 16672 36372 16724 36378
rect 16672 36314 16724 36320
rect 16670 36272 16726 36281
rect 16670 36207 16672 36216
rect 16724 36207 16726 36216
rect 16672 36178 16724 36184
rect 17052 36122 17080 43608
rect 17314 40896 17370 40905
rect 17314 40831 17370 40840
rect 17328 40225 17356 40831
rect 17314 40216 17370 40225
rect 17132 40180 17184 40186
rect 17132 40122 17184 40128
rect 17236 40174 17314 40202
rect 17144 37942 17172 40122
rect 17132 37936 17184 37942
rect 17132 37878 17184 37884
rect 17144 37806 17172 37878
rect 17132 37800 17184 37806
rect 17132 37742 17184 37748
rect 17144 37262 17172 37742
rect 17132 37256 17184 37262
rect 17132 37198 17184 37204
rect 17144 36922 17172 37198
rect 17132 36916 17184 36922
rect 17132 36858 17184 36864
rect 17236 36666 17264 40174
rect 17314 40151 17370 40160
rect 17408 38344 17460 38350
rect 17408 38286 17460 38292
rect 17420 38049 17448 38286
rect 17406 38040 17462 38049
rect 17406 37975 17408 37984
rect 17460 37975 17462 37984
rect 17408 37946 17460 37952
rect 17314 37496 17370 37505
rect 17314 37431 17370 37440
rect 17328 37330 17356 37431
rect 17316 37324 17368 37330
rect 17316 37266 17368 37272
rect 17236 36638 17356 36666
rect 17420 36650 17448 37946
rect 17130 36408 17186 36417
rect 17130 36343 17186 36352
rect 16764 36100 16816 36106
rect 16764 36042 16816 36048
rect 16868 36094 17080 36122
rect 16670 35864 16726 35873
rect 16776 35834 16804 36042
rect 16670 35799 16672 35808
rect 16724 35799 16726 35808
rect 16764 35828 16816 35834
rect 16672 35770 16724 35776
rect 16764 35770 16816 35776
rect 16762 35728 16818 35737
rect 16762 35663 16818 35672
rect 16578 35592 16634 35601
rect 16578 35527 16634 35536
rect 16592 35306 16620 35527
rect 16592 35278 16712 35306
rect 16578 35184 16634 35193
rect 16578 35119 16634 35128
rect 16592 34746 16620 35119
rect 16580 34740 16632 34746
rect 16580 34682 16632 34688
rect 16580 33992 16632 33998
rect 16580 33934 16632 33940
rect 16592 33454 16620 33934
rect 16580 33448 16632 33454
rect 16580 33390 16632 33396
rect 16580 33312 16632 33318
rect 16580 33254 16632 33260
rect 16592 33046 16620 33254
rect 16580 33040 16632 33046
rect 16580 32982 16632 32988
rect 16592 32366 16620 32982
rect 16684 32774 16712 35278
rect 16776 34513 16804 35663
rect 16762 34504 16818 34513
rect 16762 34439 16818 34448
rect 16776 33046 16804 34439
rect 16868 34134 16896 36094
rect 16948 36032 17000 36038
rect 16948 35974 17000 35980
rect 16960 34202 16988 35974
rect 17144 35465 17172 36343
rect 17224 36304 17276 36310
rect 17224 36246 17276 36252
rect 17130 35456 17186 35465
rect 17052 35414 17130 35442
rect 16948 34196 17000 34202
rect 16948 34138 17000 34144
rect 16856 34128 16908 34134
rect 16856 34070 16908 34076
rect 16854 33824 16910 33833
rect 16854 33759 16910 33768
rect 16868 33658 16896 33759
rect 16856 33652 16908 33658
rect 16856 33594 16908 33600
rect 16960 33454 16988 34138
rect 16948 33448 17000 33454
rect 16948 33390 17000 33396
rect 16856 33380 16908 33386
rect 16856 33322 16908 33328
rect 16764 33040 16816 33046
rect 16764 32982 16816 32988
rect 16672 32768 16724 32774
rect 16672 32710 16724 32716
rect 16776 32570 16804 32982
rect 16764 32564 16816 32570
rect 16764 32506 16816 32512
rect 16580 32360 16632 32366
rect 16580 32302 16632 32308
rect 16580 32224 16632 32230
rect 16578 32192 16580 32201
rect 16632 32192 16634 32201
rect 16634 32150 16712 32178
rect 16578 32127 16634 32136
rect 16684 32026 16712 32150
rect 16672 32020 16724 32026
rect 16672 31962 16724 31968
rect 16764 31884 16816 31890
rect 16764 31826 16816 31832
rect 16580 31816 16632 31822
rect 16580 31758 16632 31764
rect 16592 31346 16620 31758
rect 16672 31680 16724 31686
rect 16776 31657 16804 31826
rect 16672 31622 16724 31628
rect 16762 31648 16818 31657
rect 16580 31340 16632 31346
rect 16580 31282 16632 31288
rect 16580 31136 16632 31142
rect 16684 31124 16712 31622
rect 16762 31583 16818 31592
rect 16868 31521 16896 33322
rect 16960 32978 16988 33390
rect 16948 32972 17000 32978
rect 16948 32914 17000 32920
rect 16854 31512 16910 31521
rect 16854 31447 16910 31456
rect 16764 31204 16816 31210
rect 16764 31146 16816 31152
rect 16632 31096 16712 31124
rect 16580 31078 16632 31084
rect 16592 30598 16620 31078
rect 16776 30920 16804 31146
rect 16684 30892 16804 30920
rect 16580 30592 16632 30598
rect 16580 30534 16632 30540
rect 16684 30410 16712 30892
rect 16856 30864 16908 30870
rect 16856 30806 16908 30812
rect 16764 30796 16816 30802
rect 16764 30738 16816 30744
rect 16592 30382 16712 30410
rect 16592 29782 16620 30382
rect 16672 30048 16724 30054
rect 16776 30025 16804 30738
rect 16672 29990 16724 29996
rect 16762 30016 16818 30025
rect 16684 29850 16712 29990
rect 16762 29951 16818 29960
rect 16672 29844 16724 29850
rect 16672 29786 16724 29792
rect 16580 29776 16632 29782
rect 16580 29718 16632 29724
rect 16578 29472 16634 29481
rect 16578 29407 16634 29416
rect 16592 29170 16620 29407
rect 16684 29306 16712 29786
rect 16672 29300 16724 29306
rect 16672 29242 16724 29248
rect 16580 29164 16632 29170
rect 16580 29106 16632 29112
rect 16592 27452 16620 29106
rect 16672 29096 16724 29102
rect 16672 29038 16724 29044
rect 16684 28937 16712 29038
rect 16670 28928 16726 28937
rect 16670 28863 16726 28872
rect 16764 28620 16816 28626
rect 16764 28562 16816 28568
rect 16672 28416 16724 28422
rect 16672 28358 16724 28364
rect 16684 28014 16712 28358
rect 16776 28150 16804 28562
rect 16764 28144 16816 28150
rect 16764 28086 16816 28092
rect 16672 28008 16724 28014
rect 16724 27968 16804 27996
rect 16672 27950 16724 27956
rect 16592 27424 16712 27452
rect 16578 27024 16634 27033
rect 16578 26959 16580 26968
rect 16632 26959 16634 26968
rect 16580 26930 16632 26936
rect 16592 25922 16620 26930
rect 16684 26926 16712 27424
rect 16776 27130 16804 27968
rect 16868 27606 16896 30806
rect 16960 30666 16988 32914
rect 16948 30660 17000 30666
rect 16948 30602 17000 30608
rect 17052 30546 17080 35414
rect 17130 35391 17186 35400
rect 17132 34944 17184 34950
rect 17132 34886 17184 34892
rect 17144 30802 17172 34886
rect 17236 31210 17264 36246
rect 17328 32570 17356 36638
rect 17408 36644 17460 36650
rect 17408 36586 17460 36592
rect 17420 36242 17448 36586
rect 17408 36236 17460 36242
rect 17408 36178 17460 36184
rect 17420 35834 17448 36178
rect 17408 35828 17460 35834
rect 17408 35770 17460 35776
rect 17408 35080 17460 35086
rect 17408 35022 17460 35028
rect 17420 33862 17448 35022
rect 17408 33856 17460 33862
rect 17408 33798 17460 33804
rect 17316 32564 17368 32570
rect 17316 32506 17368 32512
rect 17316 32428 17368 32434
rect 17316 32370 17368 32376
rect 17328 31278 17356 32370
rect 17408 32224 17460 32230
rect 17408 32166 17460 32172
rect 17316 31272 17368 31278
rect 17316 31214 17368 31220
rect 17224 31204 17276 31210
rect 17224 31146 17276 31152
rect 17132 30796 17184 30802
rect 17132 30738 17184 30744
rect 17052 30518 17356 30546
rect 17222 30424 17278 30433
rect 17222 30359 17278 30368
rect 17040 30116 17092 30122
rect 17040 30058 17092 30064
rect 17132 30116 17184 30122
rect 17132 30058 17184 30064
rect 16948 29640 17000 29646
rect 16948 29582 17000 29588
rect 16856 27600 16908 27606
rect 16856 27542 16908 27548
rect 16856 27328 16908 27334
rect 16856 27270 16908 27276
rect 16764 27124 16816 27130
rect 16764 27066 16816 27072
rect 16672 26920 16724 26926
rect 16672 26862 16724 26868
rect 16672 26580 16724 26586
rect 16672 26522 16724 26528
rect 16684 26450 16712 26522
rect 16672 26444 16724 26450
rect 16672 26386 16724 26392
rect 16684 26042 16712 26386
rect 16776 26217 16804 27066
rect 16868 26450 16896 27270
rect 16960 27033 16988 29582
rect 17052 29306 17080 30058
rect 17040 29300 17092 29306
rect 17040 29242 17092 29248
rect 17144 29238 17172 30058
rect 17132 29232 17184 29238
rect 17132 29174 17184 29180
rect 17130 29064 17186 29073
rect 17130 28999 17132 29008
rect 17184 28999 17186 29008
rect 17132 28970 17184 28976
rect 17038 28928 17094 28937
rect 17038 28863 17094 28872
rect 17052 27878 17080 28863
rect 17236 28744 17264 30359
rect 17144 28716 17264 28744
rect 17040 27872 17092 27878
rect 17040 27814 17092 27820
rect 16946 27024 17002 27033
rect 16946 26959 17002 26968
rect 16856 26444 16908 26450
rect 16856 26386 16908 26392
rect 16762 26208 16818 26217
rect 16762 26143 16818 26152
rect 16672 26036 16724 26042
rect 16672 25978 16724 25984
rect 16592 25894 16896 25922
rect 16580 25832 16632 25838
rect 16580 25774 16632 25780
rect 16488 25492 16540 25498
rect 16488 25434 16540 25440
rect 16500 25158 16528 25189
rect 16488 25152 16540 25158
rect 16486 25120 16488 25129
rect 16540 25120 16542 25129
rect 16486 25055 16542 25064
rect 16500 24750 16528 25055
rect 16488 24744 16540 24750
rect 16488 24686 16540 24692
rect 16396 24608 16448 24614
rect 16396 24550 16448 24556
rect 16396 24268 16448 24274
rect 16396 24210 16448 24216
rect 16408 23526 16436 24210
rect 16592 24138 16620 25774
rect 16672 25356 16724 25362
rect 16672 25298 16724 25304
rect 16684 24585 16712 25298
rect 16762 24848 16818 24857
rect 16762 24783 16818 24792
rect 16776 24750 16804 24783
rect 16764 24744 16816 24750
rect 16764 24686 16816 24692
rect 16670 24576 16726 24585
rect 16670 24511 16726 24520
rect 16672 24268 16724 24274
rect 16672 24210 16724 24216
rect 16580 24132 16632 24138
rect 16580 24074 16632 24080
rect 16684 23798 16712 24210
rect 16776 23866 16804 24686
rect 16764 23860 16816 23866
rect 16764 23802 16816 23808
rect 16672 23792 16724 23798
rect 16868 23746 16896 25894
rect 16948 25492 17000 25498
rect 16948 25434 17000 25440
rect 16960 25362 16988 25434
rect 16948 25356 17000 25362
rect 16948 25298 17000 25304
rect 17040 25356 17092 25362
rect 17040 25298 17092 25304
rect 16948 24880 17000 24886
rect 17052 24857 17080 25298
rect 16948 24822 17000 24828
rect 17038 24848 17094 24857
rect 16960 24410 16988 24822
rect 17038 24783 17094 24792
rect 16948 24404 17000 24410
rect 16948 24346 17000 24352
rect 17144 24290 17172 28716
rect 17224 28076 17276 28082
rect 17224 28018 17276 28024
rect 17236 26586 17264 28018
rect 17328 27674 17356 30518
rect 17420 30326 17448 32166
rect 17408 30320 17460 30326
rect 17408 30262 17460 30268
rect 17408 29300 17460 29306
rect 17408 29242 17460 29248
rect 17316 27668 17368 27674
rect 17316 27610 17368 27616
rect 17420 27606 17448 29242
rect 17408 27600 17460 27606
rect 17408 27542 17460 27548
rect 17420 27130 17448 27542
rect 17408 27124 17460 27130
rect 17328 27084 17408 27112
rect 17224 26580 17276 26586
rect 17224 26522 17276 26528
rect 17328 26518 17356 27084
rect 17408 27066 17460 27072
rect 17316 26512 17368 26518
rect 17316 26454 17368 26460
rect 17316 26376 17368 26382
rect 17316 26318 17368 26324
rect 17224 26308 17276 26314
rect 17224 26250 17276 26256
rect 17236 25362 17264 26250
rect 17328 25945 17356 26318
rect 17314 25936 17370 25945
rect 17314 25871 17370 25880
rect 17224 25356 17276 25362
rect 17224 25298 17276 25304
rect 17236 25265 17264 25298
rect 17222 25256 17278 25265
rect 17222 25191 17278 25200
rect 17328 25106 17356 25871
rect 17512 25480 17540 46378
rect 17592 37188 17644 37194
rect 17592 37130 17644 37136
rect 17604 36650 17632 37130
rect 17592 36644 17644 36650
rect 17592 36586 17644 36592
rect 17696 36310 17724 76842
rect 19340 76832 19392 76838
rect 19340 76774 19392 76780
rect 17776 76424 17828 76430
rect 17776 76366 17828 76372
rect 17788 75750 17816 76366
rect 17868 76288 17920 76294
rect 17868 76230 17920 76236
rect 17880 76022 17908 76230
rect 17868 76016 17920 76022
rect 17868 75958 17920 75964
rect 19352 75954 19380 76774
rect 19248 75948 19300 75954
rect 19248 75890 19300 75896
rect 19340 75948 19392 75954
rect 19340 75890 19392 75896
rect 17776 75744 17828 75750
rect 17776 75686 17828 75692
rect 17788 75041 17816 75686
rect 19260 75206 19288 75890
rect 19248 75200 19300 75206
rect 19248 75142 19300 75148
rect 17774 75032 17830 75041
rect 17774 74967 17830 74976
rect 19260 73114 19288 75142
rect 19444 74662 19472 76894
rect 19580 76732 19876 76752
rect 19636 76730 19660 76732
rect 19716 76730 19740 76732
rect 19796 76730 19820 76732
rect 19658 76678 19660 76730
rect 19722 76678 19734 76730
rect 19796 76678 19798 76730
rect 19636 76676 19660 76678
rect 19716 76676 19740 76678
rect 19796 76676 19820 76678
rect 19580 76656 19876 76676
rect 20076 75744 20128 75750
rect 20076 75686 20128 75692
rect 19580 75644 19876 75664
rect 19636 75642 19660 75644
rect 19716 75642 19740 75644
rect 19796 75642 19820 75644
rect 19658 75590 19660 75642
rect 19722 75590 19734 75642
rect 19796 75590 19798 75642
rect 19636 75588 19660 75590
rect 19716 75588 19740 75590
rect 19796 75588 19820 75590
rect 19580 75568 19876 75588
rect 19982 75168 20038 75177
rect 19982 75103 20038 75112
rect 19892 74792 19944 74798
rect 19892 74734 19944 74740
rect 19432 74656 19484 74662
rect 19432 74598 19484 74604
rect 19580 74556 19876 74576
rect 19636 74554 19660 74556
rect 19716 74554 19740 74556
rect 19796 74554 19820 74556
rect 19658 74502 19660 74554
rect 19722 74502 19734 74554
rect 19796 74502 19798 74554
rect 19636 74500 19660 74502
rect 19716 74500 19740 74502
rect 19796 74500 19820 74502
rect 19580 74480 19876 74500
rect 19904 74390 19932 74734
rect 19892 74384 19944 74390
rect 19892 74326 19944 74332
rect 19580 73468 19876 73488
rect 19636 73466 19660 73468
rect 19716 73466 19740 73468
rect 19796 73466 19820 73468
rect 19658 73414 19660 73466
rect 19722 73414 19734 73466
rect 19796 73414 19798 73466
rect 19636 73412 19660 73414
rect 19716 73412 19740 73414
rect 19796 73412 19820 73414
rect 19580 73392 19876 73412
rect 19260 73086 19472 73114
rect 19340 73024 19392 73030
rect 19338 72992 19340 73001
rect 19392 72992 19394 73001
rect 19338 72927 19394 72936
rect 19444 72622 19472 73086
rect 19432 72616 19484 72622
rect 19338 72584 19394 72593
rect 19432 72558 19484 72564
rect 19338 72519 19340 72528
rect 19392 72519 19394 72528
rect 19340 72490 19392 72496
rect 19444 72162 19472 72558
rect 19580 72380 19876 72400
rect 19636 72378 19660 72380
rect 19716 72378 19740 72380
rect 19796 72378 19820 72380
rect 19658 72326 19660 72378
rect 19722 72326 19734 72378
rect 19796 72326 19798 72378
rect 19636 72324 19660 72326
rect 19716 72324 19740 72326
rect 19796 72324 19820 72326
rect 19580 72304 19876 72324
rect 19444 72134 19564 72162
rect 19536 71942 19564 72134
rect 19524 71936 19576 71942
rect 19522 71904 19524 71913
rect 19576 71904 19578 71913
rect 19522 71839 19578 71848
rect 18234 71496 18290 71505
rect 18234 71431 18290 71440
rect 18052 60104 18104 60110
rect 18052 60046 18104 60052
rect 17866 59800 17922 59809
rect 17866 59735 17868 59744
rect 17920 59735 17922 59744
rect 17868 59706 17920 59712
rect 17958 59392 18014 59401
rect 17958 59327 18014 59336
rect 17868 59016 17920 59022
rect 17868 58958 17920 58964
rect 17776 58880 17828 58886
rect 17776 58822 17828 58828
rect 17788 56409 17816 58822
rect 17880 57594 17908 58958
rect 17868 57588 17920 57594
rect 17868 57530 17920 57536
rect 17868 57316 17920 57322
rect 17868 57258 17920 57264
rect 17880 56846 17908 57258
rect 17868 56840 17920 56846
rect 17866 56808 17868 56817
rect 17920 56808 17922 56817
rect 17866 56743 17922 56752
rect 17866 56536 17922 56545
rect 17866 56471 17868 56480
rect 17920 56471 17922 56480
rect 17868 56442 17920 56448
rect 17774 56400 17830 56409
rect 17774 56335 17830 56344
rect 17788 54262 17816 56335
rect 17868 55276 17920 55282
rect 17868 55218 17920 55224
rect 17776 54256 17828 54262
rect 17776 54198 17828 54204
rect 17788 53038 17816 54198
rect 17880 53553 17908 55218
rect 17866 53544 17922 53553
rect 17972 53514 18000 59327
rect 18064 59022 18092 60046
rect 18144 59424 18196 59430
rect 18144 59366 18196 59372
rect 18052 59016 18104 59022
rect 18052 58958 18104 58964
rect 18052 58880 18104 58886
rect 18156 58868 18184 59366
rect 18104 58840 18184 58868
rect 18052 58822 18104 58828
rect 18156 58342 18184 58840
rect 18144 58336 18196 58342
rect 18144 58278 18196 58284
rect 18052 57928 18104 57934
rect 18052 57870 18104 57876
rect 18064 57372 18092 57870
rect 18156 57526 18184 58278
rect 18144 57520 18196 57526
rect 18144 57462 18196 57468
rect 18144 57384 18196 57390
rect 18064 57344 18144 57372
rect 18144 57326 18196 57332
rect 18052 57248 18104 57254
rect 18052 57190 18104 57196
rect 18064 56438 18092 57190
rect 18156 56817 18184 57326
rect 18142 56808 18198 56817
rect 18142 56743 18144 56752
rect 18196 56743 18198 56752
rect 18144 56714 18196 56720
rect 18052 56432 18104 56438
rect 18052 56374 18104 56380
rect 18052 55140 18104 55146
rect 18052 55082 18104 55088
rect 18064 54806 18092 55082
rect 18052 54800 18104 54806
rect 18052 54742 18104 54748
rect 18064 54330 18092 54742
rect 18052 54324 18104 54330
rect 18052 54266 18104 54272
rect 17866 53479 17922 53488
rect 17960 53508 18012 53514
rect 17960 53450 18012 53456
rect 18248 53174 18276 71431
rect 19580 71292 19876 71312
rect 19636 71290 19660 71292
rect 19716 71290 19740 71292
rect 19796 71290 19820 71292
rect 19658 71238 19660 71290
rect 19722 71238 19734 71290
rect 19796 71238 19798 71290
rect 19636 71236 19660 71238
rect 19716 71236 19740 71238
rect 19796 71236 19820 71238
rect 19580 71216 19876 71236
rect 19580 70204 19876 70224
rect 19636 70202 19660 70204
rect 19716 70202 19740 70204
rect 19796 70202 19820 70204
rect 19658 70150 19660 70202
rect 19722 70150 19734 70202
rect 19796 70150 19798 70202
rect 19636 70148 19660 70150
rect 19716 70148 19740 70150
rect 19796 70148 19820 70150
rect 19580 70128 19876 70148
rect 19580 69116 19876 69136
rect 19636 69114 19660 69116
rect 19716 69114 19740 69116
rect 19796 69114 19820 69116
rect 19658 69062 19660 69114
rect 19722 69062 19734 69114
rect 19796 69062 19798 69114
rect 19636 69060 19660 69062
rect 19716 69060 19740 69062
rect 19796 69060 19820 69062
rect 19580 69040 19876 69060
rect 19580 68028 19876 68048
rect 19636 68026 19660 68028
rect 19716 68026 19740 68028
rect 19796 68026 19820 68028
rect 19658 67974 19660 68026
rect 19722 67974 19734 68026
rect 19796 67974 19798 68026
rect 19636 67972 19660 67974
rect 19716 67972 19740 67974
rect 19796 67972 19820 67974
rect 19580 67952 19876 67972
rect 19340 67924 19392 67930
rect 19340 67866 19392 67872
rect 19352 67833 19380 67866
rect 19338 67824 19394 67833
rect 19338 67759 19394 67768
rect 19580 66940 19876 66960
rect 19636 66938 19660 66940
rect 19716 66938 19740 66940
rect 19796 66938 19820 66940
rect 19658 66886 19660 66938
rect 19722 66886 19734 66938
rect 19796 66886 19798 66938
rect 19636 66884 19660 66886
rect 19716 66884 19740 66886
rect 19796 66884 19820 66886
rect 19580 66864 19876 66884
rect 19580 65852 19876 65872
rect 19636 65850 19660 65852
rect 19716 65850 19740 65852
rect 19796 65850 19820 65852
rect 19658 65798 19660 65850
rect 19722 65798 19734 65850
rect 19796 65798 19798 65850
rect 19636 65796 19660 65798
rect 19716 65796 19740 65798
rect 19796 65796 19820 65798
rect 19580 65776 19876 65796
rect 19580 64764 19876 64784
rect 19636 64762 19660 64764
rect 19716 64762 19740 64764
rect 19796 64762 19820 64764
rect 19658 64710 19660 64762
rect 19722 64710 19734 64762
rect 19796 64710 19798 64762
rect 19636 64708 19660 64710
rect 19716 64708 19740 64710
rect 19796 64708 19820 64710
rect 19580 64688 19876 64708
rect 19580 63676 19876 63696
rect 19636 63674 19660 63676
rect 19716 63674 19740 63676
rect 19796 63674 19820 63676
rect 19658 63622 19660 63674
rect 19722 63622 19734 63674
rect 19796 63622 19798 63674
rect 19636 63620 19660 63622
rect 19716 63620 19740 63622
rect 19796 63620 19820 63622
rect 19580 63600 19876 63620
rect 18604 63232 18656 63238
rect 18604 63174 18656 63180
rect 18880 63232 18932 63238
rect 18880 63174 18932 63180
rect 18616 62762 18644 63174
rect 18892 62898 18920 63174
rect 18880 62892 18932 62898
rect 18880 62834 18932 62840
rect 18604 62756 18656 62762
rect 18604 62698 18656 62704
rect 18616 62642 18644 62698
rect 18524 62614 18644 62642
rect 18524 62354 18552 62614
rect 18892 62354 18920 62834
rect 19580 62588 19876 62608
rect 19636 62586 19660 62588
rect 19716 62586 19740 62588
rect 19796 62586 19820 62588
rect 19658 62534 19660 62586
rect 19722 62534 19734 62586
rect 19796 62534 19798 62586
rect 19636 62532 19660 62534
rect 19716 62532 19740 62534
rect 19796 62532 19820 62534
rect 19580 62512 19876 62532
rect 18512 62348 18564 62354
rect 18512 62290 18564 62296
rect 18880 62348 18932 62354
rect 18880 62290 18932 62296
rect 18420 62280 18472 62286
rect 18420 62222 18472 62228
rect 18432 62121 18460 62222
rect 18418 62112 18474 62121
rect 18418 62047 18474 62056
rect 18432 61946 18460 62047
rect 18420 61940 18472 61946
rect 18420 61882 18472 61888
rect 18432 60858 18460 61882
rect 18524 61606 18552 62290
rect 18892 61606 18920 62290
rect 19996 62257 20024 75103
rect 20088 74866 20116 75686
rect 20076 74860 20128 74866
rect 20076 74802 20128 74808
rect 20076 74656 20128 74662
rect 20076 74598 20128 74604
rect 20088 62898 20116 74598
rect 20272 74497 20300 79200
rect 21192 77926 21220 79200
rect 21180 77920 21232 77926
rect 21180 77862 21232 77868
rect 21088 76968 21140 76974
rect 21088 76910 21140 76916
rect 20904 76832 20956 76838
rect 20904 76774 20956 76780
rect 20536 76356 20588 76362
rect 20536 76298 20588 76304
rect 20548 74798 20576 76298
rect 20536 74792 20588 74798
rect 20536 74734 20588 74740
rect 20812 74656 20864 74662
rect 20812 74598 20864 74604
rect 20258 74488 20314 74497
rect 20258 74423 20314 74432
rect 20718 68368 20774 68377
rect 20718 68303 20774 68312
rect 20352 63436 20404 63442
rect 20352 63378 20404 63384
rect 20364 63034 20392 63378
rect 20352 63028 20404 63034
rect 20352 62970 20404 62976
rect 20076 62892 20128 62898
rect 20076 62834 20128 62840
rect 19062 62248 19118 62257
rect 19062 62183 19064 62192
rect 19116 62183 19118 62192
rect 19982 62248 20038 62257
rect 19982 62183 20038 62192
rect 19064 62154 19116 62160
rect 18512 61600 18564 61606
rect 18512 61542 18564 61548
rect 18880 61600 18932 61606
rect 18880 61542 18932 61548
rect 20076 61600 20128 61606
rect 20076 61542 20128 61548
rect 18420 60852 18472 60858
rect 18420 60794 18472 60800
rect 18328 58880 18380 58886
rect 18328 58822 18380 58828
rect 18340 58041 18368 58822
rect 18326 58032 18382 58041
rect 18326 57967 18382 57976
rect 18328 56908 18380 56914
rect 18328 56850 18380 56856
rect 18340 56234 18368 56850
rect 18328 56228 18380 56234
rect 18328 56170 18380 56176
rect 18340 55826 18368 56170
rect 18418 55992 18474 56001
rect 18418 55927 18474 55936
rect 18328 55820 18380 55826
rect 18328 55762 18380 55768
rect 18432 55758 18460 55927
rect 18420 55752 18472 55758
rect 18420 55694 18472 55700
rect 18524 54602 18552 61542
rect 18604 59968 18656 59974
rect 18604 59910 18656 59916
rect 18616 59566 18644 59910
rect 18604 59560 18656 59566
rect 18602 59528 18604 59537
rect 18656 59528 18658 59537
rect 18602 59463 18658 59472
rect 18696 56840 18748 56846
rect 18696 56782 18748 56788
rect 18708 55962 18736 56782
rect 18696 55956 18748 55962
rect 18696 55898 18748 55904
rect 18788 54664 18840 54670
rect 18788 54606 18840 54612
rect 18512 54596 18564 54602
rect 18512 54538 18564 54544
rect 18326 53952 18382 53961
rect 18326 53887 18382 53896
rect 18236 53168 18288 53174
rect 18236 53110 18288 53116
rect 17776 53032 17828 53038
rect 17776 52974 17828 52980
rect 18144 53032 18196 53038
rect 18144 52974 18196 52980
rect 17868 52896 17920 52902
rect 17868 52838 17920 52844
rect 17776 52488 17828 52494
rect 17776 52430 17828 52436
rect 17788 51950 17816 52430
rect 17776 51944 17828 51950
rect 17776 51886 17828 51892
rect 17788 51542 17816 51886
rect 17880 51882 17908 52838
rect 17960 52556 18012 52562
rect 17960 52498 18012 52504
rect 17972 52086 18000 52498
rect 18156 52358 18184 52974
rect 18340 52698 18368 53887
rect 18524 53038 18552 54538
rect 18800 54126 18828 54606
rect 18604 54120 18656 54126
rect 18604 54062 18656 54068
rect 18788 54120 18840 54126
rect 18788 54062 18840 54068
rect 18616 53718 18644 54062
rect 18604 53712 18656 53718
rect 18604 53654 18656 53660
rect 18616 53446 18644 53654
rect 18604 53440 18656 53446
rect 18602 53408 18604 53417
rect 18656 53408 18658 53417
rect 18602 53343 18658 53352
rect 18616 53242 18644 53343
rect 18604 53236 18656 53242
rect 18604 53178 18656 53184
rect 18512 53032 18564 53038
rect 18512 52974 18564 52980
rect 18328 52692 18380 52698
rect 18328 52634 18380 52640
rect 18144 52352 18196 52358
rect 18144 52294 18196 52300
rect 17960 52080 18012 52086
rect 17960 52022 18012 52028
rect 17868 51876 17920 51882
rect 17868 51818 17920 51824
rect 17776 51536 17828 51542
rect 17774 51504 17776 51513
rect 17828 51504 17830 51513
rect 17774 51439 17830 51448
rect 17868 51468 17920 51474
rect 17788 51413 17816 51439
rect 17972 51456 18000 52022
rect 18340 52018 18368 52634
rect 18328 52012 18380 52018
rect 18328 51954 18380 51960
rect 18420 51876 18472 51882
rect 18420 51818 18472 51824
rect 17972 51428 18092 51456
rect 17868 51410 17920 51416
rect 17880 50930 17908 51410
rect 17960 51332 18012 51338
rect 17960 51274 18012 51280
rect 17868 50924 17920 50930
rect 17868 50866 17920 50872
rect 17880 50522 17908 50866
rect 17972 50726 18000 51274
rect 17960 50720 18012 50726
rect 17960 50662 18012 50668
rect 17868 50516 17920 50522
rect 17868 50458 17920 50464
rect 17960 50380 18012 50386
rect 17960 50322 18012 50328
rect 17972 50266 18000 50322
rect 18064 50318 18092 51428
rect 18432 51241 18460 51818
rect 18418 51232 18474 51241
rect 18418 51167 18474 51176
rect 18418 50824 18474 50833
rect 18236 50788 18288 50794
rect 18418 50759 18474 50768
rect 18236 50730 18288 50736
rect 18144 50720 18196 50726
rect 18144 50662 18196 50668
rect 17880 50238 18000 50266
rect 18052 50312 18104 50318
rect 18052 50254 18104 50260
rect 17880 49434 17908 50238
rect 18156 49994 18184 50662
rect 18064 49966 18184 49994
rect 18248 49978 18276 50730
rect 18236 49972 18288 49978
rect 17868 49428 17920 49434
rect 17868 49370 17920 49376
rect 17868 49224 17920 49230
rect 17868 49166 17920 49172
rect 17776 49088 17828 49094
rect 17776 49030 17828 49036
rect 17788 44441 17816 49030
rect 17880 48890 17908 49166
rect 17868 48884 17920 48890
rect 17868 48826 17920 48832
rect 18064 46073 18092 49966
rect 18236 49914 18288 49920
rect 18144 49904 18196 49910
rect 18144 49846 18196 49852
rect 18050 46064 18106 46073
rect 18050 45999 18106 46008
rect 17774 44432 17830 44441
rect 17774 44367 17830 44376
rect 17776 43852 17828 43858
rect 17776 43794 17828 43800
rect 17788 43450 17816 43794
rect 17776 43444 17828 43450
rect 17776 43386 17828 43392
rect 17866 40624 17922 40633
rect 17866 40559 17868 40568
rect 17920 40559 17922 40568
rect 17868 40530 17920 40536
rect 17776 40520 17828 40526
rect 17776 40462 17828 40468
rect 17788 39438 17816 40462
rect 17880 40186 17908 40530
rect 17868 40180 17920 40186
rect 17868 40122 17920 40128
rect 17868 39976 17920 39982
rect 17866 39944 17868 39953
rect 17920 39944 17922 39953
rect 17866 39879 17922 39888
rect 17776 39432 17828 39438
rect 17776 39374 17828 39380
rect 17788 39098 17816 39374
rect 18052 39364 18104 39370
rect 18052 39306 18104 39312
rect 17776 39092 17828 39098
rect 17776 39034 17828 39040
rect 17788 36922 17816 39034
rect 18064 38962 18092 39306
rect 18052 38956 18104 38962
rect 18052 38898 18104 38904
rect 18052 38480 18104 38486
rect 18052 38422 18104 38428
rect 17868 38344 17920 38350
rect 17868 38286 17920 38292
rect 17880 38010 17908 38286
rect 17868 38004 17920 38010
rect 17868 37946 17920 37952
rect 17960 37664 18012 37670
rect 17880 37612 17960 37618
rect 17880 37606 18012 37612
rect 17880 37590 18000 37606
rect 17776 36916 17828 36922
rect 17776 36858 17828 36864
rect 17880 36378 17908 37590
rect 18064 37466 18092 38422
rect 18052 37460 18104 37466
rect 18052 37402 18104 37408
rect 17960 37392 18012 37398
rect 17960 37334 18012 37340
rect 17868 36372 17920 36378
rect 17868 36314 17920 36320
rect 17684 36304 17736 36310
rect 17684 36246 17736 36252
rect 17866 36272 17922 36281
rect 17866 36207 17868 36216
rect 17920 36207 17922 36216
rect 17868 36178 17920 36184
rect 17684 36100 17736 36106
rect 17684 36042 17736 36048
rect 17592 35284 17644 35290
rect 17592 35226 17644 35232
rect 17604 34542 17632 35226
rect 17696 35222 17724 36042
rect 17972 35834 18000 37334
rect 18050 36136 18106 36145
rect 18050 36071 18106 36080
rect 17960 35828 18012 35834
rect 17960 35770 18012 35776
rect 17960 35692 18012 35698
rect 17960 35634 18012 35640
rect 17972 35290 18000 35634
rect 17960 35284 18012 35290
rect 17960 35226 18012 35232
rect 18064 35222 18092 36071
rect 17684 35216 17736 35222
rect 17684 35158 17736 35164
rect 18052 35216 18104 35222
rect 18052 35158 18104 35164
rect 17960 35080 18012 35086
rect 17960 35022 18012 35028
rect 17592 34536 17644 34542
rect 17592 34478 17644 34484
rect 17774 34504 17830 34513
rect 17604 32994 17632 34478
rect 17774 34439 17830 34448
rect 17684 33992 17736 33998
rect 17684 33934 17736 33940
rect 17696 33386 17724 33934
rect 17684 33380 17736 33386
rect 17684 33322 17736 33328
rect 17696 33114 17724 33322
rect 17684 33108 17736 33114
rect 17684 33050 17736 33056
rect 17788 33046 17816 34439
rect 17972 34377 18000 35022
rect 17958 34368 18014 34377
rect 17958 34303 18014 34312
rect 17960 34128 18012 34134
rect 17958 34096 17960 34105
rect 18012 34096 18014 34105
rect 17958 34031 18014 34040
rect 17868 33924 17920 33930
rect 17868 33866 17920 33872
rect 17776 33040 17828 33046
rect 17682 33008 17738 33017
rect 17604 32966 17682 32994
rect 17776 32982 17828 32988
rect 17682 32943 17738 32952
rect 17592 32904 17644 32910
rect 17592 32846 17644 32852
rect 17604 32366 17632 32846
rect 17592 32360 17644 32366
rect 17592 32302 17644 32308
rect 17592 32224 17644 32230
rect 17592 32166 17644 32172
rect 17604 31278 17632 32166
rect 17696 31414 17724 32943
rect 17776 32904 17828 32910
rect 17776 32846 17828 32852
rect 17684 31408 17736 31414
rect 17684 31350 17736 31356
rect 17592 31272 17644 31278
rect 17592 31214 17644 31220
rect 17604 30433 17632 31214
rect 17682 30560 17738 30569
rect 17682 30495 17738 30504
rect 17590 30424 17646 30433
rect 17590 30359 17646 30368
rect 17592 30320 17644 30326
rect 17592 30262 17644 30268
rect 17604 28529 17632 30262
rect 17590 28520 17646 28529
rect 17590 28455 17646 28464
rect 17592 28416 17644 28422
rect 17592 28358 17644 28364
rect 17604 27713 17632 28358
rect 17590 27704 17646 27713
rect 17590 27639 17646 27648
rect 17592 27532 17644 27538
rect 17592 27474 17644 27480
rect 17604 27305 17632 27474
rect 17590 27296 17646 27305
rect 17590 27231 17646 27240
rect 17592 27056 17644 27062
rect 17592 26998 17644 27004
rect 17604 26450 17632 26998
rect 17592 26444 17644 26450
rect 17592 26386 17644 26392
rect 17604 25702 17632 26386
rect 17592 25696 17644 25702
rect 17592 25638 17644 25644
rect 16672 23734 16724 23740
rect 16776 23718 16896 23746
rect 16960 24262 17172 24290
rect 17236 25078 17356 25106
rect 17420 25452 17540 25480
rect 16580 23656 16632 23662
rect 16580 23598 16632 23604
rect 16396 23520 16448 23526
rect 16396 23462 16448 23468
rect 16304 23316 16356 23322
rect 16304 23258 16356 23264
rect 16408 22710 16436 23462
rect 16592 23322 16620 23598
rect 16580 23316 16632 23322
rect 16580 23258 16632 23264
rect 16396 22704 16448 22710
rect 16396 22646 16448 22652
rect 16304 22568 16356 22574
rect 16304 22510 16356 22516
rect 16316 22098 16344 22510
rect 16672 22432 16724 22438
rect 16672 22374 16724 22380
rect 16304 22092 16356 22098
rect 16304 22034 16356 22040
rect 16316 21690 16344 22034
rect 16684 21876 16712 22374
rect 16592 21848 16712 21876
rect 16304 21684 16356 21690
rect 16304 21626 16356 21632
rect 16316 19922 16344 21626
rect 16396 21548 16448 21554
rect 16396 21490 16448 21496
rect 16408 21146 16436 21490
rect 16396 21140 16448 21146
rect 16396 21082 16448 21088
rect 16304 19916 16356 19922
rect 16304 19858 16356 19864
rect 16212 19848 16264 19854
rect 16212 19790 16264 19796
rect 16028 19508 16080 19514
rect 16028 19450 16080 19456
rect 16592 19310 16620 21848
rect 16672 21480 16724 21486
rect 16672 21422 16724 21428
rect 16684 20913 16712 21422
rect 16670 20904 16726 20913
rect 16670 20839 16726 20848
rect 16776 19718 16804 23718
rect 16856 22160 16908 22166
rect 16856 22102 16908 22108
rect 16868 21146 16896 22102
rect 16856 21140 16908 21146
rect 16856 21082 16908 21088
rect 16960 20398 16988 24262
rect 17236 24154 17264 25078
rect 17316 24744 17368 24750
rect 17316 24686 17368 24692
rect 17144 24126 17264 24154
rect 17038 23216 17094 23225
rect 17038 23151 17094 23160
rect 17052 23050 17080 23151
rect 17040 23044 17092 23050
rect 17040 22986 17092 22992
rect 17144 22930 17172 24126
rect 17328 24041 17356 24686
rect 17314 24032 17370 24041
rect 17314 23967 17370 23976
rect 17224 23180 17276 23186
rect 17224 23122 17276 23128
rect 17052 22902 17172 22930
rect 17052 22234 17080 22902
rect 17040 22228 17092 22234
rect 17040 22170 17092 22176
rect 17236 22166 17264 23122
rect 17328 22166 17356 23967
rect 17224 22160 17276 22166
rect 17224 22102 17276 22108
rect 17316 22160 17368 22166
rect 17316 22102 17368 22108
rect 16948 20392 17000 20398
rect 16948 20334 17000 20340
rect 17316 20392 17368 20398
rect 17316 20334 17368 20340
rect 16764 19712 16816 19718
rect 16764 19654 16816 19660
rect 16580 19304 16632 19310
rect 16580 19246 16632 19252
rect 16592 18970 16620 19246
rect 16672 19168 16724 19174
rect 16672 19110 16724 19116
rect 16580 18964 16632 18970
rect 16580 18906 16632 18912
rect 16302 18864 16358 18873
rect 15936 18828 15988 18834
rect 16302 18799 16304 18808
rect 15936 18770 15988 18776
rect 16356 18799 16358 18808
rect 16304 18770 16356 18776
rect 15948 18426 15976 18770
rect 15936 18420 15988 18426
rect 15936 18362 15988 18368
rect 16316 18358 16344 18770
rect 16396 18760 16448 18766
rect 16396 18702 16448 18708
rect 16304 18352 16356 18358
rect 16304 18294 16356 18300
rect 16408 18154 16436 18702
rect 16396 18148 16448 18154
rect 16396 18090 16448 18096
rect 16684 18034 16712 19110
rect 16408 18006 16712 18034
rect 16408 17134 16436 18006
rect 16488 17536 16540 17542
rect 16488 17478 16540 17484
rect 16500 17134 16528 17478
rect 15844 17128 15896 17134
rect 15844 17070 15896 17076
rect 16396 17128 16448 17134
rect 16396 17070 16448 17076
rect 16488 17128 16540 17134
rect 16488 17070 16540 17076
rect 15856 16794 15884 17070
rect 15844 16788 15896 16794
rect 15844 16730 15896 16736
rect 16776 16590 16804 19654
rect 16960 17678 16988 20334
rect 17328 19718 17356 20334
rect 17316 19712 17368 19718
rect 17316 19654 17368 19660
rect 17314 19408 17370 19417
rect 17314 19343 17370 19352
rect 17328 18834 17356 19343
rect 17316 18828 17368 18834
rect 17316 18770 17368 18776
rect 17328 18426 17356 18770
rect 17316 18420 17368 18426
rect 17316 18362 17368 18368
rect 17040 18148 17092 18154
rect 17040 18090 17092 18096
rect 17052 17746 17080 18090
rect 17040 17740 17092 17746
rect 17040 17682 17092 17688
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 17052 17490 17080 17682
rect 16960 17462 17080 17490
rect 16960 17202 16988 17462
rect 17420 17252 17448 25452
rect 17500 25356 17552 25362
rect 17500 25298 17552 25304
rect 17512 24886 17540 25298
rect 17604 25265 17632 25638
rect 17696 25498 17724 30495
rect 17788 30258 17816 32846
rect 17880 32774 17908 33866
rect 18052 33856 18104 33862
rect 18052 33798 18104 33804
rect 17958 33008 18014 33017
rect 17958 32943 17960 32952
rect 18012 32943 18014 32952
rect 17960 32914 18012 32920
rect 18064 32881 18092 33798
rect 18050 32872 18106 32881
rect 18050 32807 18106 32816
rect 17868 32768 17920 32774
rect 17868 32710 17920 32716
rect 17960 32292 18012 32298
rect 17960 32234 18012 32240
rect 17972 31822 18000 32234
rect 17960 31816 18012 31822
rect 17960 31758 18012 31764
rect 18064 31210 18092 32807
rect 18052 31204 18104 31210
rect 18052 31146 18104 31152
rect 17960 31136 18012 31142
rect 17880 31084 17960 31090
rect 17880 31078 18012 31084
rect 17880 31062 18000 31078
rect 17776 30252 17828 30258
rect 17776 30194 17828 30200
rect 17880 30122 17908 31062
rect 17960 30796 18012 30802
rect 17960 30738 18012 30744
rect 17868 30116 17920 30122
rect 17868 30058 17920 30064
rect 17868 29844 17920 29850
rect 17972 29832 18000 30738
rect 18064 30433 18092 31146
rect 18050 30424 18106 30433
rect 18050 30359 18106 30368
rect 18064 30258 18092 30359
rect 18052 30252 18104 30258
rect 18052 30194 18104 30200
rect 17920 29804 18000 29832
rect 17868 29786 17920 29792
rect 18052 29708 18104 29714
rect 18052 29650 18104 29656
rect 17776 29640 17828 29646
rect 17776 29582 17828 29588
rect 17788 29306 17816 29582
rect 17776 29300 17828 29306
rect 17776 29242 17828 29248
rect 18064 29170 18092 29650
rect 18052 29164 18104 29170
rect 18052 29106 18104 29112
rect 18052 28960 18104 28966
rect 18052 28902 18104 28908
rect 17776 28620 17828 28626
rect 17776 28562 17828 28568
rect 17788 28529 17816 28562
rect 17774 28520 17830 28529
rect 17774 28455 17830 28464
rect 17788 28218 17816 28455
rect 17960 28416 18012 28422
rect 17960 28358 18012 28364
rect 17776 28212 17828 28218
rect 17776 28154 17828 28160
rect 17972 28150 18000 28358
rect 17960 28144 18012 28150
rect 17960 28086 18012 28092
rect 18064 27606 18092 28902
rect 17776 27600 17828 27606
rect 17776 27542 17828 27548
rect 18052 27600 18104 27606
rect 18052 27542 18104 27548
rect 17788 26382 17816 27542
rect 17868 27532 17920 27538
rect 17868 27474 17920 27480
rect 17776 26376 17828 26382
rect 17776 26318 17828 26324
rect 17880 26314 17908 27474
rect 18052 27464 18104 27470
rect 18050 27432 18052 27441
rect 18104 27432 18106 27441
rect 18050 27367 18106 27376
rect 17868 26308 17920 26314
rect 17868 26250 17920 26256
rect 17880 26042 17908 26250
rect 17868 26036 17920 26042
rect 17868 25978 17920 25984
rect 17684 25492 17736 25498
rect 17684 25434 17736 25440
rect 17868 25356 17920 25362
rect 17920 25316 18000 25344
rect 17868 25298 17920 25304
rect 17590 25256 17646 25265
rect 17590 25191 17646 25200
rect 17868 25220 17920 25226
rect 17868 25162 17920 25168
rect 17500 24880 17552 24886
rect 17500 24822 17552 24828
rect 17682 24712 17738 24721
rect 17682 24647 17738 24656
rect 17500 24608 17552 24614
rect 17500 24550 17552 24556
rect 17512 24342 17540 24550
rect 17500 24336 17552 24342
rect 17500 24278 17552 24284
rect 17590 24304 17646 24313
rect 17590 24239 17592 24248
rect 17644 24239 17646 24248
rect 17592 24210 17644 24216
rect 17592 23792 17644 23798
rect 17592 23734 17644 23740
rect 17500 23180 17552 23186
rect 17500 23122 17552 23128
rect 17512 22681 17540 23122
rect 17604 22778 17632 23734
rect 17592 22772 17644 22778
rect 17592 22714 17644 22720
rect 17498 22672 17554 22681
rect 17498 22607 17554 22616
rect 17696 22506 17724 24647
rect 17776 24608 17828 24614
rect 17776 24550 17828 24556
rect 17788 24177 17816 24550
rect 17880 24274 17908 25162
rect 17972 24410 18000 25316
rect 18052 25220 18104 25226
rect 18052 25162 18104 25168
rect 18064 24682 18092 25162
rect 18052 24676 18104 24682
rect 18052 24618 18104 24624
rect 17960 24404 18012 24410
rect 17960 24346 18012 24352
rect 17868 24268 17920 24274
rect 17868 24210 17920 24216
rect 17774 24168 17830 24177
rect 17774 24103 17830 24112
rect 17774 24032 17830 24041
rect 17774 23967 17830 23976
rect 17684 22500 17736 22506
rect 17684 22442 17736 22448
rect 17684 22228 17736 22234
rect 17684 22170 17736 22176
rect 17500 22092 17552 22098
rect 17500 22034 17552 22040
rect 17512 21690 17540 22034
rect 17592 21888 17644 21894
rect 17592 21830 17644 21836
rect 17500 21684 17552 21690
rect 17500 21626 17552 21632
rect 17604 20466 17632 21830
rect 17696 21010 17724 22170
rect 17788 21554 17816 23967
rect 17880 23866 17908 24210
rect 17960 24064 18012 24070
rect 17960 24006 18012 24012
rect 17868 23860 17920 23866
rect 17868 23802 17920 23808
rect 17972 23730 18000 24006
rect 17960 23724 18012 23730
rect 17960 23666 18012 23672
rect 17868 23112 17920 23118
rect 18064 23066 18092 24618
rect 17920 23060 18092 23066
rect 17868 23054 18092 23060
rect 17880 23038 18092 23054
rect 17868 22568 17920 22574
rect 17868 22510 17920 22516
rect 17880 22098 17908 22510
rect 17868 22092 17920 22098
rect 17868 22034 17920 22040
rect 17972 21962 18000 23038
rect 18052 22500 18104 22506
rect 18052 22442 18104 22448
rect 18064 22234 18092 22442
rect 18052 22228 18104 22234
rect 18052 22170 18104 22176
rect 18052 22024 18104 22030
rect 18052 21966 18104 21972
rect 17960 21956 18012 21962
rect 17960 21898 18012 21904
rect 17972 21554 18000 21898
rect 17776 21548 17828 21554
rect 17776 21490 17828 21496
rect 17960 21548 18012 21554
rect 17960 21490 18012 21496
rect 18064 21146 18092 21966
rect 18156 21842 18184 49846
rect 18248 49774 18276 49914
rect 18236 49768 18288 49774
rect 18236 49710 18288 49716
rect 18234 48920 18290 48929
rect 18234 48855 18236 48864
rect 18288 48855 18290 48864
rect 18236 48826 18288 48832
rect 18432 48278 18460 50759
rect 18524 50454 18552 52974
rect 18788 52896 18840 52902
rect 18788 52838 18840 52844
rect 18696 52556 18748 52562
rect 18696 52498 18748 52504
rect 18708 52465 18736 52498
rect 18694 52456 18750 52465
rect 18694 52391 18750 52400
rect 18708 52154 18736 52391
rect 18800 52358 18828 52838
rect 18788 52352 18840 52358
rect 18788 52294 18840 52300
rect 18696 52148 18748 52154
rect 18696 52090 18748 52096
rect 18604 51944 18656 51950
rect 18604 51886 18656 51892
rect 18616 51610 18644 51886
rect 18800 51610 18828 52294
rect 18892 52057 18920 61542
rect 19580 61500 19876 61520
rect 19636 61498 19660 61500
rect 19716 61498 19740 61500
rect 19796 61498 19820 61500
rect 19658 61446 19660 61498
rect 19722 61446 19734 61498
rect 19796 61446 19798 61498
rect 19636 61444 19660 61446
rect 19716 61444 19740 61446
rect 19796 61444 19820 61446
rect 19580 61424 19876 61444
rect 19340 61260 19392 61266
rect 19340 61202 19392 61208
rect 19352 60518 19380 61202
rect 20088 61062 20116 61542
rect 20364 61402 20392 62970
rect 20626 62384 20682 62393
rect 20626 62319 20682 62328
rect 20352 61396 20404 61402
rect 20352 61338 20404 61344
rect 20260 61124 20312 61130
rect 20260 61066 20312 61072
rect 20076 61056 20128 61062
rect 20076 60998 20128 61004
rect 20088 60722 20116 60998
rect 20076 60716 20128 60722
rect 20076 60658 20128 60664
rect 20272 60654 20300 61066
rect 19984 60648 20036 60654
rect 19984 60590 20036 60596
rect 20260 60648 20312 60654
rect 20260 60590 20312 60596
rect 19432 60580 19484 60586
rect 19432 60522 19484 60528
rect 19340 60512 19392 60518
rect 19340 60454 19392 60460
rect 19248 60172 19300 60178
rect 19248 60114 19300 60120
rect 19260 59158 19288 60114
rect 19248 59152 19300 59158
rect 19246 59120 19248 59129
rect 19300 59120 19302 59129
rect 19246 59055 19302 59064
rect 18972 59016 19024 59022
rect 18972 58958 19024 58964
rect 18984 58478 19012 58958
rect 19064 58880 19116 58886
rect 19064 58822 19116 58828
rect 19076 58682 19104 58822
rect 19064 58676 19116 58682
rect 19064 58618 19116 58624
rect 18972 58472 19024 58478
rect 18972 58414 19024 58420
rect 18984 57934 19012 58414
rect 18972 57928 19024 57934
rect 18972 57870 19024 57876
rect 18984 57798 19012 57870
rect 19076 57866 19104 58618
rect 19156 58608 19208 58614
rect 19208 58556 19288 58562
rect 19156 58550 19288 58556
rect 19168 58534 19288 58550
rect 19156 58404 19208 58410
rect 19156 58346 19208 58352
rect 19168 58002 19196 58346
rect 19156 57996 19208 58002
rect 19156 57938 19208 57944
rect 19064 57860 19116 57866
rect 19064 57802 19116 57808
rect 18972 57792 19024 57798
rect 18972 57734 19024 57740
rect 18984 57254 19012 57734
rect 19076 57594 19104 57802
rect 19064 57588 19116 57594
rect 19064 57530 19116 57536
rect 18972 57248 19024 57254
rect 18972 57190 19024 57196
rect 19076 57050 19104 57530
rect 19168 57322 19196 57938
rect 19260 57338 19288 58534
rect 19352 58138 19380 60454
rect 19444 58682 19472 60522
rect 19580 60412 19876 60432
rect 19636 60410 19660 60412
rect 19716 60410 19740 60412
rect 19796 60410 19820 60412
rect 19658 60358 19660 60410
rect 19722 60358 19734 60410
rect 19796 60358 19798 60410
rect 19636 60356 19660 60358
rect 19716 60356 19740 60358
rect 19796 60356 19820 60358
rect 19580 60336 19876 60356
rect 19708 60172 19760 60178
rect 19708 60114 19760 60120
rect 19524 59968 19576 59974
rect 19524 59910 19576 59916
rect 19536 59498 19564 59910
rect 19720 59498 19748 60114
rect 19892 59968 19944 59974
rect 19892 59910 19944 59916
rect 19904 59770 19932 59910
rect 19892 59764 19944 59770
rect 19892 59706 19944 59712
rect 19996 59702 20024 60590
rect 20076 60580 20128 60586
rect 20076 60522 20128 60528
rect 19984 59696 20036 59702
rect 19984 59638 20036 59644
rect 19524 59492 19576 59498
rect 19524 59434 19576 59440
rect 19708 59492 19760 59498
rect 19708 59434 19760 59440
rect 19580 59324 19876 59344
rect 19636 59322 19660 59324
rect 19716 59322 19740 59324
rect 19796 59322 19820 59324
rect 19658 59270 19660 59322
rect 19722 59270 19734 59322
rect 19796 59270 19798 59322
rect 19636 59268 19660 59270
rect 19716 59268 19740 59270
rect 19796 59268 19820 59270
rect 19580 59248 19876 59268
rect 19996 59158 20024 59638
rect 19984 59152 20036 59158
rect 19984 59094 20036 59100
rect 19984 58948 20036 58954
rect 19984 58890 20036 58896
rect 19892 58880 19944 58886
rect 19892 58822 19944 58828
rect 19432 58676 19484 58682
rect 19432 58618 19484 58624
rect 19580 58236 19876 58256
rect 19636 58234 19660 58236
rect 19716 58234 19740 58236
rect 19796 58234 19820 58236
rect 19658 58182 19660 58234
rect 19722 58182 19734 58234
rect 19796 58182 19798 58234
rect 19636 58180 19660 58182
rect 19716 58180 19740 58182
rect 19796 58180 19820 58182
rect 19580 58160 19876 58180
rect 19340 58132 19392 58138
rect 19340 58074 19392 58080
rect 19432 57792 19484 57798
rect 19432 57734 19484 57740
rect 19614 57760 19670 57769
rect 19444 57526 19472 57734
rect 19614 57695 19670 57704
rect 19628 57594 19656 57695
rect 19616 57588 19668 57594
rect 19616 57530 19668 57536
rect 19432 57520 19484 57526
rect 19432 57462 19484 57468
rect 19432 57384 19484 57390
rect 19156 57316 19208 57322
rect 19260 57310 19380 57338
rect 19432 57326 19484 57332
rect 19156 57258 19208 57264
rect 19248 57248 19300 57254
rect 19248 57190 19300 57196
rect 19064 57044 19116 57050
rect 19064 56986 19116 56992
rect 18972 56840 19024 56846
rect 18972 56782 19024 56788
rect 18984 56438 19012 56782
rect 19076 56710 19104 56986
rect 19156 56976 19208 56982
rect 19156 56918 19208 56924
rect 19064 56704 19116 56710
rect 19064 56646 19116 56652
rect 18972 56432 19024 56438
rect 18972 56374 19024 56380
rect 18984 55457 19012 56374
rect 19076 55962 19104 56646
rect 19168 56438 19196 56918
rect 19156 56432 19208 56438
rect 19156 56374 19208 56380
rect 19260 56386 19288 57190
rect 19352 56982 19380 57310
rect 19340 56976 19392 56982
rect 19340 56918 19392 56924
rect 19352 56778 19380 56918
rect 19444 56846 19472 57326
rect 19580 57148 19876 57168
rect 19636 57146 19660 57148
rect 19716 57146 19740 57148
rect 19796 57146 19820 57148
rect 19658 57094 19660 57146
rect 19722 57094 19734 57146
rect 19796 57094 19798 57146
rect 19636 57092 19660 57094
rect 19716 57092 19740 57094
rect 19796 57092 19820 57094
rect 19580 57072 19876 57092
rect 19432 56840 19484 56846
rect 19432 56782 19484 56788
rect 19340 56772 19392 56778
rect 19340 56714 19392 56720
rect 19444 56506 19472 56782
rect 19524 56704 19576 56710
rect 19522 56672 19524 56681
rect 19576 56672 19578 56681
rect 19522 56607 19578 56616
rect 19432 56500 19484 56506
rect 19432 56442 19484 56448
rect 19524 56500 19576 56506
rect 19524 56442 19576 56448
rect 19064 55956 19116 55962
rect 19064 55898 19116 55904
rect 19064 55820 19116 55826
rect 19064 55762 19116 55768
rect 18970 55448 19026 55457
rect 18970 55383 19026 55392
rect 19076 55214 19104 55762
rect 19168 55690 19196 56374
rect 19260 56370 19380 56386
rect 19260 56364 19392 56370
rect 19260 56358 19340 56364
rect 19340 56306 19392 56312
rect 19536 56250 19564 56442
rect 19616 56432 19668 56438
rect 19614 56400 19616 56409
rect 19904 56409 19932 58822
rect 19996 58342 20024 58890
rect 19984 58336 20036 58342
rect 19984 58278 20036 58284
rect 19996 56506 20024 58278
rect 19984 56500 20036 56506
rect 19984 56442 20036 56448
rect 19668 56400 19670 56409
rect 19614 56335 19670 56344
rect 19890 56400 19946 56409
rect 19890 56335 19946 56344
rect 20088 56250 20116 60522
rect 20272 60194 20300 60590
rect 20364 60314 20392 61338
rect 20640 60790 20668 62319
rect 20732 61130 20760 68303
rect 20720 61124 20772 61130
rect 20720 61066 20772 61072
rect 20628 60784 20680 60790
rect 20628 60726 20680 60732
rect 20536 60648 20588 60654
rect 20536 60590 20588 60596
rect 20352 60308 20404 60314
rect 20352 60250 20404 60256
rect 20180 60178 20300 60194
rect 20168 60172 20300 60178
rect 20220 60166 20300 60172
rect 20168 60114 20220 60120
rect 20168 60036 20220 60042
rect 20168 59978 20220 59984
rect 20180 59673 20208 59978
rect 20166 59664 20222 59673
rect 20166 59599 20222 59608
rect 20180 59566 20208 59599
rect 20168 59560 20220 59566
rect 20168 59502 20220 59508
rect 20168 57928 20220 57934
rect 20168 57870 20220 57876
rect 20180 57050 20208 57870
rect 20272 57474 20300 60166
rect 20364 59566 20392 60250
rect 20444 60104 20496 60110
rect 20444 60046 20496 60052
rect 20352 59560 20404 59566
rect 20352 59502 20404 59508
rect 20456 59022 20484 60046
rect 20548 59634 20576 60590
rect 20626 59800 20682 59809
rect 20626 59735 20682 59744
rect 20640 59634 20668 59735
rect 20536 59628 20588 59634
rect 20536 59570 20588 59576
rect 20628 59628 20680 59634
rect 20628 59570 20680 59576
rect 20536 59424 20588 59430
rect 20536 59366 20588 59372
rect 20444 59016 20496 59022
rect 20444 58958 20496 58964
rect 20272 57446 20392 57474
rect 20456 57458 20484 58958
rect 20548 58886 20576 59366
rect 20536 58880 20588 58886
rect 20536 58822 20588 58828
rect 20548 58342 20576 58822
rect 20536 58336 20588 58342
rect 20536 58278 20588 58284
rect 20168 57044 20220 57050
rect 20168 56986 20220 56992
rect 20180 56302 20208 56986
rect 20260 56432 20312 56438
rect 20260 56374 20312 56380
rect 19352 56222 19564 56250
rect 19904 56222 20116 56250
rect 20168 56296 20220 56302
rect 20168 56238 20220 56244
rect 19352 56166 19380 56222
rect 19340 56160 19392 56166
rect 19340 56102 19392 56108
rect 19432 56160 19484 56166
rect 19432 56102 19484 56108
rect 19352 55842 19380 56102
rect 19260 55814 19380 55842
rect 19156 55684 19208 55690
rect 19156 55626 19208 55632
rect 19064 55208 19116 55214
rect 19064 55150 19116 55156
rect 19064 54868 19116 54874
rect 19064 54810 19116 54816
rect 18972 53644 19024 53650
rect 18972 53586 19024 53592
rect 18984 53038 19012 53586
rect 19076 53514 19104 54810
rect 19260 54806 19288 55814
rect 19340 55752 19392 55758
rect 19340 55694 19392 55700
rect 19352 55078 19380 55694
rect 19444 55321 19472 56102
rect 19580 56060 19876 56080
rect 19636 56058 19660 56060
rect 19716 56058 19740 56060
rect 19796 56058 19820 56060
rect 19658 56006 19660 56058
rect 19722 56006 19734 56058
rect 19796 56006 19798 56058
rect 19636 56004 19660 56006
rect 19716 56004 19740 56006
rect 19796 56004 19820 56006
rect 19580 55984 19876 56004
rect 19524 55616 19576 55622
rect 19524 55558 19576 55564
rect 19430 55312 19486 55321
rect 19430 55247 19486 55256
rect 19536 55162 19564 55558
rect 19616 55208 19668 55214
rect 19444 55134 19564 55162
rect 19614 55176 19616 55185
rect 19668 55176 19670 55185
rect 19444 55078 19472 55134
rect 19614 55111 19670 55120
rect 19340 55072 19392 55078
rect 19340 55014 19392 55020
rect 19432 55072 19484 55078
rect 19432 55014 19484 55020
rect 19248 54800 19300 54806
rect 19248 54742 19300 54748
rect 19352 54738 19380 55014
rect 19444 54806 19472 55014
rect 19580 54972 19876 54992
rect 19636 54970 19660 54972
rect 19716 54970 19740 54972
rect 19796 54970 19820 54972
rect 19658 54918 19660 54970
rect 19722 54918 19734 54970
rect 19796 54918 19798 54970
rect 19636 54916 19660 54918
rect 19716 54916 19740 54918
rect 19796 54916 19820 54918
rect 19580 54896 19876 54916
rect 19432 54800 19484 54806
rect 19432 54742 19484 54748
rect 19340 54732 19392 54738
rect 19340 54674 19392 54680
rect 19616 54732 19668 54738
rect 19616 54674 19668 54680
rect 19246 54632 19302 54641
rect 19246 54567 19302 54576
rect 19260 53802 19288 54567
rect 19352 54369 19380 54674
rect 19338 54360 19394 54369
rect 19338 54295 19340 54304
rect 19392 54295 19394 54304
rect 19340 54266 19392 54272
rect 19352 54235 19380 54266
rect 19628 54262 19656 54674
rect 19616 54256 19668 54262
rect 19616 54198 19668 54204
rect 19432 54188 19484 54194
rect 19432 54130 19484 54136
rect 19340 53984 19392 53990
rect 19444 53961 19472 54130
rect 19628 54058 19656 54198
rect 19616 54052 19668 54058
rect 19616 53994 19668 54000
rect 19340 53926 19392 53932
rect 19430 53952 19486 53961
rect 19352 53802 19380 53926
rect 19430 53887 19486 53896
rect 19580 53884 19876 53904
rect 19636 53882 19660 53884
rect 19716 53882 19740 53884
rect 19796 53882 19820 53884
rect 19658 53830 19660 53882
rect 19722 53830 19734 53882
rect 19796 53830 19798 53882
rect 19636 53828 19660 53830
rect 19716 53828 19740 53830
rect 19796 53828 19820 53830
rect 19580 53808 19876 53828
rect 19168 53786 19380 53802
rect 19168 53780 19392 53786
rect 19168 53774 19340 53780
rect 19064 53508 19116 53514
rect 19064 53450 19116 53456
rect 18972 53032 19024 53038
rect 18972 52974 19024 52980
rect 18972 52420 19024 52426
rect 18972 52362 19024 52368
rect 18878 52048 18934 52057
rect 18878 51983 18934 51992
rect 18984 51814 19012 52362
rect 19064 52148 19116 52154
rect 19064 52090 19116 52096
rect 19076 52057 19104 52090
rect 19062 52048 19118 52057
rect 19062 51983 19118 51992
rect 19168 51950 19196 53774
rect 19340 53722 19392 53728
rect 19616 53712 19668 53718
rect 19614 53680 19616 53689
rect 19668 53680 19670 53689
rect 19614 53615 19670 53624
rect 19432 53576 19484 53582
rect 19432 53518 19484 53524
rect 19444 52562 19472 53518
rect 19522 53272 19578 53281
rect 19522 53207 19524 53216
rect 19576 53207 19578 53216
rect 19524 53178 19576 53184
rect 19580 52796 19876 52816
rect 19636 52794 19660 52796
rect 19716 52794 19740 52796
rect 19796 52794 19820 52796
rect 19658 52742 19660 52794
rect 19722 52742 19734 52794
rect 19796 52742 19798 52794
rect 19636 52740 19660 52742
rect 19716 52740 19740 52742
rect 19796 52740 19820 52742
rect 19580 52720 19876 52740
rect 19904 52562 19932 56222
rect 19982 56128 20038 56137
rect 19982 56063 20038 56072
rect 19996 55894 20024 56063
rect 19984 55888 20036 55894
rect 19984 55830 20036 55836
rect 19982 55448 20038 55457
rect 20180 55418 20208 56238
rect 20272 55962 20300 56374
rect 20260 55956 20312 55962
rect 20260 55898 20312 55904
rect 20260 55684 20312 55690
rect 20260 55626 20312 55632
rect 20272 55457 20300 55626
rect 20258 55448 20314 55457
rect 19982 55383 20038 55392
rect 20168 55412 20220 55418
rect 19996 53786 20024 55383
rect 20258 55383 20314 55392
rect 20168 55354 20220 55360
rect 20272 55282 20300 55383
rect 20260 55276 20312 55282
rect 20260 55218 20312 55224
rect 20168 54732 20220 54738
rect 20168 54674 20220 54680
rect 20076 54052 20128 54058
rect 20076 53994 20128 54000
rect 19984 53780 20036 53786
rect 19984 53722 20036 53728
rect 19996 53174 20024 53722
rect 19984 53168 20036 53174
rect 19984 53110 20036 53116
rect 19432 52556 19484 52562
rect 19432 52498 19484 52504
rect 19892 52556 19944 52562
rect 19892 52498 19944 52504
rect 19340 52420 19392 52426
rect 19340 52362 19392 52368
rect 19156 51944 19208 51950
rect 19156 51886 19208 51892
rect 19248 51876 19300 51882
rect 19248 51818 19300 51824
rect 18972 51808 19024 51814
rect 18972 51750 19024 51756
rect 18604 51604 18656 51610
rect 18604 51546 18656 51552
rect 18788 51604 18840 51610
rect 18788 51546 18840 51552
rect 18604 51060 18656 51066
rect 18604 51002 18656 51008
rect 18512 50448 18564 50454
rect 18512 50390 18564 50396
rect 18616 49774 18644 51002
rect 18800 50862 18828 51546
rect 18972 51400 19024 51406
rect 18972 51342 19024 51348
rect 18880 50992 18932 50998
rect 18880 50934 18932 50940
rect 18788 50856 18840 50862
rect 18788 50798 18840 50804
rect 18604 49768 18656 49774
rect 18604 49710 18656 49716
rect 18616 49230 18644 49710
rect 18604 49224 18656 49230
rect 18604 49166 18656 49172
rect 18696 49156 18748 49162
rect 18696 49098 18748 49104
rect 18420 48272 18472 48278
rect 18420 48214 18472 48220
rect 18604 48272 18656 48278
rect 18604 48214 18656 48220
rect 18616 47802 18644 48214
rect 18604 47796 18656 47802
rect 18604 47738 18656 47744
rect 18236 40928 18288 40934
rect 18236 40870 18288 40876
rect 18248 40089 18276 40870
rect 18234 40080 18290 40089
rect 18234 40015 18290 40024
rect 18604 39840 18656 39846
rect 18602 39808 18604 39817
rect 18656 39808 18658 39817
rect 18602 39743 18658 39752
rect 18236 39500 18288 39506
rect 18236 39442 18288 39448
rect 18248 38282 18276 39442
rect 18420 38956 18472 38962
rect 18420 38898 18472 38904
rect 18236 38276 18288 38282
rect 18236 38218 18288 38224
rect 18326 37904 18382 37913
rect 18326 37839 18382 37848
rect 18236 37800 18288 37806
rect 18236 37742 18288 37748
rect 18248 37330 18276 37742
rect 18236 37324 18288 37330
rect 18236 37266 18288 37272
rect 18248 36718 18276 37266
rect 18236 36712 18288 36718
rect 18236 36654 18288 36660
rect 18248 36378 18276 36654
rect 18236 36372 18288 36378
rect 18236 36314 18288 36320
rect 18340 36310 18368 37839
rect 18432 37806 18460 38898
rect 18708 38729 18736 49098
rect 18892 42401 18920 50934
rect 18984 50386 19012 51342
rect 19260 50862 19288 51818
rect 19248 50856 19300 50862
rect 19248 50798 19300 50804
rect 19352 50402 19380 52362
rect 18972 50380 19024 50386
rect 18972 50322 19024 50328
rect 19260 50374 19380 50402
rect 18984 49298 19012 50322
rect 19260 49858 19288 50374
rect 19340 50312 19392 50318
rect 19340 50254 19392 50260
rect 19352 49978 19380 50254
rect 19340 49972 19392 49978
rect 19340 49914 19392 49920
rect 19260 49830 19380 49858
rect 18972 49292 19024 49298
rect 18972 49234 19024 49240
rect 18984 48346 19012 49234
rect 19246 49056 19302 49065
rect 19246 48991 19302 49000
rect 19260 48754 19288 48991
rect 19248 48748 19300 48754
rect 19248 48690 19300 48696
rect 18972 48340 19024 48346
rect 18972 48282 19024 48288
rect 19062 48240 19118 48249
rect 19062 48175 19064 48184
rect 19116 48175 19118 48184
rect 19064 48146 19116 48152
rect 19076 47802 19104 48146
rect 19064 47796 19116 47802
rect 19064 47738 19116 47744
rect 19352 46209 19380 49830
rect 19444 49434 19472 52498
rect 19580 51708 19876 51728
rect 19636 51706 19660 51708
rect 19716 51706 19740 51708
rect 19796 51706 19820 51708
rect 19658 51654 19660 51706
rect 19722 51654 19734 51706
rect 19796 51654 19798 51706
rect 19636 51652 19660 51654
rect 19716 51652 19740 51654
rect 19796 51652 19820 51654
rect 19580 51632 19876 51652
rect 19524 51400 19576 51406
rect 19524 51342 19576 51348
rect 19536 50833 19564 51342
rect 19800 51332 19852 51338
rect 19800 51274 19852 51280
rect 19812 51066 19840 51274
rect 19800 51060 19852 51066
rect 19800 51002 19852 51008
rect 19522 50824 19578 50833
rect 19522 50759 19578 50768
rect 19580 50620 19876 50640
rect 19636 50618 19660 50620
rect 19716 50618 19740 50620
rect 19796 50618 19820 50620
rect 19658 50566 19660 50618
rect 19722 50566 19734 50618
rect 19796 50566 19798 50618
rect 19636 50564 19660 50566
rect 19716 50564 19740 50566
rect 19796 50564 19820 50566
rect 19580 50544 19876 50564
rect 19904 50017 19932 52498
rect 19996 52494 20024 53110
rect 19984 52488 20036 52494
rect 19984 52430 20036 52436
rect 19984 51944 20036 51950
rect 19984 51886 20036 51892
rect 19996 51785 20024 51886
rect 19982 51776 20038 51785
rect 19982 51711 20038 51720
rect 20088 51542 20116 53994
rect 20076 51536 20128 51542
rect 19982 51504 20038 51513
rect 20076 51478 20128 51484
rect 19982 51439 20038 51448
rect 19996 51406 20024 51439
rect 19984 51400 20036 51406
rect 19984 51342 20036 51348
rect 19996 50726 20024 51342
rect 20180 50969 20208 54674
rect 20260 54596 20312 54602
rect 20260 54538 20312 54544
rect 20272 53990 20300 54538
rect 20260 53984 20312 53990
rect 20260 53926 20312 53932
rect 20272 53174 20300 53926
rect 20364 53582 20392 57446
rect 20444 57452 20496 57458
rect 20444 57394 20496 57400
rect 20444 57248 20496 57254
rect 20444 57190 20496 57196
rect 20456 56914 20484 57190
rect 20444 56908 20496 56914
rect 20444 56850 20496 56856
rect 20444 55072 20496 55078
rect 20442 55040 20444 55049
rect 20496 55040 20498 55049
rect 20442 54975 20498 54984
rect 20442 54904 20498 54913
rect 20548 54890 20576 58278
rect 20628 57792 20680 57798
rect 20628 57734 20680 57740
rect 20640 57254 20668 57734
rect 20720 57384 20772 57390
rect 20720 57326 20772 57332
rect 20628 57248 20680 57254
rect 20628 57190 20680 57196
rect 20732 57050 20760 57326
rect 20720 57044 20772 57050
rect 20720 56986 20772 56992
rect 20720 55820 20772 55826
rect 20720 55762 20772 55768
rect 20732 55622 20760 55762
rect 20720 55616 20772 55622
rect 20718 55584 20720 55593
rect 20772 55584 20774 55593
rect 20718 55519 20774 55528
rect 20720 55276 20772 55282
rect 20498 54862 20576 54890
rect 20640 55236 20720 55264
rect 20442 54839 20498 54848
rect 20456 53990 20484 54839
rect 20640 54806 20668 55236
rect 20720 55218 20772 55224
rect 20628 54800 20680 54806
rect 20628 54742 20680 54748
rect 20720 54528 20772 54534
rect 20720 54470 20772 54476
rect 20628 54188 20680 54194
rect 20628 54130 20680 54136
rect 20444 53984 20496 53990
rect 20444 53926 20496 53932
rect 20456 53786 20484 53926
rect 20640 53786 20668 54130
rect 20732 54058 20760 54470
rect 20720 54052 20772 54058
rect 20720 53994 20772 54000
rect 20444 53780 20496 53786
rect 20444 53722 20496 53728
rect 20628 53780 20680 53786
rect 20628 53722 20680 53728
rect 20352 53576 20404 53582
rect 20352 53518 20404 53524
rect 20260 53168 20312 53174
rect 20260 53110 20312 53116
rect 20272 52494 20300 53110
rect 20536 53032 20588 53038
rect 20536 52974 20588 52980
rect 20444 52624 20496 52630
rect 20444 52566 20496 52572
rect 20260 52488 20312 52494
rect 20260 52430 20312 52436
rect 20456 51950 20484 52566
rect 20548 52562 20576 52974
rect 20640 52873 20668 53722
rect 20732 53718 20760 53994
rect 20720 53712 20772 53718
rect 20720 53654 20772 53660
rect 20732 53145 20760 53654
rect 20718 53136 20774 53145
rect 20718 53071 20720 53080
rect 20772 53071 20774 53080
rect 20720 53042 20772 53048
rect 20626 52864 20682 52873
rect 20626 52799 20682 52808
rect 20628 52692 20680 52698
rect 20628 52634 20680 52640
rect 20536 52556 20588 52562
rect 20536 52498 20588 52504
rect 20260 51944 20312 51950
rect 20444 51944 20496 51950
rect 20260 51886 20312 51892
rect 20350 51912 20406 51921
rect 20272 51610 20300 51886
rect 20444 51886 20496 51892
rect 20350 51847 20406 51856
rect 20260 51604 20312 51610
rect 20260 51546 20312 51552
rect 20364 51066 20392 51847
rect 20536 51604 20588 51610
rect 20536 51546 20588 51552
rect 20352 51060 20404 51066
rect 20352 51002 20404 51008
rect 20166 50960 20222 50969
rect 20166 50895 20222 50904
rect 20444 50788 20496 50794
rect 20444 50730 20496 50736
rect 19984 50720 20036 50726
rect 20352 50720 20404 50726
rect 19984 50662 20036 50668
rect 20074 50688 20130 50697
rect 20352 50662 20404 50668
rect 20074 50623 20130 50632
rect 19890 50008 19946 50017
rect 19890 49943 19946 49952
rect 20088 49774 20116 50623
rect 20168 50312 20220 50318
rect 20168 50254 20220 50260
rect 20076 49768 20128 49774
rect 20076 49710 20128 49716
rect 19580 49532 19876 49552
rect 19636 49530 19660 49532
rect 19716 49530 19740 49532
rect 19796 49530 19820 49532
rect 19658 49478 19660 49530
rect 19722 49478 19734 49530
rect 19796 49478 19798 49530
rect 19636 49476 19660 49478
rect 19716 49476 19740 49478
rect 19796 49476 19820 49478
rect 19580 49456 19876 49476
rect 19432 49428 19484 49434
rect 19432 49370 19484 49376
rect 19444 48686 19472 49370
rect 19708 49224 19760 49230
rect 19708 49166 19760 49172
rect 19524 48748 19576 48754
rect 19720 48736 19748 49166
rect 20076 48884 20128 48890
rect 20076 48826 20128 48832
rect 19982 48784 20038 48793
rect 19720 48708 19840 48736
rect 19982 48719 20038 48728
rect 19524 48690 19576 48696
rect 19432 48680 19484 48686
rect 19536 48657 19564 48690
rect 19432 48622 19484 48628
rect 19522 48648 19578 48657
rect 19444 48210 19472 48622
rect 19522 48583 19578 48592
rect 19812 48600 19840 48708
rect 19996 48686 20024 48719
rect 19984 48680 20036 48686
rect 19984 48622 20036 48628
rect 19812 48572 19932 48600
rect 19580 48444 19876 48464
rect 19636 48442 19660 48444
rect 19716 48442 19740 48444
rect 19796 48442 19820 48444
rect 19658 48390 19660 48442
rect 19722 48390 19734 48442
rect 19796 48390 19798 48442
rect 19636 48388 19660 48390
rect 19716 48388 19740 48390
rect 19796 48388 19820 48390
rect 19580 48368 19876 48388
rect 19432 48204 19484 48210
rect 19432 48146 19484 48152
rect 19444 47802 19472 48146
rect 19904 48074 19932 48572
rect 19996 48278 20024 48622
rect 19984 48272 20036 48278
rect 19984 48214 20036 48220
rect 19984 48136 20036 48142
rect 19984 48078 20036 48084
rect 19892 48068 19944 48074
rect 19892 48010 19944 48016
rect 19432 47796 19484 47802
rect 19432 47738 19484 47744
rect 19444 47258 19472 47738
rect 19580 47356 19876 47376
rect 19636 47354 19660 47356
rect 19716 47354 19740 47356
rect 19796 47354 19820 47356
rect 19658 47302 19660 47354
rect 19722 47302 19734 47354
rect 19796 47302 19798 47354
rect 19636 47300 19660 47302
rect 19716 47300 19740 47302
rect 19796 47300 19820 47302
rect 19580 47280 19876 47300
rect 19432 47252 19484 47258
rect 19432 47194 19484 47200
rect 19904 47122 19932 48010
rect 19892 47116 19944 47122
rect 19892 47058 19944 47064
rect 19904 46714 19932 47058
rect 19996 47025 20024 48078
rect 20088 47802 20116 48826
rect 20076 47796 20128 47802
rect 20076 47738 20128 47744
rect 20076 47456 20128 47462
rect 20076 47398 20128 47404
rect 19982 47016 20038 47025
rect 19982 46951 20038 46960
rect 20088 46889 20116 47398
rect 20074 46880 20130 46889
rect 20074 46815 20130 46824
rect 19892 46708 19944 46714
rect 19892 46650 19944 46656
rect 19580 46268 19876 46288
rect 19636 46266 19660 46268
rect 19716 46266 19740 46268
rect 19796 46266 19820 46268
rect 19658 46214 19660 46266
rect 19722 46214 19734 46266
rect 19796 46214 19798 46266
rect 19636 46212 19660 46214
rect 19716 46212 19740 46214
rect 19796 46212 19820 46214
rect 19338 46200 19394 46209
rect 19580 46192 19876 46212
rect 19338 46135 19394 46144
rect 19580 45180 19876 45200
rect 19636 45178 19660 45180
rect 19716 45178 19740 45180
rect 19796 45178 19820 45180
rect 19658 45126 19660 45178
rect 19722 45126 19734 45178
rect 19796 45126 19798 45178
rect 19636 45124 19660 45126
rect 19716 45124 19740 45126
rect 19796 45124 19820 45126
rect 19580 45104 19876 45124
rect 19580 44092 19876 44112
rect 19636 44090 19660 44092
rect 19716 44090 19740 44092
rect 19796 44090 19820 44092
rect 19658 44038 19660 44090
rect 19722 44038 19734 44090
rect 19796 44038 19798 44090
rect 19636 44036 19660 44038
rect 19716 44036 19740 44038
rect 19796 44036 19820 44038
rect 19580 44016 19876 44036
rect 19246 43208 19302 43217
rect 19246 43143 19302 43152
rect 18878 42392 18934 42401
rect 18878 42327 18934 42336
rect 19064 42016 19116 42022
rect 19064 41958 19116 41964
rect 19076 41614 19104 41958
rect 19064 41608 19116 41614
rect 19064 41550 19116 41556
rect 18972 40928 19024 40934
rect 18972 40870 19024 40876
rect 18984 40594 19012 40870
rect 19260 40769 19288 43143
rect 19580 43004 19876 43024
rect 19636 43002 19660 43004
rect 19716 43002 19740 43004
rect 19796 43002 19820 43004
rect 19658 42950 19660 43002
rect 19722 42950 19734 43002
rect 19796 42950 19798 43002
rect 19636 42948 19660 42950
rect 19716 42948 19740 42950
rect 19796 42948 19820 42950
rect 19580 42928 19876 42948
rect 19708 42560 19760 42566
rect 19708 42502 19760 42508
rect 19720 42158 19748 42502
rect 19708 42152 19760 42158
rect 19760 42100 19932 42106
rect 19708 42094 19932 42100
rect 19720 42078 19932 42094
rect 19340 42016 19392 42022
rect 19340 41958 19392 41964
rect 19352 41070 19380 41958
rect 19580 41916 19876 41936
rect 19636 41914 19660 41916
rect 19716 41914 19740 41916
rect 19796 41914 19820 41916
rect 19658 41862 19660 41914
rect 19722 41862 19734 41914
rect 19796 41862 19798 41914
rect 19636 41860 19660 41862
rect 19716 41860 19740 41862
rect 19796 41860 19820 41862
rect 19580 41840 19876 41860
rect 19904 41682 19932 42078
rect 19892 41676 19944 41682
rect 19892 41618 19944 41624
rect 19524 41608 19576 41614
rect 19524 41550 19576 41556
rect 19432 41472 19484 41478
rect 19432 41414 19484 41420
rect 19340 41064 19392 41070
rect 19340 41006 19392 41012
rect 19246 40760 19302 40769
rect 19246 40695 19302 40704
rect 19444 40610 19472 41414
rect 19536 41002 19564 41550
rect 19904 41206 19932 41618
rect 19892 41200 19944 41206
rect 19892 41142 19944 41148
rect 19904 41070 19932 41142
rect 19892 41064 19944 41070
rect 19892 41006 19944 41012
rect 19524 40996 19576 41002
rect 19524 40938 19576 40944
rect 19580 40828 19876 40848
rect 19636 40826 19660 40828
rect 19716 40826 19740 40828
rect 19796 40826 19820 40828
rect 19658 40774 19660 40826
rect 19722 40774 19734 40826
rect 19796 40774 19798 40826
rect 19636 40772 19660 40774
rect 19716 40772 19740 40774
rect 19796 40772 19820 40774
rect 19580 40752 19876 40772
rect 19352 40594 19472 40610
rect 18972 40588 19024 40594
rect 18972 40530 19024 40536
rect 19340 40588 19472 40594
rect 19392 40582 19472 40588
rect 19708 40588 19760 40594
rect 19340 40530 19392 40536
rect 19708 40530 19760 40536
rect 19984 40588 20036 40594
rect 19984 40530 20036 40536
rect 20076 40588 20128 40594
rect 20076 40530 20128 40536
rect 19720 40458 19748 40530
rect 19708 40452 19760 40458
rect 19708 40394 19760 40400
rect 19340 40384 19392 40390
rect 19340 40326 19392 40332
rect 19062 39672 19118 39681
rect 19062 39607 19064 39616
rect 19116 39607 19118 39616
rect 19064 39578 19116 39584
rect 19076 38962 19104 39578
rect 19352 39098 19380 40326
rect 19720 39953 19748 40394
rect 19706 39944 19762 39953
rect 19706 39879 19762 39888
rect 19580 39740 19876 39760
rect 19636 39738 19660 39740
rect 19716 39738 19740 39740
rect 19796 39738 19820 39740
rect 19658 39686 19660 39738
rect 19722 39686 19734 39738
rect 19796 39686 19798 39738
rect 19636 39684 19660 39686
rect 19716 39684 19740 39686
rect 19796 39684 19820 39686
rect 19580 39664 19876 39684
rect 19996 39574 20024 40530
rect 20088 40050 20116 40530
rect 20076 40044 20128 40050
rect 20076 39986 20128 39992
rect 19984 39568 20036 39574
rect 19984 39510 20036 39516
rect 19892 39500 19944 39506
rect 19892 39442 19944 39448
rect 19340 39092 19392 39098
rect 19340 39034 19392 39040
rect 19064 38956 19116 38962
rect 19064 38898 19116 38904
rect 19156 38888 19208 38894
rect 19156 38830 19208 38836
rect 18694 38720 18750 38729
rect 18694 38655 18750 38664
rect 19168 38418 19196 38830
rect 19904 38826 19932 39442
rect 19984 39024 20036 39030
rect 19984 38966 20036 38972
rect 19892 38820 19944 38826
rect 19892 38762 19944 38768
rect 19580 38652 19876 38672
rect 19636 38650 19660 38652
rect 19716 38650 19740 38652
rect 19796 38650 19820 38652
rect 19658 38598 19660 38650
rect 19722 38598 19734 38650
rect 19796 38598 19798 38650
rect 19636 38596 19660 38598
rect 19716 38596 19740 38598
rect 19796 38596 19820 38598
rect 19580 38576 19876 38596
rect 19996 38554 20024 38966
rect 20088 38894 20116 39986
rect 20076 38888 20128 38894
rect 20076 38830 20128 38836
rect 19340 38548 19392 38554
rect 19340 38490 19392 38496
rect 19984 38548 20036 38554
rect 19984 38490 20036 38496
rect 19064 38412 19116 38418
rect 19064 38354 19116 38360
rect 19156 38412 19208 38418
rect 19156 38354 19208 38360
rect 18786 38312 18842 38321
rect 18786 38247 18842 38256
rect 18800 38214 18828 38247
rect 18788 38208 18840 38214
rect 18788 38150 18840 38156
rect 18602 37904 18658 37913
rect 18602 37839 18658 37848
rect 18420 37800 18472 37806
rect 18420 37742 18472 37748
rect 18432 37618 18460 37742
rect 18432 37590 18552 37618
rect 18524 37466 18552 37590
rect 18420 37460 18472 37466
rect 18420 37402 18472 37408
rect 18512 37460 18564 37466
rect 18512 37402 18564 37408
rect 18432 37369 18460 37402
rect 18418 37360 18474 37369
rect 18418 37295 18474 37304
rect 18616 37176 18644 37839
rect 18800 37806 18828 38150
rect 19076 37806 19104 38354
rect 18788 37800 18840 37806
rect 18788 37742 18840 37748
rect 18880 37800 18932 37806
rect 19064 37800 19116 37806
rect 18880 37742 18932 37748
rect 18970 37768 19026 37777
rect 18432 37148 18644 37176
rect 18328 36304 18380 36310
rect 18328 36246 18380 36252
rect 18236 36032 18288 36038
rect 18236 35974 18288 35980
rect 18248 34066 18276 35974
rect 18328 35624 18380 35630
rect 18328 35566 18380 35572
rect 18340 34746 18368 35566
rect 18328 34740 18380 34746
rect 18328 34682 18380 34688
rect 18326 34640 18382 34649
rect 18326 34575 18382 34584
rect 18340 34134 18368 34575
rect 18328 34128 18380 34134
rect 18328 34070 18380 34076
rect 18236 34060 18288 34066
rect 18236 34002 18288 34008
rect 18248 33658 18276 34002
rect 18236 33652 18288 33658
rect 18236 33594 18288 33600
rect 18248 33318 18276 33594
rect 18326 33552 18382 33561
rect 18326 33487 18382 33496
rect 18236 33312 18288 33318
rect 18236 33254 18288 33260
rect 18340 32910 18368 33487
rect 18328 32904 18380 32910
rect 18328 32846 18380 32852
rect 18328 32768 18380 32774
rect 18328 32710 18380 32716
rect 18340 32473 18368 32710
rect 18326 32464 18382 32473
rect 18326 32399 18382 32408
rect 18432 32366 18460 37148
rect 18786 37088 18842 37097
rect 18786 37023 18842 37032
rect 18512 36576 18564 36582
rect 18512 36518 18564 36524
rect 18420 32360 18472 32366
rect 18420 32302 18472 32308
rect 18420 32224 18472 32230
rect 18420 32166 18472 32172
rect 18326 31920 18382 31929
rect 18326 31855 18328 31864
rect 18380 31855 18382 31864
rect 18328 31826 18380 31832
rect 18432 31793 18460 32166
rect 18234 31784 18290 31793
rect 18234 31719 18290 31728
rect 18418 31784 18474 31793
rect 18418 31719 18474 31728
rect 18248 30734 18276 31719
rect 18524 31634 18552 36518
rect 18602 36272 18658 36281
rect 18602 36207 18658 36216
rect 18616 33114 18644 36207
rect 18696 34944 18748 34950
rect 18696 34886 18748 34892
rect 18708 34678 18736 34886
rect 18696 34672 18748 34678
rect 18696 34614 18748 34620
rect 18708 34202 18736 34614
rect 18800 34354 18828 37023
rect 18892 36718 18920 37742
rect 19064 37742 19116 37748
rect 18970 37703 19026 37712
rect 18984 37330 19012 37703
rect 19156 37664 19208 37670
rect 19156 37606 19208 37612
rect 19168 37330 19196 37606
rect 18972 37324 19024 37330
rect 18972 37266 19024 37272
rect 19156 37324 19208 37330
rect 19156 37266 19208 37272
rect 18880 36712 18932 36718
rect 18880 36654 18932 36660
rect 18984 36378 19012 37266
rect 19064 36576 19116 36582
rect 19352 36530 19380 38490
rect 19798 38040 19854 38049
rect 19798 37975 19800 37984
rect 19852 37975 19854 37984
rect 19800 37946 19852 37952
rect 20076 37800 20128 37806
rect 20076 37742 20128 37748
rect 19984 37732 20036 37738
rect 19984 37674 20036 37680
rect 19580 37564 19876 37584
rect 19636 37562 19660 37564
rect 19716 37562 19740 37564
rect 19796 37562 19820 37564
rect 19658 37510 19660 37562
rect 19722 37510 19734 37562
rect 19796 37510 19798 37562
rect 19636 37508 19660 37510
rect 19716 37508 19740 37510
rect 19796 37508 19820 37510
rect 19580 37488 19876 37508
rect 19996 37398 20024 37674
rect 20088 37641 20116 37742
rect 20074 37632 20130 37641
rect 20074 37567 20130 37576
rect 19984 37392 20036 37398
rect 19984 37334 20036 37340
rect 19996 36922 20024 37334
rect 19984 36916 20036 36922
rect 19984 36858 20036 36864
rect 19064 36518 19116 36524
rect 18972 36372 19024 36378
rect 18972 36314 19024 36320
rect 18880 36236 18932 36242
rect 18880 36178 18932 36184
rect 18892 35494 18920 36178
rect 18880 35488 18932 35494
rect 18880 35430 18932 35436
rect 18892 35154 18920 35430
rect 18880 35148 18932 35154
rect 18880 35090 18932 35096
rect 18892 34542 18920 35090
rect 18880 34536 18932 34542
rect 18880 34478 18932 34484
rect 18800 34326 19012 34354
rect 18696 34196 18748 34202
rect 18696 34138 18748 34144
rect 18694 33688 18750 33697
rect 18694 33623 18750 33632
rect 18708 33454 18736 33623
rect 18696 33448 18748 33454
rect 18696 33390 18748 33396
rect 18788 33380 18840 33386
rect 18788 33322 18840 33328
rect 18604 33108 18656 33114
rect 18604 33050 18656 33056
rect 18694 33008 18750 33017
rect 18694 32943 18750 32952
rect 18432 31606 18552 31634
rect 18328 30932 18380 30938
rect 18328 30874 18380 30880
rect 18236 30728 18288 30734
rect 18236 30670 18288 30676
rect 18248 30394 18276 30670
rect 18236 30388 18288 30394
rect 18236 30330 18288 30336
rect 18234 30288 18290 30297
rect 18234 30223 18290 30232
rect 18248 28218 18276 30223
rect 18340 30054 18368 30874
rect 18432 30569 18460 31606
rect 18510 31512 18566 31521
rect 18510 31447 18566 31456
rect 18418 30560 18474 30569
rect 18418 30495 18474 30504
rect 18420 30116 18472 30122
rect 18420 30058 18472 30064
rect 18328 30048 18380 30054
rect 18328 29990 18380 29996
rect 18432 29782 18460 30058
rect 18420 29776 18472 29782
rect 18420 29718 18472 29724
rect 18420 29028 18472 29034
rect 18420 28970 18472 28976
rect 18432 28801 18460 28970
rect 18418 28792 18474 28801
rect 18418 28727 18474 28736
rect 18328 28620 18380 28626
rect 18328 28562 18380 28568
rect 18236 28212 18288 28218
rect 18236 28154 18288 28160
rect 18340 27674 18368 28562
rect 18328 27668 18380 27674
rect 18328 27610 18380 27616
rect 18236 26240 18288 26246
rect 18236 26182 18288 26188
rect 18248 25906 18276 26182
rect 18236 25900 18288 25906
rect 18236 25842 18288 25848
rect 18234 24168 18290 24177
rect 18234 24103 18290 24112
rect 18248 22030 18276 24103
rect 18340 23905 18368 27610
rect 18524 26586 18552 31447
rect 18604 31204 18656 31210
rect 18604 31146 18656 31152
rect 18616 30802 18644 31146
rect 18708 30938 18736 32943
rect 18800 32881 18828 33322
rect 18786 32872 18842 32881
rect 18786 32807 18788 32816
rect 18840 32807 18842 32816
rect 18788 32778 18840 32784
rect 18800 32747 18828 32778
rect 18880 32768 18932 32774
rect 18880 32710 18932 32716
rect 18786 32600 18842 32609
rect 18786 32535 18842 32544
rect 18800 32065 18828 32535
rect 18892 32502 18920 32710
rect 18880 32496 18932 32502
rect 18880 32438 18932 32444
rect 18786 32056 18842 32065
rect 18984 32026 19012 34326
rect 19076 32774 19104 36518
rect 19168 36502 19380 36530
rect 19984 36576 20036 36582
rect 19984 36518 20036 36524
rect 19168 36038 19196 36502
rect 19580 36476 19876 36496
rect 19636 36474 19660 36476
rect 19716 36474 19740 36476
rect 19796 36474 19820 36476
rect 19658 36422 19660 36474
rect 19722 36422 19734 36474
rect 19796 36422 19798 36474
rect 19636 36420 19660 36422
rect 19716 36420 19740 36422
rect 19796 36420 19820 36422
rect 19338 36408 19394 36417
rect 19580 36400 19876 36420
rect 19338 36343 19394 36352
rect 19352 36242 19380 36343
rect 19340 36236 19392 36242
rect 19340 36178 19392 36184
rect 19248 36100 19300 36106
rect 19248 36042 19300 36048
rect 19156 36032 19208 36038
rect 19156 35974 19208 35980
rect 19154 35864 19210 35873
rect 19154 35799 19210 35808
rect 19168 35154 19196 35799
rect 19260 35630 19288 36042
rect 19432 36032 19484 36038
rect 19338 36000 19394 36009
rect 19432 35974 19484 35980
rect 19338 35935 19394 35944
rect 19248 35624 19300 35630
rect 19248 35566 19300 35572
rect 19352 35290 19380 35935
rect 19444 35698 19472 35974
rect 19432 35692 19484 35698
rect 19432 35634 19484 35640
rect 19340 35284 19392 35290
rect 19340 35226 19392 35232
rect 19444 35222 19472 35634
rect 19892 35556 19944 35562
rect 19892 35498 19944 35504
rect 19580 35388 19876 35408
rect 19636 35386 19660 35388
rect 19716 35386 19740 35388
rect 19796 35386 19820 35388
rect 19658 35334 19660 35386
rect 19722 35334 19734 35386
rect 19796 35334 19798 35386
rect 19636 35332 19660 35334
rect 19716 35332 19740 35334
rect 19796 35332 19820 35334
rect 19580 35312 19876 35332
rect 19432 35216 19484 35222
rect 19338 35184 19394 35193
rect 19156 35148 19208 35154
rect 19432 35158 19484 35164
rect 19338 35119 19340 35128
rect 19156 35090 19208 35096
rect 19392 35119 19394 35128
rect 19340 35090 19392 35096
rect 19340 35012 19392 35018
rect 19340 34954 19392 34960
rect 19352 34241 19380 34954
rect 19616 34944 19668 34950
rect 19616 34886 19668 34892
rect 19628 34785 19656 34886
rect 19614 34776 19670 34785
rect 19904 34746 19932 35498
rect 19614 34711 19670 34720
rect 19892 34740 19944 34746
rect 19628 34542 19656 34711
rect 19892 34682 19944 34688
rect 19616 34536 19668 34542
rect 19616 34478 19668 34484
rect 19432 34468 19484 34474
rect 19432 34410 19484 34416
rect 19338 34232 19394 34241
rect 19338 34167 19394 34176
rect 19248 34128 19300 34134
rect 19248 34070 19300 34076
rect 19156 33856 19208 33862
rect 19156 33798 19208 33804
rect 19168 33386 19196 33798
rect 19156 33380 19208 33386
rect 19156 33322 19208 33328
rect 19154 33280 19210 33289
rect 19260 33266 19288 34070
rect 19444 33969 19472 34410
rect 19580 34300 19876 34320
rect 19636 34298 19660 34300
rect 19716 34298 19740 34300
rect 19796 34298 19820 34300
rect 19658 34246 19660 34298
rect 19722 34246 19734 34298
rect 19796 34246 19798 34298
rect 19636 34244 19660 34246
rect 19716 34244 19740 34246
rect 19796 34244 19820 34246
rect 19580 34224 19876 34244
rect 19430 33960 19486 33969
rect 19430 33895 19486 33904
rect 19614 33960 19670 33969
rect 19614 33895 19670 33904
rect 19340 33856 19392 33862
rect 19340 33798 19392 33804
rect 19210 33238 19288 33266
rect 19154 33215 19210 33224
rect 19064 32768 19116 32774
rect 19064 32710 19116 32716
rect 19064 32292 19116 32298
rect 19064 32234 19116 32240
rect 18786 31991 18842 32000
rect 18972 32020 19024 32026
rect 18800 31906 18828 31991
rect 18972 31962 19024 31968
rect 18800 31878 19012 31906
rect 18880 31816 18932 31822
rect 18880 31758 18932 31764
rect 18892 31385 18920 31758
rect 18878 31376 18934 31385
rect 18878 31311 18934 31320
rect 18696 30932 18748 30938
rect 18696 30874 18748 30880
rect 18604 30796 18656 30802
rect 18604 30738 18656 30744
rect 18616 30705 18644 30738
rect 18602 30696 18658 30705
rect 18602 30631 18658 30640
rect 18788 30592 18840 30598
rect 18788 30534 18840 30540
rect 18800 30161 18828 30534
rect 18984 30190 19012 31878
rect 19076 31346 19104 32234
rect 19064 31340 19116 31346
rect 19064 31282 19116 31288
rect 19062 30696 19118 30705
rect 19062 30631 19118 30640
rect 19076 30326 19104 30631
rect 19064 30320 19116 30326
rect 19064 30262 19116 30268
rect 18972 30184 19024 30190
rect 18786 30152 18842 30161
rect 18972 30126 19024 30132
rect 18786 30087 18788 30096
rect 18840 30087 18842 30096
rect 18788 30058 18840 30064
rect 18880 30048 18932 30054
rect 18880 29990 18932 29996
rect 18696 29844 18748 29850
rect 18696 29786 18748 29792
rect 18604 29028 18656 29034
rect 18604 28970 18656 28976
rect 18616 28558 18644 28970
rect 18708 28966 18736 29786
rect 18788 29504 18840 29510
rect 18788 29446 18840 29452
rect 18800 29102 18828 29446
rect 18788 29096 18840 29102
rect 18788 29038 18840 29044
rect 18696 28960 18748 28966
rect 18696 28902 18748 28908
rect 18708 28762 18736 28902
rect 18892 28762 18920 29990
rect 19064 29640 19116 29646
rect 19064 29582 19116 29588
rect 18970 29472 19026 29481
rect 18970 29407 19026 29416
rect 18696 28756 18748 28762
rect 18696 28698 18748 28704
rect 18880 28756 18932 28762
rect 18880 28698 18932 28704
rect 18604 28552 18656 28558
rect 18604 28494 18656 28500
rect 18616 28422 18644 28494
rect 18604 28416 18656 28422
rect 18604 28358 18656 28364
rect 18616 27674 18644 28358
rect 18604 27668 18656 27674
rect 18604 27610 18656 27616
rect 18708 27305 18736 28698
rect 18984 28694 19012 29407
rect 18972 28688 19024 28694
rect 18878 28656 18934 28665
rect 18972 28630 19024 28636
rect 18878 28591 18880 28600
rect 18932 28591 18934 28600
rect 18880 28562 18932 28568
rect 18972 28552 19024 28558
rect 18972 28494 19024 28500
rect 18878 28384 18934 28393
rect 18878 28319 18934 28328
rect 18892 28218 18920 28319
rect 18880 28212 18932 28218
rect 18880 28154 18932 28160
rect 18786 28112 18842 28121
rect 18786 28047 18842 28056
rect 18694 27296 18750 27305
rect 18694 27231 18750 27240
rect 18800 27130 18828 28047
rect 18892 28014 18920 28154
rect 18880 28008 18932 28014
rect 18880 27950 18932 27956
rect 18984 27538 19012 28494
rect 18972 27532 19024 27538
rect 18972 27474 19024 27480
rect 18984 27441 19012 27474
rect 18970 27432 19026 27441
rect 18970 27367 19026 27376
rect 18788 27124 18840 27130
rect 18788 27066 18840 27072
rect 18800 26926 18828 27066
rect 18788 26920 18840 26926
rect 18788 26862 18840 26868
rect 18880 26784 18932 26790
rect 18880 26726 18932 26732
rect 18512 26580 18564 26586
rect 18512 26522 18564 26528
rect 18512 26444 18564 26450
rect 18512 26386 18564 26392
rect 18524 25974 18552 26386
rect 18604 26376 18656 26382
rect 18604 26318 18656 26324
rect 18512 25968 18564 25974
rect 18512 25910 18564 25916
rect 18524 25430 18552 25910
rect 18512 25424 18564 25430
rect 18512 25366 18564 25372
rect 18326 23896 18382 23905
rect 18326 23831 18328 23840
rect 18380 23831 18382 23840
rect 18328 23802 18380 23808
rect 18340 23771 18368 23802
rect 18512 23656 18564 23662
rect 18512 23598 18564 23604
rect 18524 23322 18552 23598
rect 18512 23316 18564 23322
rect 18512 23258 18564 23264
rect 18616 22982 18644 26318
rect 18696 25832 18748 25838
rect 18694 25800 18696 25809
rect 18788 25832 18840 25838
rect 18748 25800 18750 25809
rect 18788 25774 18840 25780
rect 18694 25735 18750 25744
rect 18800 25673 18828 25774
rect 18786 25664 18842 25673
rect 18786 25599 18842 25608
rect 18800 25158 18828 25599
rect 18788 25152 18840 25158
rect 18788 25094 18840 25100
rect 18694 24984 18750 24993
rect 18694 24919 18750 24928
rect 18708 24750 18736 24919
rect 18696 24744 18748 24750
rect 18696 24686 18748 24692
rect 18800 24596 18828 25094
rect 18708 24568 18828 24596
rect 18604 22976 18656 22982
rect 18604 22918 18656 22924
rect 18420 22704 18472 22710
rect 18420 22646 18472 22652
rect 18326 22536 18382 22545
rect 18326 22471 18328 22480
rect 18380 22471 18382 22480
rect 18328 22442 18380 22448
rect 18236 22024 18288 22030
rect 18432 22001 18460 22646
rect 18616 22574 18644 22918
rect 18604 22568 18656 22574
rect 18604 22510 18656 22516
rect 18512 22500 18564 22506
rect 18512 22442 18564 22448
rect 18524 22409 18552 22442
rect 18510 22400 18566 22409
rect 18510 22335 18566 22344
rect 18602 22128 18658 22137
rect 18602 22063 18658 22072
rect 18236 21966 18288 21972
rect 18418 21992 18474 22001
rect 18418 21927 18474 21936
rect 18156 21814 18552 21842
rect 18052 21140 18104 21146
rect 18052 21082 18104 21088
rect 17684 21004 17736 21010
rect 17684 20946 17736 20952
rect 17696 20602 17724 20946
rect 18328 20936 18380 20942
rect 18328 20878 18380 20884
rect 17960 20800 18012 20806
rect 17960 20742 18012 20748
rect 17684 20596 17736 20602
rect 17684 20538 17736 20544
rect 17868 20596 17920 20602
rect 17972 20584 18000 20742
rect 17920 20556 18000 20584
rect 17868 20538 17920 20544
rect 17592 20460 17644 20466
rect 17592 20402 17644 20408
rect 17684 19984 17736 19990
rect 17684 19926 17736 19932
rect 17696 19174 17724 19926
rect 17776 19848 17828 19854
rect 17776 19790 17828 19796
rect 17684 19168 17736 19174
rect 17684 19110 17736 19116
rect 17788 18970 17816 19790
rect 17776 18964 17828 18970
rect 17776 18906 17828 18912
rect 17500 18624 17552 18630
rect 17500 18566 17552 18572
rect 17512 17746 17540 18566
rect 17880 17814 17908 20538
rect 18340 19922 18368 20878
rect 17960 19916 18012 19922
rect 17960 19858 18012 19864
rect 18144 19916 18196 19922
rect 18144 19858 18196 19864
rect 18328 19916 18380 19922
rect 18328 19858 18380 19864
rect 17972 19174 18000 19858
rect 18156 19825 18184 19858
rect 18142 19816 18198 19825
rect 18142 19751 18198 19760
rect 18156 19310 18184 19751
rect 18144 19304 18196 19310
rect 18144 19246 18196 19252
rect 17960 19168 18012 19174
rect 17960 19110 18012 19116
rect 17960 18964 18012 18970
rect 17960 18906 18012 18912
rect 17972 18465 18000 18906
rect 17958 18456 18014 18465
rect 18156 18426 18184 19246
rect 18420 19236 18472 19242
rect 18420 19178 18472 19184
rect 18432 18834 18460 19178
rect 18420 18828 18472 18834
rect 18420 18770 18472 18776
rect 17958 18391 18014 18400
rect 18144 18420 18196 18426
rect 18144 18362 18196 18368
rect 17960 18148 18012 18154
rect 17960 18090 18012 18096
rect 17868 17808 17920 17814
rect 17868 17750 17920 17756
rect 17500 17740 17552 17746
rect 17500 17682 17552 17688
rect 17512 17338 17540 17682
rect 17500 17332 17552 17338
rect 17500 17274 17552 17280
rect 17052 17224 17448 17252
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 16396 16584 16448 16590
rect 16396 16526 16448 16532
rect 16764 16584 16816 16590
rect 16764 16526 16816 16532
rect 16408 15978 16436 16526
rect 16396 15972 16448 15978
rect 16396 15914 16448 15920
rect 15844 15360 15896 15366
rect 15844 15302 15896 15308
rect 15856 14958 15884 15302
rect 16856 15156 16908 15162
rect 16856 15098 16908 15104
rect 16028 15088 16080 15094
rect 16028 15030 16080 15036
rect 15844 14952 15896 14958
rect 15844 14894 15896 14900
rect 15856 14550 15884 14894
rect 15844 14544 15896 14550
rect 15844 14486 15896 14492
rect 15936 12912 15988 12918
rect 15936 12854 15988 12860
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15752 12096 15804 12102
rect 15752 12038 15804 12044
rect 15304 11694 15332 12038
rect 15948 11898 15976 12854
rect 15936 11892 15988 11898
rect 15936 11834 15988 11840
rect 15292 11688 15344 11694
rect 15292 11630 15344 11636
rect 15304 11286 15332 11630
rect 15292 11280 15344 11286
rect 15292 11222 15344 11228
rect 15304 10810 15332 11222
rect 15844 11076 15896 11082
rect 15844 11018 15896 11024
rect 15292 10804 15344 10810
rect 15292 10746 15344 10752
rect 15566 8528 15622 8537
rect 15566 8463 15622 8472
rect 14832 3188 14884 3194
rect 14832 3130 14884 3136
rect 15580 898 15608 8463
rect 15856 4049 15884 11018
rect 16040 5273 16068 15030
rect 16868 14958 16896 15098
rect 16856 14952 16908 14958
rect 16856 14894 16908 14900
rect 16486 13424 16542 13433
rect 16486 13359 16542 13368
rect 16764 13388 16816 13394
rect 16500 13326 16528 13359
rect 16764 13330 16816 13336
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 16488 13320 16540 13326
rect 16488 13262 16540 13268
rect 16580 13320 16632 13326
rect 16580 13262 16632 13268
rect 16592 12986 16620 13262
rect 16580 12980 16632 12986
rect 16580 12922 16632 12928
rect 16776 12850 16804 13330
rect 16960 12986 16988 13330
rect 16948 12980 17000 12986
rect 16948 12922 17000 12928
rect 16764 12844 16816 12850
rect 16764 12786 16816 12792
rect 16396 12232 16448 12238
rect 16396 12174 16448 12180
rect 16408 11898 16436 12174
rect 16396 11892 16448 11898
rect 16396 11834 16448 11840
rect 16212 11552 16264 11558
rect 16212 11494 16264 11500
rect 16224 11218 16252 11494
rect 16776 11234 16804 12786
rect 16212 11212 16264 11218
rect 16212 11154 16264 11160
rect 16408 11206 16804 11234
rect 16224 10810 16252 11154
rect 16408 11150 16436 11206
rect 16396 11144 16448 11150
rect 16396 11086 16448 11092
rect 16488 11144 16540 11150
rect 16488 11086 16540 11092
rect 16212 10804 16264 10810
rect 16212 10746 16264 10752
rect 16408 10742 16436 11086
rect 16396 10736 16448 10742
rect 16396 10678 16448 10684
rect 16500 10674 16528 11086
rect 16488 10668 16540 10674
rect 16488 10610 16540 10616
rect 17052 9761 17080 17224
rect 17512 17134 17540 17274
rect 17880 17270 17908 17750
rect 17972 17746 18000 18090
rect 18432 17882 18460 18770
rect 18420 17876 18472 17882
rect 18340 17836 18420 17864
rect 17960 17740 18012 17746
rect 17960 17682 18012 17688
rect 17868 17264 17920 17270
rect 17868 17206 17920 17212
rect 17500 17128 17552 17134
rect 17500 17070 17552 17076
rect 17316 17060 17368 17066
rect 17316 17002 17368 17008
rect 17328 13394 17356 17002
rect 17512 16658 17540 17070
rect 18340 16658 18368 17836
rect 18420 17818 18472 17824
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 17500 16652 17552 16658
rect 17500 16594 17552 16600
rect 17684 16652 17736 16658
rect 17684 16594 17736 16600
rect 18328 16652 18380 16658
rect 18328 16594 18380 16600
rect 17512 16250 17540 16594
rect 17500 16244 17552 16250
rect 17500 16186 17552 16192
rect 17696 16182 17724 16594
rect 17960 16448 18012 16454
rect 17960 16390 18012 16396
rect 17684 16176 17736 16182
rect 17684 16118 17736 16124
rect 17972 15706 18000 16390
rect 18050 15736 18106 15745
rect 17960 15700 18012 15706
rect 18050 15671 18106 15680
rect 17960 15642 18012 15648
rect 17972 15026 18000 15642
rect 18064 15638 18092 15671
rect 18052 15632 18104 15638
rect 18052 15574 18104 15580
rect 17960 15020 18012 15026
rect 17960 14962 18012 14968
rect 17972 14482 18000 14962
rect 18064 14958 18092 15574
rect 18326 15192 18382 15201
rect 18326 15127 18328 15136
rect 18380 15127 18382 15136
rect 18328 15098 18380 15104
rect 18052 14952 18104 14958
rect 18052 14894 18104 14900
rect 17960 14476 18012 14482
rect 17960 14418 18012 14424
rect 17500 14408 17552 14414
rect 17500 14350 17552 14356
rect 17316 13388 17368 13394
rect 17316 13330 17368 13336
rect 17132 12980 17184 12986
rect 17132 12922 17184 12928
rect 17144 12442 17172 12922
rect 17328 12918 17356 13330
rect 17316 12912 17368 12918
rect 17316 12854 17368 12860
rect 17132 12436 17184 12442
rect 17132 12378 17184 12384
rect 17512 12306 17540 14350
rect 17972 14074 18000 14418
rect 17960 14068 18012 14074
rect 17960 14010 18012 14016
rect 18064 13546 18092 14894
rect 18340 14414 18368 14445
rect 18328 14408 18380 14414
rect 18326 14376 18328 14385
rect 18380 14376 18382 14385
rect 18326 14311 18382 14320
rect 18340 14074 18368 14311
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 17880 13518 18092 13546
rect 17880 13462 17908 13518
rect 17868 13456 17920 13462
rect 17868 13398 17920 13404
rect 17500 12300 17552 12306
rect 17500 12242 17552 12248
rect 17512 11898 17540 12242
rect 18064 12238 18092 13518
rect 18432 12374 18460 17478
rect 18420 12368 18472 12374
rect 18420 12310 18472 12316
rect 18052 12232 18104 12238
rect 18052 12174 18104 12180
rect 18328 12232 18380 12238
rect 18328 12174 18380 12180
rect 17868 12096 17920 12102
rect 17868 12038 17920 12044
rect 17500 11892 17552 11898
rect 17500 11834 17552 11840
rect 17512 11150 17540 11834
rect 17880 11150 17908 12038
rect 18340 11898 18368 12174
rect 18432 12102 18460 12310
rect 18420 12096 18472 12102
rect 18420 12038 18472 12044
rect 18328 11892 18380 11898
rect 18328 11834 18380 11840
rect 17500 11144 17552 11150
rect 17500 11086 17552 11092
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17512 10742 17540 11086
rect 17880 10810 17908 11086
rect 17868 10804 17920 10810
rect 17868 10746 17920 10752
rect 17500 10736 17552 10742
rect 17500 10678 17552 10684
rect 18236 10736 18288 10742
rect 18236 10678 18288 10684
rect 16118 9752 16174 9761
rect 16118 9687 16174 9696
rect 17038 9752 17094 9761
rect 17038 9687 17094 9696
rect 16026 5264 16082 5273
rect 16026 5199 16082 5208
rect 15842 4040 15898 4049
rect 15842 3975 15898 3984
rect 15580 870 15700 898
rect 15672 800 15700 870
rect 16132 800 16160 9687
rect 17960 4140 18012 4146
rect 17960 4082 18012 4088
rect 17038 4040 17094 4049
rect 17038 3975 17094 3984
rect 17052 800 17080 3975
rect 17972 800 18000 4082
rect 18248 3369 18276 10678
rect 18524 9081 18552 21814
rect 18616 21146 18644 22063
rect 18708 21894 18736 24568
rect 18788 24336 18840 24342
rect 18892 24324 18920 26726
rect 18972 26512 19024 26518
rect 18970 26480 18972 26489
rect 19024 26480 19026 26489
rect 18970 26415 19026 26424
rect 19076 26042 19104 29582
rect 19168 29306 19196 33215
rect 19248 32360 19300 32366
rect 19248 32302 19300 32308
rect 19260 30938 19288 32302
rect 19352 31822 19380 33798
rect 19444 33658 19472 33895
rect 19432 33652 19484 33658
rect 19432 33594 19484 33600
rect 19628 33522 19656 33895
rect 19616 33516 19668 33522
rect 19616 33458 19668 33464
rect 19432 33448 19484 33454
rect 19432 33390 19484 33396
rect 19444 32978 19472 33390
rect 19580 33212 19876 33232
rect 19636 33210 19660 33212
rect 19716 33210 19740 33212
rect 19796 33210 19820 33212
rect 19658 33158 19660 33210
rect 19722 33158 19734 33210
rect 19796 33158 19798 33210
rect 19636 33156 19660 33158
rect 19716 33156 19740 33158
rect 19796 33156 19820 33158
rect 19580 33136 19876 33156
rect 19432 32972 19484 32978
rect 19432 32914 19484 32920
rect 19616 32836 19668 32842
rect 19616 32778 19668 32784
rect 19432 32768 19484 32774
rect 19432 32710 19484 32716
rect 19340 31816 19392 31822
rect 19340 31758 19392 31764
rect 19340 31680 19392 31686
rect 19340 31622 19392 31628
rect 19352 31482 19380 31622
rect 19340 31476 19392 31482
rect 19340 31418 19392 31424
rect 19352 31346 19380 31418
rect 19340 31340 19392 31346
rect 19340 31282 19392 31288
rect 19248 30932 19300 30938
rect 19248 30874 19300 30880
rect 19352 30818 19380 31282
rect 19444 31142 19472 32710
rect 19628 32298 19656 32778
rect 19904 32570 19932 34682
rect 19996 34377 20024 36518
rect 20074 35048 20130 35057
rect 20074 34983 20076 34992
rect 20128 34983 20130 34992
rect 20076 34954 20128 34960
rect 20074 34912 20130 34921
rect 20074 34847 20130 34856
rect 19982 34368 20038 34377
rect 19982 34303 20038 34312
rect 20088 33590 20116 34847
rect 20076 33584 20128 33590
rect 20076 33526 20128 33532
rect 19984 33516 20036 33522
rect 19984 33458 20036 33464
rect 19892 32564 19944 32570
rect 19892 32506 19944 32512
rect 19892 32428 19944 32434
rect 19892 32370 19944 32376
rect 19616 32292 19668 32298
rect 19616 32234 19668 32240
rect 19580 32124 19876 32144
rect 19636 32122 19660 32124
rect 19716 32122 19740 32124
rect 19796 32122 19820 32124
rect 19658 32070 19660 32122
rect 19722 32070 19734 32122
rect 19796 32070 19798 32122
rect 19636 32068 19660 32070
rect 19716 32068 19740 32070
rect 19796 32068 19820 32070
rect 19580 32048 19876 32068
rect 19904 31958 19932 32370
rect 19616 31952 19668 31958
rect 19616 31894 19668 31900
rect 19892 31952 19944 31958
rect 19892 31894 19944 31900
rect 19628 31249 19656 31894
rect 19892 31748 19944 31754
rect 19892 31690 19944 31696
rect 19904 31521 19932 31690
rect 19890 31512 19946 31521
rect 19890 31447 19946 31456
rect 19904 31346 19932 31447
rect 19892 31340 19944 31346
rect 19892 31282 19944 31288
rect 19614 31240 19670 31249
rect 19614 31175 19670 31184
rect 19890 31240 19946 31249
rect 19890 31175 19946 31184
rect 19432 31136 19484 31142
rect 19432 31078 19484 31084
rect 19580 31036 19876 31056
rect 19636 31034 19660 31036
rect 19716 31034 19740 31036
rect 19796 31034 19820 31036
rect 19658 30982 19660 31034
rect 19722 30982 19734 31034
rect 19796 30982 19798 31034
rect 19636 30980 19660 30982
rect 19716 30980 19740 30982
rect 19796 30980 19820 30982
rect 19580 30960 19876 30980
rect 19260 30790 19380 30818
rect 19260 30297 19288 30790
rect 19340 30592 19392 30598
rect 19340 30534 19392 30540
rect 19246 30288 19302 30297
rect 19246 30223 19302 30232
rect 19248 30048 19300 30054
rect 19248 29990 19300 29996
rect 19156 29300 19208 29306
rect 19156 29242 19208 29248
rect 19154 29200 19210 29209
rect 19154 29135 19156 29144
rect 19208 29135 19210 29144
rect 19156 29106 19208 29112
rect 19156 29028 19208 29034
rect 19156 28970 19208 28976
rect 19168 27402 19196 28970
rect 19260 28937 19288 29990
rect 19246 28928 19302 28937
rect 19246 28863 19302 28872
rect 19352 28558 19380 30534
rect 19580 29948 19876 29968
rect 19636 29946 19660 29948
rect 19716 29946 19740 29948
rect 19796 29946 19820 29948
rect 19658 29894 19660 29946
rect 19722 29894 19734 29946
rect 19796 29894 19798 29946
rect 19636 29892 19660 29894
rect 19716 29892 19740 29894
rect 19796 29892 19820 29894
rect 19580 29872 19876 29892
rect 19904 29730 19932 31175
rect 19996 30841 20024 33458
rect 20076 32564 20128 32570
rect 20076 32506 20128 32512
rect 19982 30832 20038 30841
rect 19982 30767 20038 30776
rect 19996 30734 20024 30767
rect 19984 30728 20036 30734
rect 19984 30670 20036 30676
rect 20088 30326 20116 32506
rect 20076 30320 20128 30326
rect 20076 30262 20128 30268
rect 19984 30252 20036 30258
rect 19984 30194 20036 30200
rect 19524 29708 19576 29714
rect 19524 29650 19576 29656
rect 19812 29702 19932 29730
rect 19536 29209 19564 29650
rect 19708 29640 19760 29646
rect 19708 29582 19760 29588
rect 19720 29306 19748 29582
rect 19812 29306 19840 29702
rect 19996 29345 20024 30194
rect 20076 30184 20128 30190
rect 20076 30126 20128 30132
rect 20088 30025 20116 30126
rect 20074 30016 20130 30025
rect 20074 29951 20130 29960
rect 20088 29850 20116 29951
rect 20076 29844 20128 29850
rect 20076 29786 20128 29792
rect 19982 29336 20038 29345
rect 19708 29300 19760 29306
rect 19708 29242 19760 29248
rect 19800 29300 19852 29306
rect 19982 29271 20038 29280
rect 19800 29242 19852 29248
rect 19522 29200 19578 29209
rect 19720 29186 19748 29242
rect 19720 29158 19932 29186
rect 19522 29135 19578 29144
rect 19580 28860 19876 28880
rect 19636 28858 19660 28860
rect 19716 28858 19740 28860
rect 19796 28858 19820 28860
rect 19658 28806 19660 28858
rect 19722 28806 19734 28858
rect 19796 28806 19798 28858
rect 19636 28804 19660 28806
rect 19716 28804 19740 28806
rect 19796 28804 19820 28806
rect 19580 28784 19876 28804
rect 19340 28552 19392 28558
rect 19340 28494 19392 28500
rect 19156 27396 19208 27402
rect 19156 27338 19208 27344
rect 19064 26036 19116 26042
rect 19064 25978 19116 25984
rect 19168 25945 19196 27338
rect 19248 27328 19300 27334
rect 19248 27270 19300 27276
rect 19260 26382 19288 27270
rect 19248 26376 19300 26382
rect 19248 26318 19300 26324
rect 19352 26246 19380 28494
rect 19800 28484 19852 28490
rect 19800 28426 19852 28432
rect 19812 28218 19840 28426
rect 19904 28393 19932 29158
rect 19984 28688 20036 28694
rect 19984 28630 20036 28636
rect 19890 28384 19946 28393
rect 19890 28319 19946 28328
rect 19996 28234 20024 28630
rect 19800 28212 19852 28218
rect 19800 28154 19852 28160
rect 19904 28206 20024 28234
rect 19812 28014 19840 28154
rect 19800 28008 19852 28014
rect 19800 27950 19852 27956
rect 19580 27772 19876 27792
rect 19636 27770 19660 27772
rect 19716 27770 19740 27772
rect 19796 27770 19820 27772
rect 19658 27718 19660 27770
rect 19722 27718 19734 27770
rect 19796 27718 19798 27770
rect 19636 27716 19660 27718
rect 19716 27716 19740 27718
rect 19796 27716 19820 27718
rect 19430 27704 19486 27713
rect 19580 27696 19876 27716
rect 19430 27639 19486 27648
rect 19444 27606 19472 27639
rect 19432 27600 19484 27606
rect 19904 27554 19932 28206
rect 20076 27872 20128 27878
rect 20076 27814 20128 27820
rect 19432 27542 19484 27548
rect 19524 27532 19576 27538
rect 19524 27474 19576 27480
rect 19812 27526 19932 27554
rect 19984 27600 20036 27606
rect 19984 27542 20036 27548
rect 19430 27160 19486 27169
rect 19430 27095 19486 27104
rect 19444 26926 19472 27095
rect 19432 26920 19484 26926
rect 19430 26888 19432 26897
rect 19484 26888 19486 26897
rect 19430 26823 19486 26832
rect 19536 26772 19564 27474
rect 19444 26744 19564 26772
rect 19812 26772 19840 27526
rect 19996 26926 20024 27542
rect 19984 26920 20036 26926
rect 19984 26862 20036 26868
rect 19812 26744 20024 26772
rect 19340 26240 19392 26246
rect 19340 26182 19392 26188
rect 19444 26194 19472 26744
rect 19580 26684 19876 26704
rect 19636 26682 19660 26684
rect 19716 26682 19740 26684
rect 19796 26682 19820 26684
rect 19658 26630 19660 26682
rect 19722 26630 19734 26682
rect 19796 26630 19798 26682
rect 19636 26628 19660 26630
rect 19716 26628 19740 26630
rect 19796 26628 19820 26630
rect 19580 26608 19876 26628
rect 19616 26376 19668 26382
rect 19616 26318 19668 26324
rect 19628 26217 19656 26318
rect 19614 26208 19670 26217
rect 19352 26058 19380 26182
rect 19444 26166 19564 26194
rect 19352 26030 19472 26058
rect 19154 25936 19210 25945
rect 19154 25871 19210 25880
rect 19340 25900 19392 25906
rect 19340 25842 19392 25848
rect 19352 25362 19380 25842
rect 19444 25838 19472 26030
rect 19432 25832 19484 25838
rect 19432 25774 19484 25780
rect 19536 25684 19564 26166
rect 19614 26143 19670 26152
rect 19892 25968 19944 25974
rect 19892 25910 19944 25916
rect 19444 25656 19564 25684
rect 19444 25430 19472 25656
rect 19580 25596 19876 25616
rect 19636 25594 19660 25596
rect 19716 25594 19740 25596
rect 19796 25594 19820 25596
rect 19658 25542 19660 25594
rect 19722 25542 19734 25594
rect 19796 25542 19798 25594
rect 19636 25540 19660 25542
rect 19716 25540 19740 25542
rect 19796 25540 19820 25542
rect 19580 25520 19876 25540
rect 19432 25424 19484 25430
rect 19432 25366 19484 25372
rect 19616 25424 19668 25430
rect 19616 25366 19668 25372
rect 19248 25356 19300 25362
rect 19248 25298 19300 25304
rect 19340 25356 19392 25362
rect 19340 25298 19392 25304
rect 19260 24750 19288 25298
rect 19064 24744 19116 24750
rect 19064 24686 19116 24692
rect 19248 24744 19300 24750
rect 19248 24686 19300 24692
rect 19076 24614 19104 24686
rect 19064 24608 19116 24614
rect 19064 24550 19116 24556
rect 19352 24410 19380 25298
rect 19524 25220 19576 25226
rect 19444 25180 19524 25208
rect 19340 24404 19392 24410
rect 19340 24346 19392 24352
rect 18972 24336 19024 24342
rect 18892 24296 18972 24324
rect 18788 24278 18840 24284
rect 19444 24313 19472 25180
rect 19524 25162 19576 25168
rect 19628 24954 19656 25366
rect 19798 25256 19854 25265
rect 19798 25191 19854 25200
rect 19616 24948 19668 24954
rect 19616 24890 19668 24896
rect 19812 24682 19840 25191
rect 19800 24676 19852 24682
rect 19800 24618 19852 24624
rect 19580 24508 19876 24528
rect 19636 24506 19660 24508
rect 19716 24506 19740 24508
rect 19796 24506 19820 24508
rect 19658 24454 19660 24506
rect 19722 24454 19734 24506
rect 19796 24454 19798 24506
rect 19636 24452 19660 24454
rect 19716 24452 19740 24454
rect 19796 24452 19820 24454
rect 19580 24432 19876 24452
rect 18972 24278 19024 24284
rect 19430 24304 19486 24313
rect 18800 23254 18828 24278
rect 18880 23588 18932 23594
rect 18880 23530 18932 23536
rect 18788 23248 18840 23254
rect 18788 23190 18840 23196
rect 18892 22642 18920 23530
rect 18880 22636 18932 22642
rect 18880 22578 18932 22584
rect 18786 22264 18842 22273
rect 18786 22199 18842 22208
rect 18800 22030 18828 22199
rect 18880 22092 18932 22098
rect 18984 22080 19012 24278
rect 19430 24239 19486 24248
rect 19340 24132 19392 24138
rect 19340 24074 19392 24080
rect 19246 23896 19302 23905
rect 19246 23831 19302 23840
rect 19156 23656 19208 23662
rect 19156 23598 19208 23604
rect 19168 23089 19196 23598
rect 19260 23526 19288 23831
rect 19248 23520 19300 23526
rect 19248 23462 19300 23468
rect 19352 23338 19380 24074
rect 19444 23662 19472 24239
rect 19524 23792 19576 23798
rect 19524 23734 19576 23740
rect 19432 23656 19484 23662
rect 19432 23598 19484 23604
rect 19536 23508 19564 23734
rect 19260 23310 19380 23338
rect 19444 23480 19564 23508
rect 19154 23080 19210 23089
rect 19154 23015 19210 23024
rect 19064 22568 19116 22574
rect 19064 22510 19116 22516
rect 18932 22052 19012 22080
rect 18880 22034 18932 22040
rect 18788 22024 18840 22030
rect 18788 21966 18840 21972
rect 18696 21888 18748 21894
rect 18696 21830 18748 21836
rect 18800 21729 18828 21966
rect 18786 21720 18842 21729
rect 18892 21690 18920 22034
rect 18786 21655 18842 21664
rect 18880 21684 18932 21690
rect 18880 21626 18932 21632
rect 18788 21480 18840 21486
rect 18788 21422 18840 21428
rect 18604 21140 18656 21146
rect 18604 21082 18656 21088
rect 18800 21049 18828 21422
rect 19076 21078 19104 22510
rect 19156 22500 19208 22506
rect 19156 22442 19208 22448
rect 19168 21593 19196 22442
rect 19260 22234 19288 23310
rect 19444 23186 19472 23480
rect 19580 23420 19876 23440
rect 19636 23418 19660 23420
rect 19716 23418 19740 23420
rect 19796 23418 19820 23420
rect 19658 23366 19660 23418
rect 19722 23366 19734 23418
rect 19796 23366 19798 23418
rect 19636 23364 19660 23366
rect 19716 23364 19740 23366
rect 19796 23364 19820 23366
rect 19580 23344 19876 23364
rect 19904 23304 19932 25910
rect 19996 24750 20024 26744
rect 20088 25906 20116 27814
rect 20076 25900 20128 25906
rect 20076 25842 20128 25848
rect 20088 25498 20116 25842
rect 20076 25492 20128 25498
rect 20076 25434 20128 25440
rect 20088 24954 20116 25434
rect 20076 24948 20128 24954
rect 20076 24890 20128 24896
rect 20076 24812 20128 24818
rect 20076 24754 20128 24760
rect 19984 24744 20036 24750
rect 19984 24686 20036 24692
rect 19984 24608 20036 24614
rect 19984 24550 20036 24556
rect 19996 24410 20024 24550
rect 19984 24404 20036 24410
rect 19984 24346 20036 24352
rect 19996 24274 20024 24346
rect 19984 24268 20036 24274
rect 19984 24210 20036 24216
rect 20088 24041 20116 24754
rect 20074 24032 20130 24041
rect 20074 23967 20130 23976
rect 19904 23276 20024 23304
rect 19432 23180 19484 23186
rect 19432 23122 19484 23128
rect 19800 23180 19852 23186
rect 19800 23122 19852 23128
rect 19892 23180 19944 23186
rect 19892 23122 19944 23128
rect 19340 23112 19392 23118
rect 19340 23054 19392 23060
rect 19248 22228 19300 22234
rect 19248 22170 19300 22176
rect 19154 21584 19210 21593
rect 19154 21519 19210 21528
rect 19064 21072 19116 21078
rect 18786 21040 18842 21049
rect 19064 21014 19116 21020
rect 19156 21072 19208 21078
rect 19156 21014 19208 21020
rect 18786 20975 18842 20984
rect 18800 19310 18828 20975
rect 18970 20904 19026 20913
rect 18970 20839 19026 20848
rect 18984 19310 19012 20839
rect 19076 20602 19104 21014
rect 19064 20596 19116 20602
rect 19064 20538 19116 20544
rect 19168 20058 19196 21014
rect 19352 20992 19380 23054
rect 19444 22166 19472 23122
rect 19812 22778 19840 23122
rect 19800 22772 19852 22778
rect 19800 22714 19852 22720
rect 19580 22332 19876 22352
rect 19636 22330 19660 22332
rect 19716 22330 19740 22332
rect 19796 22330 19820 22332
rect 19658 22278 19660 22330
rect 19722 22278 19734 22330
rect 19796 22278 19798 22330
rect 19636 22276 19660 22278
rect 19716 22276 19740 22278
rect 19796 22276 19820 22278
rect 19580 22256 19876 22276
rect 19432 22160 19484 22166
rect 19432 22102 19484 22108
rect 19904 22001 19932 23122
rect 19996 23118 20024 23276
rect 19984 23112 20036 23118
rect 19984 23054 20036 23060
rect 20074 23080 20130 23089
rect 19996 22710 20024 23054
rect 20074 23015 20130 23024
rect 19984 22704 20036 22710
rect 19984 22646 20036 22652
rect 19984 22432 20036 22438
rect 19984 22374 20036 22380
rect 19890 21992 19946 22001
rect 19890 21927 19946 21936
rect 19904 21622 19932 21927
rect 19892 21616 19944 21622
rect 19614 21584 19670 21593
rect 19892 21558 19944 21564
rect 19614 21519 19616 21528
rect 19668 21519 19670 21528
rect 19616 21490 19668 21496
rect 19432 21344 19484 21350
rect 19432 21286 19484 21292
rect 19444 21060 19472 21286
rect 19580 21244 19876 21264
rect 19636 21242 19660 21244
rect 19716 21242 19740 21244
rect 19796 21242 19820 21244
rect 19658 21190 19660 21242
rect 19722 21190 19734 21242
rect 19796 21190 19798 21242
rect 19636 21188 19660 21190
rect 19716 21188 19740 21190
rect 19796 21188 19820 21190
rect 19580 21168 19876 21188
rect 19996 21146 20024 22374
rect 19984 21140 20036 21146
rect 19984 21082 20036 21088
rect 19444 21032 19564 21060
rect 19352 20964 19472 20992
rect 19340 20868 19392 20874
rect 19340 20810 19392 20816
rect 19352 20602 19380 20810
rect 19340 20596 19392 20602
rect 19340 20538 19392 20544
rect 19444 20466 19472 20964
rect 19536 20505 19564 21032
rect 19708 21004 19760 21010
rect 19708 20946 19760 20952
rect 19720 20806 19748 20946
rect 19708 20800 19760 20806
rect 19708 20742 19760 20748
rect 19522 20496 19578 20505
rect 19432 20460 19484 20466
rect 19522 20431 19578 20440
rect 19432 20402 19484 20408
rect 19444 20058 19472 20402
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 19580 20156 19876 20176
rect 19636 20154 19660 20156
rect 19716 20154 19740 20156
rect 19796 20154 19820 20156
rect 19658 20102 19660 20154
rect 19722 20102 19734 20154
rect 19796 20102 19798 20154
rect 19636 20100 19660 20102
rect 19716 20100 19740 20102
rect 19796 20100 19820 20102
rect 19580 20080 19876 20100
rect 19156 20052 19208 20058
rect 19156 19994 19208 20000
rect 19432 20052 19484 20058
rect 19432 19994 19484 20000
rect 19444 19310 19472 19994
rect 19996 19990 20024 20198
rect 19984 19984 20036 19990
rect 19984 19926 20036 19932
rect 20088 19514 20116 23015
rect 20076 19508 20128 19514
rect 20076 19450 20128 19456
rect 18788 19304 18840 19310
rect 18788 19246 18840 19252
rect 18972 19304 19024 19310
rect 19156 19304 19208 19310
rect 18972 19246 19024 19252
rect 19154 19272 19156 19281
rect 19432 19304 19484 19310
rect 19208 19272 19210 19281
rect 18800 18834 18828 19246
rect 18984 19174 19012 19246
rect 19432 19246 19484 19252
rect 19154 19207 19210 19216
rect 18972 19168 19024 19174
rect 18972 19110 19024 19116
rect 18788 18828 18840 18834
rect 18788 18770 18840 18776
rect 18800 18086 18828 18770
rect 18984 18426 19012 19110
rect 19168 18970 19196 19207
rect 19580 19068 19876 19088
rect 19636 19066 19660 19068
rect 19716 19066 19740 19068
rect 19796 19066 19820 19068
rect 19658 19014 19660 19066
rect 19722 19014 19734 19066
rect 19796 19014 19798 19066
rect 19636 19012 19660 19014
rect 19716 19012 19740 19014
rect 19796 19012 19820 19014
rect 19580 18992 19876 19012
rect 19156 18964 19208 18970
rect 19156 18906 19208 18912
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 18972 18420 19024 18426
rect 18972 18362 19024 18368
rect 18788 18080 18840 18086
rect 18788 18022 18840 18028
rect 19248 17876 19300 17882
rect 19352 17864 19380 18770
rect 19580 17980 19876 18000
rect 19636 17978 19660 17980
rect 19716 17978 19740 17980
rect 19796 17978 19820 17980
rect 19658 17926 19660 17978
rect 19722 17926 19734 17978
rect 19796 17926 19798 17978
rect 19636 17924 19660 17926
rect 19716 17924 19740 17926
rect 19796 17924 19820 17926
rect 19580 17904 19876 17924
rect 20074 17912 20130 17921
rect 19300 17836 19380 17864
rect 20074 17847 20130 17856
rect 19248 17818 19300 17824
rect 20088 17746 20116 17847
rect 19156 17740 19208 17746
rect 19156 17682 19208 17688
rect 20076 17740 20128 17746
rect 20076 17682 20128 17688
rect 18604 17604 18656 17610
rect 18604 17546 18656 17552
rect 18616 17338 18644 17546
rect 19168 17338 19196 17682
rect 18604 17332 18656 17338
rect 18604 17274 18656 17280
rect 19156 17332 19208 17338
rect 19156 17274 19208 17280
rect 19580 16892 19876 16912
rect 19636 16890 19660 16892
rect 19716 16890 19740 16892
rect 19796 16890 19820 16892
rect 19658 16838 19660 16890
rect 19722 16838 19734 16890
rect 19796 16838 19798 16890
rect 19636 16836 19660 16838
rect 19716 16836 19740 16838
rect 19796 16836 19820 16838
rect 19580 16816 19876 16836
rect 19154 16552 19210 16561
rect 19154 16487 19210 16496
rect 18604 15088 18656 15094
rect 18604 15030 18656 15036
rect 18616 12170 18644 15030
rect 18972 14884 19024 14890
rect 18972 14826 19024 14832
rect 18984 14618 19012 14826
rect 18972 14612 19024 14618
rect 18972 14554 19024 14560
rect 18970 14512 19026 14521
rect 18970 14447 19026 14456
rect 18604 12164 18656 12170
rect 18604 12106 18656 12112
rect 18616 11558 18644 12106
rect 18880 12096 18932 12102
rect 18880 12038 18932 12044
rect 18604 11552 18656 11558
rect 18604 11494 18656 11500
rect 18616 11218 18644 11494
rect 18604 11212 18656 11218
rect 18604 11154 18656 11160
rect 18604 11076 18656 11082
rect 18604 11018 18656 11024
rect 18616 10742 18644 11018
rect 18604 10736 18656 10742
rect 18604 10678 18656 10684
rect 18892 9081 18920 12038
rect 18510 9072 18566 9081
rect 18510 9007 18566 9016
rect 18878 9072 18934 9081
rect 18878 9007 18934 9016
rect 18984 4842 19012 14447
rect 18892 4814 19012 4842
rect 18234 3360 18290 3369
rect 18234 3295 18290 3304
rect 18248 2514 18276 3295
rect 18236 2508 18288 2514
rect 18236 2450 18288 2456
rect 18892 800 18920 4814
rect 19168 4146 19196 16487
rect 19580 15804 19876 15824
rect 19636 15802 19660 15804
rect 19716 15802 19740 15804
rect 19796 15802 19820 15804
rect 19658 15750 19660 15802
rect 19722 15750 19734 15802
rect 19796 15750 19798 15802
rect 19636 15748 19660 15750
rect 19716 15748 19740 15750
rect 19796 15748 19820 15750
rect 19580 15728 19876 15748
rect 20180 15473 20208 50254
rect 20260 49700 20312 49706
rect 20260 49642 20312 49648
rect 20272 49434 20300 49642
rect 20260 49428 20312 49434
rect 20260 49370 20312 49376
rect 20364 48929 20392 50662
rect 20350 48920 20406 48929
rect 20350 48855 20406 48864
rect 20352 48680 20404 48686
rect 20352 48622 20404 48628
rect 20258 48376 20314 48385
rect 20258 48311 20314 48320
rect 20272 48074 20300 48311
rect 20260 48068 20312 48074
rect 20260 48010 20312 48016
rect 20364 46986 20392 48622
rect 20456 48278 20484 50730
rect 20444 48272 20496 48278
rect 20444 48214 20496 48220
rect 20548 48124 20576 51546
rect 20640 50386 20668 52634
rect 20720 52488 20772 52494
rect 20720 52430 20772 52436
rect 20732 51649 20760 52430
rect 20718 51640 20774 51649
rect 20718 51575 20774 51584
rect 20720 50856 20772 50862
rect 20720 50798 20772 50804
rect 20628 50380 20680 50386
rect 20628 50322 20680 50328
rect 20732 49434 20760 50798
rect 20720 49428 20772 49434
rect 20720 49370 20772 49376
rect 20628 49292 20680 49298
rect 20628 49234 20680 49240
rect 20640 49201 20668 49234
rect 20626 49192 20682 49201
rect 20626 49127 20682 49136
rect 20640 48890 20668 49127
rect 20628 48884 20680 48890
rect 20628 48826 20680 48832
rect 20720 48136 20772 48142
rect 20548 48096 20720 48124
rect 20720 48078 20772 48084
rect 20352 46980 20404 46986
rect 20352 46922 20404 46928
rect 20260 40928 20312 40934
rect 20260 40870 20312 40876
rect 20272 40594 20300 40870
rect 20260 40588 20312 40594
rect 20260 40530 20312 40536
rect 20272 40458 20300 40530
rect 20260 40452 20312 40458
rect 20260 40394 20312 40400
rect 20272 39302 20300 40394
rect 20364 39914 20392 46922
rect 20444 42084 20496 42090
rect 20444 42026 20496 42032
rect 20352 39908 20404 39914
rect 20352 39850 20404 39856
rect 20260 39296 20312 39302
rect 20260 39238 20312 39244
rect 20272 38962 20300 39238
rect 20260 38956 20312 38962
rect 20260 38898 20312 38904
rect 20456 38418 20484 42026
rect 20720 40724 20772 40730
rect 20720 40666 20772 40672
rect 20732 40633 20760 40666
rect 20718 40624 20774 40633
rect 20718 40559 20774 40568
rect 20536 39908 20588 39914
rect 20536 39850 20588 39856
rect 20444 38412 20496 38418
rect 20444 38354 20496 38360
rect 20352 37732 20404 37738
rect 20352 37674 20404 37680
rect 20364 37466 20392 37674
rect 20444 37664 20496 37670
rect 20444 37606 20496 37612
rect 20352 37460 20404 37466
rect 20352 37402 20404 37408
rect 20258 37224 20314 37233
rect 20258 37159 20314 37168
rect 20272 36922 20300 37159
rect 20260 36916 20312 36922
rect 20260 36858 20312 36864
rect 20352 35012 20404 35018
rect 20352 34954 20404 34960
rect 20364 34626 20392 34954
rect 20272 34598 20392 34626
rect 20272 34134 20300 34598
rect 20352 34536 20404 34542
rect 20352 34478 20404 34484
rect 20364 34406 20392 34478
rect 20352 34400 20404 34406
rect 20352 34342 20404 34348
rect 20364 34241 20392 34342
rect 20350 34232 20406 34241
rect 20350 34167 20406 34176
rect 20260 34128 20312 34134
rect 20260 34070 20312 34076
rect 20352 34060 20404 34066
rect 20352 34002 20404 34008
rect 20260 33380 20312 33386
rect 20260 33322 20312 33328
rect 20272 33114 20300 33322
rect 20364 33318 20392 34002
rect 20352 33312 20404 33318
rect 20352 33254 20404 33260
rect 20260 33108 20312 33114
rect 20260 33050 20312 33056
rect 20272 32026 20300 33050
rect 20364 32910 20392 33254
rect 20352 32904 20404 32910
rect 20352 32846 20404 32852
rect 20260 32020 20312 32026
rect 20260 31962 20312 31968
rect 20260 31884 20312 31890
rect 20260 31826 20312 31832
rect 20272 28082 20300 31826
rect 20364 31770 20392 32846
rect 20456 31890 20484 37606
rect 20548 34513 20576 39850
rect 20824 39386 20852 74598
rect 20916 69737 20944 76774
rect 21100 76378 21128 76910
rect 22112 76514 22140 79200
rect 21916 76492 21968 76498
rect 21916 76434 21968 76440
rect 22020 76486 22140 76514
rect 21178 76392 21234 76401
rect 21100 76350 21178 76378
rect 21178 76327 21180 76336
rect 21232 76327 21234 76336
rect 21180 76298 21232 76304
rect 21928 75970 21956 76434
rect 22020 76430 22048 76486
rect 22008 76424 22060 76430
rect 22008 76366 22060 76372
rect 22020 76090 22048 76366
rect 22928 76288 22980 76294
rect 22928 76230 22980 76236
rect 22008 76084 22060 76090
rect 22008 76026 22060 76032
rect 21928 75942 22048 75970
rect 22020 75750 22048 75942
rect 22008 75744 22060 75750
rect 22008 75686 22060 75692
rect 21362 75304 21418 75313
rect 21362 75239 21418 75248
rect 21270 74488 21326 74497
rect 21270 74423 21326 74432
rect 21088 72480 21140 72486
rect 21088 72422 21140 72428
rect 21100 71913 21128 72422
rect 21086 71904 21142 71913
rect 21086 71839 21142 71848
rect 20902 69728 20958 69737
rect 20902 69663 20958 69672
rect 20902 67960 20958 67969
rect 20902 67895 20904 67904
rect 20956 67895 20958 67904
rect 20904 67866 20956 67872
rect 21088 63368 21140 63374
rect 21088 63310 21140 63316
rect 21100 62830 21128 63310
rect 21088 62824 21140 62830
rect 21088 62766 21140 62772
rect 21180 62144 21232 62150
rect 21180 62086 21232 62092
rect 21088 60104 21140 60110
rect 21088 60046 21140 60052
rect 20904 59424 20956 59430
rect 20904 59366 20956 59372
rect 20916 59129 20944 59366
rect 20902 59120 20958 59129
rect 20902 59055 20904 59064
rect 20956 59055 20958 59064
rect 20904 59026 20956 59032
rect 20916 58070 20944 59026
rect 20904 58064 20956 58070
rect 20904 58006 20956 58012
rect 20904 57860 20956 57866
rect 20904 57802 20956 57808
rect 20916 57254 20944 57802
rect 20904 57248 20956 57254
rect 20904 57190 20956 57196
rect 20916 56438 20944 57190
rect 21100 56778 21128 60046
rect 21192 58546 21220 62086
rect 21180 58540 21232 58546
rect 21180 58482 21232 58488
rect 21180 57792 21232 57798
rect 21180 57734 21232 57740
rect 21192 57594 21220 57734
rect 21180 57588 21232 57594
rect 21180 57530 21232 57536
rect 21088 56772 21140 56778
rect 21088 56714 21140 56720
rect 20904 56432 20956 56438
rect 20904 56374 20956 56380
rect 20902 56264 20958 56273
rect 20902 56199 20904 56208
rect 20956 56199 20958 56208
rect 20904 56170 20956 56176
rect 21088 55820 21140 55826
rect 21088 55762 21140 55768
rect 20996 55616 21048 55622
rect 20996 55558 21048 55564
rect 20902 54224 20958 54233
rect 20902 54159 20958 54168
rect 20916 52562 20944 54159
rect 21008 52630 21036 55558
rect 21100 55282 21128 55762
rect 21180 55752 21232 55758
rect 21180 55694 21232 55700
rect 21088 55276 21140 55282
rect 21088 55218 21140 55224
rect 21192 55214 21220 55694
rect 21180 55208 21232 55214
rect 21180 55150 21232 55156
rect 21088 55140 21140 55146
rect 21088 55082 21140 55088
rect 21100 54534 21128 55082
rect 21088 54528 21140 54534
rect 21088 54470 21140 54476
rect 21100 54058 21128 54470
rect 21192 54194 21220 55150
rect 21180 54188 21232 54194
rect 21180 54130 21232 54136
rect 21088 54052 21140 54058
rect 21088 53994 21140 54000
rect 20996 52624 21048 52630
rect 21048 52572 21128 52578
rect 20996 52566 21128 52572
rect 20904 52556 20956 52562
rect 21008 52550 21128 52566
rect 20904 52498 20956 52504
rect 20916 52154 20944 52498
rect 20994 52456 21050 52465
rect 20994 52391 21050 52400
rect 20904 52148 20956 52154
rect 20904 52090 20956 52096
rect 20902 51912 20958 51921
rect 20902 51847 20958 51856
rect 20916 51474 20944 51847
rect 20904 51468 20956 51474
rect 20904 51410 20956 51416
rect 20902 50824 20958 50833
rect 20902 50759 20958 50768
rect 20916 50726 20944 50759
rect 20904 50720 20956 50726
rect 20904 50662 20956 50668
rect 21008 48890 21036 52391
rect 21100 50454 21128 52550
rect 21180 51536 21232 51542
rect 21180 51478 21232 51484
rect 21192 50726 21220 51478
rect 21180 50720 21232 50726
rect 21180 50662 21232 50668
rect 21088 50448 21140 50454
rect 21088 50390 21140 50396
rect 21100 49910 21128 50390
rect 21088 49904 21140 49910
rect 21088 49846 21140 49852
rect 21088 49768 21140 49774
rect 21086 49736 21088 49745
rect 21140 49736 21142 49745
rect 21086 49671 21142 49680
rect 21178 48920 21234 48929
rect 20996 48884 21048 48890
rect 21178 48855 21234 48864
rect 20996 48826 21048 48832
rect 20904 48544 20956 48550
rect 20904 48486 20956 48492
rect 20916 46714 20944 48486
rect 21192 48210 21220 48855
rect 21180 48204 21232 48210
rect 21180 48146 21232 48152
rect 21088 48068 21140 48074
rect 21088 48010 21140 48016
rect 21100 47598 21128 48010
rect 21192 47802 21220 48146
rect 21180 47796 21232 47802
rect 21180 47738 21232 47744
rect 21088 47592 21140 47598
rect 21088 47534 21140 47540
rect 20994 47288 21050 47297
rect 20994 47223 21050 47232
rect 21180 47252 21232 47258
rect 20904 46708 20956 46714
rect 20904 46650 20956 46656
rect 21008 46510 21036 47223
rect 21180 47194 21232 47200
rect 21192 47161 21220 47194
rect 21178 47152 21234 47161
rect 21178 47087 21234 47096
rect 20996 46504 21048 46510
rect 20996 46446 21048 46452
rect 21180 46028 21232 46034
rect 21180 45970 21232 45976
rect 21192 45286 21220 45970
rect 21180 45280 21232 45286
rect 21180 45222 21232 45228
rect 20904 43852 20956 43858
rect 20904 43794 20956 43800
rect 20916 43382 20944 43794
rect 21192 43790 21220 45222
rect 21180 43784 21232 43790
rect 21180 43726 21232 43732
rect 21192 43450 21220 43726
rect 21180 43444 21232 43450
rect 21180 43386 21232 43392
rect 20904 43376 20956 43382
rect 20904 43318 20956 43324
rect 20916 42770 20944 43318
rect 20904 42764 20956 42770
rect 20904 42706 20956 42712
rect 20996 42764 21048 42770
rect 20996 42706 21048 42712
rect 20916 42294 20944 42706
rect 21008 42362 21036 42706
rect 20996 42356 21048 42362
rect 20996 42298 21048 42304
rect 20904 42288 20956 42294
rect 20904 42230 20956 42236
rect 20916 41818 20944 42230
rect 20904 41812 20956 41818
rect 20904 41754 20956 41760
rect 20916 41070 20944 41754
rect 20904 41064 20956 41070
rect 20904 41006 20956 41012
rect 21180 41064 21232 41070
rect 21180 41006 21232 41012
rect 21192 40730 21220 41006
rect 21180 40724 21232 40730
rect 21180 40666 21232 40672
rect 21088 40588 21140 40594
rect 21088 40530 21140 40536
rect 20996 39840 21048 39846
rect 20996 39782 21048 39788
rect 20824 39358 20944 39386
rect 20812 37800 20864 37806
rect 20812 37742 20864 37748
rect 20824 37505 20852 37742
rect 20810 37496 20866 37505
rect 20810 37431 20812 37440
rect 20864 37431 20866 37440
rect 20812 37402 20864 37408
rect 20824 37371 20852 37402
rect 20916 37233 20944 39358
rect 21008 39098 21036 39782
rect 21100 39642 21128 40530
rect 21192 39982 21220 40666
rect 21180 39976 21232 39982
rect 21180 39918 21232 39924
rect 21088 39636 21140 39642
rect 21088 39578 21140 39584
rect 21192 39506 21220 39918
rect 21180 39500 21232 39506
rect 21180 39442 21232 39448
rect 20996 39092 21048 39098
rect 20996 39034 21048 39040
rect 21008 38826 21036 39034
rect 20996 38820 21048 38826
rect 20996 38762 21048 38768
rect 21008 38554 21036 38762
rect 21192 38554 21220 39442
rect 20996 38548 21048 38554
rect 20996 38490 21048 38496
rect 21180 38548 21232 38554
rect 21180 38490 21232 38496
rect 20996 38412 21048 38418
rect 20996 38354 21048 38360
rect 21008 37913 21036 38354
rect 21088 38344 21140 38350
rect 21086 38312 21088 38321
rect 21140 38312 21142 38321
rect 21086 38247 21142 38256
rect 20994 37904 21050 37913
rect 20994 37839 21050 37848
rect 21100 37670 21128 38247
rect 21088 37664 21140 37670
rect 21088 37606 21140 37612
rect 20902 37224 20958 37233
rect 20902 37159 20958 37168
rect 20904 36576 20956 36582
rect 20904 36518 20956 36524
rect 21180 36576 21232 36582
rect 21180 36518 21232 36524
rect 20916 36281 20944 36518
rect 20902 36272 20958 36281
rect 21192 36242 21220 36518
rect 20902 36207 20958 36216
rect 21180 36236 21232 36242
rect 21180 36178 21232 36184
rect 21192 36038 21220 36178
rect 21088 36032 21140 36038
rect 21088 35974 21140 35980
rect 21180 36032 21232 36038
rect 21180 35974 21232 35980
rect 21100 35737 21128 35974
rect 21086 35728 21142 35737
rect 21086 35663 21142 35672
rect 20994 35592 21050 35601
rect 20628 35556 20680 35562
rect 20994 35527 21050 35536
rect 20628 35498 20680 35504
rect 20640 35442 20668 35498
rect 20640 35414 20760 35442
rect 20534 34504 20590 34513
rect 20534 34439 20590 34448
rect 20732 34202 20760 35414
rect 20902 34912 20958 34921
rect 20902 34847 20958 34856
rect 20812 34672 20864 34678
rect 20810 34640 20812 34649
rect 20864 34640 20866 34649
rect 20810 34575 20866 34584
rect 20916 34513 20944 34847
rect 21008 34678 21036 35527
rect 21100 35154 21128 35663
rect 21192 35630 21220 35974
rect 21180 35624 21232 35630
rect 21180 35566 21232 35572
rect 21088 35148 21140 35154
rect 21088 35090 21140 35096
rect 21100 34746 21128 35090
rect 21088 34740 21140 34746
rect 21088 34682 21140 34688
rect 20996 34672 21048 34678
rect 20996 34614 21048 34620
rect 21088 34536 21140 34542
rect 20902 34504 20958 34513
rect 21088 34478 21140 34484
rect 20902 34439 20958 34448
rect 20720 34196 20772 34202
rect 20720 34138 20772 34144
rect 20904 34060 20956 34066
rect 20904 34002 20956 34008
rect 20996 34060 21048 34066
rect 20996 34002 21048 34008
rect 20628 33992 20680 33998
rect 20628 33934 20680 33940
rect 20534 33280 20590 33289
rect 20534 33215 20590 33224
rect 20548 32842 20576 33215
rect 20536 32836 20588 32842
rect 20536 32778 20588 32784
rect 20640 32201 20668 33934
rect 20720 33856 20772 33862
rect 20720 33798 20772 33804
rect 20732 33697 20760 33798
rect 20718 33688 20774 33697
rect 20916 33658 20944 34002
rect 20718 33623 20774 33632
rect 20904 33652 20956 33658
rect 20904 33594 20956 33600
rect 21008 33538 21036 34002
rect 20916 33510 21036 33538
rect 20916 33454 20944 33510
rect 20904 33448 20956 33454
rect 20824 33408 20904 33436
rect 20824 33266 20852 33408
rect 20904 33390 20956 33396
rect 20994 33416 21050 33425
rect 20994 33351 21050 33360
rect 20824 33238 20944 33266
rect 20718 33144 20774 33153
rect 20718 33079 20774 33088
rect 20732 32774 20760 33079
rect 20812 32904 20864 32910
rect 20812 32846 20864 32852
rect 20720 32768 20772 32774
rect 20824 32745 20852 32846
rect 20720 32710 20772 32716
rect 20810 32736 20866 32745
rect 20626 32192 20682 32201
rect 20626 32127 20682 32136
rect 20536 31952 20588 31958
rect 20536 31894 20588 31900
rect 20732 31906 20760 32710
rect 20810 32671 20866 32680
rect 20812 32360 20864 32366
rect 20812 32302 20864 32308
rect 20824 32026 20852 32302
rect 20916 32230 20944 33238
rect 21008 32298 21036 33351
rect 21100 32570 21128 34478
rect 21192 33130 21220 35566
rect 21284 35290 21312 74423
rect 21376 67561 21404 75239
rect 21822 73264 21878 73273
rect 21822 73199 21878 73208
rect 21362 67552 21418 67561
rect 21362 67487 21418 67496
rect 21730 63472 21786 63481
rect 21640 63436 21692 63442
rect 21730 63407 21786 63416
rect 21640 63378 21692 63384
rect 21652 63186 21680 63378
rect 21744 63306 21772 63407
rect 21732 63300 21784 63306
rect 21732 63242 21784 63248
rect 21652 63158 21772 63186
rect 21744 62830 21772 63158
rect 21456 62824 21508 62830
rect 21456 62766 21508 62772
rect 21732 62824 21784 62830
rect 21732 62766 21784 62772
rect 21468 61962 21496 62766
rect 21744 62150 21772 62766
rect 21732 62144 21784 62150
rect 21732 62086 21784 62092
rect 21468 61934 21772 61962
rect 21364 61192 21416 61198
rect 21364 61134 21416 61140
rect 21376 60858 21404 61134
rect 21364 60852 21416 60858
rect 21364 60794 21416 60800
rect 21548 60580 21600 60586
rect 21548 60522 21600 60528
rect 21560 60314 21588 60522
rect 21640 60512 21692 60518
rect 21640 60454 21692 60460
rect 21548 60308 21600 60314
rect 21548 60250 21600 60256
rect 21546 59528 21602 59537
rect 21546 59463 21602 59472
rect 21560 59226 21588 59463
rect 21548 59220 21600 59226
rect 21548 59162 21600 59168
rect 21652 58478 21680 60454
rect 21640 58472 21692 58478
rect 21640 58414 21692 58420
rect 21454 58304 21510 58313
rect 21454 58239 21510 58248
rect 21364 57792 21416 57798
rect 21364 57734 21416 57740
rect 21376 57390 21404 57734
rect 21364 57384 21416 57390
rect 21364 57326 21416 57332
rect 21468 56982 21496 58239
rect 21652 57905 21680 58414
rect 21638 57896 21694 57905
rect 21638 57831 21694 57840
rect 21456 56976 21508 56982
rect 21456 56918 21508 56924
rect 21548 56908 21600 56914
rect 21548 56850 21600 56856
rect 21362 56808 21418 56817
rect 21362 56743 21418 56752
rect 21376 56506 21404 56743
rect 21454 56672 21510 56681
rect 21454 56607 21510 56616
rect 21468 56506 21496 56607
rect 21560 56545 21588 56850
rect 21546 56536 21602 56545
rect 21364 56500 21416 56506
rect 21364 56442 21416 56448
rect 21456 56500 21508 56506
rect 21546 56471 21602 56480
rect 21456 56442 21508 56448
rect 21456 56364 21508 56370
rect 21456 56306 21508 56312
rect 21364 56228 21416 56234
rect 21364 56170 21416 56176
rect 21376 55185 21404 56170
rect 21468 55729 21496 56306
rect 21454 55720 21510 55729
rect 21454 55655 21510 55664
rect 21362 55176 21418 55185
rect 21362 55111 21418 55120
rect 21376 54097 21404 55111
rect 21652 55078 21680 57831
rect 21640 55072 21692 55078
rect 21640 55014 21692 55020
rect 21456 54732 21508 54738
rect 21456 54674 21508 54680
rect 21640 54732 21692 54738
rect 21640 54674 21692 54680
rect 21468 54194 21496 54674
rect 21546 54632 21602 54641
rect 21546 54567 21602 54576
rect 21456 54188 21508 54194
rect 21456 54130 21508 54136
rect 21362 54088 21418 54097
rect 21362 54023 21418 54032
rect 21560 53718 21588 54567
rect 21652 54126 21680 54674
rect 21640 54120 21692 54126
rect 21640 54062 21692 54068
rect 21652 53961 21680 54062
rect 21638 53952 21694 53961
rect 21638 53887 21694 53896
rect 21548 53712 21600 53718
rect 21548 53654 21600 53660
rect 21640 53644 21692 53650
rect 21640 53586 21692 53592
rect 21364 53576 21416 53582
rect 21364 53518 21416 53524
rect 21376 53038 21404 53518
rect 21364 53032 21416 53038
rect 21364 52974 21416 52980
rect 21376 51610 21404 52974
rect 21652 52698 21680 53586
rect 21640 52692 21692 52698
rect 21640 52634 21692 52640
rect 21548 51944 21600 51950
rect 21546 51912 21548 51921
rect 21600 51912 21602 51921
rect 21546 51847 21602 51856
rect 21640 51876 21692 51882
rect 21640 51818 21692 51824
rect 21456 51808 21508 51814
rect 21456 51750 21508 51756
rect 21364 51604 21416 51610
rect 21364 51546 21416 51552
rect 21364 51400 21416 51406
rect 21364 51342 21416 51348
rect 21376 50862 21404 51342
rect 21364 50856 21416 50862
rect 21364 50798 21416 50804
rect 21376 50522 21404 50798
rect 21364 50516 21416 50522
rect 21364 50458 21416 50464
rect 21468 48210 21496 51750
rect 21546 51640 21602 51649
rect 21546 51575 21602 51584
rect 21560 49434 21588 51575
rect 21652 50930 21680 51818
rect 21744 51474 21772 61934
rect 21836 60110 21864 73199
rect 22020 71074 22048 75686
rect 22020 71058 22140 71074
rect 22020 71052 22152 71058
rect 22020 71046 22100 71052
rect 22100 70994 22152 71000
rect 22744 71052 22796 71058
rect 22744 70994 22796 71000
rect 22756 70650 22784 70994
rect 22744 70644 22796 70650
rect 22744 70586 22796 70592
rect 22756 68814 22784 70586
rect 22834 69864 22890 69873
rect 22834 69799 22890 69808
rect 22848 68882 22876 69799
rect 22836 68876 22888 68882
rect 22836 68818 22888 68824
rect 22560 68808 22612 68814
rect 22560 68750 22612 68756
rect 22744 68808 22796 68814
rect 22744 68750 22796 68756
rect 22572 68270 22600 68750
rect 22848 68474 22876 68818
rect 22836 68468 22888 68474
rect 22836 68410 22888 68416
rect 22560 68264 22612 68270
rect 22560 68206 22612 68212
rect 22190 67552 22246 67561
rect 22190 67487 22246 67496
rect 22008 62688 22060 62694
rect 22008 62630 22060 62636
rect 22020 62150 22048 62630
rect 22008 62144 22060 62150
rect 22006 62112 22008 62121
rect 22060 62112 22062 62121
rect 22006 62047 22062 62056
rect 21916 61600 21968 61606
rect 21916 61542 21968 61548
rect 21928 61266 21956 61542
rect 22020 61418 22048 62047
rect 22020 61390 22140 61418
rect 21916 61260 21968 61266
rect 21916 61202 21968 61208
rect 22008 61192 22060 61198
rect 22008 61134 22060 61140
rect 22020 60353 22048 61134
rect 22112 61062 22140 61390
rect 22100 61056 22152 61062
rect 22100 60998 22152 61004
rect 22100 60648 22152 60654
rect 22100 60590 22152 60596
rect 22006 60344 22062 60353
rect 22006 60279 22062 60288
rect 21824 60104 21876 60110
rect 21824 60046 21876 60052
rect 21824 59968 21876 59974
rect 21824 59910 21876 59916
rect 21836 59566 21864 59910
rect 22112 59673 22140 60590
rect 22204 59702 22232 67487
rect 22282 66736 22338 66745
rect 22282 66671 22338 66680
rect 22296 62898 22324 66671
rect 22284 62892 22336 62898
rect 22284 62834 22336 62840
rect 22466 62248 22522 62257
rect 22466 62183 22522 62192
rect 22376 60648 22428 60654
rect 22376 60590 22428 60596
rect 22388 60518 22416 60590
rect 22376 60512 22428 60518
rect 22376 60454 22428 60460
rect 22388 59809 22416 60454
rect 22374 59800 22430 59809
rect 22374 59735 22430 59744
rect 22192 59696 22244 59702
rect 22098 59664 22154 59673
rect 22192 59638 22244 59644
rect 22098 59599 22154 59608
rect 21824 59560 21876 59566
rect 22112 59548 22140 59599
rect 22376 59560 22428 59566
rect 22112 59520 22232 59548
rect 21824 59502 21876 59508
rect 21836 59158 21864 59502
rect 22100 59220 22152 59226
rect 22100 59162 22152 59168
rect 21824 59152 21876 59158
rect 21824 59094 21876 59100
rect 21836 58478 21864 59094
rect 21916 58880 21968 58886
rect 22112 58834 22140 59162
rect 21916 58822 21968 58828
rect 21928 58546 21956 58822
rect 22020 58806 22140 58834
rect 21916 58540 21968 58546
rect 21916 58482 21968 58488
rect 21824 58472 21876 58478
rect 21824 58414 21876 58420
rect 22020 57882 22048 58806
rect 21928 57854 22048 57882
rect 21928 57458 21956 57854
rect 22008 57792 22060 57798
rect 22008 57734 22060 57740
rect 22020 57526 22048 57734
rect 22008 57520 22060 57526
rect 22008 57462 22060 57468
rect 21916 57452 21968 57458
rect 21916 57394 21968 57400
rect 22204 57338 22232 59520
rect 22376 59502 22428 59508
rect 22388 59226 22416 59502
rect 22376 59220 22428 59226
rect 22376 59162 22428 59168
rect 22376 58472 22428 58478
rect 22376 58414 22428 58420
rect 22388 57798 22416 58414
rect 22480 57866 22508 62183
rect 22560 61056 22612 61062
rect 22560 60998 22612 61004
rect 22572 60654 22600 60998
rect 22560 60648 22612 60654
rect 22560 60590 22612 60596
rect 22836 60172 22888 60178
rect 22836 60114 22888 60120
rect 22558 59800 22614 59809
rect 22848 59770 22876 60114
rect 22558 59735 22614 59744
rect 22836 59764 22888 59770
rect 22468 57860 22520 57866
rect 22468 57802 22520 57808
rect 22376 57792 22428 57798
rect 22376 57734 22428 57740
rect 22388 57390 22416 57734
rect 21836 57310 22232 57338
rect 22284 57384 22336 57390
rect 22284 57326 22336 57332
rect 22376 57384 22428 57390
rect 22376 57326 22428 57332
rect 21836 53174 21864 57310
rect 22100 56908 22152 56914
rect 22100 56850 22152 56856
rect 22008 56772 22060 56778
rect 22008 56714 22060 56720
rect 21914 56672 21970 56681
rect 21914 56607 21970 56616
rect 21928 56438 21956 56607
rect 21916 56432 21968 56438
rect 21916 56374 21968 56380
rect 21916 56296 21968 56302
rect 21916 56238 21968 56244
rect 21928 54874 21956 56238
rect 21916 54868 21968 54874
rect 21916 54810 21968 54816
rect 21928 54210 21956 54810
rect 22020 54330 22048 56714
rect 22112 56166 22140 56850
rect 22296 56302 22324 57326
rect 22388 56710 22416 57326
rect 22572 56846 22600 59735
rect 22836 59706 22888 59712
rect 22744 59628 22796 59634
rect 22744 59570 22796 59576
rect 22756 59022 22784 59570
rect 22940 59072 22968 76230
rect 23032 70961 23060 79200
rect 23952 73273 23980 79200
rect 24412 78010 24440 79200
rect 24228 77982 24440 78010
rect 24228 77178 24256 77982
rect 24308 77920 24360 77926
rect 24308 77862 24360 77868
rect 24320 77586 24348 77862
rect 24308 77580 24360 77586
rect 24308 77522 24360 77528
rect 24216 77172 24268 77178
rect 24216 77114 24268 77120
rect 24320 77110 24348 77522
rect 24676 77376 24728 77382
rect 24676 77318 24728 77324
rect 24398 77208 24454 77217
rect 24398 77143 24400 77152
rect 24452 77143 24454 77152
rect 24400 77114 24452 77120
rect 24308 77104 24360 77110
rect 24308 77046 24360 77052
rect 24688 76974 24716 77318
rect 24676 76968 24728 76974
rect 24676 76910 24728 76916
rect 24122 76392 24178 76401
rect 24122 76327 24178 76336
rect 24136 76294 24164 76327
rect 24688 76294 24716 76910
rect 24124 76288 24176 76294
rect 24124 76230 24176 76236
rect 24676 76288 24728 76294
rect 24676 76230 24728 76236
rect 24688 76129 24716 76230
rect 24674 76120 24730 76129
rect 24674 76055 24730 76064
rect 25332 75886 25360 79200
rect 25870 76120 25926 76129
rect 25870 76055 25926 76064
rect 25884 75886 25912 76055
rect 25320 75880 25372 75886
rect 25320 75822 25372 75828
rect 25872 75880 25924 75886
rect 25924 75828 26004 75834
rect 25872 75822 26004 75828
rect 25884 75806 26004 75822
rect 25976 75206 26004 75806
rect 25964 75200 26016 75206
rect 25964 75142 26016 75148
rect 24766 74488 24822 74497
rect 24766 74423 24822 74432
rect 23938 73264 23994 73273
rect 23938 73199 23994 73208
rect 23204 71052 23256 71058
rect 23204 70994 23256 71000
rect 23018 70952 23074 70961
rect 23018 70887 23074 70896
rect 23216 70514 23244 70994
rect 24308 70984 24360 70990
rect 24306 70952 24308 70961
rect 24360 70952 24362 70961
rect 24306 70887 24362 70896
rect 23388 70644 23440 70650
rect 23388 70586 23440 70592
rect 23204 70508 23256 70514
rect 23204 70450 23256 70456
rect 23020 60852 23072 60858
rect 23020 60794 23072 60800
rect 23032 60042 23060 60794
rect 23020 60036 23072 60042
rect 23020 59978 23072 59984
rect 23032 59090 23060 59978
rect 22848 59044 22968 59072
rect 23020 59084 23072 59090
rect 22744 59016 22796 59022
rect 22744 58958 22796 58964
rect 22756 58342 22784 58958
rect 22744 58336 22796 58342
rect 22744 58278 22796 58284
rect 22650 58032 22706 58041
rect 22650 57967 22706 57976
rect 22560 56840 22612 56846
rect 22560 56782 22612 56788
rect 22376 56704 22428 56710
rect 22376 56646 22428 56652
rect 22284 56296 22336 56302
rect 22284 56238 22336 56244
rect 22100 56160 22152 56166
rect 22100 56102 22152 56108
rect 22112 56001 22140 56102
rect 22098 55992 22154 56001
rect 22098 55927 22154 55936
rect 22284 54664 22336 54670
rect 22284 54606 22336 54612
rect 22008 54324 22060 54330
rect 22008 54266 22060 54272
rect 22192 54324 22244 54330
rect 22192 54266 22244 54272
rect 21928 54182 22048 54210
rect 22020 54126 22048 54182
rect 22008 54120 22060 54126
rect 22008 54062 22060 54068
rect 21916 54052 21968 54058
rect 21916 53994 21968 54000
rect 21824 53168 21876 53174
rect 21824 53110 21876 53116
rect 21928 52714 21956 53994
rect 21928 52686 22140 52714
rect 22112 52630 22140 52686
rect 22100 52624 22152 52630
rect 22100 52566 22152 52572
rect 22112 52358 22140 52566
rect 22204 52562 22232 54266
rect 22296 53632 22324 54606
rect 22388 54194 22416 56646
rect 22572 56166 22600 56782
rect 22560 56160 22612 56166
rect 22560 56102 22612 56108
rect 22468 55752 22520 55758
rect 22466 55720 22468 55729
rect 22520 55720 22522 55729
rect 22466 55655 22522 55664
rect 22572 55622 22600 56102
rect 22560 55616 22612 55622
rect 22560 55558 22612 55564
rect 22468 54664 22520 54670
rect 22468 54606 22520 54612
rect 22480 54505 22508 54606
rect 22466 54496 22522 54505
rect 22466 54431 22522 54440
rect 22376 54188 22428 54194
rect 22376 54130 22428 54136
rect 22376 54052 22428 54058
rect 22376 53994 22428 54000
rect 22388 53786 22416 53994
rect 22376 53780 22428 53786
rect 22376 53722 22428 53728
rect 22376 53644 22428 53650
rect 22296 53604 22376 53632
rect 22376 53586 22428 53592
rect 22284 53032 22336 53038
rect 22282 53000 22284 53009
rect 22336 53000 22338 53009
rect 22388 52970 22416 53586
rect 22282 52935 22338 52944
rect 22376 52964 22428 52970
rect 22376 52906 22428 52912
rect 22388 52601 22416 52906
rect 22374 52592 22430 52601
rect 22192 52556 22244 52562
rect 22374 52527 22430 52536
rect 22192 52498 22244 52504
rect 22100 52352 22152 52358
rect 22100 52294 22152 52300
rect 21822 52048 21878 52057
rect 21822 51983 21878 51992
rect 21836 51610 21864 51983
rect 21824 51604 21876 51610
rect 21824 51546 21876 51552
rect 22008 51604 22060 51610
rect 22008 51546 22060 51552
rect 22020 51474 22048 51546
rect 21732 51468 21784 51474
rect 21732 51410 21784 51416
rect 22008 51468 22060 51474
rect 22008 51410 22060 51416
rect 22112 51406 22140 52294
rect 22204 51814 22232 52498
rect 22282 52184 22338 52193
rect 22282 52119 22338 52128
rect 22296 52086 22324 52119
rect 22284 52080 22336 52086
rect 22284 52022 22336 52028
rect 22388 51950 22416 52527
rect 22376 51944 22428 51950
rect 22376 51886 22428 51892
rect 22192 51808 22244 51814
rect 22192 51750 22244 51756
rect 22388 51542 22416 51886
rect 22376 51536 22428 51542
rect 22376 51478 22428 51484
rect 22100 51400 22152 51406
rect 22100 51342 22152 51348
rect 21732 51264 21784 51270
rect 21732 51206 21784 51212
rect 21744 51105 21772 51206
rect 21730 51096 21786 51105
rect 21730 51031 21786 51040
rect 22008 51060 22060 51066
rect 21640 50924 21692 50930
rect 21640 50866 21692 50872
rect 21744 50386 21772 51031
rect 22112 51048 22140 51342
rect 22284 51332 22336 51338
rect 22284 51274 22336 51280
rect 22296 51066 22324 51274
rect 22284 51060 22336 51066
rect 22060 51020 22140 51048
rect 22204 51020 22284 51048
rect 22008 51002 22060 51008
rect 22006 50960 22062 50969
rect 22006 50895 22008 50904
rect 22060 50895 22062 50904
rect 22008 50866 22060 50872
rect 21822 50824 21878 50833
rect 21822 50759 21878 50768
rect 21732 50380 21784 50386
rect 21732 50322 21784 50328
rect 21744 49978 21772 50322
rect 21732 49972 21784 49978
rect 21732 49914 21784 49920
rect 21548 49428 21600 49434
rect 21548 49370 21600 49376
rect 21456 48204 21508 48210
rect 21456 48146 21508 48152
rect 21362 47832 21418 47841
rect 21362 47767 21418 47776
rect 21376 43382 21404 47767
rect 21468 47258 21496 48146
rect 21640 47592 21692 47598
rect 21640 47534 21692 47540
rect 21456 47252 21508 47258
rect 21456 47194 21508 47200
rect 21652 45898 21680 47534
rect 21640 45892 21692 45898
rect 21640 45834 21692 45840
rect 21364 43376 21416 43382
rect 21364 43318 21416 43324
rect 21364 41064 21416 41070
rect 21362 41032 21364 41041
rect 21416 41032 21418 41041
rect 21362 40967 21418 40976
rect 21364 40384 21416 40390
rect 21364 40326 21416 40332
rect 21376 40050 21404 40326
rect 21364 40044 21416 40050
rect 21364 39986 21416 39992
rect 21376 39642 21404 39986
rect 21364 39636 21416 39642
rect 21364 39578 21416 39584
rect 21732 39432 21784 39438
rect 21732 39374 21784 39380
rect 21638 38856 21694 38865
rect 21744 38826 21772 39374
rect 21638 38791 21694 38800
rect 21732 38820 21784 38826
rect 21652 38758 21680 38791
rect 21732 38762 21784 38768
rect 21640 38752 21692 38758
rect 21640 38694 21692 38700
rect 21638 38040 21694 38049
rect 21638 37975 21694 37984
rect 21546 37904 21602 37913
rect 21546 37839 21548 37848
rect 21600 37839 21602 37848
rect 21548 37810 21600 37816
rect 21652 37369 21680 37975
rect 21638 37360 21694 37369
rect 21638 37295 21694 37304
rect 21652 36922 21680 37295
rect 21640 36916 21692 36922
rect 21640 36858 21692 36864
rect 21272 35284 21324 35290
rect 21272 35226 21324 35232
rect 21362 34640 21418 34649
rect 21362 34575 21418 34584
rect 21376 34474 21404 34575
rect 21364 34468 21416 34474
rect 21364 34410 21416 34416
rect 21548 33924 21600 33930
rect 21548 33866 21600 33872
rect 21272 33856 21324 33862
rect 21272 33798 21324 33804
rect 21284 33318 21312 33798
rect 21364 33448 21416 33454
rect 21364 33390 21416 33396
rect 21272 33312 21324 33318
rect 21272 33254 21324 33260
rect 21192 33102 21312 33130
rect 21178 32736 21234 32745
rect 21178 32671 21234 32680
rect 21088 32564 21140 32570
rect 21088 32506 21140 32512
rect 21100 32434 21128 32506
rect 21088 32428 21140 32434
rect 21088 32370 21140 32376
rect 21192 32298 21220 32671
rect 20996 32292 21048 32298
rect 20996 32234 21048 32240
rect 21180 32292 21232 32298
rect 21180 32234 21232 32240
rect 20904 32224 20956 32230
rect 20904 32166 20956 32172
rect 20994 32192 21050 32201
rect 20812 32020 20864 32026
rect 20812 31962 20864 31968
rect 20444 31884 20496 31890
rect 20444 31826 20496 31832
rect 20364 31742 20484 31770
rect 20352 31204 20404 31210
rect 20352 31146 20404 31152
rect 20364 31113 20392 31146
rect 20350 31104 20406 31113
rect 20350 31039 20406 31048
rect 20364 30870 20392 31039
rect 20352 30864 20404 30870
rect 20352 30806 20404 30812
rect 20352 30660 20404 30666
rect 20352 30602 20404 30608
rect 20364 29560 20392 30602
rect 20456 30394 20484 31742
rect 20444 30388 20496 30394
rect 20444 30330 20496 30336
rect 20444 30184 20496 30190
rect 20444 30126 20496 30132
rect 20456 29782 20484 30126
rect 20444 29776 20496 29782
rect 20444 29718 20496 29724
rect 20444 29572 20496 29578
rect 20364 29532 20444 29560
rect 20444 29514 20496 29520
rect 20456 28966 20484 29514
rect 20444 28960 20496 28966
rect 20444 28902 20496 28908
rect 20456 28762 20484 28902
rect 20444 28756 20496 28762
rect 20444 28698 20496 28704
rect 20444 28552 20496 28558
rect 20444 28494 20496 28500
rect 20260 28076 20312 28082
rect 20260 28018 20312 28024
rect 20258 27976 20314 27985
rect 20456 27962 20484 28494
rect 20258 27911 20314 27920
rect 20364 27934 20484 27962
rect 20272 27878 20300 27911
rect 20260 27872 20312 27878
rect 20260 27814 20312 27820
rect 20258 27704 20314 27713
rect 20364 27674 20392 27934
rect 20444 27872 20496 27878
rect 20444 27814 20496 27820
rect 20258 27639 20260 27648
rect 20312 27639 20314 27648
rect 20352 27668 20404 27674
rect 20260 27610 20312 27616
rect 20352 27610 20404 27616
rect 20260 26988 20312 26994
rect 20260 26930 20312 26936
rect 20272 20754 20300 26930
rect 20352 26920 20404 26926
rect 20352 26862 20404 26868
rect 20364 26450 20392 26862
rect 20456 26586 20484 27814
rect 20444 26580 20496 26586
rect 20444 26522 20496 26528
rect 20352 26444 20404 26450
rect 20352 26386 20404 26392
rect 20352 25764 20404 25770
rect 20352 25706 20404 25712
rect 20364 22137 20392 25706
rect 20444 25152 20496 25158
rect 20444 25094 20496 25100
rect 20456 24993 20484 25094
rect 20442 24984 20498 24993
rect 20442 24919 20498 24928
rect 20444 24812 20496 24818
rect 20444 24754 20496 24760
rect 20456 24721 20484 24754
rect 20442 24712 20498 24721
rect 20442 24647 20498 24656
rect 20444 22636 20496 22642
rect 20444 22578 20496 22584
rect 20456 22273 20484 22578
rect 20442 22264 20498 22273
rect 20442 22199 20498 22208
rect 20456 22166 20484 22199
rect 20444 22160 20496 22166
rect 20350 22128 20406 22137
rect 20444 22102 20496 22108
rect 20548 22114 20576 31894
rect 20732 31878 20852 31906
rect 20720 31816 20772 31822
rect 20720 31758 20772 31764
rect 20732 30938 20760 31758
rect 20824 31686 20852 31878
rect 20812 31680 20864 31686
rect 20812 31622 20864 31628
rect 20720 30932 20772 30938
rect 20720 30874 20772 30880
rect 20720 30728 20772 30734
rect 20720 30670 20772 30676
rect 20732 30433 20760 30670
rect 20718 30424 20774 30433
rect 20718 30359 20774 30368
rect 20720 30320 20772 30326
rect 20720 30262 20772 30268
rect 20732 30122 20760 30262
rect 20720 30116 20772 30122
rect 20720 30058 20772 30064
rect 20732 29850 20760 30058
rect 20824 30054 20852 31622
rect 20812 30048 20864 30054
rect 20812 29990 20864 29996
rect 20810 29880 20866 29889
rect 20720 29844 20772 29850
rect 20810 29815 20866 29824
rect 20720 29786 20772 29792
rect 20628 29504 20680 29510
rect 20628 29446 20680 29452
rect 20640 29102 20668 29446
rect 20628 29096 20680 29102
rect 20680 29056 20760 29084
rect 20628 29038 20680 29044
rect 20732 28694 20760 29056
rect 20720 28688 20772 28694
rect 20720 28630 20772 28636
rect 20732 28529 20760 28630
rect 20718 28520 20774 28529
rect 20718 28455 20774 28464
rect 20628 28212 20680 28218
rect 20680 28172 20760 28200
rect 20628 28154 20680 28160
rect 20628 27600 20680 27606
rect 20628 27542 20680 27548
rect 20640 26994 20668 27542
rect 20628 26988 20680 26994
rect 20628 26930 20680 26936
rect 20626 26888 20682 26897
rect 20626 26823 20628 26832
rect 20680 26823 20682 26832
rect 20628 26794 20680 26800
rect 20628 26376 20680 26382
rect 20628 26318 20680 26324
rect 20640 25974 20668 26318
rect 20628 25968 20680 25974
rect 20628 25910 20680 25916
rect 20640 24410 20668 25910
rect 20628 24404 20680 24410
rect 20628 24346 20680 24352
rect 20640 23186 20668 24346
rect 20732 24274 20760 28172
rect 20824 28150 20852 29815
rect 20916 29306 20944 32166
rect 20994 32127 21050 32136
rect 21008 31793 21036 32127
rect 20994 31784 21050 31793
rect 20994 31719 21050 31728
rect 21008 29850 21036 31719
rect 21088 30932 21140 30938
rect 21088 30874 21140 30880
rect 20996 29844 21048 29850
rect 20996 29786 21048 29792
rect 20904 29300 20956 29306
rect 20904 29242 20956 29248
rect 21008 29238 21036 29786
rect 21100 29628 21128 30874
rect 21192 30394 21220 32234
rect 21284 32026 21312 33102
rect 21272 32020 21324 32026
rect 21272 31962 21324 31968
rect 21376 31890 21404 33390
rect 21456 33312 21508 33318
rect 21456 33254 21508 33260
rect 21468 33153 21496 33254
rect 21454 33144 21510 33153
rect 21454 33079 21510 33088
rect 21560 32994 21588 33866
rect 21730 33824 21786 33833
rect 21730 33759 21786 33768
rect 21638 33688 21694 33697
rect 21638 33623 21694 33632
rect 21652 33386 21680 33623
rect 21744 33522 21772 33759
rect 21732 33516 21784 33522
rect 21732 33458 21784 33464
rect 21640 33380 21692 33386
rect 21640 33322 21692 33328
rect 21468 32966 21588 32994
rect 21652 32994 21680 33322
rect 21744 33114 21772 33458
rect 21732 33108 21784 33114
rect 21732 33050 21784 33056
rect 21652 32966 21772 32994
rect 21468 32434 21496 32966
rect 21640 32904 21692 32910
rect 21640 32846 21692 32852
rect 21456 32428 21508 32434
rect 21456 32370 21508 32376
rect 21546 32328 21602 32337
rect 21468 32286 21546 32314
rect 21468 31890 21496 32286
rect 21546 32263 21602 32272
rect 21548 32224 21600 32230
rect 21548 32166 21600 32172
rect 21560 32026 21588 32166
rect 21548 32020 21600 32026
rect 21548 31962 21600 31968
rect 21364 31884 21416 31890
rect 21364 31826 21416 31832
rect 21456 31884 21508 31890
rect 21456 31826 21508 31832
rect 21272 31680 21324 31686
rect 21272 31622 21324 31628
rect 21284 30870 21312 31622
rect 21376 30938 21404 31826
rect 21468 31482 21496 31826
rect 21456 31476 21508 31482
rect 21456 31418 21508 31424
rect 21454 31376 21510 31385
rect 21454 31311 21510 31320
rect 21468 31278 21496 31311
rect 21456 31272 21508 31278
rect 21456 31214 21508 31220
rect 21456 31136 21508 31142
rect 21456 31078 21508 31084
rect 21364 30932 21416 30938
rect 21364 30874 21416 30880
rect 21272 30864 21324 30870
rect 21272 30806 21324 30812
rect 21284 30433 21312 30806
rect 21364 30796 21416 30802
rect 21364 30738 21416 30744
rect 21376 30705 21404 30738
rect 21362 30696 21418 30705
rect 21362 30631 21418 30640
rect 21270 30424 21326 30433
rect 21180 30388 21232 30394
rect 21376 30394 21404 30631
rect 21468 30569 21496 31078
rect 21454 30560 21510 30569
rect 21454 30495 21510 30504
rect 21270 30359 21326 30368
rect 21364 30388 21416 30394
rect 21180 30330 21232 30336
rect 21364 30330 21416 30336
rect 21272 30320 21324 30326
rect 21272 30262 21324 30268
rect 21180 30184 21232 30190
rect 21180 30126 21232 30132
rect 21192 29753 21220 30126
rect 21178 29744 21234 29753
rect 21178 29679 21234 29688
rect 21180 29640 21232 29646
rect 21100 29600 21180 29628
rect 21180 29582 21232 29588
rect 21192 29510 21220 29582
rect 21180 29504 21232 29510
rect 21180 29446 21232 29452
rect 20996 29232 21048 29238
rect 20996 29174 21048 29180
rect 21088 29028 21140 29034
rect 21088 28970 21140 28976
rect 20904 28688 20956 28694
rect 20904 28630 20956 28636
rect 20812 28144 20864 28150
rect 20812 28086 20864 28092
rect 20812 28008 20864 28014
rect 20810 27976 20812 27985
rect 20864 27976 20866 27985
rect 20916 27946 20944 28630
rect 20994 28520 21050 28529
rect 20994 28455 21050 28464
rect 21008 28218 21036 28455
rect 20996 28212 21048 28218
rect 20996 28154 21048 28160
rect 20996 28076 21048 28082
rect 20996 28018 21048 28024
rect 20810 27911 20866 27920
rect 20904 27940 20956 27946
rect 20904 27882 20956 27888
rect 20812 27872 20864 27878
rect 20812 27814 20864 27820
rect 20824 26790 20852 27814
rect 20904 27328 20956 27334
rect 20904 27270 20956 27276
rect 20916 26994 20944 27270
rect 20904 26988 20956 26994
rect 20904 26930 20956 26936
rect 20904 26852 20956 26858
rect 20904 26794 20956 26800
rect 20812 26784 20864 26790
rect 20812 26726 20864 26732
rect 20812 26512 20864 26518
rect 20916 26489 20944 26794
rect 20812 26454 20864 26460
rect 20902 26480 20958 26489
rect 20824 25922 20852 26454
rect 20902 26415 20958 26424
rect 20904 26308 20956 26314
rect 20904 26250 20956 26256
rect 20916 26081 20944 26250
rect 20902 26072 20958 26081
rect 20902 26007 20958 26016
rect 21008 25956 21036 28018
rect 21100 27538 21128 28970
rect 21192 28762 21220 29446
rect 21180 28756 21232 28762
rect 21180 28698 21232 28704
rect 21284 28665 21312 30262
rect 21560 29782 21588 31962
rect 21652 31822 21680 32846
rect 21744 32609 21772 32966
rect 21730 32600 21786 32609
rect 21730 32535 21786 32544
rect 21732 32496 21784 32502
rect 21732 32438 21784 32444
rect 21640 31816 21692 31822
rect 21640 31758 21692 31764
rect 21640 31340 21692 31346
rect 21640 31282 21692 31288
rect 21652 31142 21680 31282
rect 21640 31136 21692 31142
rect 21640 31078 21692 31084
rect 21652 29850 21680 31078
rect 21744 30870 21772 32438
rect 21732 30864 21784 30870
rect 21732 30806 21784 30812
rect 21732 30184 21784 30190
rect 21732 30126 21784 30132
rect 21640 29844 21692 29850
rect 21640 29786 21692 29792
rect 21548 29776 21600 29782
rect 21548 29718 21600 29724
rect 21744 29646 21772 30126
rect 21364 29640 21416 29646
rect 21732 29640 21784 29646
rect 21364 29582 21416 29588
rect 21546 29608 21602 29617
rect 21270 28656 21326 28665
rect 21180 28620 21232 28626
rect 21270 28591 21326 28600
rect 21180 28562 21232 28568
rect 21192 27878 21220 28562
rect 21284 28558 21312 28591
rect 21272 28552 21324 28558
rect 21272 28494 21324 28500
rect 21272 28416 21324 28422
rect 21272 28358 21324 28364
rect 21180 27872 21232 27878
rect 21180 27814 21232 27820
rect 21178 27704 21234 27713
rect 21284 27674 21312 28358
rect 21178 27639 21234 27648
rect 21272 27668 21324 27674
rect 21088 27532 21140 27538
rect 21088 27474 21140 27480
rect 21100 27130 21128 27474
rect 21088 27124 21140 27130
rect 21088 27066 21140 27072
rect 21088 26988 21140 26994
rect 21088 26930 21140 26936
rect 21100 26382 21128 26930
rect 21192 26790 21220 27639
rect 21272 27610 21324 27616
rect 21270 27568 21326 27577
rect 21270 27503 21326 27512
rect 21284 27470 21312 27503
rect 21272 27464 21324 27470
rect 21272 27406 21324 27412
rect 21180 26784 21232 26790
rect 21180 26726 21232 26732
rect 21192 26518 21220 26726
rect 21284 26586 21312 27406
rect 21272 26580 21324 26586
rect 21272 26522 21324 26528
rect 21180 26512 21232 26518
rect 21180 26454 21232 26460
rect 21088 26376 21140 26382
rect 21088 26318 21140 26324
rect 21100 26081 21128 26318
rect 21180 26308 21232 26314
rect 21180 26250 21232 26256
rect 21086 26072 21142 26081
rect 21086 26007 21142 26016
rect 21008 25928 21128 25956
rect 20824 25894 20944 25922
rect 20812 25764 20864 25770
rect 20812 25706 20864 25712
rect 20824 25673 20852 25706
rect 20810 25664 20866 25673
rect 20810 25599 20866 25608
rect 20810 24848 20866 24857
rect 20810 24783 20866 24792
rect 20824 24750 20852 24783
rect 20812 24744 20864 24750
rect 20812 24686 20864 24692
rect 20812 24608 20864 24614
rect 20812 24550 20864 24556
rect 20720 24268 20772 24274
rect 20720 24210 20772 24216
rect 20720 23724 20772 23730
rect 20720 23666 20772 23672
rect 20628 23180 20680 23186
rect 20628 23122 20680 23128
rect 20732 22658 20760 23666
rect 20824 23254 20852 24550
rect 20916 24206 20944 25894
rect 20994 25800 21050 25809
rect 20994 25735 21050 25744
rect 21008 24596 21036 25735
rect 21100 25362 21128 25928
rect 21088 25356 21140 25362
rect 21088 25298 21140 25304
rect 21192 24954 21220 26250
rect 21272 26036 21324 26042
rect 21272 25978 21324 25984
rect 21284 25537 21312 25978
rect 21376 25838 21404 29582
rect 21732 29582 21784 29588
rect 21546 29543 21602 29552
rect 21560 29510 21588 29543
rect 21548 29504 21600 29510
rect 21548 29446 21600 29452
rect 21548 29232 21600 29238
rect 21548 29174 21600 29180
rect 21456 28688 21508 28694
rect 21456 28630 21508 28636
rect 21468 27849 21496 28630
rect 21454 27840 21510 27849
rect 21454 27775 21510 27784
rect 21560 27418 21588 29174
rect 21640 28552 21692 28558
rect 21640 28494 21692 28500
rect 21652 27606 21680 28494
rect 21730 28112 21786 28121
rect 21730 28047 21732 28056
rect 21784 28047 21786 28056
rect 21732 28018 21784 28024
rect 21732 27940 21784 27946
rect 21732 27882 21784 27888
rect 21640 27600 21692 27606
rect 21640 27542 21692 27548
rect 21744 27538 21772 27882
rect 21732 27532 21784 27538
rect 21732 27474 21784 27480
rect 21560 27390 21680 27418
rect 21548 27328 21600 27334
rect 21548 27270 21600 27276
rect 21456 26920 21508 26926
rect 21456 26862 21508 26868
rect 21468 26761 21496 26862
rect 21454 26752 21510 26761
rect 21454 26687 21510 26696
rect 21454 26480 21510 26489
rect 21454 26415 21456 26424
rect 21508 26415 21510 26424
rect 21456 26386 21508 26392
rect 21468 26042 21496 26386
rect 21456 26036 21508 26042
rect 21456 25978 21508 25984
rect 21456 25900 21508 25906
rect 21456 25842 21508 25848
rect 21364 25832 21416 25838
rect 21364 25774 21416 25780
rect 21270 25528 21326 25537
rect 21270 25463 21326 25472
rect 21272 25356 21324 25362
rect 21272 25298 21324 25304
rect 21180 24948 21232 24954
rect 21180 24890 21232 24896
rect 21088 24744 21140 24750
rect 21086 24712 21088 24721
rect 21140 24712 21142 24721
rect 21086 24647 21142 24656
rect 21008 24568 21128 24596
rect 20904 24200 20956 24206
rect 20904 24142 20956 24148
rect 20904 23656 20956 23662
rect 20904 23598 20956 23604
rect 20812 23248 20864 23254
rect 20812 23190 20864 23196
rect 20916 22982 20944 23598
rect 20996 23588 21048 23594
rect 20996 23530 21048 23536
rect 20904 22976 20956 22982
rect 20904 22918 20956 22924
rect 20812 22772 20864 22778
rect 20812 22714 20864 22720
rect 20640 22630 20760 22658
rect 20640 22574 20668 22630
rect 20628 22568 20680 22574
rect 20628 22510 20680 22516
rect 20640 22234 20668 22510
rect 20628 22228 20680 22234
rect 20628 22170 20680 22176
rect 20548 22086 20668 22114
rect 20350 22063 20406 22072
rect 20640 22080 20668 22086
rect 20640 22052 20760 22080
rect 20444 21888 20496 21894
rect 20444 21830 20496 21836
rect 20456 21486 20484 21830
rect 20352 21480 20404 21486
rect 20444 21480 20496 21486
rect 20352 21422 20404 21428
rect 20442 21448 20444 21457
rect 20496 21448 20498 21457
rect 20364 21010 20392 21422
rect 20442 21383 20498 21392
rect 20456 21078 20484 21383
rect 20628 21140 20680 21146
rect 20628 21082 20680 21088
rect 20444 21072 20496 21078
rect 20444 21014 20496 21020
rect 20352 21004 20404 21010
rect 20352 20946 20404 20952
rect 20536 20936 20588 20942
rect 20536 20878 20588 20884
rect 20272 20726 20484 20754
rect 20260 20392 20312 20398
rect 20260 20334 20312 20340
rect 20272 20058 20300 20334
rect 20260 20052 20312 20058
rect 20260 19994 20312 20000
rect 20272 18902 20300 19994
rect 20260 18896 20312 18902
rect 20260 18838 20312 18844
rect 20456 18834 20484 20726
rect 20548 20466 20576 20878
rect 20536 20460 20588 20466
rect 20536 20402 20588 20408
rect 20548 20058 20576 20402
rect 20640 20380 20668 21082
rect 20732 20534 20760 22052
rect 20824 20874 20852 22714
rect 20916 22642 20944 22918
rect 20904 22636 20956 22642
rect 20904 22578 20956 22584
rect 21008 22098 21036 23530
rect 20996 22092 21048 22098
rect 20996 22034 21048 22040
rect 21008 21690 21036 22034
rect 21100 21894 21128 24568
rect 21192 23225 21220 24890
rect 21178 23216 21234 23225
rect 21178 23151 21234 23160
rect 21180 22976 21232 22982
rect 21180 22918 21232 22924
rect 21192 22545 21220 22918
rect 21178 22536 21234 22545
rect 21178 22471 21234 22480
rect 21178 22400 21234 22409
rect 21178 22335 21234 22344
rect 21088 21888 21140 21894
rect 21088 21830 21140 21836
rect 20996 21684 21048 21690
rect 20996 21626 21048 21632
rect 21088 21140 21140 21146
rect 21088 21082 21140 21088
rect 21100 21049 21128 21082
rect 21086 21040 21142 21049
rect 21192 21010 21220 22335
rect 21284 21554 21312 25298
rect 21468 25242 21496 25842
rect 21376 25214 21496 25242
rect 21376 23186 21404 25214
rect 21456 25152 21508 25158
rect 21456 25094 21508 25100
rect 21468 24886 21496 25094
rect 21456 24880 21508 24886
rect 21456 24822 21508 24828
rect 21456 24744 21508 24750
rect 21456 24686 21508 24692
rect 21468 24410 21496 24686
rect 21560 24682 21588 27270
rect 21652 25906 21680 27390
rect 21730 27296 21786 27305
rect 21730 27231 21786 27240
rect 21744 26790 21772 27231
rect 21732 26784 21784 26790
rect 21732 26726 21784 26732
rect 21732 26580 21784 26586
rect 21732 26522 21784 26528
rect 21744 25974 21772 26522
rect 21732 25968 21784 25974
rect 21732 25910 21784 25916
rect 21640 25900 21692 25906
rect 21640 25842 21692 25848
rect 21732 25832 21784 25838
rect 21732 25774 21784 25780
rect 21640 25696 21692 25702
rect 21640 25638 21692 25644
rect 21548 24676 21600 24682
rect 21548 24618 21600 24624
rect 21560 24410 21588 24618
rect 21456 24404 21508 24410
rect 21456 24346 21508 24352
rect 21548 24404 21600 24410
rect 21548 24346 21600 24352
rect 21548 24268 21600 24274
rect 21548 24210 21600 24216
rect 21454 24168 21510 24177
rect 21454 24103 21510 24112
rect 21468 23730 21496 24103
rect 21560 24041 21588 24210
rect 21546 24032 21602 24041
rect 21546 23967 21602 23976
rect 21560 23866 21588 23967
rect 21548 23860 21600 23866
rect 21548 23802 21600 23808
rect 21652 23798 21680 25638
rect 21640 23792 21692 23798
rect 21640 23734 21692 23740
rect 21456 23724 21508 23730
rect 21456 23666 21508 23672
rect 21364 23180 21416 23186
rect 21364 23122 21416 23128
rect 21376 22778 21404 23122
rect 21364 22772 21416 22778
rect 21364 22714 21416 22720
rect 21468 22681 21496 23666
rect 21548 23656 21600 23662
rect 21546 23624 21548 23633
rect 21600 23624 21602 23633
rect 21546 23559 21602 23568
rect 21560 23526 21588 23559
rect 21548 23520 21600 23526
rect 21548 23462 21600 23468
rect 21548 23248 21600 23254
rect 21548 23190 21600 23196
rect 21560 22953 21588 23190
rect 21652 23168 21680 23734
rect 21744 23322 21772 25774
rect 21732 23316 21784 23322
rect 21732 23258 21784 23264
rect 21652 23140 21772 23168
rect 21638 23080 21694 23089
rect 21638 23015 21694 23024
rect 21546 22944 21602 22953
rect 21546 22879 21602 22888
rect 21454 22672 21510 22681
rect 21454 22607 21510 22616
rect 21560 22166 21588 22879
rect 21548 22160 21600 22166
rect 21548 22102 21600 22108
rect 21362 21720 21418 21729
rect 21362 21655 21418 21664
rect 21272 21548 21324 21554
rect 21272 21490 21324 21496
rect 21376 21146 21404 21655
rect 21364 21140 21416 21146
rect 21364 21082 21416 21088
rect 21086 20975 21142 20984
rect 21180 21004 21232 21010
rect 21180 20946 21232 20952
rect 21364 21004 21416 21010
rect 21364 20946 21416 20952
rect 20812 20868 20864 20874
rect 20812 20810 20864 20816
rect 20720 20528 20772 20534
rect 20720 20470 20772 20476
rect 20720 20392 20772 20398
rect 20640 20352 20720 20380
rect 20720 20334 20772 20340
rect 21376 20058 21404 20946
rect 20536 20052 20588 20058
rect 20536 19994 20588 20000
rect 21364 20052 21416 20058
rect 21364 19994 21416 20000
rect 20996 19916 21048 19922
rect 20996 19858 21048 19864
rect 21008 19514 21036 19858
rect 21086 19816 21142 19825
rect 21086 19751 21088 19760
rect 21140 19751 21142 19760
rect 21088 19722 21140 19728
rect 20996 19508 21048 19514
rect 20996 19450 21048 19456
rect 20444 18828 20496 18834
rect 20444 18770 20496 18776
rect 21178 15600 21234 15609
rect 21178 15535 21180 15544
rect 21232 15535 21234 15544
rect 21180 15506 21232 15512
rect 20166 15464 20222 15473
rect 20166 15399 20222 15408
rect 21192 15162 21220 15506
rect 21272 15496 21324 15502
rect 21272 15438 21324 15444
rect 21180 15156 21232 15162
rect 21180 15098 21232 15104
rect 21284 14822 21312 15438
rect 21272 14816 21324 14822
rect 21272 14758 21324 14764
rect 19580 14716 19876 14736
rect 19636 14714 19660 14716
rect 19716 14714 19740 14716
rect 19796 14714 19820 14716
rect 19658 14662 19660 14714
rect 19722 14662 19734 14714
rect 19796 14662 19798 14714
rect 19636 14660 19660 14662
rect 19716 14660 19740 14662
rect 19796 14660 19820 14662
rect 19580 14640 19876 14660
rect 21284 14385 21312 14758
rect 21270 14376 21326 14385
rect 21270 14311 21326 14320
rect 19580 13628 19876 13648
rect 19636 13626 19660 13628
rect 19716 13626 19740 13628
rect 19796 13626 19820 13628
rect 19658 13574 19660 13626
rect 19722 13574 19734 13626
rect 19796 13574 19798 13626
rect 19636 13572 19660 13574
rect 19716 13572 19740 13574
rect 19796 13572 19820 13574
rect 19580 13552 19876 13572
rect 21284 13530 21312 14311
rect 21272 13524 21324 13530
rect 21272 13466 21324 13472
rect 19580 12540 19876 12560
rect 19636 12538 19660 12540
rect 19716 12538 19740 12540
rect 19796 12538 19820 12540
rect 19658 12486 19660 12538
rect 19722 12486 19734 12538
rect 19796 12486 19798 12538
rect 19636 12484 19660 12486
rect 19716 12484 19740 12486
rect 19796 12484 19820 12486
rect 19580 12464 19876 12484
rect 19248 12300 19300 12306
rect 19248 12242 19300 12248
rect 19260 11626 19288 12242
rect 21560 11898 21588 22102
rect 21652 19553 21680 23015
rect 21744 22574 21772 23140
rect 21732 22568 21784 22574
rect 21732 22510 21784 22516
rect 21744 22234 21772 22510
rect 21732 22228 21784 22234
rect 21732 22170 21784 22176
rect 21638 19544 21694 19553
rect 21638 19479 21694 19488
rect 21548 11892 21600 11898
rect 21548 11834 21600 11840
rect 19432 11688 19484 11694
rect 19432 11630 19484 11636
rect 19984 11688 20036 11694
rect 19984 11630 20036 11636
rect 19248 11620 19300 11626
rect 19248 11562 19300 11568
rect 19260 11286 19288 11562
rect 19248 11280 19300 11286
rect 19248 11222 19300 11228
rect 19444 11082 19472 11630
rect 19580 11452 19876 11472
rect 19636 11450 19660 11452
rect 19716 11450 19740 11452
rect 19796 11450 19820 11452
rect 19658 11398 19660 11450
rect 19722 11398 19734 11450
rect 19796 11398 19798 11450
rect 19636 11396 19660 11398
rect 19716 11396 19740 11398
rect 19796 11396 19820 11398
rect 19580 11376 19876 11396
rect 19432 11076 19484 11082
rect 19432 11018 19484 11024
rect 19580 10364 19876 10384
rect 19636 10362 19660 10364
rect 19716 10362 19740 10364
rect 19796 10362 19820 10364
rect 19658 10310 19660 10362
rect 19722 10310 19734 10362
rect 19796 10310 19798 10362
rect 19636 10308 19660 10310
rect 19716 10308 19740 10310
rect 19796 10308 19820 10310
rect 19580 10288 19876 10308
rect 19996 10305 20024 11630
rect 19982 10296 20038 10305
rect 19982 10231 20038 10240
rect 19430 9480 19486 9489
rect 19430 9415 19486 9424
rect 19444 6905 19472 9415
rect 19580 9276 19876 9296
rect 19636 9274 19660 9276
rect 19716 9274 19740 9276
rect 19796 9274 19820 9276
rect 19658 9222 19660 9274
rect 19722 9222 19734 9274
rect 19796 9222 19798 9274
rect 19636 9220 19660 9222
rect 19716 9220 19740 9222
rect 19796 9220 19820 9222
rect 19580 9200 19876 9220
rect 19580 8188 19876 8208
rect 19636 8186 19660 8188
rect 19716 8186 19740 8188
rect 19796 8186 19820 8188
rect 19658 8134 19660 8186
rect 19722 8134 19734 8186
rect 19796 8134 19798 8186
rect 19636 8132 19660 8134
rect 19716 8132 19740 8134
rect 19796 8132 19820 8134
rect 19580 8112 19876 8132
rect 19580 7100 19876 7120
rect 19636 7098 19660 7100
rect 19716 7098 19740 7100
rect 19796 7098 19820 7100
rect 19658 7046 19660 7098
rect 19722 7046 19734 7098
rect 19796 7046 19798 7098
rect 19636 7044 19660 7046
rect 19716 7044 19740 7046
rect 19796 7044 19820 7046
rect 19580 7024 19876 7044
rect 19430 6896 19486 6905
rect 19430 6831 19486 6840
rect 19580 6012 19876 6032
rect 19636 6010 19660 6012
rect 19716 6010 19740 6012
rect 19796 6010 19820 6012
rect 19658 5958 19660 6010
rect 19722 5958 19734 6010
rect 19796 5958 19798 6010
rect 19636 5956 19660 5958
rect 19716 5956 19740 5958
rect 19796 5956 19820 5958
rect 19580 5936 19876 5956
rect 19580 4924 19876 4944
rect 19636 4922 19660 4924
rect 19716 4922 19740 4924
rect 19796 4922 19820 4924
rect 19658 4870 19660 4922
rect 19722 4870 19734 4922
rect 19796 4870 19798 4922
rect 19636 4868 19660 4870
rect 19716 4868 19740 4870
rect 19796 4868 19820 4870
rect 19580 4848 19876 4868
rect 21732 4820 21784 4826
rect 21732 4762 21784 4768
rect 19246 4312 19302 4321
rect 19430 4312 19486 4321
rect 19302 4270 19430 4298
rect 19246 4247 19302 4256
rect 19430 4247 19486 4256
rect 19156 4140 19208 4146
rect 19156 4082 19208 4088
rect 19432 4004 19484 4010
rect 19432 3946 19484 3952
rect 19444 3398 19472 3946
rect 19580 3836 19876 3856
rect 19636 3834 19660 3836
rect 19716 3834 19740 3836
rect 19796 3834 19820 3836
rect 19658 3782 19660 3834
rect 19722 3782 19734 3834
rect 19796 3782 19798 3834
rect 19636 3780 19660 3782
rect 19716 3780 19740 3782
rect 19796 3780 19820 3782
rect 19580 3760 19876 3780
rect 19432 3392 19484 3398
rect 19430 3360 19432 3369
rect 20812 3392 20864 3398
rect 19484 3360 19486 3369
rect 20812 3334 20864 3340
rect 19430 3295 19486 3304
rect 20720 3120 20772 3126
rect 20720 3062 20772 3068
rect 19580 2748 19876 2768
rect 19636 2746 19660 2748
rect 19716 2746 19740 2748
rect 19796 2746 19820 2748
rect 19658 2694 19660 2746
rect 19722 2694 19734 2746
rect 19796 2694 19798 2746
rect 19636 2692 19660 2694
rect 19716 2692 19740 2694
rect 19796 2692 19820 2694
rect 19580 2672 19876 2692
rect 18972 2440 19024 2446
rect 18972 2382 19024 2388
rect 18984 2281 19012 2382
rect 19800 2304 19852 2310
rect 18970 2272 19026 2281
rect 19800 2246 19852 2252
rect 18970 2207 19026 2216
rect 19812 800 19840 2246
rect 20732 800 20760 3062
rect 20824 2990 20852 3334
rect 20812 2984 20864 2990
rect 20812 2926 20864 2932
rect 20824 2650 20852 2926
rect 21744 2666 21772 4762
rect 21836 4146 21864 50759
rect 22008 50720 22060 50726
rect 22008 50662 22060 50668
rect 22020 47666 22048 50662
rect 22204 50368 22232 51020
rect 22284 51002 22336 51008
rect 22112 50340 22232 50368
rect 22284 50380 22336 50386
rect 22112 48754 22140 50340
rect 22284 50322 22336 50328
rect 22192 50244 22244 50250
rect 22192 50186 22244 50192
rect 22204 49774 22232 50186
rect 22192 49768 22244 49774
rect 22192 49710 22244 49716
rect 22296 49706 22324 50322
rect 22284 49700 22336 49706
rect 22284 49642 22336 49648
rect 22192 49632 22244 49638
rect 22192 49574 22244 49580
rect 22204 49337 22232 49574
rect 22190 49328 22246 49337
rect 22296 49298 22324 49642
rect 22190 49263 22246 49272
rect 22284 49292 22336 49298
rect 22284 49234 22336 49240
rect 22100 48748 22152 48754
rect 22100 48690 22152 48696
rect 22296 48550 22324 49234
rect 22388 49162 22416 51478
rect 22480 50182 22508 54431
rect 22560 54120 22612 54126
rect 22560 54062 22612 54068
rect 22572 53242 22600 54062
rect 22560 53236 22612 53242
rect 22560 53178 22612 53184
rect 22560 51944 22612 51950
rect 22560 51886 22612 51892
rect 22572 51542 22600 51886
rect 22560 51536 22612 51542
rect 22560 51478 22612 51484
rect 22664 51388 22692 57967
rect 22756 57934 22784 58278
rect 22848 58177 22876 59044
rect 23020 59026 23072 59032
rect 23032 58682 23060 59026
rect 23020 58676 23072 58682
rect 23020 58618 23072 58624
rect 23032 58410 23060 58618
rect 23020 58404 23072 58410
rect 23020 58346 23072 58352
rect 22834 58168 22890 58177
rect 22834 58103 22890 58112
rect 22744 57928 22796 57934
rect 22744 57870 22796 57876
rect 22836 57928 22888 57934
rect 22836 57870 22888 57876
rect 22756 57390 22784 57870
rect 22744 57384 22796 57390
rect 22744 57326 22796 57332
rect 22848 57050 22876 57870
rect 22836 57044 22888 57050
rect 22836 56986 22888 56992
rect 22848 55962 22876 56986
rect 22928 56908 22980 56914
rect 22928 56850 22980 56856
rect 22836 55956 22888 55962
rect 22836 55898 22888 55904
rect 22848 55418 22876 55898
rect 22940 55826 22968 56850
rect 23018 55992 23074 56001
rect 23018 55927 23074 55936
rect 22928 55820 22980 55826
rect 22928 55762 22980 55768
rect 22836 55412 22888 55418
rect 22836 55354 22888 55360
rect 22836 54800 22888 54806
rect 22836 54742 22888 54748
rect 22744 54732 22796 54738
rect 22744 54674 22796 54680
rect 22756 54641 22784 54674
rect 22742 54632 22798 54641
rect 22742 54567 22798 54576
rect 22848 53990 22876 54742
rect 22836 53984 22888 53990
rect 22836 53926 22888 53932
rect 22848 53632 22876 53926
rect 22940 53786 22968 55762
rect 22928 53780 22980 53786
rect 22928 53722 22980 53728
rect 22848 53604 22968 53632
rect 22940 52902 22968 53604
rect 22928 52896 22980 52902
rect 22928 52838 22980 52844
rect 22836 52420 22888 52426
rect 22836 52362 22888 52368
rect 22572 51360 22692 51388
rect 22468 50176 22520 50182
rect 22468 50118 22520 50124
rect 22376 49156 22428 49162
rect 22376 49098 22428 49104
rect 22480 49065 22508 50118
rect 22572 49978 22600 51360
rect 22652 50380 22704 50386
rect 22652 50322 22704 50328
rect 22560 49972 22612 49978
rect 22560 49914 22612 49920
rect 22560 49428 22612 49434
rect 22560 49370 22612 49376
rect 22466 49056 22522 49065
rect 22466 48991 22522 49000
rect 22376 48748 22428 48754
rect 22376 48690 22428 48696
rect 22284 48544 22336 48550
rect 22284 48486 22336 48492
rect 22388 48278 22416 48690
rect 22572 48686 22600 49370
rect 22664 49298 22692 50322
rect 22652 49292 22704 49298
rect 22652 49234 22704 49240
rect 22560 48680 22612 48686
rect 22560 48622 22612 48628
rect 22560 48544 22612 48550
rect 22560 48486 22612 48492
rect 22376 48272 22428 48278
rect 22374 48240 22376 48249
rect 22428 48240 22430 48249
rect 22572 48210 22600 48486
rect 22664 48346 22692 49234
rect 22744 48680 22796 48686
rect 22742 48648 22744 48657
rect 22796 48648 22798 48657
rect 22742 48583 22798 48592
rect 22652 48340 22704 48346
rect 22652 48282 22704 48288
rect 22374 48175 22430 48184
rect 22560 48204 22612 48210
rect 22560 48146 22612 48152
rect 22008 47660 22060 47666
rect 22008 47602 22060 47608
rect 22572 47258 22600 48146
rect 22744 47796 22796 47802
rect 22744 47738 22796 47744
rect 22560 47252 22612 47258
rect 22560 47194 22612 47200
rect 22100 47116 22152 47122
rect 22100 47058 22152 47064
rect 21914 47016 21970 47025
rect 22112 47002 22140 47058
rect 21914 46951 21916 46960
rect 21968 46951 21970 46960
rect 22020 46974 22140 47002
rect 22192 46980 22244 46986
rect 21916 46922 21968 46928
rect 21928 46510 21956 46922
rect 22020 46714 22048 46974
rect 22192 46922 22244 46928
rect 22008 46708 22060 46714
rect 22008 46650 22060 46656
rect 22204 46646 22232 46922
rect 22756 46918 22784 47738
rect 22284 46912 22336 46918
rect 22744 46912 22796 46918
rect 22284 46854 22336 46860
rect 22466 46880 22522 46889
rect 22192 46640 22244 46646
rect 22192 46582 22244 46588
rect 21916 46504 21968 46510
rect 21916 46446 21968 46452
rect 22100 46504 22152 46510
rect 22100 46446 22152 46452
rect 22112 46170 22140 46446
rect 22100 46164 22152 46170
rect 22100 46106 22152 46112
rect 22296 46034 22324 46854
rect 22744 46854 22796 46860
rect 22466 46815 22522 46824
rect 22480 46578 22508 46815
rect 22468 46572 22520 46578
rect 22468 46514 22520 46520
rect 22376 46164 22428 46170
rect 22376 46106 22428 46112
rect 22284 46028 22336 46034
rect 22284 45970 22336 45976
rect 22388 45898 22416 46106
rect 22744 46028 22796 46034
rect 22744 45970 22796 45976
rect 22376 45892 22428 45898
rect 22376 45834 22428 45840
rect 22388 44742 22416 45834
rect 22468 45348 22520 45354
rect 22468 45290 22520 45296
rect 22480 45082 22508 45290
rect 22756 45286 22784 45970
rect 22744 45280 22796 45286
rect 22744 45222 22796 45228
rect 22756 45082 22784 45222
rect 22468 45076 22520 45082
rect 22468 45018 22520 45024
rect 22744 45076 22796 45082
rect 22744 45018 22796 45024
rect 22376 44736 22428 44742
rect 22376 44678 22428 44684
rect 22388 44198 22416 44678
rect 22376 44192 22428 44198
rect 22376 44134 22428 44140
rect 22008 43648 22060 43654
rect 22008 43590 22060 43596
rect 22020 42770 22048 43590
rect 22008 42764 22060 42770
rect 22008 42706 22060 42712
rect 22388 38808 22416 44134
rect 22468 40928 22520 40934
rect 22468 40870 22520 40876
rect 22480 39302 22508 40870
rect 22468 39296 22520 39302
rect 22468 39238 22520 39244
rect 22480 39098 22508 39238
rect 22468 39092 22520 39098
rect 22468 39034 22520 39040
rect 22468 38820 22520 38826
rect 22388 38780 22468 38808
rect 22468 38762 22520 38768
rect 22282 37224 22338 37233
rect 22282 37159 22338 37168
rect 22296 34592 22324 37159
rect 22374 36136 22430 36145
rect 22374 36071 22430 36080
rect 22204 34564 22324 34592
rect 22100 34400 22152 34406
rect 22098 34368 22100 34377
rect 22152 34368 22154 34377
rect 22098 34303 22154 34312
rect 22100 34128 22152 34134
rect 22100 34070 22152 34076
rect 22008 33652 22060 33658
rect 22008 33594 22060 33600
rect 22020 33425 22048 33594
rect 22006 33416 22062 33425
rect 21928 33374 22006 33402
rect 21928 29170 21956 33374
rect 22006 33351 22062 33360
rect 22008 33312 22060 33318
rect 22008 33254 22060 33260
rect 22020 33046 22048 33254
rect 22008 33040 22060 33046
rect 22008 32982 22060 32988
rect 22112 32910 22140 34070
rect 22100 32904 22152 32910
rect 22100 32846 22152 32852
rect 22100 32564 22152 32570
rect 22100 32506 22152 32512
rect 22008 32428 22060 32434
rect 22008 32370 22060 32376
rect 22020 31346 22048 32370
rect 22008 31340 22060 31346
rect 22008 31282 22060 31288
rect 22020 30734 22048 30765
rect 22008 30728 22060 30734
rect 22006 30696 22008 30705
rect 22060 30696 22062 30705
rect 22006 30631 22062 30640
rect 22020 30326 22048 30631
rect 22008 30320 22060 30326
rect 22008 30262 22060 30268
rect 22112 30025 22140 32506
rect 22204 30258 22232 34564
rect 22388 34490 22416 36071
rect 22296 34462 22416 34490
rect 22296 30802 22324 34462
rect 22480 34354 22508 38762
rect 22742 37768 22798 37777
rect 22742 37703 22798 37712
rect 22650 35864 22706 35873
rect 22650 35799 22706 35808
rect 22560 35556 22612 35562
rect 22560 35498 22612 35504
rect 22572 35154 22600 35498
rect 22664 35290 22692 35799
rect 22652 35284 22704 35290
rect 22652 35226 22704 35232
rect 22560 35148 22612 35154
rect 22560 35090 22612 35096
rect 22572 34746 22600 35090
rect 22652 35080 22704 35086
rect 22652 35022 22704 35028
rect 22560 34740 22612 34746
rect 22560 34682 22612 34688
rect 22560 34536 22612 34542
rect 22560 34478 22612 34484
rect 22388 34326 22508 34354
rect 22284 30796 22336 30802
rect 22284 30738 22336 30744
rect 22192 30252 22244 30258
rect 22192 30194 22244 30200
rect 22192 30116 22244 30122
rect 22192 30058 22244 30064
rect 22098 30016 22154 30025
rect 22098 29951 22154 29960
rect 22008 29708 22060 29714
rect 22008 29650 22060 29656
rect 22100 29708 22152 29714
rect 22100 29650 22152 29656
rect 21916 29164 21968 29170
rect 21916 29106 21968 29112
rect 21928 28762 21956 29106
rect 21916 28756 21968 28762
rect 21916 28698 21968 28704
rect 21928 28558 21956 28698
rect 21916 28552 21968 28558
rect 21916 28494 21968 28500
rect 21928 28218 21956 28494
rect 22020 28490 22048 29650
rect 22112 28966 22140 29650
rect 22100 28960 22152 28966
rect 22100 28902 22152 28908
rect 22100 28688 22152 28694
rect 22100 28630 22152 28636
rect 22112 28529 22140 28630
rect 22098 28520 22154 28529
rect 22008 28484 22060 28490
rect 22098 28455 22154 28464
rect 22008 28426 22060 28432
rect 21916 28212 21968 28218
rect 21916 28154 21968 28160
rect 21916 27872 21968 27878
rect 21916 27814 21968 27820
rect 21928 27674 21956 27814
rect 21916 27668 21968 27674
rect 21916 27610 21968 27616
rect 22020 27554 22048 28426
rect 22204 28234 22232 30058
rect 22296 29850 22324 30738
rect 22284 29844 22336 29850
rect 22284 29786 22336 29792
rect 22282 29064 22338 29073
rect 22282 28999 22338 29008
rect 21928 27526 22048 27554
rect 22112 28206 22232 28234
rect 21928 26586 21956 27526
rect 22008 27464 22060 27470
rect 22112 27452 22140 28206
rect 22192 27940 22244 27946
rect 22192 27882 22244 27888
rect 22204 27577 22232 27882
rect 22190 27568 22246 27577
rect 22190 27503 22246 27512
rect 22296 27470 22324 28999
rect 22284 27464 22336 27470
rect 22112 27424 22232 27452
rect 22008 27406 22060 27412
rect 21916 26580 21968 26586
rect 21916 26522 21968 26528
rect 22020 26518 22048 27406
rect 22100 26784 22152 26790
rect 22100 26726 22152 26732
rect 22008 26512 22060 26518
rect 22008 26454 22060 26460
rect 22112 26450 22140 26726
rect 22100 26444 22152 26450
rect 22100 26386 22152 26392
rect 21916 26376 21968 26382
rect 21916 26318 21968 26324
rect 21928 24206 21956 26318
rect 22100 26308 22152 26314
rect 22100 26250 22152 26256
rect 22008 24676 22060 24682
rect 22008 24618 22060 24624
rect 22020 24449 22048 24618
rect 22006 24440 22062 24449
rect 22006 24375 22062 24384
rect 22008 24336 22060 24342
rect 22008 24278 22060 24284
rect 21916 24200 21968 24206
rect 21916 24142 21968 24148
rect 21916 23588 21968 23594
rect 21916 23530 21968 23536
rect 21928 23186 21956 23530
rect 21916 23180 21968 23186
rect 21916 23122 21968 23128
rect 22020 23089 22048 24278
rect 22006 23080 22062 23089
rect 22006 23015 22062 23024
rect 22008 22704 22060 22710
rect 22006 22672 22008 22681
rect 22060 22672 22062 22681
rect 22006 22607 22062 22616
rect 21916 22024 21968 22030
rect 21916 21966 21968 21972
rect 21928 21865 21956 21966
rect 21914 21856 21970 21865
rect 21914 21791 21970 21800
rect 21928 21690 21956 21791
rect 21916 21684 21968 21690
rect 21916 21626 21968 21632
rect 22112 19938 22140 26250
rect 22204 25401 22232 27424
rect 22284 27406 22336 27412
rect 22284 27328 22336 27334
rect 22284 27270 22336 27276
rect 22296 27169 22324 27270
rect 22282 27160 22338 27169
rect 22282 27095 22338 27104
rect 22284 26852 22336 26858
rect 22284 26794 22336 26800
rect 22190 25392 22246 25401
rect 22190 25327 22246 25336
rect 22192 25288 22244 25294
rect 22192 25230 22244 25236
rect 22204 25129 22232 25230
rect 22190 25120 22246 25129
rect 22190 25055 22246 25064
rect 22204 24274 22232 25055
rect 22296 24818 22324 26794
rect 22284 24812 22336 24818
rect 22284 24754 22336 24760
rect 22192 24268 22244 24274
rect 22192 24210 22244 24216
rect 22192 23520 22244 23526
rect 22192 23462 22244 23468
rect 22204 22982 22232 23462
rect 22192 22976 22244 22982
rect 22192 22918 22244 22924
rect 22192 21344 22244 21350
rect 22192 21286 22244 21292
rect 22204 20641 22232 21286
rect 22190 20632 22246 20641
rect 22190 20567 22246 20576
rect 22020 19922 22140 19938
rect 22008 19916 22140 19922
rect 22060 19910 22140 19916
rect 22008 19858 22060 19864
rect 22100 18080 22152 18086
rect 22100 18022 22152 18028
rect 22008 15496 22060 15502
rect 22008 15438 22060 15444
rect 22020 15314 22048 15438
rect 22112 15314 22140 18022
rect 22190 17912 22246 17921
rect 22190 17847 22246 17856
rect 22020 15286 22140 15314
rect 22100 14272 22152 14278
rect 21928 14220 22100 14226
rect 21928 14214 22152 14220
rect 21928 14198 22140 14214
rect 21928 13394 21956 14198
rect 22006 13968 22062 13977
rect 22006 13903 22062 13912
rect 21916 13388 21968 13394
rect 21916 13330 21968 13336
rect 21928 12986 21956 13330
rect 21916 12980 21968 12986
rect 21916 12922 21968 12928
rect 22020 4826 22048 13903
rect 22098 13560 22154 13569
rect 22098 13495 22154 13504
rect 22112 10033 22140 13495
rect 22098 10024 22154 10033
rect 22098 9959 22154 9968
rect 22008 4820 22060 4826
rect 22008 4762 22060 4768
rect 21824 4140 21876 4146
rect 21824 4082 21876 4088
rect 22204 3074 22232 17847
rect 22388 3194 22416 34326
rect 22468 33856 22520 33862
rect 22468 33798 22520 33804
rect 22480 33561 22508 33798
rect 22466 33552 22522 33561
rect 22466 33487 22522 33496
rect 22468 32904 22520 32910
rect 22468 32846 22520 32852
rect 22480 32298 22508 32846
rect 22572 32774 22600 34478
rect 22664 34474 22692 35022
rect 22652 34468 22704 34474
rect 22652 34410 22704 34416
rect 22652 32836 22704 32842
rect 22652 32778 22704 32784
rect 22560 32768 22612 32774
rect 22560 32710 22612 32716
rect 22560 32360 22612 32366
rect 22664 32348 22692 32778
rect 22612 32320 22692 32348
rect 22560 32302 22612 32308
rect 22468 32292 22520 32298
rect 22468 32234 22520 32240
rect 22468 31884 22520 31890
rect 22468 31826 22520 31832
rect 22480 31142 22508 31826
rect 22468 31136 22520 31142
rect 22468 31078 22520 31084
rect 22572 30954 22600 32302
rect 22652 31204 22704 31210
rect 22652 31146 22704 31152
rect 22480 30926 22600 30954
rect 22480 30598 22508 30926
rect 22560 30660 22612 30666
rect 22560 30602 22612 30608
rect 22468 30592 22520 30598
rect 22468 30534 22520 30540
rect 22572 30433 22600 30602
rect 22558 30424 22614 30433
rect 22558 30359 22560 30368
rect 22612 30359 22614 30368
rect 22560 30330 22612 30336
rect 22572 30299 22600 30330
rect 22560 30048 22612 30054
rect 22558 30016 22560 30025
rect 22612 30016 22614 30025
rect 22558 29951 22614 29960
rect 22468 29504 22520 29510
rect 22468 29446 22520 29452
rect 22480 29102 22508 29446
rect 22664 29170 22692 31146
rect 22652 29164 22704 29170
rect 22652 29106 22704 29112
rect 22468 29096 22520 29102
rect 22466 29064 22468 29073
rect 22520 29064 22522 29073
rect 22466 28999 22522 29008
rect 22652 29028 22704 29034
rect 22652 28970 22704 28976
rect 22468 28756 22520 28762
rect 22468 28698 22520 28704
rect 22480 27878 22508 28698
rect 22560 28552 22612 28558
rect 22560 28494 22612 28500
rect 22468 27872 22520 27878
rect 22468 27814 22520 27820
rect 22572 27674 22600 28494
rect 22560 27668 22612 27674
rect 22560 27610 22612 27616
rect 22468 27328 22520 27334
rect 22468 27270 22520 27276
rect 22480 25922 22508 27270
rect 22572 26586 22600 27610
rect 22560 26580 22612 26586
rect 22560 26522 22612 26528
rect 22558 26344 22614 26353
rect 22558 26279 22614 26288
rect 22572 26042 22600 26279
rect 22560 26036 22612 26042
rect 22560 25978 22612 25984
rect 22480 25894 22600 25922
rect 22468 25832 22520 25838
rect 22468 25774 22520 25780
rect 22480 24410 22508 25774
rect 22572 25362 22600 25894
rect 22560 25356 22612 25362
rect 22560 25298 22612 25304
rect 22468 24404 22520 24410
rect 22468 24346 22520 24352
rect 22468 24268 22520 24274
rect 22468 24210 22520 24216
rect 22560 24268 22612 24274
rect 22560 24210 22612 24216
rect 22480 24070 22508 24210
rect 22468 24064 22520 24070
rect 22468 24006 22520 24012
rect 22480 21894 22508 24006
rect 22572 23866 22600 24210
rect 22560 23860 22612 23866
rect 22560 23802 22612 23808
rect 22468 21888 22520 21894
rect 22468 21830 22520 21836
rect 22480 19961 22508 21830
rect 22664 21418 22692 28970
rect 22756 27538 22784 37703
rect 22848 36825 22876 52362
rect 22940 51785 22968 52838
rect 22926 51776 22982 51785
rect 22926 51711 22982 51720
rect 22940 50454 22968 51711
rect 22928 50448 22980 50454
rect 22928 50390 22980 50396
rect 22928 49972 22980 49978
rect 22928 49914 22980 49920
rect 22940 46510 22968 49914
rect 23032 48754 23060 55927
rect 23112 55820 23164 55826
rect 23112 55762 23164 55768
rect 23124 54670 23152 55762
rect 23112 54664 23164 54670
rect 23112 54606 23164 54612
rect 23110 53408 23166 53417
rect 23110 53343 23166 53352
rect 23124 52698 23152 53343
rect 23112 52692 23164 52698
rect 23112 52634 23164 52640
rect 23124 52154 23152 52634
rect 23112 52148 23164 52154
rect 23112 52090 23164 52096
rect 23112 51400 23164 51406
rect 23112 51342 23164 51348
rect 23020 48748 23072 48754
rect 23020 48690 23072 48696
rect 23018 48512 23074 48521
rect 23018 48447 23074 48456
rect 23032 48278 23060 48447
rect 23020 48272 23072 48278
rect 23020 48214 23072 48220
rect 23020 47184 23072 47190
rect 23020 47126 23072 47132
rect 22928 46504 22980 46510
rect 22928 46446 22980 46452
rect 22940 46102 22968 46446
rect 22928 46096 22980 46102
rect 22928 46038 22980 46044
rect 22928 45960 22980 45966
rect 22928 45902 22980 45908
rect 22940 45626 22968 45902
rect 22928 45620 22980 45626
rect 22928 45562 22980 45568
rect 23032 45082 23060 47126
rect 23020 45076 23072 45082
rect 23020 45018 23072 45024
rect 23124 38729 23152 51342
rect 23110 38720 23166 38729
rect 23110 38655 23166 38664
rect 23112 37256 23164 37262
rect 23112 37198 23164 37204
rect 22834 36816 22890 36825
rect 22834 36751 22890 36760
rect 23124 36582 23152 37198
rect 23112 36576 23164 36582
rect 23112 36518 23164 36524
rect 22836 34944 22888 34950
rect 22836 34886 22888 34892
rect 22848 32042 22876 34886
rect 23020 33992 23072 33998
rect 23020 33934 23072 33940
rect 23032 33386 23060 33934
rect 23020 33380 23072 33386
rect 23020 33322 23072 33328
rect 22928 32972 22980 32978
rect 22928 32914 22980 32920
rect 22940 32230 22968 32914
rect 22928 32224 22980 32230
rect 22926 32192 22928 32201
rect 22980 32192 22982 32201
rect 22926 32127 22982 32136
rect 22926 32056 22982 32065
rect 22848 32014 22926 32042
rect 22926 31991 22982 32000
rect 22836 31952 22888 31958
rect 22834 31920 22836 31929
rect 22888 31920 22890 31929
rect 22834 31855 22890 31864
rect 22940 31736 22968 31991
rect 22848 31708 22968 31736
rect 22848 31210 22876 31708
rect 22926 31648 22982 31657
rect 22926 31583 22982 31592
rect 22836 31204 22888 31210
rect 22836 31146 22888 31152
rect 22940 30938 22968 31583
rect 22928 30932 22980 30938
rect 22928 30874 22980 30880
rect 22836 30796 22888 30802
rect 22836 30738 22888 30744
rect 22848 30122 22876 30738
rect 22836 30116 22888 30122
rect 22836 30058 22888 30064
rect 22928 29504 22980 29510
rect 22928 29446 22980 29452
rect 22834 28384 22890 28393
rect 22834 28319 22890 28328
rect 22744 27532 22796 27538
rect 22744 27474 22796 27480
rect 22744 27328 22796 27334
rect 22744 27270 22796 27276
rect 22756 27033 22784 27270
rect 22742 27024 22798 27033
rect 22742 26959 22798 26968
rect 22756 25498 22784 26959
rect 22848 26382 22876 28319
rect 22940 27946 22968 29446
rect 22928 27940 22980 27946
rect 22928 27882 22980 27888
rect 22928 26512 22980 26518
rect 22928 26454 22980 26460
rect 22836 26376 22888 26382
rect 22834 26344 22836 26353
rect 22888 26344 22890 26353
rect 22834 26279 22890 26288
rect 22836 26240 22888 26246
rect 22836 26182 22888 26188
rect 22848 25809 22876 26182
rect 22940 25974 22968 26454
rect 22928 25968 22980 25974
rect 22928 25910 22980 25916
rect 22834 25800 22890 25809
rect 22834 25735 22890 25744
rect 22848 25702 22876 25735
rect 22836 25696 22888 25702
rect 22836 25638 22888 25644
rect 22744 25492 22796 25498
rect 22744 25434 22796 25440
rect 22848 25430 22876 25638
rect 22836 25424 22888 25430
rect 22836 25366 22888 25372
rect 22926 25392 22982 25401
rect 22926 25327 22982 25336
rect 22834 23624 22890 23633
rect 22834 23559 22890 23568
rect 22744 23180 22796 23186
rect 22744 23122 22796 23128
rect 22756 22778 22784 23122
rect 22848 23089 22876 23559
rect 22940 23118 22968 25327
rect 22928 23112 22980 23118
rect 22834 23080 22890 23089
rect 22928 23054 22980 23060
rect 22834 23015 22836 23024
rect 22888 23015 22890 23024
rect 22836 22986 22888 22992
rect 22744 22772 22796 22778
rect 22744 22714 22796 22720
rect 22940 22273 22968 23054
rect 22926 22264 22982 22273
rect 22926 22199 22982 22208
rect 22652 21412 22704 21418
rect 22652 21354 22704 21360
rect 22466 19952 22522 19961
rect 22466 19887 22522 19896
rect 22742 19136 22798 19145
rect 22742 19071 22798 19080
rect 22756 18834 22784 19071
rect 22744 18828 22796 18834
rect 22744 18770 22796 18776
rect 22468 18760 22520 18766
rect 22468 18702 22520 18708
rect 22480 18086 22508 18702
rect 22756 18426 22784 18770
rect 22744 18420 22796 18426
rect 22744 18362 22796 18368
rect 22468 18080 22520 18086
rect 22468 18022 22520 18028
rect 22650 16416 22706 16425
rect 22650 16351 22706 16360
rect 22468 15360 22520 15366
rect 22468 15302 22520 15308
rect 22480 13841 22508 15302
rect 22466 13832 22522 13841
rect 22466 13767 22522 13776
rect 22664 11257 22692 16351
rect 22650 11248 22706 11257
rect 22650 11183 22706 11192
rect 23032 5137 23060 33322
rect 23112 33312 23164 33318
rect 23110 33280 23112 33289
rect 23164 33280 23166 33289
rect 23110 33215 23166 33224
rect 23112 31884 23164 31890
rect 23112 31826 23164 31832
rect 23124 31482 23152 31826
rect 23112 31476 23164 31482
rect 23112 31418 23164 31424
rect 23124 31249 23152 31418
rect 23110 31240 23166 31249
rect 23110 31175 23166 31184
rect 23112 31136 23164 31142
rect 23112 31078 23164 31084
rect 23124 30870 23152 31078
rect 23112 30864 23164 30870
rect 23112 30806 23164 30812
rect 23112 29708 23164 29714
rect 23112 29650 23164 29656
rect 23124 29345 23152 29650
rect 23110 29336 23166 29345
rect 23110 29271 23112 29280
rect 23164 29271 23166 29280
rect 23112 29242 23164 29248
rect 23124 29211 23152 29242
rect 23110 28792 23166 28801
rect 23110 28727 23112 28736
rect 23164 28727 23166 28736
rect 23112 28698 23164 28704
rect 23112 28620 23164 28626
rect 23112 28562 23164 28568
rect 23124 28150 23152 28562
rect 23112 28144 23164 28150
rect 23110 28112 23112 28121
rect 23164 28112 23166 28121
rect 23110 28047 23166 28056
rect 23112 28008 23164 28014
rect 23112 27950 23164 27956
rect 23124 24410 23152 27950
rect 23112 24404 23164 24410
rect 23112 24346 23164 24352
rect 23112 22704 23164 22710
rect 23112 22646 23164 22652
rect 23124 22574 23152 22646
rect 23112 22568 23164 22574
rect 23110 22536 23112 22545
rect 23164 22536 23166 22545
rect 23110 22471 23166 22480
rect 23112 22024 23164 22030
rect 23112 21966 23164 21972
rect 23124 21418 23152 21966
rect 23112 21412 23164 21418
rect 23112 21354 23164 21360
rect 23112 14272 23164 14278
rect 23216 14249 23244 70450
rect 23400 69850 23428 70586
rect 24214 70000 24270 70009
rect 24214 69935 24270 69944
rect 24228 69902 24256 69935
rect 23480 69896 23532 69902
rect 23400 69844 23480 69850
rect 23400 69838 23532 69844
rect 23940 69896 23992 69902
rect 23940 69838 23992 69844
rect 24216 69896 24268 69902
rect 24216 69838 24268 69844
rect 23400 69822 23520 69838
rect 23952 69562 23980 69838
rect 23940 69556 23992 69562
rect 23940 69498 23992 69504
rect 24228 69494 24256 69838
rect 24676 69760 24728 69766
rect 24676 69702 24728 69708
rect 24216 69488 24268 69494
rect 24216 69430 24268 69436
rect 23940 68672 23992 68678
rect 23940 68614 23992 68620
rect 24032 68672 24084 68678
rect 24032 68614 24084 68620
rect 23386 61432 23442 61441
rect 23386 61367 23442 61376
rect 23296 59424 23348 59430
rect 23296 59366 23348 59372
rect 23308 59090 23336 59366
rect 23400 59106 23428 61367
rect 23846 60344 23902 60353
rect 23846 60279 23902 60288
rect 23860 59974 23888 60279
rect 23848 59968 23900 59974
rect 23848 59910 23900 59916
rect 23296 59084 23348 59090
rect 23400 59078 23520 59106
rect 23860 59090 23888 59910
rect 23952 59401 23980 68614
rect 24044 68270 24072 68614
rect 24688 68338 24716 69702
rect 24676 68332 24728 68338
rect 24676 68274 24728 68280
rect 24032 68264 24084 68270
rect 24032 68206 24084 68212
rect 24306 68232 24362 68241
rect 24044 67658 24072 68206
rect 24306 68167 24362 68176
rect 24032 67652 24084 67658
rect 24032 67594 24084 67600
rect 24320 60722 24348 68167
rect 24492 67652 24544 67658
rect 24492 67594 24544 67600
rect 24308 60716 24360 60722
rect 24308 60658 24360 60664
rect 24504 60314 24532 67594
rect 24492 60308 24544 60314
rect 24492 60250 24544 60256
rect 24308 59968 24360 59974
rect 24308 59910 24360 59916
rect 24216 59560 24268 59566
rect 24216 59502 24268 59508
rect 24320 59514 24348 59910
rect 24400 59628 24452 59634
rect 24504 59616 24532 60250
rect 24452 59588 24532 59616
rect 24400 59570 24452 59576
rect 23938 59392 23994 59401
rect 23938 59327 23994 59336
rect 23296 59026 23348 59032
rect 23386 58984 23442 58993
rect 23386 58919 23388 58928
rect 23440 58919 23442 58928
rect 23388 58890 23440 58896
rect 23492 58834 23520 59078
rect 23848 59084 23900 59090
rect 23848 59026 23900 59032
rect 24228 58886 24256 59502
rect 24320 59486 24532 59514
rect 24504 59158 24532 59486
rect 24492 59152 24544 59158
rect 24492 59094 24544 59100
rect 24308 59084 24360 59090
rect 24308 59026 24360 59032
rect 23400 58806 23520 58834
rect 24216 58880 24268 58886
rect 24216 58822 24268 58828
rect 23296 57996 23348 58002
rect 23296 57938 23348 57944
rect 23308 57254 23336 57938
rect 23296 57248 23348 57254
rect 23296 57190 23348 57196
rect 23308 56914 23336 57190
rect 23296 56908 23348 56914
rect 23296 56850 23348 56856
rect 23308 56506 23336 56850
rect 23296 56500 23348 56506
rect 23296 56442 23348 56448
rect 23296 55616 23348 55622
rect 23296 55558 23348 55564
rect 23308 53582 23336 55558
rect 23296 53576 23348 53582
rect 23296 53518 23348 53524
rect 23296 53440 23348 53446
rect 23296 53382 23348 53388
rect 23308 52154 23336 53382
rect 23296 52148 23348 52154
rect 23296 52090 23348 52096
rect 23296 51876 23348 51882
rect 23296 51818 23348 51824
rect 23308 51649 23336 51818
rect 23294 51640 23350 51649
rect 23294 51575 23296 51584
rect 23348 51575 23350 51584
rect 23296 51546 23348 51552
rect 23400 51490 23428 58806
rect 24124 58608 24176 58614
rect 24124 58550 24176 58556
rect 24032 57996 24084 58002
rect 24032 57938 24084 57944
rect 23480 57792 23532 57798
rect 23480 57734 23532 57740
rect 23492 56914 23520 57734
rect 23572 57384 23624 57390
rect 23572 57326 23624 57332
rect 23480 56908 23532 56914
rect 23480 56850 23532 56856
rect 23492 56166 23520 56850
rect 23480 56160 23532 56166
rect 23480 56102 23532 56108
rect 23584 56114 23612 57326
rect 23662 56400 23718 56409
rect 23662 56335 23718 56344
rect 23676 56302 23704 56335
rect 23664 56296 23716 56302
rect 23664 56238 23716 56244
rect 23848 56160 23900 56166
rect 23492 55978 23520 56102
rect 23584 56086 23704 56114
rect 23848 56102 23900 56108
rect 23492 55950 23612 55978
rect 23478 53952 23534 53961
rect 23478 53887 23534 53896
rect 23492 53242 23520 53887
rect 23584 53718 23612 55950
rect 23676 55622 23704 56086
rect 23664 55616 23716 55622
rect 23664 55558 23716 55564
rect 23676 55214 23704 55558
rect 23860 55214 23888 56102
rect 23940 55820 23992 55826
rect 23940 55762 23992 55768
rect 23664 55208 23716 55214
rect 23664 55150 23716 55156
rect 23848 55208 23900 55214
rect 23848 55150 23900 55156
rect 23572 53712 23624 53718
rect 23572 53654 23624 53660
rect 23676 53417 23704 55150
rect 23860 54874 23888 55150
rect 23952 55078 23980 55762
rect 23940 55072 23992 55078
rect 23940 55014 23992 55020
rect 23952 54874 23980 55014
rect 23848 54868 23900 54874
rect 23848 54810 23900 54816
rect 23940 54868 23992 54874
rect 23940 54810 23992 54816
rect 23860 54330 23888 54810
rect 23952 54738 23980 54810
rect 23940 54732 23992 54738
rect 23940 54674 23992 54680
rect 23848 54324 23900 54330
rect 23848 54266 23900 54272
rect 23860 53650 23888 54266
rect 23952 54262 23980 54674
rect 23940 54256 23992 54262
rect 23940 54198 23992 54204
rect 23848 53644 23900 53650
rect 23848 53586 23900 53592
rect 23754 53544 23810 53553
rect 23754 53479 23810 53488
rect 23848 53508 23900 53514
rect 23662 53408 23718 53417
rect 23662 53343 23718 53352
rect 23480 53236 23532 53242
rect 23480 53178 23532 53184
rect 23768 53174 23796 53479
rect 23848 53450 23900 53456
rect 23756 53168 23808 53174
rect 23756 53110 23808 53116
rect 23768 52698 23796 53110
rect 23756 52692 23808 52698
rect 23756 52634 23808 52640
rect 23480 51944 23532 51950
rect 23480 51886 23532 51892
rect 23308 51462 23428 51490
rect 23308 37262 23336 51462
rect 23388 51060 23440 51066
rect 23492 51048 23520 51886
rect 23440 51020 23520 51048
rect 23388 51002 23440 51008
rect 23860 50318 23888 53450
rect 23952 53174 23980 54198
rect 23940 53168 23992 53174
rect 23940 53110 23992 53116
rect 23952 52902 23980 52933
rect 23940 52896 23992 52902
rect 23938 52864 23940 52873
rect 23992 52864 23994 52873
rect 23938 52799 23994 52808
rect 23952 52698 23980 52799
rect 23940 52692 23992 52698
rect 23940 52634 23992 52640
rect 23952 52086 23980 52634
rect 23940 52080 23992 52086
rect 23940 52022 23992 52028
rect 23952 51474 23980 52022
rect 23940 51468 23992 51474
rect 23940 51410 23992 51416
rect 23952 50522 23980 51410
rect 23940 50516 23992 50522
rect 23940 50458 23992 50464
rect 23664 50312 23716 50318
rect 23664 50254 23716 50260
rect 23848 50312 23900 50318
rect 23848 50254 23900 50260
rect 23480 49836 23532 49842
rect 23480 49778 23532 49784
rect 23388 49768 23440 49774
rect 23388 49710 23440 49716
rect 23400 48142 23428 49710
rect 23388 48136 23440 48142
rect 23388 48078 23440 48084
rect 23400 47802 23428 48078
rect 23388 47796 23440 47802
rect 23388 47738 23440 47744
rect 23388 47592 23440 47598
rect 23492 47580 23520 49778
rect 23572 49292 23624 49298
rect 23572 49234 23624 49240
rect 23584 48822 23612 49234
rect 23572 48816 23624 48822
rect 23676 48793 23704 50254
rect 23756 49632 23808 49638
rect 23756 49574 23808 49580
rect 23572 48758 23624 48764
rect 23662 48784 23718 48793
rect 23662 48719 23718 48728
rect 23572 48272 23624 48278
rect 23572 48214 23624 48220
rect 23440 47552 23520 47580
rect 23388 47534 23440 47540
rect 23584 47530 23612 48214
rect 23664 48068 23716 48074
rect 23768 48056 23796 49574
rect 23860 49094 23888 50254
rect 23940 49904 23992 49910
rect 23940 49846 23992 49852
rect 23952 49774 23980 49846
rect 23940 49768 23992 49774
rect 23940 49710 23992 49716
rect 23848 49088 23900 49094
rect 23848 49030 23900 49036
rect 23848 48204 23900 48210
rect 23848 48146 23900 48152
rect 23716 48028 23796 48056
rect 23664 48010 23716 48016
rect 23664 47660 23716 47666
rect 23664 47602 23716 47608
rect 23572 47524 23624 47530
rect 23572 47466 23624 47472
rect 23570 47152 23626 47161
rect 23570 47087 23626 47096
rect 23584 46986 23612 47087
rect 23676 47054 23704 47602
rect 23768 47258 23796 48028
rect 23756 47252 23808 47258
rect 23756 47194 23808 47200
rect 23860 47190 23888 48146
rect 23952 47734 23980 49710
rect 24044 49434 24072 57938
rect 24136 57594 24164 58550
rect 24216 58472 24268 58478
rect 24320 58460 24348 59026
rect 24504 58478 24532 59094
rect 24584 58880 24636 58886
rect 24584 58822 24636 58828
rect 24268 58432 24348 58460
rect 24492 58472 24544 58478
rect 24216 58414 24268 58420
rect 24492 58414 24544 58420
rect 24228 57798 24256 58414
rect 24504 58313 24532 58414
rect 24490 58304 24546 58313
rect 24490 58239 24546 58248
rect 24504 58138 24532 58239
rect 24492 58132 24544 58138
rect 24492 58074 24544 58080
rect 24306 57896 24362 57905
rect 24306 57831 24308 57840
rect 24360 57831 24362 57840
rect 24308 57802 24360 57808
rect 24216 57792 24268 57798
rect 24216 57734 24268 57740
rect 24124 57588 24176 57594
rect 24124 57530 24176 57536
rect 24136 57390 24164 57530
rect 24124 57384 24176 57390
rect 24124 57326 24176 57332
rect 24308 57248 24360 57254
rect 24308 57190 24360 57196
rect 24216 55344 24268 55350
rect 24216 55286 24268 55292
rect 24124 53644 24176 53650
rect 24124 53586 24176 53592
rect 24136 53553 24164 53586
rect 24122 53544 24178 53553
rect 24122 53479 24178 53488
rect 24124 52012 24176 52018
rect 24124 51954 24176 51960
rect 24136 50386 24164 51954
rect 24228 50561 24256 55286
rect 24320 54806 24348 57190
rect 24400 56840 24452 56846
rect 24398 56808 24400 56817
rect 24452 56808 24454 56817
rect 24398 56743 24454 56752
rect 24492 56160 24544 56166
rect 24490 56128 24492 56137
rect 24544 56128 24546 56137
rect 24490 56063 24546 56072
rect 24492 55956 24544 55962
rect 24492 55898 24544 55904
rect 24504 55214 24532 55898
rect 24492 55208 24544 55214
rect 24492 55150 24544 55156
rect 24308 54800 24360 54806
rect 24308 54742 24360 54748
rect 24320 54330 24348 54742
rect 24492 54528 24544 54534
rect 24492 54470 24544 54476
rect 24308 54324 24360 54330
rect 24308 54266 24360 54272
rect 24504 54233 24532 54470
rect 24490 54224 24546 54233
rect 24490 54159 24546 54168
rect 24492 54052 24544 54058
rect 24492 53994 24544 54000
rect 24504 53961 24532 53994
rect 24490 53952 24546 53961
rect 24490 53887 24546 53896
rect 24492 53644 24544 53650
rect 24492 53586 24544 53592
rect 24400 53508 24452 53514
rect 24400 53450 24452 53456
rect 24308 51468 24360 51474
rect 24308 51410 24360 51416
rect 24320 51066 24348 51410
rect 24308 51060 24360 51066
rect 24308 51002 24360 51008
rect 24308 50720 24360 50726
rect 24308 50662 24360 50668
rect 24214 50552 24270 50561
rect 24214 50487 24270 50496
rect 24124 50380 24176 50386
rect 24124 50322 24176 50328
rect 24136 49978 24164 50322
rect 24124 49972 24176 49978
rect 24124 49914 24176 49920
rect 24320 49910 24348 50662
rect 24308 49904 24360 49910
rect 24308 49846 24360 49852
rect 24032 49428 24084 49434
rect 24032 49370 24084 49376
rect 24032 49292 24084 49298
rect 24032 49234 24084 49240
rect 24044 49065 24072 49234
rect 24030 49056 24086 49065
rect 24030 48991 24086 49000
rect 24214 48920 24270 48929
rect 24214 48855 24270 48864
rect 24124 48544 24176 48550
rect 24124 48486 24176 48492
rect 24136 48278 24164 48486
rect 24124 48272 24176 48278
rect 24124 48214 24176 48220
rect 24032 48000 24084 48006
rect 24032 47942 24084 47948
rect 23940 47728 23992 47734
rect 23940 47670 23992 47676
rect 24044 47598 24072 47942
rect 24032 47592 24084 47598
rect 23952 47552 24032 47580
rect 23848 47184 23900 47190
rect 23848 47126 23900 47132
rect 23664 47048 23716 47054
rect 23664 46990 23716 46996
rect 23754 47016 23810 47025
rect 23572 46980 23624 46986
rect 23572 46922 23624 46928
rect 23676 46170 23704 46990
rect 23754 46951 23810 46960
rect 23664 46164 23716 46170
rect 23664 46106 23716 46112
rect 23388 45892 23440 45898
rect 23388 45834 23440 45840
rect 23400 45626 23428 45834
rect 23480 45824 23532 45830
rect 23480 45766 23532 45772
rect 23388 45620 23440 45626
rect 23388 45562 23440 45568
rect 23492 45558 23520 45766
rect 23480 45552 23532 45558
rect 23480 45494 23532 45500
rect 23768 45082 23796 46951
rect 23952 45665 23980 47552
rect 24032 47534 24084 47540
rect 24044 47469 24072 47534
rect 24136 47258 24164 48214
rect 24228 47297 24256 48855
rect 24308 48136 24360 48142
rect 24308 48078 24360 48084
rect 24214 47288 24270 47297
rect 24124 47252 24176 47258
rect 24214 47223 24270 47232
rect 24124 47194 24176 47200
rect 24228 47190 24256 47223
rect 24216 47184 24268 47190
rect 24216 47126 24268 47132
rect 24320 47054 24348 48078
rect 24308 47048 24360 47054
rect 24308 46990 24360 46996
rect 24032 46912 24084 46918
rect 24032 46854 24084 46860
rect 24044 46510 24072 46854
rect 24032 46504 24084 46510
rect 24032 46446 24084 46452
rect 24032 45960 24084 45966
rect 24032 45902 24084 45908
rect 23938 45656 23994 45665
rect 23938 45591 23994 45600
rect 23952 45490 23980 45591
rect 23940 45484 23992 45490
rect 23940 45426 23992 45432
rect 23756 45076 23808 45082
rect 23756 45018 23808 45024
rect 23848 44940 23900 44946
rect 23848 44882 23900 44888
rect 23570 44432 23626 44441
rect 23570 44367 23626 44376
rect 23584 43722 23612 44367
rect 23860 44334 23888 44882
rect 24044 44334 24072 45902
rect 24308 45892 24360 45898
rect 24308 45834 24360 45840
rect 24124 45348 24176 45354
rect 24124 45290 24176 45296
rect 23848 44328 23900 44334
rect 24032 44328 24084 44334
rect 23848 44270 23900 44276
rect 24030 44296 24032 44305
rect 24084 44296 24086 44305
rect 23860 43858 23888 44270
rect 24030 44231 24086 44240
rect 23848 43852 23900 43858
rect 23848 43794 23900 43800
rect 23572 43716 23624 43722
rect 23572 43658 23624 43664
rect 23860 43110 23888 43794
rect 23848 43104 23900 43110
rect 23848 43046 23900 43052
rect 23572 41676 23624 41682
rect 23572 41618 23624 41624
rect 23386 41440 23442 41449
rect 23386 41375 23442 41384
rect 23400 40594 23428 41375
rect 23584 41206 23612 41618
rect 23768 41614 23796 41645
rect 23756 41608 23808 41614
rect 23754 41576 23756 41585
rect 23808 41576 23810 41585
rect 23754 41511 23810 41520
rect 23768 41274 23796 41511
rect 23860 41449 23888 43046
rect 24136 42770 24164 45290
rect 24320 45014 24348 45834
rect 24308 45008 24360 45014
rect 24308 44950 24360 44956
rect 24216 44328 24268 44334
rect 24216 44270 24268 44276
rect 24228 43858 24256 44270
rect 24320 43994 24348 44950
rect 24308 43988 24360 43994
rect 24308 43930 24360 43936
rect 24216 43852 24268 43858
rect 24216 43794 24268 43800
rect 24124 42764 24176 42770
rect 24124 42706 24176 42712
rect 24136 42158 24164 42706
rect 24124 42152 24176 42158
rect 24124 42094 24176 42100
rect 24308 42016 24360 42022
rect 24308 41958 24360 41964
rect 24320 41834 24348 41958
rect 24228 41818 24348 41834
rect 24216 41812 24348 41818
rect 24268 41806 24348 41812
rect 24216 41754 24268 41760
rect 23846 41440 23902 41449
rect 23846 41375 23902 41384
rect 23756 41268 23808 41274
rect 23756 41210 23808 41216
rect 23572 41200 23624 41206
rect 23572 41142 23624 41148
rect 23478 41032 23534 41041
rect 23478 40967 23534 40976
rect 23492 40730 23520 40967
rect 23480 40724 23532 40730
rect 23480 40666 23532 40672
rect 23388 40588 23440 40594
rect 23388 40530 23440 40536
rect 23400 40186 23428 40530
rect 23388 40180 23440 40186
rect 23388 40122 23440 40128
rect 23584 39982 23612 41142
rect 23572 39976 23624 39982
rect 23572 39918 23624 39924
rect 24320 38418 24348 41806
rect 24308 38412 24360 38418
rect 24308 38354 24360 38360
rect 24124 38208 24176 38214
rect 24124 38150 24176 38156
rect 23754 37632 23810 37641
rect 23754 37567 23810 37576
rect 23296 37256 23348 37262
rect 23296 37198 23348 37204
rect 23308 36922 23336 37198
rect 23296 36916 23348 36922
rect 23296 36858 23348 36864
rect 23296 36576 23348 36582
rect 23296 36518 23348 36524
rect 23308 36174 23336 36518
rect 23386 36272 23442 36281
rect 23386 36207 23388 36216
rect 23440 36207 23442 36216
rect 23388 36178 23440 36184
rect 23296 36168 23348 36174
rect 23296 36110 23348 36116
rect 23308 35698 23336 36110
rect 23400 35834 23428 36178
rect 23388 35828 23440 35834
rect 23388 35770 23440 35776
rect 23296 35692 23348 35698
rect 23296 35634 23348 35640
rect 23308 35018 23336 35634
rect 23388 35284 23440 35290
rect 23388 35226 23440 35232
rect 23296 35012 23348 35018
rect 23296 34954 23348 34960
rect 23308 34066 23336 34954
rect 23296 34060 23348 34066
rect 23296 34002 23348 34008
rect 23308 33318 23336 34002
rect 23296 33312 23348 33318
rect 23296 33254 23348 33260
rect 23296 32768 23348 32774
rect 23296 32710 23348 32716
rect 23308 32502 23336 32710
rect 23296 32496 23348 32502
rect 23296 32438 23348 32444
rect 23294 32056 23350 32065
rect 23294 31991 23296 32000
rect 23348 31991 23350 32000
rect 23296 31962 23348 31968
rect 23308 31822 23336 31962
rect 23296 31816 23348 31822
rect 23400 31804 23428 35226
rect 23480 35216 23532 35222
rect 23480 35158 23532 35164
rect 23492 34542 23520 35158
rect 23768 34762 23796 37567
rect 23848 37324 23900 37330
rect 23848 37266 23900 37272
rect 23860 36378 23888 37266
rect 23848 36372 23900 36378
rect 23848 36314 23900 36320
rect 23940 35488 23992 35494
rect 23940 35430 23992 35436
rect 23952 35018 23980 35430
rect 23940 35012 23992 35018
rect 23940 34954 23992 34960
rect 23848 34944 23900 34950
rect 23846 34912 23848 34921
rect 23900 34912 23902 34921
rect 23846 34847 23902 34856
rect 23768 34734 23888 34762
rect 23480 34536 23532 34542
rect 23480 34478 23532 34484
rect 23756 33924 23808 33930
rect 23756 33866 23808 33872
rect 23768 33454 23796 33866
rect 23756 33448 23808 33454
rect 23756 33390 23808 33396
rect 23756 33312 23808 33318
rect 23756 33254 23808 33260
rect 23768 32910 23796 33254
rect 23664 32904 23716 32910
rect 23662 32872 23664 32881
rect 23756 32904 23808 32910
rect 23716 32872 23718 32881
rect 23756 32846 23808 32852
rect 23662 32807 23718 32816
rect 23664 32360 23716 32366
rect 23768 32348 23796 32846
rect 23716 32320 23796 32348
rect 23664 32302 23716 32308
rect 23676 32201 23704 32302
rect 23662 32192 23718 32201
rect 23662 32127 23718 32136
rect 23400 31776 23612 31804
rect 23296 31758 23348 31764
rect 23308 28082 23336 31758
rect 23584 31736 23612 31776
rect 23492 31708 23612 31736
rect 23492 31278 23520 31708
rect 23570 31648 23626 31657
rect 23570 31583 23626 31592
rect 23480 31272 23532 31278
rect 23480 31214 23532 31220
rect 23388 31136 23440 31142
rect 23388 31078 23440 31084
rect 23400 30190 23428 31078
rect 23478 30288 23534 30297
rect 23478 30223 23534 30232
rect 23388 30184 23440 30190
rect 23388 30126 23440 30132
rect 23400 29782 23428 30126
rect 23492 29782 23520 30223
rect 23388 29776 23440 29782
rect 23388 29718 23440 29724
rect 23480 29776 23532 29782
rect 23480 29718 23532 29724
rect 23492 29306 23520 29718
rect 23480 29300 23532 29306
rect 23480 29242 23532 29248
rect 23480 29164 23532 29170
rect 23480 29106 23532 29112
rect 23388 28688 23440 28694
rect 23388 28630 23440 28636
rect 23296 28076 23348 28082
rect 23296 28018 23348 28024
rect 23400 27985 23428 28630
rect 23386 27976 23442 27985
rect 23386 27911 23442 27920
rect 23294 27568 23350 27577
rect 23294 27503 23350 27512
rect 23308 27169 23336 27503
rect 23400 27470 23428 27911
rect 23388 27464 23440 27470
rect 23388 27406 23440 27412
rect 23294 27160 23350 27169
rect 23294 27095 23350 27104
rect 23308 26926 23336 27095
rect 23400 26994 23428 27406
rect 23388 26988 23440 26994
rect 23388 26930 23440 26936
rect 23296 26920 23348 26926
rect 23492 26874 23520 29106
rect 23296 26862 23348 26868
rect 23400 26846 23520 26874
rect 23400 26353 23428 26846
rect 23480 26784 23532 26790
rect 23480 26726 23532 26732
rect 23492 26586 23520 26726
rect 23480 26580 23532 26586
rect 23480 26522 23532 26528
rect 23480 26376 23532 26382
rect 23386 26344 23442 26353
rect 23480 26318 23532 26324
rect 23386 26279 23442 26288
rect 23296 26240 23348 26246
rect 23492 26194 23520 26318
rect 23296 26182 23348 26188
rect 23308 25673 23336 26182
rect 23400 26166 23520 26194
rect 23294 25664 23350 25673
rect 23294 25599 23350 25608
rect 23308 23866 23336 25599
rect 23400 24274 23428 26166
rect 23480 26036 23532 26042
rect 23480 25978 23532 25984
rect 23492 24954 23520 25978
rect 23480 24948 23532 24954
rect 23480 24890 23532 24896
rect 23388 24268 23440 24274
rect 23388 24210 23440 24216
rect 23480 24268 23532 24274
rect 23480 24210 23532 24216
rect 23296 23860 23348 23866
rect 23296 23802 23348 23808
rect 23388 23180 23440 23186
rect 23492 23168 23520 24210
rect 23584 24206 23612 31583
rect 23754 31512 23810 31521
rect 23754 31447 23810 31456
rect 23768 31210 23796 31447
rect 23756 31204 23808 31210
rect 23756 31146 23808 31152
rect 23664 30932 23716 30938
rect 23664 30874 23716 30880
rect 23676 30054 23704 30874
rect 23756 30592 23808 30598
rect 23756 30534 23808 30540
rect 23664 30048 23716 30054
rect 23664 29990 23716 29996
rect 23768 29850 23796 30534
rect 23860 30326 23888 34734
rect 24032 34400 24084 34406
rect 24032 34342 24084 34348
rect 24044 34082 24072 34342
rect 24136 34202 24164 38150
rect 24320 38010 24348 38354
rect 24308 38004 24360 38010
rect 24308 37946 24360 37952
rect 24216 37120 24268 37126
rect 24216 37062 24268 37068
rect 24228 36038 24256 37062
rect 24216 36032 24268 36038
rect 24216 35974 24268 35980
rect 24216 34740 24268 34746
rect 24216 34682 24268 34688
rect 24124 34196 24176 34202
rect 24124 34138 24176 34144
rect 24044 34054 24164 34082
rect 24136 33454 24164 34054
rect 24124 33448 24176 33454
rect 24124 33390 24176 33396
rect 24136 32434 24164 33390
rect 24228 32978 24256 34682
rect 24216 32972 24268 32978
rect 24216 32914 24268 32920
rect 24124 32428 24176 32434
rect 24124 32370 24176 32376
rect 23940 32360 23992 32366
rect 23938 32328 23940 32337
rect 23992 32328 23994 32337
rect 23938 32263 23994 32272
rect 24214 32328 24270 32337
rect 24214 32263 24270 32272
rect 24228 32026 24256 32263
rect 24216 32020 24268 32026
rect 24216 31962 24268 31968
rect 24124 31952 24176 31958
rect 24124 31894 24176 31900
rect 23940 31748 23992 31754
rect 23940 31690 23992 31696
rect 23952 31634 23980 31690
rect 23952 31606 24072 31634
rect 24044 31414 24072 31606
rect 24032 31408 24084 31414
rect 24032 31350 24084 31356
rect 23940 31340 23992 31346
rect 23940 31282 23992 31288
rect 23952 30938 23980 31282
rect 23940 30932 23992 30938
rect 23940 30874 23992 30880
rect 23848 30320 23900 30326
rect 24044 30297 24072 31350
rect 23848 30262 23900 30268
rect 24030 30288 24086 30297
rect 24030 30223 24086 30232
rect 23940 30184 23992 30190
rect 24136 30138 24164 31894
rect 24308 31816 24360 31822
rect 24308 31758 24360 31764
rect 24320 30666 24348 31758
rect 24308 30660 24360 30666
rect 24308 30602 24360 30608
rect 24216 30592 24268 30598
rect 24216 30534 24268 30540
rect 24228 30190 24256 30534
rect 23940 30126 23992 30132
rect 23952 29889 23980 30126
rect 24044 30122 24164 30138
rect 24216 30184 24268 30190
rect 24216 30126 24268 30132
rect 24032 30116 24164 30122
rect 24084 30110 24164 30116
rect 24032 30058 24084 30064
rect 23938 29880 23994 29889
rect 23756 29844 23808 29850
rect 23938 29815 23994 29824
rect 23756 29786 23808 29792
rect 23846 29744 23902 29753
rect 23846 29679 23902 29688
rect 23662 29608 23718 29617
rect 23662 29543 23718 29552
rect 23676 28762 23704 29543
rect 23860 29170 23888 29679
rect 23940 29572 23992 29578
rect 23940 29514 23992 29520
rect 23848 29164 23900 29170
rect 23848 29106 23900 29112
rect 23756 29096 23808 29102
rect 23756 29038 23808 29044
rect 23768 28801 23796 29038
rect 23754 28792 23810 28801
rect 23664 28756 23716 28762
rect 23810 28750 23888 28778
rect 23952 28762 23980 29514
rect 23754 28727 23810 28736
rect 23664 28698 23716 28704
rect 23676 27606 23704 28698
rect 23860 27656 23888 28750
rect 23940 28756 23992 28762
rect 23940 28698 23992 28704
rect 23952 28422 23980 28698
rect 23940 28416 23992 28422
rect 23940 28358 23992 28364
rect 23938 28248 23994 28257
rect 24044 28234 24072 30058
rect 24124 30048 24176 30054
rect 24124 29990 24176 29996
rect 24136 28393 24164 29990
rect 24320 29850 24348 30602
rect 24308 29844 24360 29850
rect 24308 29786 24360 29792
rect 24216 28620 24268 28626
rect 24216 28562 24268 28568
rect 24122 28384 24178 28393
rect 24122 28319 24178 28328
rect 24044 28206 24164 28234
rect 23938 28183 23940 28192
rect 23992 28183 23994 28192
rect 23940 28154 23992 28160
rect 24032 28144 24084 28150
rect 24032 28086 24084 28092
rect 23940 27940 23992 27946
rect 24044 27928 24072 28086
rect 23992 27900 24072 27928
rect 23940 27882 23992 27888
rect 23768 27628 23888 27656
rect 23664 27600 23716 27606
rect 23664 27542 23716 27548
rect 23664 27464 23716 27470
rect 23664 27406 23716 27412
rect 23572 24200 23624 24206
rect 23572 24142 23624 24148
rect 23584 23186 23612 24142
rect 23676 23905 23704 27406
rect 23768 25362 23796 27628
rect 23848 27532 23900 27538
rect 23848 27474 23900 27480
rect 23860 27334 23888 27474
rect 23848 27328 23900 27334
rect 23848 27270 23900 27276
rect 23756 25356 23808 25362
rect 23756 25298 23808 25304
rect 23768 24834 23796 25298
rect 23860 25265 23888 27270
rect 23952 27062 23980 27882
rect 24136 27674 24164 28206
rect 24124 27668 24176 27674
rect 24124 27610 24176 27616
rect 24032 27600 24084 27606
rect 24032 27542 24084 27548
rect 23940 27056 23992 27062
rect 23940 26998 23992 27004
rect 23952 26518 23980 26998
rect 24044 26858 24072 27542
rect 24124 27464 24176 27470
rect 24124 27406 24176 27412
rect 24032 26852 24084 26858
rect 24032 26794 24084 26800
rect 23940 26512 23992 26518
rect 23940 26454 23992 26460
rect 23938 26344 23994 26353
rect 24136 26314 24164 27406
rect 24228 26450 24256 28562
rect 24308 28416 24360 28422
rect 24308 28358 24360 28364
rect 24320 26994 24348 28358
rect 24308 26988 24360 26994
rect 24308 26930 24360 26936
rect 24308 26784 24360 26790
rect 24308 26726 24360 26732
rect 24216 26444 24268 26450
rect 24216 26386 24268 26392
rect 24228 26353 24256 26386
rect 24214 26344 24270 26353
rect 23938 26279 23994 26288
rect 24124 26308 24176 26314
rect 23952 25906 23980 26279
rect 24214 26279 24270 26288
rect 24124 26250 24176 26256
rect 23940 25900 23992 25906
rect 23940 25842 23992 25848
rect 23952 25362 23980 25842
rect 24032 25832 24084 25838
rect 24032 25774 24084 25780
rect 24044 25362 24072 25774
rect 24124 25696 24176 25702
rect 24124 25638 24176 25644
rect 23940 25356 23992 25362
rect 23940 25298 23992 25304
rect 24032 25356 24084 25362
rect 24032 25298 24084 25304
rect 23846 25256 23902 25265
rect 23846 25191 23902 25200
rect 23768 24806 23980 24834
rect 23756 24744 23808 24750
rect 23756 24686 23808 24692
rect 23768 24585 23796 24686
rect 23754 24576 23810 24585
rect 23754 24511 23810 24520
rect 23846 24440 23902 24449
rect 23756 24404 23808 24410
rect 23846 24375 23902 24384
rect 23756 24346 23808 24352
rect 23768 24313 23796 24346
rect 23754 24304 23810 24313
rect 23754 24239 23810 24248
rect 23662 23896 23718 23905
rect 23860 23866 23888 24375
rect 23952 24138 23980 24806
rect 23940 24132 23992 24138
rect 23940 24074 23992 24080
rect 23662 23831 23718 23840
rect 23848 23860 23900 23866
rect 23848 23802 23900 23808
rect 23662 23760 23718 23769
rect 23662 23695 23718 23704
rect 23676 23662 23704 23695
rect 23952 23662 23980 24074
rect 23664 23656 23716 23662
rect 23664 23598 23716 23604
rect 23940 23656 23992 23662
rect 23940 23598 23992 23604
rect 23440 23140 23520 23168
rect 23572 23180 23624 23186
rect 23388 23122 23440 23128
rect 23572 23122 23624 23128
rect 23848 23112 23900 23118
rect 23294 23080 23350 23089
rect 23848 23054 23900 23060
rect 23294 23015 23350 23024
rect 23308 14482 23336 23015
rect 23860 22778 23888 23054
rect 24044 22817 24072 25298
rect 24030 22808 24086 22817
rect 23848 22772 23900 22778
rect 24030 22743 24086 22752
rect 23848 22714 23900 22720
rect 23860 22681 23888 22714
rect 23846 22672 23902 22681
rect 23846 22607 23902 22616
rect 23388 22024 23440 22030
rect 23386 21992 23388 22001
rect 23440 21992 23442 22001
rect 23386 21927 23442 21936
rect 23400 21690 23428 21927
rect 23388 21684 23440 21690
rect 23388 21626 23440 21632
rect 23846 19272 23902 19281
rect 23846 19207 23902 19216
rect 23860 18970 23888 19207
rect 23848 18964 23900 18970
rect 23848 18906 23900 18912
rect 24136 17241 24164 25638
rect 24216 24676 24268 24682
rect 24216 24618 24268 24624
rect 24228 24274 24256 24618
rect 24216 24268 24268 24274
rect 24216 24210 24268 24216
rect 24228 23866 24256 24210
rect 24216 23860 24268 23866
rect 24216 23802 24268 23808
rect 24320 22409 24348 26726
rect 24306 22400 24362 22409
rect 24306 22335 24362 22344
rect 24122 17232 24178 17241
rect 24122 17167 24178 17176
rect 24308 16652 24360 16658
rect 24308 16594 24360 16600
rect 23848 16584 23900 16590
rect 23848 16526 23900 16532
rect 23860 15910 23888 16526
rect 24320 15910 24348 16594
rect 23848 15904 23900 15910
rect 23848 15846 23900 15852
rect 24308 15904 24360 15910
rect 24308 15846 24360 15852
rect 23296 14476 23348 14482
rect 23296 14418 23348 14424
rect 23112 14214 23164 14220
rect 23202 14240 23258 14249
rect 23124 13977 23152 14214
rect 23202 14175 23258 14184
rect 23308 14074 23336 14418
rect 23296 14068 23348 14074
rect 23296 14010 23348 14016
rect 23110 13968 23166 13977
rect 23110 13903 23166 13912
rect 23478 13424 23534 13433
rect 23478 13359 23534 13368
rect 23492 7449 23520 13359
rect 23478 7440 23534 7449
rect 23478 7375 23534 7384
rect 23860 7313 23888 15846
rect 23938 11112 23994 11121
rect 23938 11047 23994 11056
rect 23846 7304 23902 7313
rect 23846 7239 23902 7248
rect 23018 5128 23074 5137
rect 23018 5063 23074 5072
rect 22744 4072 22796 4078
rect 22744 4014 22796 4020
rect 22376 3188 22428 3194
rect 22376 3130 22428 3136
rect 22204 3046 22600 3074
rect 20812 2644 20864 2650
rect 20812 2586 20864 2592
rect 21652 2638 21772 2666
rect 21652 800 21680 2638
rect 22572 800 22600 3046
rect 3422 776 3478 785
rect 3422 711 3478 720
rect 4158 0 4214 800
rect 5078 0 5134 800
rect 5998 0 6054 800
rect 6918 0 6974 800
rect 7838 0 7894 800
rect 8298 0 8354 800
rect 9218 0 9274 800
rect 10138 0 10194 800
rect 11058 0 11114 800
rect 11978 0 12034 800
rect 12898 0 12954 800
rect 13818 0 13874 800
rect 14738 0 14794 800
rect 15658 0 15714 800
rect 16118 0 16174 800
rect 17038 0 17094 800
rect 17958 0 18014 800
rect 18878 0 18934 800
rect 19798 0 19854 800
rect 20718 0 20774 800
rect 21638 0 21694 800
rect 22558 0 22614 800
rect 22756 241 22784 4014
rect 23754 2408 23810 2417
rect 23754 2343 23756 2352
rect 23808 2343 23810 2352
rect 23756 2314 23808 2320
rect 23480 1420 23532 1426
rect 23480 1362 23532 1368
rect 23492 800 23520 1362
rect 23952 800 23980 11047
rect 24412 7721 24440 53450
rect 24504 52494 24532 53586
rect 24492 52488 24544 52494
rect 24492 52430 24544 52436
rect 24492 50380 24544 50386
rect 24492 50322 24544 50328
rect 24504 50289 24532 50322
rect 24490 50280 24546 50289
rect 24490 50215 24546 50224
rect 24490 48240 24546 48249
rect 24490 48175 24492 48184
rect 24544 48175 24546 48184
rect 24492 48146 24544 48152
rect 24492 47592 24544 47598
rect 24492 47534 24544 47540
rect 24504 47025 24532 47534
rect 24490 47016 24546 47025
rect 24490 46951 24546 46960
rect 24492 43308 24544 43314
rect 24492 43250 24544 43256
rect 24504 42906 24532 43250
rect 24492 42900 24544 42906
rect 24492 42842 24544 42848
rect 24492 38344 24544 38350
rect 24492 38286 24544 38292
rect 24504 37369 24532 38286
rect 24490 37360 24546 37369
rect 24490 37295 24546 37304
rect 24492 34536 24544 34542
rect 24492 34478 24544 34484
rect 24504 33454 24532 34478
rect 24492 33448 24544 33454
rect 24492 33390 24544 33396
rect 24504 31482 24532 33390
rect 24492 31476 24544 31482
rect 24492 31418 24544 31424
rect 24492 31204 24544 31210
rect 24492 31146 24544 31152
rect 24504 30802 24532 31146
rect 24492 30796 24544 30802
rect 24492 30738 24544 30744
rect 24492 30660 24544 30666
rect 24492 30602 24544 30608
rect 24504 30122 24532 30602
rect 24492 30116 24544 30122
rect 24492 30058 24544 30064
rect 24492 27600 24544 27606
rect 24492 27542 24544 27548
rect 24504 26625 24532 27542
rect 24490 26616 24546 26625
rect 24490 26551 24546 26560
rect 24504 26450 24532 26551
rect 24492 26444 24544 26450
rect 24492 26386 24544 26392
rect 24490 23080 24546 23089
rect 24490 23015 24492 23024
rect 24544 23015 24546 23024
rect 24492 22986 24544 22992
rect 24492 21888 24544 21894
rect 24490 21856 24492 21865
rect 24544 21856 24546 21865
rect 24490 21791 24546 21800
rect 24398 7712 24454 7721
rect 24398 7647 24454 7656
rect 24596 1426 24624 58822
rect 24780 58546 24808 74423
rect 25686 73944 25742 73953
rect 25686 73879 25742 73888
rect 25228 69284 25280 69290
rect 25228 69226 25280 69232
rect 25240 68882 25268 69226
rect 25228 68876 25280 68882
rect 25228 68818 25280 68824
rect 25240 67658 25268 68818
rect 25318 68232 25374 68241
rect 25318 68167 25374 68176
rect 25228 67652 25280 67658
rect 25228 67594 25280 67600
rect 25332 64410 25360 68167
rect 25240 64382 25360 64410
rect 24950 61296 25006 61305
rect 24950 61231 25006 61240
rect 24768 58540 24820 58546
rect 24768 58482 24820 58488
rect 24768 57792 24820 57798
rect 24768 57734 24820 57740
rect 24676 56840 24728 56846
rect 24676 56782 24728 56788
rect 24688 55729 24716 56782
rect 24780 56710 24808 57734
rect 24860 56908 24912 56914
rect 24860 56850 24912 56856
rect 24768 56704 24820 56710
rect 24768 56646 24820 56652
rect 24872 56522 24900 56850
rect 24780 56494 24900 56522
rect 24780 56166 24808 56494
rect 24964 56370 24992 61231
rect 25042 59392 25098 59401
rect 25042 59327 25098 59336
rect 25056 57338 25084 59327
rect 25136 59016 25188 59022
rect 25136 58958 25188 58964
rect 25148 58682 25176 58958
rect 25240 58954 25268 64382
rect 25504 60648 25556 60654
rect 25318 60616 25374 60625
rect 25504 60590 25556 60596
rect 25318 60551 25374 60560
rect 25332 60314 25360 60551
rect 25320 60308 25372 60314
rect 25320 60250 25372 60256
rect 25516 59770 25544 60590
rect 25504 59764 25556 59770
rect 25504 59706 25556 59712
rect 25228 58948 25280 58954
rect 25228 58890 25280 58896
rect 25136 58676 25188 58682
rect 25136 58618 25188 58624
rect 25148 57594 25176 58618
rect 25228 58404 25280 58410
rect 25228 58346 25280 58352
rect 25240 58002 25268 58346
rect 25320 58336 25372 58342
rect 25320 58278 25372 58284
rect 25228 57996 25280 58002
rect 25228 57938 25280 57944
rect 25136 57588 25188 57594
rect 25136 57530 25188 57536
rect 25240 57526 25268 57938
rect 25228 57520 25280 57526
rect 25228 57462 25280 57468
rect 25056 57310 25268 57338
rect 25136 56704 25188 56710
rect 25136 56646 25188 56652
rect 24952 56364 25004 56370
rect 24952 56306 25004 56312
rect 25148 56302 25176 56646
rect 25136 56296 25188 56302
rect 25136 56238 25188 56244
rect 24768 56160 24820 56166
rect 24768 56102 24820 56108
rect 24952 55820 25004 55826
rect 24952 55762 25004 55768
rect 24674 55720 24730 55729
rect 24674 55655 24730 55664
rect 24688 55570 24716 55655
rect 24860 55616 24912 55622
rect 24688 55564 24860 55570
rect 24688 55558 24912 55564
rect 24688 55542 24900 55558
rect 24688 53650 24716 55542
rect 24964 55418 24992 55762
rect 24952 55412 25004 55418
rect 24952 55354 25004 55360
rect 24768 54256 24820 54262
rect 24964 54210 24992 55354
rect 25136 54800 25188 54806
rect 25136 54742 25188 54748
rect 25044 54732 25096 54738
rect 25044 54674 25096 54680
rect 24768 54198 24820 54204
rect 24676 53644 24728 53650
rect 24676 53586 24728 53592
rect 24780 53242 24808 54198
rect 24872 54182 24992 54210
rect 24768 53236 24820 53242
rect 24768 53178 24820 53184
rect 24768 52896 24820 52902
rect 24768 52838 24820 52844
rect 24676 52556 24728 52562
rect 24676 52498 24728 52504
rect 24688 51814 24716 52498
rect 24676 51808 24728 51814
rect 24676 51750 24728 51756
rect 24688 50833 24716 51750
rect 24780 51406 24808 52838
rect 24872 52018 24900 54182
rect 25056 54126 25084 54674
rect 24952 54120 25004 54126
rect 24952 54062 25004 54068
rect 25044 54120 25096 54126
rect 25044 54062 25096 54068
rect 24964 53446 24992 54062
rect 24952 53440 25004 53446
rect 24952 53382 25004 53388
rect 24964 52630 24992 53382
rect 25042 53000 25098 53009
rect 25042 52935 25098 52944
rect 24952 52624 25004 52630
rect 24952 52566 25004 52572
rect 24952 52420 25004 52426
rect 24952 52362 25004 52368
rect 24860 52012 24912 52018
rect 24860 51954 24912 51960
rect 24858 51912 24914 51921
rect 24858 51847 24914 51856
rect 24872 51610 24900 51847
rect 24860 51604 24912 51610
rect 24860 51546 24912 51552
rect 24964 51474 24992 52362
rect 25056 51474 25084 52935
rect 25148 52154 25176 54742
rect 25240 53666 25268 57310
rect 25332 56545 25360 58278
rect 25596 57316 25648 57322
rect 25596 57258 25648 57264
rect 25504 56704 25556 56710
rect 25502 56672 25504 56681
rect 25556 56672 25558 56681
rect 25502 56607 25558 56616
rect 25318 56536 25374 56545
rect 25318 56471 25374 56480
rect 25320 56296 25372 56302
rect 25320 56238 25372 56244
rect 25332 53802 25360 56238
rect 25608 55826 25636 57258
rect 25596 55820 25648 55826
rect 25596 55762 25648 55768
rect 25504 54664 25556 54670
rect 25504 54606 25556 54612
rect 25412 54596 25464 54602
rect 25412 54538 25464 54544
rect 25424 54194 25452 54538
rect 25412 54188 25464 54194
rect 25412 54130 25464 54136
rect 25424 53938 25452 54130
rect 25516 54126 25544 54606
rect 25608 54194 25636 55762
rect 25596 54188 25648 54194
rect 25596 54130 25648 54136
rect 25504 54120 25556 54126
rect 25504 54062 25556 54068
rect 25424 53910 25544 53938
rect 25332 53774 25452 53802
rect 25240 53638 25360 53666
rect 25228 53508 25280 53514
rect 25228 53450 25280 53456
rect 25240 53038 25268 53450
rect 25228 53032 25280 53038
rect 25228 52974 25280 52980
rect 25226 52184 25282 52193
rect 25136 52148 25188 52154
rect 25226 52119 25282 52128
rect 25136 52090 25188 52096
rect 24952 51468 25004 51474
rect 24952 51410 25004 51416
rect 25044 51468 25096 51474
rect 25044 51410 25096 51416
rect 24768 51400 24820 51406
rect 24768 51342 24820 51348
rect 24858 51368 24914 51377
rect 24858 51303 24914 51312
rect 24872 51066 24900 51303
rect 24950 51232 25006 51241
rect 24950 51167 25006 51176
rect 24860 51060 24912 51066
rect 24860 51002 24912 51008
rect 24768 50992 24820 50998
rect 24768 50934 24820 50940
rect 24674 50824 24730 50833
rect 24674 50759 24730 50768
rect 24674 49736 24730 49745
rect 24674 49671 24730 49680
rect 24688 48385 24716 49671
rect 24780 49434 24808 50934
rect 24860 50856 24912 50862
rect 24860 50798 24912 50804
rect 24768 49428 24820 49434
rect 24768 49370 24820 49376
rect 24768 49224 24820 49230
rect 24768 49166 24820 49172
rect 24674 48376 24730 48385
rect 24674 48311 24730 48320
rect 24688 48142 24716 48311
rect 24676 48136 24728 48142
rect 24676 48078 24728 48084
rect 24676 47592 24728 47598
rect 24676 47534 24728 47540
rect 24688 46578 24716 47534
rect 24676 46572 24728 46578
rect 24676 46514 24728 46520
rect 24676 45960 24728 45966
rect 24676 45902 24728 45908
rect 24688 45558 24716 45902
rect 24676 45552 24728 45558
rect 24676 45494 24728 45500
rect 24688 44946 24716 45494
rect 24676 44940 24728 44946
rect 24676 44882 24728 44888
rect 24688 44538 24716 44882
rect 24676 44532 24728 44538
rect 24676 44474 24728 44480
rect 24674 44024 24730 44033
rect 24674 43959 24730 43968
rect 24688 43314 24716 43959
rect 24676 43308 24728 43314
rect 24676 43250 24728 43256
rect 24674 43208 24730 43217
rect 24674 43143 24676 43152
rect 24728 43143 24730 43152
rect 24676 43114 24728 43120
rect 24780 40905 24808 49166
rect 24872 47841 24900 50798
rect 24964 48890 24992 51167
rect 25240 50153 25268 52119
rect 25332 52034 25360 53638
rect 25424 52193 25452 53774
rect 25516 53446 25544 53910
rect 25504 53440 25556 53446
rect 25504 53382 25556 53388
rect 25410 52184 25466 52193
rect 25516 52154 25544 53382
rect 25596 53100 25648 53106
rect 25596 53042 25648 53048
rect 25410 52119 25466 52128
rect 25504 52148 25556 52154
rect 25504 52090 25556 52096
rect 25332 52006 25452 52034
rect 25320 51808 25372 51814
rect 25320 51750 25372 51756
rect 25332 51474 25360 51750
rect 25320 51468 25372 51474
rect 25320 51410 25372 51416
rect 25332 50182 25360 51410
rect 25320 50176 25372 50182
rect 25226 50144 25282 50153
rect 25320 50118 25372 50124
rect 25226 50079 25282 50088
rect 25136 49836 25188 49842
rect 25136 49778 25188 49784
rect 25044 49428 25096 49434
rect 25044 49370 25096 49376
rect 24952 48884 25004 48890
rect 24952 48826 25004 48832
rect 25056 48686 25084 49370
rect 25044 48680 25096 48686
rect 25044 48622 25096 48628
rect 24952 48544 25004 48550
rect 24952 48486 25004 48492
rect 24964 48226 24992 48486
rect 25056 48346 25084 48622
rect 25044 48340 25096 48346
rect 25044 48282 25096 48288
rect 25148 48226 25176 49778
rect 25240 49706 25268 50079
rect 25228 49700 25280 49706
rect 25228 49642 25280 49648
rect 25424 49042 25452 52006
rect 25502 51096 25558 51105
rect 25502 51031 25558 51040
rect 25516 50862 25544 51031
rect 25608 50969 25636 53042
rect 25594 50960 25650 50969
rect 25594 50895 25650 50904
rect 25504 50856 25556 50862
rect 25504 50798 25556 50804
rect 25596 50176 25648 50182
rect 25596 50118 25648 50124
rect 25608 49774 25636 50118
rect 25596 49768 25648 49774
rect 25596 49710 25648 49716
rect 25504 49700 25556 49706
rect 25504 49642 25556 49648
rect 25240 49014 25452 49042
rect 25240 48618 25268 49014
rect 25412 48884 25464 48890
rect 25412 48826 25464 48832
rect 25228 48612 25280 48618
rect 25228 48554 25280 48560
rect 25240 48385 25268 48554
rect 25226 48376 25282 48385
rect 25226 48311 25282 48320
rect 24964 48198 25176 48226
rect 24858 47832 24914 47841
rect 24858 47767 24914 47776
rect 24964 47666 24992 48198
rect 24952 47660 25004 47666
rect 24952 47602 25004 47608
rect 25240 47410 25268 48311
rect 25320 47524 25372 47530
rect 25320 47466 25372 47472
rect 25332 47433 25360 47466
rect 25148 47382 25268 47410
rect 25318 47424 25374 47433
rect 24860 46504 24912 46510
rect 24860 46446 24912 46452
rect 24872 46034 24900 46446
rect 24860 46028 24912 46034
rect 24860 45970 24912 45976
rect 24872 45286 24900 45970
rect 25044 45416 25096 45422
rect 25044 45358 25096 45364
rect 24860 45280 24912 45286
rect 24860 45222 24912 45228
rect 24872 44928 24900 45222
rect 24952 44940 25004 44946
rect 24872 44900 24952 44928
rect 24872 43994 24900 44900
rect 24952 44882 25004 44888
rect 24952 44260 25004 44266
rect 24952 44202 25004 44208
rect 24860 43988 24912 43994
rect 24860 43930 24912 43936
rect 24860 41472 24912 41478
rect 24858 41440 24860 41449
rect 24912 41440 24914 41449
rect 24858 41375 24914 41384
rect 24766 40896 24822 40905
rect 24766 40831 24822 40840
rect 24766 40760 24822 40769
rect 24766 40695 24822 40704
rect 24674 34776 24730 34785
rect 24674 34711 24676 34720
rect 24728 34711 24730 34720
rect 24676 34682 24728 34688
rect 24676 33856 24728 33862
rect 24676 33798 24728 33804
rect 24688 33454 24716 33798
rect 24780 33658 24808 40695
rect 24964 37330 24992 44202
rect 25056 43722 25084 45358
rect 25044 43716 25096 43722
rect 25044 43658 25096 43664
rect 25056 39506 25084 43658
rect 25148 43246 25176 47382
rect 25318 47359 25374 47368
rect 25226 47288 25282 47297
rect 25226 47223 25282 47232
rect 25240 47122 25268 47223
rect 25228 47116 25280 47122
rect 25228 47058 25280 47064
rect 25240 46714 25268 47058
rect 25228 46708 25280 46714
rect 25228 46650 25280 46656
rect 25240 44742 25268 46650
rect 25228 44736 25280 44742
rect 25228 44678 25280 44684
rect 25228 43852 25280 43858
rect 25228 43794 25280 43800
rect 25136 43240 25188 43246
rect 25136 43182 25188 43188
rect 25148 42906 25176 43182
rect 25136 42900 25188 42906
rect 25136 42842 25188 42848
rect 25240 42566 25268 43794
rect 25228 42560 25280 42566
rect 25228 42502 25280 42508
rect 25136 39976 25188 39982
rect 25136 39918 25188 39924
rect 25148 39642 25176 39918
rect 25136 39636 25188 39642
rect 25136 39578 25188 39584
rect 25044 39500 25096 39506
rect 25044 39442 25096 39448
rect 25056 38554 25084 39442
rect 25148 38962 25176 39578
rect 25136 38956 25188 38962
rect 25136 38898 25188 38904
rect 25044 38548 25096 38554
rect 25044 38490 25096 38496
rect 24952 37324 25004 37330
rect 24952 37266 25004 37272
rect 25042 34640 25098 34649
rect 25042 34575 25098 34584
rect 24860 34468 24912 34474
rect 24860 34410 24912 34416
rect 24768 33652 24820 33658
rect 24768 33594 24820 33600
rect 24872 33454 24900 34410
rect 25056 34202 25084 34575
rect 25044 34196 25096 34202
rect 25044 34138 25096 34144
rect 24676 33448 24728 33454
rect 24676 33390 24728 33396
rect 24860 33448 24912 33454
rect 24860 33390 24912 33396
rect 25042 33416 25098 33425
rect 24688 33266 24716 33390
rect 25042 33351 25098 33360
rect 24688 33238 24900 33266
rect 24872 32570 24900 33238
rect 24952 32836 25004 32842
rect 24952 32778 25004 32784
rect 24860 32564 24912 32570
rect 24860 32506 24912 32512
rect 24858 32464 24914 32473
rect 24858 32399 24914 32408
rect 24872 32026 24900 32399
rect 24860 32020 24912 32026
rect 24860 31962 24912 31968
rect 24964 31890 24992 32778
rect 25056 32026 25084 33351
rect 25044 32020 25096 32026
rect 25044 31962 25096 31968
rect 24768 31884 24820 31890
rect 24768 31826 24820 31832
rect 24952 31884 25004 31890
rect 24952 31826 25004 31832
rect 24780 31210 24808 31826
rect 24952 31476 25004 31482
rect 24952 31418 25004 31424
rect 24964 31260 24992 31418
rect 25056 31385 25084 31962
rect 25136 31816 25188 31822
rect 25136 31758 25188 31764
rect 25042 31376 25098 31385
rect 25042 31311 25098 31320
rect 24964 31232 25084 31260
rect 24768 31204 24820 31210
rect 24768 31146 24820 31152
rect 24952 31136 25004 31142
rect 24858 31104 24914 31113
rect 24952 31078 25004 31084
rect 24858 31039 24914 31048
rect 24872 30938 24900 31039
rect 24860 30932 24912 30938
rect 24860 30874 24912 30880
rect 24860 30796 24912 30802
rect 24860 30738 24912 30744
rect 24676 30728 24728 30734
rect 24676 30670 24728 30676
rect 24688 30054 24716 30670
rect 24768 30252 24820 30258
rect 24768 30194 24820 30200
rect 24676 30048 24728 30054
rect 24674 30016 24676 30025
rect 24728 30016 24730 30025
rect 24674 29951 24730 29960
rect 24780 29889 24808 30194
rect 24766 29880 24822 29889
rect 24872 29850 24900 30738
rect 24964 30598 24992 31078
rect 24952 30592 25004 30598
rect 24952 30534 25004 30540
rect 24950 30288 25006 30297
rect 24950 30223 25006 30232
rect 24964 30054 24992 30223
rect 24952 30048 25004 30054
rect 24952 29990 25004 29996
rect 24766 29815 24822 29824
rect 24860 29844 24912 29850
rect 24780 29782 24808 29815
rect 24860 29786 24912 29792
rect 24768 29776 24820 29782
rect 24768 29718 24820 29724
rect 24964 29594 24992 29990
rect 24780 29566 24992 29594
rect 24780 28422 24808 29566
rect 24860 28756 24912 28762
rect 24860 28698 24912 28704
rect 24768 28416 24820 28422
rect 24768 28358 24820 28364
rect 24872 28014 24900 28698
rect 25056 28422 25084 31232
rect 25044 28416 25096 28422
rect 25044 28358 25096 28364
rect 24676 28008 24728 28014
rect 24676 27950 24728 27956
rect 24860 28008 24912 28014
rect 24860 27950 24912 27956
rect 24688 27674 24716 27950
rect 24872 27690 24900 27950
rect 25044 27872 25096 27878
rect 25044 27814 25096 27820
rect 24676 27668 24728 27674
rect 24872 27662 24992 27690
rect 24676 27610 24728 27616
rect 24676 27532 24728 27538
rect 24728 27492 24808 27520
rect 24676 27474 24728 27480
rect 24676 26920 24728 26926
rect 24676 26862 24728 26868
rect 24688 26625 24716 26862
rect 24780 26790 24808 27492
rect 24860 27328 24912 27334
rect 24860 27270 24912 27276
rect 24768 26784 24820 26790
rect 24766 26752 24768 26761
rect 24820 26752 24822 26761
rect 24766 26687 24822 26696
rect 24674 26616 24730 26625
rect 24674 26551 24730 26560
rect 24688 26518 24716 26551
rect 24676 26512 24728 26518
rect 24676 26454 24728 26460
rect 24872 25945 24900 27270
rect 24858 25936 24914 25945
rect 24964 25906 24992 27662
rect 25056 27130 25084 27814
rect 25044 27124 25096 27130
rect 25044 27066 25096 27072
rect 25042 27024 25098 27033
rect 25042 26959 25098 26968
rect 25056 26466 25084 26959
rect 25148 26586 25176 31758
rect 25136 26580 25188 26586
rect 25136 26522 25188 26528
rect 25056 26438 25176 26466
rect 25044 26308 25096 26314
rect 25044 26250 25096 26256
rect 25056 26217 25084 26250
rect 25042 26208 25098 26217
rect 25042 26143 25098 26152
rect 24858 25871 24914 25880
rect 24952 25900 25004 25906
rect 24952 25842 25004 25848
rect 24860 25832 24912 25838
rect 24860 25774 24912 25780
rect 24768 25288 24820 25294
rect 24768 25230 24820 25236
rect 24674 24848 24730 24857
rect 24674 24783 24676 24792
rect 24728 24783 24730 24792
rect 24676 24754 24728 24760
rect 24780 24426 24808 25230
rect 24872 25158 24900 25774
rect 24860 25152 24912 25158
rect 24860 25094 24912 25100
rect 24688 24410 24808 24426
rect 24872 24410 24900 25094
rect 24964 24818 24992 25842
rect 24952 24812 25004 24818
rect 24952 24754 25004 24760
rect 25044 24744 25096 24750
rect 25044 24686 25096 24692
rect 24676 24404 24808 24410
rect 24728 24398 24808 24404
rect 24860 24404 24912 24410
rect 24676 24346 24728 24352
rect 24860 24346 24912 24352
rect 25056 24342 25084 24686
rect 25148 24426 25176 26438
rect 25240 24800 25268 42502
rect 25332 38486 25360 47359
rect 25424 47258 25452 48826
rect 25412 47252 25464 47258
rect 25412 47194 25464 47200
rect 25412 45824 25464 45830
rect 25410 45792 25412 45801
rect 25464 45792 25466 45801
rect 25410 45727 25466 45736
rect 25424 45490 25452 45727
rect 25412 45484 25464 45490
rect 25412 45426 25464 45432
rect 25516 44266 25544 49642
rect 25596 49632 25648 49638
rect 25596 49574 25648 49580
rect 25608 49434 25636 49574
rect 25596 49428 25648 49434
rect 25596 49370 25648 49376
rect 25596 48340 25648 48346
rect 25596 48282 25648 48288
rect 25608 47598 25636 48282
rect 25596 47592 25648 47598
rect 25596 47534 25648 47540
rect 25596 47456 25648 47462
rect 25596 47398 25648 47404
rect 25608 47190 25636 47398
rect 25596 47184 25648 47190
rect 25596 47126 25648 47132
rect 25594 47016 25650 47025
rect 25594 46951 25650 46960
rect 25504 44260 25556 44266
rect 25504 44202 25556 44208
rect 25502 44160 25558 44169
rect 25502 44095 25558 44104
rect 25516 43314 25544 44095
rect 25608 43858 25636 46951
rect 25596 43852 25648 43858
rect 25596 43794 25648 43800
rect 25504 43308 25556 43314
rect 25504 43250 25556 43256
rect 25410 40080 25466 40089
rect 25410 40015 25466 40024
rect 25424 38894 25452 40015
rect 25412 38888 25464 38894
rect 25412 38830 25464 38836
rect 25320 38480 25372 38486
rect 25320 38422 25372 38428
rect 25424 37806 25452 38830
rect 25516 38350 25544 43250
rect 25700 42294 25728 73879
rect 25976 69562 26004 75142
rect 26252 74746 26280 79200
rect 26976 76832 27028 76838
rect 26976 76774 27028 76780
rect 26252 74718 26832 74746
rect 26332 73908 26384 73914
rect 26332 73850 26384 73856
rect 26146 69592 26202 69601
rect 25964 69556 26016 69562
rect 26146 69527 26202 69536
rect 25964 69498 26016 69504
rect 25872 68196 25924 68202
rect 25872 68138 25924 68144
rect 25778 64152 25834 64161
rect 25778 64087 25834 64096
rect 25792 62286 25820 64087
rect 25780 62280 25832 62286
rect 25780 62222 25832 62228
rect 25780 56704 25832 56710
rect 25780 56646 25832 56652
rect 25792 56302 25820 56646
rect 25780 56296 25832 56302
rect 25780 56238 25832 56244
rect 25780 55616 25832 55622
rect 25780 55558 25832 55564
rect 25792 54534 25820 55558
rect 25780 54528 25832 54534
rect 25780 54470 25832 54476
rect 25792 54097 25820 54470
rect 25778 54088 25834 54097
rect 25778 54023 25834 54032
rect 25778 53136 25834 53145
rect 25778 53071 25834 53080
rect 25792 52970 25820 53071
rect 25780 52964 25832 52970
rect 25780 52906 25832 52912
rect 25792 52698 25820 52906
rect 25780 52692 25832 52698
rect 25780 52634 25832 52640
rect 25778 52592 25834 52601
rect 25778 52527 25780 52536
rect 25832 52527 25834 52536
rect 25780 52498 25832 52504
rect 25780 51876 25832 51882
rect 25780 51818 25832 51824
rect 25792 50017 25820 51818
rect 25778 50008 25834 50017
rect 25778 49943 25834 49952
rect 25780 48544 25832 48550
rect 25780 48486 25832 48492
rect 25792 47258 25820 48486
rect 25780 47252 25832 47258
rect 25780 47194 25832 47200
rect 25780 46368 25832 46374
rect 25778 46336 25780 46345
rect 25832 46336 25834 46345
rect 25778 46271 25834 46280
rect 25780 44736 25832 44742
rect 25780 44678 25832 44684
rect 25792 42770 25820 44678
rect 25780 42764 25832 42770
rect 25780 42706 25832 42712
rect 25688 42288 25740 42294
rect 25688 42230 25740 42236
rect 25688 42152 25740 42158
rect 25688 42094 25740 42100
rect 25700 41818 25728 42094
rect 25688 41812 25740 41818
rect 25688 41754 25740 41760
rect 25688 40384 25740 40390
rect 25688 40326 25740 40332
rect 25700 40050 25728 40326
rect 25688 40044 25740 40050
rect 25688 39986 25740 39992
rect 25780 39908 25832 39914
rect 25780 39850 25832 39856
rect 25792 38894 25820 39850
rect 25780 38888 25832 38894
rect 25778 38856 25780 38865
rect 25832 38856 25834 38865
rect 25778 38791 25834 38800
rect 25504 38344 25556 38350
rect 25504 38286 25556 38292
rect 25516 38010 25544 38286
rect 25504 38004 25556 38010
rect 25504 37946 25556 37952
rect 25412 37800 25464 37806
rect 25412 37742 25464 37748
rect 25688 37800 25740 37806
rect 25688 37742 25740 37748
rect 25700 37466 25728 37742
rect 25688 37460 25740 37466
rect 25688 37402 25740 37408
rect 25412 36712 25464 36718
rect 25688 36712 25740 36718
rect 25412 36654 25464 36660
rect 25686 36680 25688 36689
rect 25740 36680 25742 36689
rect 25424 36174 25452 36654
rect 25686 36615 25742 36624
rect 25412 36168 25464 36174
rect 25412 36110 25464 36116
rect 25884 34785 25912 68138
rect 25976 62370 26004 69498
rect 25976 62354 26096 62370
rect 25976 62348 26108 62354
rect 25976 62342 26056 62348
rect 26056 62290 26108 62296
rect 25964 62280 26016 62286
rect 25964 62222 26016 62228
rect 25976 55842 26004 62222
rect 26056 61056 26108 61062
rect 26056 60998 26108 61004
rect 26068 60654 26096 60998
rect 26056 60648 26108 60654
rect 26056 60590 26108 60596
rect 26054 56400 26110 56409
rect 26054 56335 26056 56344
rect 26108 56335 26110 56344
rect 26056 56306 26108 56312
rect 25976 55814 26096 55842
rect 25964 54732 26016 54738
rect 25964 54674 26016 54680
rect 25976 53990 26004 54674
rect 25964 53984 26016 53990
rect 25964 53926 26016 53932
rect 25976 49842 26004 53926
rect 25964 49836 26016 49842
rect 25964 49778 26016 49784
rect 25964 49632 26016 49638
rect 25964 49574 26016 49580
rect 25976 49094 26004 49574
rect 25964 49088 26016 49094
rect 25964 49030 26016 49036
rect 25976 48793 26004 49030
rect 25962 48784 26018 48793
rect 25962 48719 26018 48728
rect 25976 48550 26004 48719
rect 25964 48544 26016 48550
rect 25964 48486 26016 48492
rect 25964 47524 26016 47530
rect 25964 47466 26016 47472
rect 25976 46170 26004 47466
rect 25964 46164 26016 46170
rect 25964 46106 26016 46112
rect 25976 45626 26004 46106
rect 25964 45620 26016 45626
rect 25964 45562 26016 45568
rect 25964 44736 26016 44742
rect 25962 44704 25964 44713
rect 26016 44704 26018 44713
rect 25962 44639 26018 44648
rect 25976 44402 26004 44639
rect 25964 44396 26016 44402
rect 25964 44338 26016 44344
rect 25962 44296 26018 44305
rect 25962 44231 26018 44240
rect 25976 43994 26004 44231
rect 25964 43988 26016 43994
rect 25964 43930 26016 43936
rect 25964 42560 26016 42566
rect 25964 42502 26016 42508
rect 25976 42158 26004 42502
rect 25964 42152 26016 42158
rect 25964 42094 26016 42100
rect 26068 38962 26096 55814
rect 26160 44334 26188 69527
rect 26344 65521 26372 73850
rect 26424 67584 26476 67590
rect 26424 67526 26476 67532
rect 26436 67386 26464 67526
rect 26424 67380 26476 67386
rect 26424 67322 26476 67328
rect 26330 65512 26386 65521
rect 26330 65447 26386 65456
rect 26804 62354 26832 74718
rect 26516 62348 26568 62354
rect 26516 62290 26568 62296
rect 26792 62348 26844 62354
rect 26792 62290 26844 62296
rect 26528 61878 26556 62290
rect 26804 61946 26832 62290
rect 26792 61940 26844 61946
rect 26792 61882 26844 61888
rect 26516 61872 26568 61878
rect 26516 61814 26568 61820
rect 26240 60648 26292 60654
rect 26238 60616 26240 60625
rect 26292 60616 26294 60625
rect 26238 60551 26294 60560
rect 26516 60580 26568 60586
rect 26516 60522 26568 60528
rect 26528 59498 26556 60522
rect 26608 60104 26660 60110
rect 26608 60046 26660 60052
rect 26620 59634 26648 60046
rect 26608 59628 26660 59634
rect 26608 59570 26660 59576
rect 26516 59492 26568 59498
rect 26516 59434 26568 59440
rect 26528 59158 26556 59434
rect 26620 59158 26648 59570
rect 26792 59560 26844 59566
rect 26792 59502 26844 59508
rect 26516 59152 26568 59158
rect 26516 59094 26568 59100
rect 26608 59152 26660 59158
rect 26608 59094 26660 59100
rect 26620 58138 26648 59094
rect 26804 58342 26832 59502
rect 26884 58472 26936 58478
rect 26884 58414 26936 58420
rect 26792 58336 26844 58342
rect 26792 58278 26844 58284
rect 26608 58132 26660 58138
rect 26608 58074 26660 58080
rect 26896 57798 26924 58414
rect 26884 57792 26936 57798
rect 26884 57734 26936 57740
rect 26700 57384 26752 57390
rect 26700 57326 26752 57332
rect 26712 57050 26740 57326
rect 26700 57044 26752 57050
rect 26700 56986 26752 56992
rect 26516 56908 26568 56914
rect 26516 56850 26568 56856
rect 26332 56228 26384 56234
rect 26332 56170 26384 56176
rect 26344 55321 26372 56170
rect 26528 56166 26556 56850
rect 26516 56160 26568 56166
rect 26516 56102 26568 56108
rect 26528 55865 26556 56102
rect 26514 55856 26570 55865
rect 26988 55842 27016 76774
rect 27172 73914 27200 79200
rect 28092 77466 28120 79200
rect 28000 77438 28120 77466
rect 27528 75812 27580 75818
rect 27528 75754 27580 75760
rect 27160 73908 27212 73914
rect 27160 73850 27212 73856
rect 27434 72856 27490 72865
rect 27434 72791 27490 72800
rect 27250 67280 27306 67289
rect 27250 67215 27306 67224
rect 27068 67040 27120 67046
rect 27068 66982 27120 66988
rect 27080 60353 27108 66982
rect 27158 64016 27214 64025
rect 27158 63951 27214 63960
rect 27066 60344 27122 60353
rect 27066 60279 27122 60288
rect 27068 59016 27120 59022
rect 27068 58958 27120 58964
rect 27080 55962 27108 58958
rect 27068 55956 27120 55962
rect 27068 55898 27120 55904
rect 26988 55814 27108 55842
rect 26514 55791 26570 55800
rect 26516 55752 26568 55758
rect 26516 55694 26568 55700
rect 26528 55350 26556 55694
rect 26516 55344 26568 55350
rect 26330 55312 26386 55321
rect 26240 55276 26292 55282
rect 26516 55286 26568 55292
rect 26330 55247 26386 55256
rect 26240 55218 26292 55224
rect 26252 54806 26280 55218
rect 26344 55078 26372 55247
rect 26332 55072 26384 55078
rect 26332 55014 26384 55020
rect 26240 54800 26292 54806
rect 26240 54742 26292 54748
rect 26238 54632 26294 54641
rect 26238 54567 26294 54576
rect 26252 54194 26280 54567
rect 26240 54188 26292 54194
rect 26240 54130 26292 54136
rect 26240 54052 26292 54058
rect 26240 53994 26292 54000
rect 26252 53446 26280 53994
rect 26332 53984 26384 53990
rect 26332 53926 26384 53932
rect 26344 53582 26372 53926
rect 26332 53576 26384 53582
rect 26332 53518 26384 53524
rect 26240 53440 26292 53446
rect 26240 53382 26292 53388
rect 26252 53038 26280 53382
rect 26240 53032 26292 53038
rect 26240 52974 26292 52980
rect 26344 52902 26372 53518
rect 26528 53038 26556 55286
rect 26608 55140 26660 55146
rect 26608 55082 26660 55088
rect 26516 53032 26568 53038
rect 26516 52974 26568 52980
rect 26240 52896 26292 52902
rect 26240 52838 26292 52844
rect 26332 52896 26384 52902
rect 26332 52838 26384 52844
rect 26252 52358 26280 52838
rect 26240 52352 26292 52358
rect 26240 52294 26292 52300
rect 26240 51808 26292 51814
rect 26240 51750 26292 51756
rect 26252 49910 26280 51750
rect 26344 51270 26372 52838
rect 26332 51264 26384 51270
rect 26332 51206 26384 51212
rect 26344 49910 26372 51206
rect 26424 50788 26476 50794
rect 26424 50730 26476 50736
rect 26240 49904 26292 49910
rect 26240 49846 26292 49852
rect 26332 49904 26384 49910
rect 26332 49846 26384 49852
rect 26332 49700 26384 49706
rect 26332 49642 26384 49648
rect 26240 49088 26292 49094
rect 26240 49030 26292 49036
rect 26252 48754 26280 49030
rect 26240 48748 26292 48754
rect 26240 48690 26292 48696
rect 26344 48618 26372 49642
rect 26332 48612 26384 48618
rect 26332 48554 26384 48560
rect 26344 48498 26372 48554
rect 26252 48470 26372 48498
rect 26252 48006 26280 48470
rect 26436 48278 26464 50730
rect 26424 48272 26476 48278
rect 26424 48214 26476 48220
rect 26240 48000 26292 48006
rect 26436 47977 26464 48214
rect 26240 47942 26292 47948
rect 26422 47968 26478 47977
rect 26252 45937 26280 47942
rect 26422 47903 26478 47912
rect 26332 47660 26384 47666
rect 26332 47602 26384 47608
rect 26238 45928 26294 45937
rect 26238 45863 26294 45872
rect 26344 45082 26372 47602
rect 26528 46578 26556 52974
rect 26620 48278 26648 55082
rect 26792 55072 26844 55078
rect 26792 55014 26844 55020
rect 26804 54913 26832 55014
rect 26790 54904 26846 54913
rect 26790 54839 26846 54848
rect 26804 54126 26832 54839
rect 26884 54528 26936 54534
rect 26884 54470 26936 54476
rect 26700 54120 26752 54126
rect 26700 54062 26752 54068
rect 26792 54120 26844 54126
rect 26792 54062 26844 54068
rect 26712 53446 26740 54062
rect 26896 54058 26924 54470
rect 26884 54052 26936 54058
rect 26884 53994 26936 54000
rect 26700 53440 26752 53446
rect 26700 53382 26752 53388
rect 26712 53281 26740 53382
rect 26698 53272 26754 53281
rect 26698 53207 26754 53216
rect 26792 52964 26844 52970
rect 26896 52952 26924 53994
rect 26844 52924 26924 52952
rect 26792 52906 26844 52912
rect 26792 52352 26844 52358
rect 26792 52294 26844 52300
rect 26884 52352 26936 52358
rect 26884 52294 26936 52300
rect 26804 51950 26832 52294
rect 26896 51950 26924 52294
rect 26792 51944 26844 51950
rect 26792 51886 26844 51892
rect 26884 51944 26936 51950
rect 26884 51886 26936 51892
rect 26804 50130 26832 51886
rect 26896 51610 26924 51886
rect 26884 51604 26936 51610
rect 26884 51546 26936 51552
rect 26976 51468 27028 51474
rect 26976 51410 27028 51416
rect 26884 51400 26936 51406
rect 26884 51342 26936 51348
rect 26896 50726 26924 51342
rect 26884 50720 26936 50726
rect 26882 50688 26884 50697
rect 26936 50688 26938 50697
rect 26882 50623 26938 50632
rect 26712 50102 26832 50130
rect 26712 49434 26740 50102
rect 26790 50008 26846 50017
rect 26790 49943 26846 49952
rect 26700 49428 26752 49434
rect 26700 49370 26752 49376
rect 26804 49366 26832 49943
rect 26792 49360 26844 49366
rect 26792 49302 26844 49308
rect 26700 49292 26752 49298
rect 26700 49234 26752 49240
rect 26712 48890 26740 49234
rect 26700 48884 26752 48890
rect 26700 48826 26752 48832
rect 26804 48550 26832 49302
rect 26792 48544 26844 48550
rect 26792 48486 26844 48492
rect 26608 48272 26660 48278
rect 26608 48214 26660 48220
rect 26620 47841 26648 48214
rect 26792 48204 26844 48210
rect 26792 48146 26844 48152
rect 26606 47832 26662 47841
rect 26606 47767 26662 47776
rect 26804 47462 26832 48146
rect 26792 47456 26844 47462
rect 26792 47398 26844 47404
rect 26804 47002 26832 47398
rect 26896 47190 26924 50623
rect 26988 50522 27016 51410
rect 27080 50862 27108 55814
rect 27172 53632 27200 63951
rect 27264 59702 27292 67215
rect 27252 59696 27304 59702
rect 27252 59638 27304 59644
rect 27252 59084 27304 59090
rect 27252 59026 27304 59032
rect 27264 58614 27292 59026
rect 27252 58608 27304 58614
rect 27252 58550 27304 58556
rect 27264 57526 27292 58550
rect 27344 57928 27396 57934
rect 27344 57870 27396 57876
rect 27252 57520 27304 57526
rect 27252 57462 27304 57468
rect 27356 56982 27384 57870
rect 27344 56976 27396 56982
rect 27344 56918 27396 56924
rect 27356 56506 27384 56918
rect 27344 56500 27396 56506
rect 27344 56442 27396 56448
rect 27344 53644 27396 53650
rect 27172 53604 27292 53632
rect 27160 53508 27212 53514
rect 27160 53450 27212 53456
rect 27172 53038 27200 53450
rect 27160 53032 27212 53038
rect 27160 52974 27212 52980
rect 27160 52896 27212 52902
rect 27160 52838 27212 52844
rect 27172 52494 27200 52838
rect 27160 52488 27212 52494
rect 27160 52430 27212 52436
rect 27264 51542 27292 53604
rect 27344 53586 27396 53592
rect 27356 52902 27384 53586
rect 27344 52896 27396 52902
rect 27344 52838 27396 52844
rect 27356 52018 27384 52838
rect 27448 52630 27476 72791
rect 27540 69057 27568 75754
rect 28000 74497 28028 77438
rect 28080 77376 28132 77382
rect 28080 77318 28132 77324
rect 28908 77376 28960 77382
rect 28908 77318 28960 77324
rect 27986 74488 28042 74497
rect 27986 74423 28042 74432
rect 27526 69048 27582 69057
rect 27526 68983 27582 68992
rect 27804 62144 27856 62150
rect 27804 62086 27856 62092
rect 27816 60178 27844 62086
rect 27804 60172 27856 60178
rect 27804 60114 27856 60120
rect 27712 58608 27764 58614
rect 27712 58550 27764 58556
rect 27620 58472 27672 58478
rect 27540 58432 27620 58460
rect 27540 57458 27568 58432
rect 27724 58449 27752 58550
rect 27620 58414 27672 58420
rect 27710 58440 27766 58449
rect 27710 58375 27766 58384
rect 27620 58336 27672 58342
rect 27620 58278 27672 58284
rect 27528 57452 27580 57458
rect 27528 57394 27580 57400
rect 27632 56914 27660 58278
rect 28092 57633 28120 77318
rect 28816 76968 28868 76974
rect 28816 76910 28868 76916
rect 28828 76430 28856 76910
rect 28816 76424 28868 76430
rect 28816 76366 28868 76372
rect 28828 76129 28856 76366
rect 28814 76120 28870 76129
rect 28814 76055 28870 76064
rect 28828 76022 28856 76055
rect 28816 76016 28868 76022
rect 28816 75958 28868 75964
rect 28816 73024 28868 73030
rect 28814 72992 28816 73001
rect 28868 72992 28870 73001
rect 28814 72927 28870 72936
rect 28920 70666 28948 77318
rect 29012 76430 29040 79200
rect 29092 77512 29144 77518
rect 29092 77454 29144 77460
rect 29104 77178 29132 77454
rect 29460 77376 29512 77382
rect 29460 77318 29512 77324
rect 29092 77172 29144 77178
rect 29092 77114 29144 77120
rect 29472 76974 29500 77318
rect 29460 76968 29512 76974
rect 29460 76910 29512 76916
rect 29000 76424 29052 76430
rect 29000 76366 29052 76372
rect 29012 76090 29040 76366
rect 29000 76084 29052 76090
rect 29000 76026 29052 76032
rect 29826 75576 29882 75585
rect 29826 75511 29882 75520
rect 29840 75478 29868 75511
rect 29828 75472 29880 75478
rect 29828 75414 29880 75420
rect 29368 75336 29420 75342
rect 29368 75278 29420 75284
rect 29380 74662 29408 75278
rect 29368 74656 29420 74662
rect 29368 74598 29420 74604
rect 28828 70638 28948 70666
rect 28828 70122 28856 70638
rect 28828 70094 28948 70122
rect 28920 62830 28948 70094
rect 28724 62824 28776 62830
rect 28724 62766 28776 62772
rect 28908 62824 28960 62830
rect 28908 62766 28960 62772
rect 28172 60172 28224 60178
rect 28172 60114 28224 60120
rect 28184 59430 28212 60114
rect 28172 59424 28224 59430
rect 28172 59366 28224 59372
rect 28078 57624 28134 57633
rect 28078 57559 28134 57568
rect 27620 56908 27672 56914
rect 27620 56850 27672 56856
rect 27528 56840 27580 56846
rect 27528 56782 27580 56788
rect 27540 56506 27568 56782
rect 27528 56500 27580 56506
rect 27528 56442 27580 56448
rect 27804 56296 27856 56302
rect 27804 56238 27856 56244
rect 27816 55622 27844 56238
rect 27804 55616 27856 55622
rect 27804 55558 27856 55564
rect 27528 54664 27580 54670
rect 27528 54606 27580 54612
rect 27540 53650 27568 54606
rect 27816 53972 27844 55558
rect 27986 55448 28042 55457
rect 27986 55383 28042 55392
rect 28000 55214 28028 55383
rect 27988 55208 28040 55214
rect 27988 55150 28040 55156
rect 27894 55040 27950 55049
rect 27894 54975 27950 54984
rect 27908 54330 27936 54975
rect 28092 54874 28120 57559
rect 28080 54868 28132 54874
rect 28080 54810 28132 54816
rect 27896 54324 27948 54330
rect 27896 54266 27948 54272
rect 27908 54126 27936 54266
rect 27896 54120 27948 54126
rect 27896 54062 27948 54068
rect 27816 53944 27936 53972
rect 27528 53644 27580 53650
rect 27528 53586 27580 53592
rect 27618 53544 27674 53553
rect 27618 53479 27674 53488
rect 27436 52624 27488 52630
rect 27436 52566 27488 52572
rect 27528 52556 27580 52562
rect 27528 52498 27580 52504
rect 27344 52012 27396 52018
rect 27344 51954 27396 51960
rect 27540 51882 27568 52498
rect 27632 52086 27660 53479
rect 27712 52148 27764 52154
rect 27712 52090 27764 52096
rect 27620 52080 27672 52086
rect 27620 52022 27672 52028
rect 27528 51876 27580 51882
rect 27528 51818 27580 51824
rect 27252 51536 27304 51542
rect 27252 51478 27304 51484
rect 27068 50856 27120 50862
rect 27068 50798 27120 50804
rect 26976 50516 27028 50522
rect 26976 50458 27028 50464
rect 26988 49842 27016 50458
rect 27080 50454 27108 50798
rect 27068 50448 27120 50454
rect 27068 50390 27120 50396
rect 27264 50386 27292 51478
rect 27528 51264 27580 51270
rect 27528 51206 27580 51212
rect 27344 50924 27396 50930
rect 27344 50866 27396 50872
rect 27252 50380 27304 50386
rect 27252 50322 27304 50328
rect 26976 49836 27028 49842
rect 26976 49778 27028 49784
rect 27264 49434 27292 50322
rect 27252 49428 27304 49434
rect 27252 49370 27304 49376
rect 27068 49224 27120 49230
rect 27068 49166 27120 49172
rect 27080 48210 27108 49166
rect 27158 49056 27214 49065
rect 27158 48991 27214 49000
rect 27172 48686 27200 48991
rect 27160 48680 27212 48686
rect 27160 48622 27212 48628
rect 27068 48204 27120 48210
rect 27068 48146 27120 48152
rect 27080 47802 27108 48146
rect 27356 48113 27384 50866
rect 27540 50726 27568 51206
rect 27620 50992 27672 50998
rect 27620 50934 27672 50940
rect 27528 50720 27580 50726
rect 27528 50662 27580 50668
rect 27528 50516 27580 50522
rect 27528 50458 27580 50464
rect 27540 49774 27568 50458
rect 27528 49768 27580 49774
rect 27632 49745 27660 50934
rect 27724 50454 27752 52090
rect 27804 50720 27856 50726
rect 27804 50662 27856 50668
rect 27712 50448 27764 50454
rect 27712 50390 27764 50396
rect 27528 49710 27580 49716
rect 27618 49736 27674 49745
rect 27618 49671 27674 49680
rect 27724 49450 27752 50390
rect 27816 50250 27844 50662
rect 27804 50244 27856 50250
rect 27804 50186 27856 50192
rect 27908 49881 27936 53944
rect 28184 53650 28212 59366
rect 28736 58070 28764 62766
rect 29090 62112 29146 62121
rect 29090 62047 29146 62056
rect 29000 59560 29052 59566
rect 29000 59502 29052 59508
rect 29012 59242 29040 59502
rect 28920 59214 29040 59242
rect 28724 58064 28776 58070
rect 28724 58006 28776 58012
rect 28448 57996 28500 58002
rect 28448 57938 28500 57944
rect 28816 57996 28868 58002
rect 28816 57938 28868 57944
rect 28356 57792 28408 57798
rect 28356 57734 28408 57740
rect 28368 57390 28396 57734
rect 28460 57458 28488 57938
rect 28540 57928 28592 57934
rect 28540 57870 28592 57876
rect 28632 57928 28684 57934
rect 28632 57870 28684 57876
rect 28448 57452 28500 57458
rect 28448 57394 28500 57400
rect 28356 57384 28408 57390
rect 28356 57326 28408 57332
rect 28264 56908 28316 56914
rect 28264 56850 28316 56856
rect 28276 56250 28304 56850
rect 28368 56370 28396 57326
rect 28460 56778 28488 57394
rect 28552 57254 28580 57870
rect 28644 57458 28672 57870
rect 28632 57452 28684 57458
rect 28632 57394 28684 57400
rect 28540 57248 28592 57254
rect 28540 57190 28592 57196
rect 28448 56772 28500 56778
rect 28448 56714 28500 56720
rect 28356 56364 28408 56370
rect 28356 56306 28408 56312
rect 28276 56222 28396 56250
rect 28368 56166 28396 56222
rect 28356 56160 28408 56166
rect 28356 56102 28408 56108
rect 28264 55820 28316 55826
rect 28264 55762 28316 55768
rect 28276 55282 28304 55762
rect 28264 55276 28316 55282
rect 28264 55218 28316 55224
rect 28172 53644 28224 53650
rect 28172 53586 28224 53592
rect 28368 53530 28396 56102
rect 28460 55842 28488 56714
rect 28552 55962 28580 57190
rect 28644 56846 28672 57394
rect 28724 57316 28776 57322
rect 28724 57258 28776 57264
rect 28632 56840 28684 56846
rect 28632 56782 28684 56788
rect 28540 55956 28592 55962
rect 28540 55898 28592 55904
rect 28460 55814 28580 55842
rect 28184 53502 28396 53530
rect 28080 51944 28132 51950
rect 28080 51886 28132 51892
rect 27988 51604 28040 51610
rect 27988 51546 28040 51552
rect 28000 50794 28028 51546
rect 28092 51066 28120 51886
rect 28080 51060 28132 51066
rect 28080 51002 28132 51008
rect 28184 50946 28212 53502
rect 28264 52488 28316 52494
rect 28264 52430 28316 52436
rect 28276 52154 28304 52430
rect 28356 52420 28408 52426
rect 28356 52362 28408 52368
rect 28264 52148 28316 52154
rect 28264 52090 28316 52096
rect 28264 51808 28316 51814
rect 28368 51796 28396 52362
rect 28316 51768 28396 51796
rect 28264 51750 28316 51756
rect 28368 51406 28396 51768
rect 28356 51400 28408 51406
rect 28356 51342 28408 51348
rect 28448 51400 28500 51406
rect 28448 51342 28500 51348
rect 28368 51066 28396 51342
rect 28460 51241 28488 51342
rect 28446 51232 28502 51241
rect 28446 51167 28502 51176
rect 28356 51060 28408 51066
rect 28356 51002 28408 51008
rect 28184 50918 28488 50946
rect 27988 50788 28040 50794
rect 27988 50730 28040 50736
rect 28172 50788 28224 50794
rect 28172 50730 28224 50736
rect 27894 49872 27950 49881
rect 27894 49807 27950 49816
rect 27908 49774 27936 49807
rect 27804 49768 27856 49774
rect 27804 49710 27856 49716
rect 27896 49768 27948 49774
rect 27896 49710 27948 49716
rect 27540 49422 27752 49450
rect 27540 49366 27568 49422
rect 27528 49360 27580 49366
rect 27528 49302 27580 49308
rect 27620 48816 27672 48822
rect 27620 48758 27672 48764
rect 27436 48544 27488 48550
rect 27436 48486 27488 48492
rect 27342 48104 27398 48113
rect 27342 48039 27398 48048
rect 27068 47796 27120 47802
rect 27068 47738 27120 47744
rect 27080 47258 27108 47738
rect 27068 47252 27120 47258
rect 27068 47194 27120 47200
rect 26884 47184 26936 47190
rect 26884 47126 26936 47132
rect 26884 47048 26936 47054
rect 26804 46996 26884 47002
rect 26804 46990 26936 46996
rect 26804 46974 26924 46990
rect 26516 46572 26568 46578
rect 26516 46514 26568 46520
rect 26424 46436 26476 46442
rect 26424 46378 26476 46384
rect 26436 45830 26464 46378
rect 26424 45824 26476 45830
rect 26424 45766 26476 45772
rect 26332 45076 26384 45082
rect 26332 45018 26384 45024
rect 26436 44334 26464 45766
rect 26528 45626 26556 46514
rect 26608 46504 26660 46510
rect 26608 46446 26660 46452
rect 26516 45620 26568 45626
rect 26516 45562 26568 45568
rect 26620 45490 26648 46446
rect 26896 46345 26924 46974
rect 27080 46510 27108 47194
rect 27158 47152 27214 47161
rect 27158 47087 27160 47096
rect 27212 47087 27214 47096
rect 27160 47058 27212 47064
rect 27172 46714 27200 47058
rect 27448 47054 27476 48486
rect 27632 48278 27660 48758
rect 27620 48272 27672 48278
rect 27620 48214 27672 48220
rect 27528 48204 27580 48210
rect 27528 48146 27580 48152
rect 27540 47530 27568 48146
rect 27724 47682 27752 49422
rect 27816 48210 27844 49710
rect 28000 49337 28028 50730
rect 28184 50522 28212 50730
rect 28356 50720 28408 50726
rect 28356 50662 28408 50668
rect 28172 50516 28224 50522
rect 28172 50458 28224 50464
rect 28078 50416 28134 50425
rect 28368 50386 28396 50662
rect 28078 50351 28134 50360
rect 28356 50380 28408 50386
rect 27986 49328 28042 49337
rect 27986 49263 28042 49272
rect 27988 49224 28040 49230
rect 27988 49166 28040 49172
rect 28000 48550 28028 49166
rect 27988 48544 28040 48550
rect 27986 48512 27988 48521
rect 28040 48512 28042 48521
rect 27986 48447 28042 48456
rect 28092 48362 28120 50351
rect 28356 50322 28408 50328
rect 28264 50312 28316 50318
rect 28264 50254 28316 50260
rect 28172 48680 28224 48686
rect 28172 48622 28224 48628
rect 27908 48334 28120 48362
rect 28184 48346 28212 48622
rect 28172 48340 28224 48346
rect 27804 48204 27856 48210
rect 27804 48146 27856 48152
rect 27632 47654 27752 47682
rect 27528 47524 27580 47530
rect 27528 47466 27580 47472
rect 27540 47122 27568 47466
rect 27528 47116 27580 47122
rect 27528 47058 27580 47064
rect 27436 47048 27488 47054
rect 27540 47025 27568 47058
rect 27436 46990 27488 46996
rect 27526 47016 27582 47025
rect 27250 46880 27306 46889
rect 27250 46815 27306 46824
rect 27160 46708 27212 46714
rect 27160 46650 27212 46656
rect 27068 46504 27120 46510
rect 27068 46446 27120 46452
rect 26882 46336 26938 46345
rect 26882 46271 26938 46280
rect 26608 45484 26660 45490
rect 26608 45426 26660 45432
rect 26516 45416 26568 45422
rect 26516 45358 26568 45364
rect 26148 44328 26200 44334
rect 26424 44328 26476 44334
rect 26148 44270 26200 44276
rect 26422 44296 26424 44305
rect 26476 44296 26478 44305
rect 26422 44231 26478 44240
rect 26330 44024 26386 44033
rect 26330 43959 26332 43968
rect 26384 43959 26386 43968
rect 26332 43930 26384 43936
rect 26344 43246 26372 43930
rect 26528 43858 26556 45358
rect 26620 44402 26648 45426
rect 26896 45422 26924 46271
rect 27264 46170 27292 46815
rect 27448 46170 27476 46990
rect 27526 46951 27582 46960
rect 27252 46164 27304 46170
rect 27436 46164 27488 46170
rect 27252 46106 27304 46112
rect 27356 46124 27436 46152
rect 27356 45422 27384 46124
rect 27632 46152 27660 47654
rect 27816 47598 27844 48146
rect 27712 47592 27764 47598
rect 27712 47534 27764 47540
rect 27804 47592 27856 47598
rect 27804 47534 27856 47540
rect 27724 47054 27752 47534
rect 27712 47048 27764 47054
rect 27712 46990 27764 46996
rect 27804 46368 27856 46374
rect 27804 46310 27856 46316
rect 27632 46124 27752 46152
rect 27436 46106 27488 46112
rect 27434 46064 27490 46073
rect 27434 45999 27490 46008
rect 27528 46028 27580 46034
rect 26792 45416 26844 45422
rect 26792 45358 26844 45364
rect 26884 45416 26936 45422
rect 26884 45358 26936 45364
rect 27344 45416 27396 45422
rect 27344 45358 27396 45364
rect 26700 44872 26752 44878
rect 26700 44814 26752 44820
rect 26712 44538 26740 44814
rect 26804 44742 26832 45358
rect 26896 44810 26924 45358
rect 27448 45082 27476 45999
rect 27528 45970 27580 45976
rect 27620 46028 27672 46034
rect 27620 45970 27672 45976
rect 27540 45937 27568 45970
rect 27526 45928 27582 45937
rect 27526 45863 27582 45872
rect 27632 45626 27660 45970
rect 27620 45620 27672 45626
rect 27620 45562 27672 45568
rect 27436 45076 27488 45082
rect 27436 45018 27488 45024
rect 27620 44940 27672 44946
rect 27620 44882 27672 44888
rect 26884 44804 26936 44810
rect 26884 44746 26936 44752
rect 26792 44736 26844 44742
rect 26792 44678 26844 44684
rect 26896 44538 26924 44746
rect 27252 44736 27304 44742
rect 27252 44678 27304 44684
rect 26700 44532 26752 44538
rect 26700 44474 26752 44480
rect 26884 44532 26936 44538
rect 26884 44474 26936 44480
rect 26608 44396 26660 44402
rect 26608 44338 26660 44344
rect 26608 43988 26660 43994
rect 26608 43930 26660 43936
rect 26516 43852 26568 43858
rect 26516 43794 26568 43800
rect 26332 43240 26384 43246
rect 26332 43182 26384 43188
rect 26528 43110 26556 43794
rect 26620 43761 26648 43930
rect 26606 43752 26662 43761
rect 26606 43687 26662 43696
rect 26516 43104 26568 43110
rect 26516 43046 26568 43052
rect 26528 42514 26556 43046
rect 26620 42838 26648 43687
rect 27158 43344 27214 43353
rect 26700 43308 26752 43314
rect 27158 43279 27214 43288
rect 26700 43250 26752 43256
rect 26608 42832 26660 42838
rect 26608 42774 26660 42780
rect 26528 42486 26648 42514
rect 26620 42022 26648 42486
rect 26712 42226 26740 43250
rect 27172 43246 27200 43279
rect 27160 43240 27212 43246
rect 27160 43182 27212 43188
rect 27068 43172 27120 43178
rect 27068 43114 27120 43120
rect 26976 42764 27028 42770
rect 26976 42706 27028 42712
rect 26988 42362 27016 42706
rect 26976 42356 27028 42362
rect 26976 42298 27028 42304
rect 26700 42220 26752 42226
rect 26700 42162 26752 42168
rect 26608 42016 26660 42022
rect 26608 41958 26660 41964
rect 26516 40044 26568 40050
rect 26516 39986 26568 39992
rect 26528 39574 26556 39986
rect 26516 39568 26568 39574
rect 26516 39510 26568 39516
rect 26528 38962 26556 39510
rect 26620 39506 26648 41958
rect 26884 39976 26936 39982
rect 26884 39918 26936 39924
rect 26608 39500 26660 39506
rect 26608 39442 26660 39448
rect 26620 39098 26648 39442
rect 26608 39092 26660 39098
rect 26608 39034 26660 39040
rect 26056 38956 26108 38962
rect 26056 38898 26108 38904
rect 26516 38956 26568 38962
rect 26516 38898 26568 38904
rect 26896 38894 26924 39918
rect 26884 38888 26936 38894
rect 26884 38830 26936 38836
rect 26974 38856 27030 38865
rect 26792 38820 26844 38826
rect 26792 38762 26844 38768
rect 26146 38720 26202 38729
rect 26146 38655 26202 38664
rect 25964 37732 26016 37738
rect 25964 37674 26016 37680
rect 25870 34776 25926 34785
rect 25870 34711 25926 34720
rect 25318 33960 25374 33969
rect 25318 33895 25374 33904
rect 25332 33386 25360 33895
rect 25594 33688 25650 33697
rect 25594 33623 25596 33632
rect 25648 33623 25650 33632
rect 25596 33594 25648 33600
rect 25504 33448 25556 33454
rect 25504 33390 25556 33396
rect 25320 33380 25372 33386
rect 25320 33322 25372 33328
rect 25332 32910 25360 33322
rect 25320 32904 25372 32910
rect 25320 32846 25372 32852
rect 25332 31278 25360 32846
rect 25320 31272 25372 31278
rect 25320 31214 25372 31220
rect 25412 31136 25464 31142
rect 25318 31104 25374 31113
rect 25412 31078 25464 31084
rect 25318 31039 25374 31048
rect 25332 30122 25360 31039
rect 25424 30705 25452 31078
rect 25516 30954 25544 33390
rect 25594 33008 25650 33017
rect 25594 32943 25650 32952
rect 25608 32570 25636 32943
rect 25596 32564 25648 32570
rect 25596 32506 25648 32512
rect 25780 32496 25832 32502
rect 25780 32438 25832 32444
rect 25688 32224 25740 32230
rect 25688 32166 25740 32172
rect 25596 31952 25648 31958
rect 25594 31920 25596 31929
rect 25648 31920 25650 31929
rect 25594 31855 25650 31864
rect 25700 31226 25728 32166
rect 25792 31754 25820 32438
rect 25780 31748 25832 31754
rect 25780 31690 25832 31696
rect 25780 31340 25832 31346
rect 25832 31300 25912 31328
rect 25780 31282 25832 31288
rect 25700 31198 25820 31226
rect 25516 30926 25636 30954
rect 25410 30696 25466 30705
rect 25410 30631 25466 30640
rect 25412 30592 25464 30598
rect 25412 30534 25464 30540
rect 25424 30410 25452 30534
rect 25424 30382 25544 30410
rect 25320 30116 25372 30122
rect 25320 30058 25372 30064
rect 25332 29782 25360 30058
rect 25516 30054 25544 30382
rect 25504 30048 25556 30054
rect 25504 29990 25556 29996
rect 25320 29776 25372 29782
rect 25320 29718 25372 29724
rect 25332 29306 25360 29718
rect 25320 29300 25372 29306
rect 25320 29242 25372 29248
rect 25320 29028 25372 29034
rect 25320 28970 25372 28976
rect 25332 27606 25360 28970
rect 25516 27962 25544 29990
rect 25608 28762 25636 30926
rect 25686 30152 25742 30161
rect 25686 30087 25742 30096
rect 25700 29850 25728 30087
rect 25688 29844 25740 29850
rect 25688 29786 25740 29792
rect 25688 29708 25740 29714
rect 25688 29650 25740 29656
rect 25596 28756 25648 28762
rect 25596 28698 25648 28704
rect 25596 28416 25648 28422
rect 25596 28358 25648 28364
rect 25608 28082 25636 28358
rect 25596 28076 25648 28082
rect 25596 28018 25648 28024
rect 25424 27934 25544 27962
rect 25320 27600 25372 27606
rect 25320 27542 25372 27548
rect 25320 27328 25372 27334
rect 25320 27270 25372 27276
rect 25332 27062 25360 27270
rect 25320 27056 25372 27062
rect 25424 27033 25452 27934
rect 25320 26998 25372 27004
rect 25410 27024 25466 27033
rect 25410 26959 25466 26968
rect 25502 26480 25558 26489
rect 25502 26415 25558 26424
rect 25516 26314 25544 26415
rect 25504 26308 25556 26314
rect 25504 26250 25556 26256
rect 25318 26072 25374 26081
rect 25318 26007 25320 26016
rect 25372 26007 25374 26016
rect 25320 25978 25372 25984
rect 25318 25528 25374 25537
rect 25318 25463 25320 25472
rect 25372 25463 25374 25472
rect 25320 25434 25372 25440
rect 25608 25362 25636 28018
rect 25700 26518 25728 29650
rect 25792 26897 25820 31198
rect 25884 30394 25912 31300
rect 25872 30388 25924 30394
rect 25872 30330 25924 30336
rect 25870 30152 25926 30161
rect 25870 30087 25872 30096
rect 25924 30087 25926 30096
rect 25872 30058 25924 30064
rect 25884 29714 25912 30058
rect 25872 29708 25924 29714
rect 25872 29650 25924 29656
rect 25872 29300 25924 29306
rect 25872 29242 25924 29248
rect 25884 28422 25912 29242
rect 25872 28416 25924 28422
rect 25872 28358 25924 28364
rect 25884 28218 25912 28358
rect 25872 28212 25924 28218
rect 25872 28154 25924 28160
rect 25884 27674 25912 28154
rect 25872 27668 25924 27674
rect 25872 27610 25924 27616
rect 25884 27130 25912 27610
rect 25872 27124 25924 27130
rect 25872 27066 25924 27072
rect 25884 26926 25912 27066
rect 25872 26920 25924 26926
rect 25778 26888 25834 26897
rect 25872 26862 25924 26868
rect 25778 26823 25834 26832
rect 25872 26784 25924 26790
rect 25872 26726 25924 26732
rect 25778 26616 25834 26625
rect 25778 26551 25834 26560
rect 25688 26512 25740 26518
rect 25688 26454 25740 26460
rect 25596 25356 25648 25362
rect 25596 25298 25648 25304
rect 25792 24818 25820 26551
rect 25884 26314 25912 26726
rect 25872 26308 25924 26314
rect 25872 26250 25924 26256
rect 25872 25832 25924 25838
rect 25870 25800 25872 25809
rect 25924 25800 25926 25809
rect 25870 25735 25926 25744
rect 25780 24812 25832 24818
rect 25240 24772 25360 24800
rect 25226 24712 25282 24721
rect 25226 24647 25282 24656
rect 25240 24614 25268 24647
rect 25228 24608 25280 24614
rect 25228 24550 25280 24556
rect 25148 24398 25268 24426
rect 25044 24336 25096 24342
rect 25044 24278 25096 24284
rect 25240 24274 25268 24398
rect 25228 24268 25280 24274
rect 25228 24210 25280 24216
rect 25044 23656 25096 23662
rect 25044 23598 25096 23604
rect 24674 23216 24730 23225
rect 24674 23151 24676 23160
rect 24728 23151 24730 23160
rect 24676 23122 24728 23128
rect 24688 22778 24716 23122
rect 24676 22772 24728 22778
rect 24676 22714 24728 22720
rect 24952 21412 25004 21418
rect 24952 21354 25004 21360
rect 24676 21344 24728 21350
rect 24676 21286 24728 21292
rect 24688 7857 24716 21286
rect 24964 20806 24992 21354
rect 24952 20800 25004 20806
rect 24952 20742 25004 20748
rect 24964 18601 24992 20742
rect 24950 18592 25006 18601
rect 24950 18527 25006 18536
rect 24768 15904 24820 15910
rect 24964 15858 24992 18527
rect 24820 15852 24992 15858
rect 24768 15846 24992 15852
rect 24780 15830 24992 15846
rect 24858 15464 24914 15473
rect 24858 15399 24914 15408
rect 24674 7848 24730 7857
rect 24674 7783 24730 7792
rect 24584 1420 24636 1426
rect 24584 1362 24636 1368
rect 24872 800 24900 15399
rect 24964 14006 24992 15830
rect 24952 14000 25004 14006
rect 24952 13942 25004 13948
rect 24964 6905 24992 13942
rect 25056 7585 25084 23598
rect 25240 22982 25268 24210
rect 25228 22976 25280 22982
rect 25228 22918 25280 22924
rect 25240 22642 25268 22918
rect 25228 22636 25280 22642
rect 25228 22578 25280 22584
rect 25228 21480 25280 21486
rect 25228 21422 25280 21428
rect 25240 21350 25268 21422
rect 25228 21344 25280 21350
rect 25228 21286 25280 21292
rect 25332 16726 25360 24772
rect 25780 24754 25832 24760
rect 25596 24132 25648 24138
rect 25596 24074 25648 24080
rect 25412 24064 25464 24070
rect 25410 24032 25412 24041
rect 25464 24032 25466 24041
rect 25410 23967 25466 23976
rect 25608 23322 25636 24074
rect 25596 23316 25648 23322
rect 25596 23258 25648 23264
rect 25320 16720 25372 16726
rect 25320 16662 25372 16668
rect 25134 13968 25190 13977
rect 25134 13903 25190 13912
rect 25148 13870 25176 13903
rect 25136 13864 25188 13870
rect 25136 13806 25188 13812
rect 25778 7712 25834 7721
rect 25778 7647 25834 7656
rect 25042 7576 25098 7585
rect 25042 7511 25098 7520
rect 24950 6896 25006 6905
rect 24950 6831 25006 6840
rect 25792 800 25820 7647
rect 25976 6361 26004 37674
rect 26054 33688 26110 33697
rect 26054 33623 26110 33632
rect 26068 31482 26096 33623
rect 26056 31476 26108 31482
rect 26056 31418 26108 31424
rect 26160 31328 26188 38655
rect 26804 37806 26832 38762
rect 26896 38554 26924 38830
rect 26974 38791 27030 38800
rect 26884 38548 26936 38554
rect 26884 38490 26936 38496
rect 26792 37800 26844 37806
rect 26792 37742 26844 37748
rect 26884 37664 26936 37670
rect 26884 37606 26936 37612
rect 26790 37496 26846 37505
rect 26790 37431 26846 37440
rect 26804 36922 26832 37431
rect 26792 36916 26844 36922
rect 26792 36858 26844 36864
rect 26700 34604 26752 34610
rect 26700 34546 26752 34552
rect 26240 34536 26292 34542
rect 26240 34478 26292 34484
rect 26252 33862 26280 34478
rect 26332 33924 26384 33930
rect 26332 33866 26384 33872
rect 26240 33856 26292 33862
rect 26240 33798 26292 33804
rect 26252 33318 26280 33798
rect 26240 33312 26292 33318
rect 26240 33254 26292 33260
rect 26252 33114 26280 33254
rect 26240 33108 26292 33114
rect 26240 33050 26292 33056
rect 26344 32570 26372 33866
rect 26332 32564 26384 32570
rect 26332 32506 26384 32512
rect 26424 32360 26476 32366
rect 26424 32302 26476 32308
rect 26240 32292 26292 32298
rect 26240 32234 26292 32240
rect 26068 31300 26188 31328
rect 26068 30954 26096 31300
rect 26252 31278 26280 32234
rect 26436 32230 26464 32302
rect 26332 32224 26384 32230
rect 26332 32166 26384 32172
rect 26424 32224 26476 32230
rect 26424 32166 26476 32172
rect 26344 32065 26372 32166
rect 26330 32056 26386 32065
rect 26330 31991 26386 32000
rect 26436 31793 26464 32166
rect 26422 31784 26478 31793
rect 26422 31719 26478 31728
rect 26240 31272 26292 31278
rect 26240 31214 26292 31220
rect 26068 30926 26188 30954
rect 26056 28960 26108 28966
rect 26056 28902 26108 28908
rect 26068 28762 26096 28902
rect 26056 28756 26108 28762
rect 26056 28698 26108 28704
rect 26054 27432 26110 27441
rect 26054 27367 26110 27376
rect 26068 27130 26096 27367
rect 26056 27124 26108 27130
rect 26056 27066 26108 27072
rect 26056 26240 26108 26246
rect 26056 26182 26108 26188
rect 26068 25838 26096 26182
rect 26056 25832 26108 25838
rect 26056 25774 26108 25780
rect 26056 25288 26108 25294
rect 26056 25230 26108 25236
rect 26068 24018 26096 25230
rect 26160 24177 26188 30926
rect 26252 30297 26280 31214
rect 26332 31204 26384 31210
rect 26332 31146 26384 31152
rect 26238 30288 26294 30297
rect 26238 30223 26294 30232
rect 26240 30048 26292 30054
rect 26240 29990 26292 29996
rect 26252 29889 26280 29990
rect 26238 29880 26294 29889
rect 26238 29815 26294 29824
rect 26344 29782 26372 31146
rect 26436 30598 26464 31719
rect 26514 31376 26570 31385
rect 26514 31311 26570 31320
rect 26424 30592 26476 30598
rect 26424 30534 26476 30540
rect 26332 29776 26384 29782
rect 26436 29753 26464 30534
rect 26332 29718 26384 29724
rect 26422 29744 26478 29753
rect 26344 29510 26372 29718
rect 26528 29714 26556 31311
rect 26606 30832 26662 30841
rect 26606 30767 26662 30776
rect 26620 30326 26648 30767
rect 26608 30320 26660 30326
rect 26608 30262 26660 30268
rect 26608 30184 26660 30190
rect 26608 30126 26660 30132
rect 26422 29679 26478 29688
rect 26516 29708 26568 29714
rect 26516 29650 26568 29656
rect 26332 29504 26384 29510
rect 26332 29446 26384 29452
rect 26528 29306 26556 29650
rect 26620 29578 26648 30126
rect 26608 29572 26660 29578
rect 26608 29514 26660 29520
rect 26516 29300 26568 29306
rect 26516 29242 26568 29248
rect 26240 29164 26292 29170
rect 26240 29106 26292 29112
rect 26252 28762 26280 29106
rect 26514 29064 26570 29073
rect 26332 29028 26384 29034
rect 26514 28999 26570 29008
rect 26332 28970 26384 28976
rect 26240 28756 26292 28762
rect 26240 28698 26292 28704
rect 26240 26784 26292 26790
rect 26240 26726 26292 26732
rect 26252 24857 26280 26726
rect 26238 24848 26294 24857
rect 26238 24783 26294 24792
rect 26146 24168 26202 24177
rect 26146 24103 26202 24112
rect 26068 23990 26280 24018
rect 26252 23866 26280 23990
rect 26240 23860 26292 23866
rect 26240 23802 26292 23808
rect 26344 14521 26372 28970
rect 26422 28520 26478 28529
rect 26528 28490 26556 28999
rect 26608 28688 26660 28694
rect 26608 28630 26660 28636
rect 26422 28455 26478 28464
rect 26516 28484 26568 28490
rect 26436 26586 26464 28455
rect 26516 28426 26568 28432
rect 26620 28218 26648 28630
rect 26608 28212 26660 28218
rect 26608 28154 26660 28160
rect 26516 27872 26568 27878
rect 26516 27814 26568 27820
rect 26424 26580 26476 26586
rect 26424 26522 26476 26528
rect 26424 25764 26476 25770
rect 26424 25706 26476 25712
rect 26436 23769 26464 25706
rect 26422 23760 26478 23769
rect 26422 23695 26478 23704
rect 26422 23352 26478 23361
rect 26422 23287 26478 23296
rect 26436 21690 26464 23287
rect 26424 21684 26476 21690
rect 26424 21626 26476 21632
rect 26330 14512 26386 14521
rect 26330 14447 26386 14456
rect 26528 7857 26556 27814
rect 26712 26926 26740 34546
rect 26804 32337 26832 36858
rect 26790 32328 26846 32337
rect 26790 32263 26846 32272
rect 26792 31884 26844 31890
rect 26792 31826 26844 31832
rect 26804 31482 26832 31826
rect 26792 31476 26844 31482
rect 26792 31418 26844 31424
rect 26792 31136 26844 31142
rect 26792 31078 26844 31084
rect 26804 29102 26832 31078
rect 26792 29096 26844 29102
rect 26792 29038 26844 29044
rect 26804 28694 26832 29038
rect 26792 28688 26844 28694
rect 26792 28630 26844 28636
rect 26792 28552 26844 28558
rect 26792 28494 26844 28500
rect 26804 28393 26832 28494
rect 26790 28384 26846 28393
rect 26790 28319 26846 28328
rect 26804 27674 26832 28319
rect 26792 27668 26844 27674
rect 26792 27610 26844 27616
rect 26700 26920 26752 26926
rect 26700 26862 26752 26868
rect 26804 26858 26832 27610
rect 26792 26852 26844 26858
rect 26792 26794 26844 26800
rect 26700 26784 26752 26790
rect 26700 26726 26752 26732
rect 26712 25906 26740 26726
rect 26790 26344 26846 26353
rect 26790 26279 26846 26288
rect 26700 25900 26752 25906
rect 26700 25842 26752 25848
rect 26804 25430 26832 26279
rect 26792 25424 26844 25430
rect 26792 25366 26844 25372
rect 26608 25356 26660 25362
rect 26608 25298 26660 25304
rect 26620 24954 26648 25298
rect 26608 24948 26660 24954
rect 26608 24890 26660 24896
rect 26620 22681 26648 24890
rect 26606 22672 26662 22681
rect 26606 22607 26662 22616
rect 26896 10577 26924 37606
rect 26988 35714 27016 38791
rect 27080 35873 27108 43114
rect 27172 41818 27200 43182
rect 27264 42770 27292 44678
rect 27528 44396 27580 44402
rect 27528 44338 27580 44344
rect 27344 44260 27396 44266
rect 27344 44202 27396 44208
rect 27356 43858 27384 44202
rect 27540 43858 27568 44338
rect 27632 44266 27660 44882
rect 27724 44810 27752 46124
rect 27816 45393 27844 46310
rect 27802 45384 27858 45393
rect 27908 45370 27936 48334
rect 28172 48282 28224 48288
rect 28170 48240 28226 48249
rect 28170 48175 28226 48184
rect 28080 48068 28132 48074
rect 28080 48010 28132 48016
rect 27988 47592 28040 47598
rect 27988 47534 28040 47540
rect 28000 45490 28028 47534
rect 28092 46374 28120 48010
rect 28184 46646 28212 48175
rect 28172 46640 28224 46646
rect 28172 46582 28224 46588
rect 28172 46504 28224 46510
rect 28172 46446 28224 46452
rect 28080 46368 28132 46374
rect 28080 46310 28132 46316
rect 28078 45928 28134 45937
rect 28078 45863 28134 45872
rect 28092 45558 28120 45863
rect 28184 45626 28212 46446
rect 28172 45620 28224 45626
rect 28172 45562 28224 45568
rect 28080 45552 28132 45558
rect 28080 45494 28132 45500
rect 27988 45484 28040 45490
rect 27988 45426 28040 45432
rect 28184 45422 28212 45562
rect 28172 45416 28224 45422
rect 27908 45342 28120 45370
rect 28172 45358 28224 45364
rect 27802 45319 27858 45328
rect 27988 45280 28040 45286
rect 27988 45222 28040 45228
rect 28092 45234 28120 45342
rect 27712 44804 27764 44810
rect 27712 44746 27764 44752
rect 27804 44736 27856 44742
rect 27804 44678 27856 44684
rect 27712 44396 27764 44402
rect 27712 44338 27764 44344
rect 27620 44260 27672 44266
rect 27620 44202 27672 44208
rect 27344 43852 27396 43858
rect 27344 43794 27396 43800
rect 27528 43852 27580 43858
rect 27528 43794 27580 43800
rect 27356 42906 27384 43794
rect 27436 43716 27488 43722
rect 27436 43658 27488 43664
rect 27448 43314 27476 43658
rect 27436 43308 27488 43314
rect 27436 43250 27488 43256
rect 27344 42900 27396 42906
rect 27344 42842 27396 42848
rect 27632 42770 27660 44202
rect 27252 42764 27304 42770
rect 27252 42706 27304 42712
rect 27620 42764 27672 42770
rect 27620 42706 27672 42712
rect 27528 42696 27580 42702
rect 27528 42638 27580 42644
rect 27540 42378 27568 42638
rect 27724 42378 27752 44338
rect 27540 42362 27752 42378
rect 27528 42356 27752 42362
rect 27580 42350 27752 42356
rect 27528 42298 27580 42304
rect 27540 42242 27568 42298
rect 27448 42214 27568 42242
rect 27160 41812 27212 41818
rect 27160 41754 27212 41760
rect 27252 41608 27304 41614
rect 27252 41550 27304 41556
rect 27264 41449 27292 41550
rect 27250 41440 27306 41449
rect 27250 41375 27306 41384
rect 27252 39024 27304 39030
rect 27252 38966 27304 38972
rect 27160 38956 27212 38962
rect 27160 38898 27212 38904
rect 27172 38554 27200 38898
rect 27160 38548 27212 38554
rect 27160 38490 27212 38496
rect 27264 37874 27292 38966
rect 27252 37868 27304 37874
rect 27252 37810 27304 37816
rect 27264 37466 27292 37810
rect 27252 37460 27304 37466
rect 27252 37402 27304 37408
rect 27448 37330 27476 42214
rect 27526 41712 27582 41721
rect 27526 41647 27582 41656
rect 27540 41614 27568 41647
rect 27528 41608 27580 41614
rect 27528 41550 27580 41556
rect 27540 41274 27568 41550
rect 27710 41440 27766 41449
rect 27710 41375 27766 41384
rect 27724 41274 27752 41375
rect 27528 41268 27580 41274
rect 27528 41210 27580 41216
rect 27712 41268 27764 41274
rect 27712 41210 27764 41216
rect 27712 38208 27764 38214
rect 27712 38150 27764 38156
rect 27724 37806 27752 38150
rect 27712 37800 27764 37806
rect 27712 37742 27764 37748
rect 27436 37324 27488 37330
rect 27436 37266 27488 37272
rect 27448 36922 27476 37266
rect 27436 36916 27488 36922
rect 27436 36858 27488 36864
rect 27448 36417 27476 36858
rect 27434 36408 27490 36417
rect 27434 36343 27490 36352
rect 27066 35864 27122 35873
rect 27066 35799 27122 35808
rect 26988 35686 27108 35714
rect 26974 32328 27030 32337
rect 26974 32263 27030 32272
rect 26988 31482 27016 32263
rect 26976 31476 27028 31482
rect 26976 31418 27028 31424
rect 26976 29776 27028 29782
rect 26976 29718 27028 29724
rect 26988 29510 27016 29718
rect 26976 29504 27028 29510
rect 26974 29472 26976 29481
rect 27028 29472 27030 29481
rect 26974 29407 27030 29416
rect 26988 29381 27016 29407
rect 27080 29238 27108 35686
rect 27618 34232 27674 34241
rect 27618 34167 27674 34176
rect 27632 34066 27660 34167
rect 27620 34060 27672 34066
rect 27620 34002 27672 34008
rect 27434 33824 27490 33833
rect 27434 33759 27490 33768
rect 27344 32972 27396 32978
rect 27344 32914 27396 32920
rect 27160 32360 27212 32366
rect 27160 32302 27212 32308
rect 27172 31657 27200 32302
rect 27356 31822 27384 32914
rect 27344 31816 27396 31822
rect 27344 31758 27396 31764
rect 27158 31648 27214 31657
rect 27158 31583 27214 31592
rect 27250 31376 27306 31385
rect 27250 31311 27306 31320
rect 27264 31278 27292 31311
rect 27252 31272 27304 31278
rect 27252 31214 27304 31220
rect 27356 30734 27384 31758
rect 27448 31482 27476 33759
rect 27632 33658 27660 34002
rect 27712 33856 27764 33862
rect 27712 33798 27764 33804
rect 27620 33652 27672 33658
rect 27620 33594 27672 33600
rect 27724 32026 27752 33798
rect 27712 32020 27764 32026
rect 27712 31962 27764 31968
rect 27620 31816 27672 31822
rect 27620 31758 27672 31764
rect 27526 31648 27582 31657
rect 27526 31583 27582 31592
rect 27436 31476 27488 31482
rect 27436 31418 27488 31424
rect 27540 30818 27568 31583
rect 27448 30790 27568 30818
rect 27344 30728 27396 30734
rect 27344 30670 27396 30676
rect 27344 30116 27396 30122
rect 27344 30058 27396 30064
rect 27250 30016 27306 30025
rect 27250 29951 27306 29960
rect 27264 29782 27292 29951
rect 27252 29776 27304 29782
rect 27252 29718 27304 29724
rect 27252 29572 27304 29578
rect 27252 29514 27304 29520
rect 27068 29232 27120 29238
rect 27068 29174 27120 29180
rect 27160 28416 27212 28422
rect 27160 28358 27212 28364
rect 27068 28076 27120 28082
rect 27068 28018 27120 28024
rect 27080 27674 27108 28018
rect 27068 27668 27120 27674
rect 27068 27610 27120 27616
rect 27068 27532 27120 27538
rect 27068 27474 27120 27480
rect 27080 27130 27108 27474
rect 27068 27124 27120 27130
rect 27068 27066 27120 27072
rect 27068 26920 27120 26926
rect 27068 26862 27120 26868
rect 26976 26376 27028 26382
rect 26976 26318 27028 26324
rect 26988 26042 27016 26318
rect 26976 26036 27028 26042
rect 26976 25978 27028 25984
rect 27080 17921 27108 26862
rect 27172 21457 27200 28358
rect 27264 26874 27292 29514
rect 27356 28762 27384 30058
rect 27448 29152 27476 30790
rect 27528 30728 27580 30734
rect 27632 30716 27660 31758
rect 27712 31680 27764 31686
rect 27712 31622 27764 31628
rect 27580 30688 27660 30716
rect 27528 30670 27580 30676
rect 27528 30388 27580 30394
rect 27528 30330 27580 30336
rect 27540 29730 27568 30330
rect 27632 30326 27660 30688
rect 27620 30320 27672 30326
rect 27620 30262 27672 30268
rect 27724 29850 27752 31622
rect 27712 29844 27764 29850
rect 27712 29786 27764 29792
rect 27540 29702 27752 29730
rect 27620 29640 27672 29646
rect 27620 29582 27672 29588
rect 27448 29124 27568 29152
rect 27436 29028 27488 29034
rect 27436 28970 27488 28976
rect 27344 28756 27396 28762
rect 27344 28698 27396 28704
rect 27344 28484 27396 28490
rect 27344 28426 27396 28432
rect 27356 27606 27384 28426
rect 27448 28218 27476 28970
rect 27436 28212 27488 28218
rect 27436 28154 27488 28160
rect 27344 27600 27396 27606
rect 27344 27542 27396 27548
rect 27264 26846 27384 26874
rect 27252 26784 27304 26790
rect 27252 26726 27304 26732
rect 27264 25702 27292 26726
rect 27252 25696 27304 25702
rect 27252 25638 27304 25644
rect 27356 25498 27384 26846
rect 27540 26568 27568 29124
rect 27632 28490 27660 29582
rect 27724 28762 27752 29702
rect 27712 28756 27764 28762
rect 27712 28698 27764 28704
rect 27620 28484 27672 28490
rect 27620 28426 27672 28432
rect 27816 27441 27844 44678
rect 27894 44568 27950 44577
rect 27894 44503 27950 44512
rect 27908 44470 27936 44503
rect 28000 44470 28028 45222
rect 28092 45206 28212 45234
rect 28080 44804 28132 44810
rect 28080 44746 28132 44752
rect 27896 44464 27948 44470
rect 27896 44406 27948 44412
rect 27988 44464 28040 44470
rect 27988 44406 28040 44412
rect 27908 43450 27936 44406
rect 28000 43994 28028 44406
rect 27988 43988 28040 43994
rect 27988 43930 28040 43936
rect 27988 43852 28040 43858
rect 27988 43794 28040 43800
rect 27896 43444 27948 43450
rect 27896 43386 27948 43392
rect 28000 42294 28028 43794
rect 28092 43450 28120 44746
rect 28080 43444 28132 43450
rect 28080 43386 28132 43392
rect 28184 43194 28212 45206
rect 28276 43330 28304 50254
rect 28368 49978 28396 50322
rect 28356 49972 28408 49978
rect 28356 49914 28408 49920
rect 28460 49858 28488 50918
rect 28552 50425 28580 55814
rect 28736 50930 28764 57258
rect 28828 54670 28856 57938
rect 28920 56982 28948 59214
rect 29104 59158 29132 62047
rect 29274 61160 29330 61169
rect 29274 61095 29330 61104
rect 29184 60172 29236 60178
rect 29184 60114 29236 60120
rect 29196 59430 29224 60114
rect 29184 59424 29236 59430
rect 29184 59366 29236 59372
rect 29092 59152 29144 59158
rect 29092 59094 29144 59100
rect 29000 59016 29052 59022
rect 29000 58958 29052 58964
rect 29012 58478 29040 58958
rect 29000 58472 29052 58478
rect 29000 58414 29052 58420
rect 28998 57624 29054 57633
rect 28998 57559 29000 57568
rect 29052 57559 29054 57568
rect 29000 57530 29052 57536
rect 29012 57390 29040 57530
rect 29000 57384 29052 57390
rect 29000 57326 29052 57332
rect 28908 56976 28960 56982
rect 28908 56918 28960 56924
rect 28908 56772 28960 56778
rect 28908 56714 28960 56720
rect 28816 54664 28868 54670
rect 28816 54606 28868 54612
rect 28828 54330 28856 54606
rect 28816 54324 28868 54330
rect 28816 54266 28868 54272
rect 28920 54097 28948 56714
rect 29000 54732 29052 54738
rect 29000 54674 29052 54680
rect 29012 54330 29040 54674
rect 29092 54528 29144 54534
rect 29092 54470 29144 54476
rect 29000 54324 29052 54330
rect 29000 54266 29052 54272
rect 28906 54088 28962 54097
rect 28906 54023 28962 54032
rect 28998 53408 29054 53417
rect 28998 53343 29054 53352
rect 29012 51814 29040 53343
rect 29104 52698 29132 54470
rect 29196 52737 29224 59366
rect 29182 52728 29238 52737
rect 29092 52692 29144 52698
rect 29182 52663 29238 52672
rect 29092 52634 29144 52640
rect 29092 51944 29144 51950
rect 29092 51886 29144 51892
rect 29000 51808 29052 51814
rect 29000 51750 29052 51756
rect 29104 51542 29132 51886
rect 29092 51536 29144 51542
rect 29092 51478 29144 51484
rect 28908 51264 28960 51270
rect 28908 51206 28960 51212
rect 28724 50924 28776 50930
rect 28724 50866 28776 50872
rect 28538 50416 28594 50425
rect 28538 50351 28594 50360
rect 28540 50244 28592 50250
rect 28540 50186 28592 50192
rect 28368 49830 28488 49858
rect 28368 47705 28396 49830
rect 28552 48550 28580 50186
rect 28632 49768 28684 49774
rect 28632 49710 28684 49716
rect 28540 48544 28592 48550
rect 28540 48486 28592 48492
rect 28448 48272 28500 48278
rect 28448 48214 28500 48220
rect 28354 47696 28410 47705
rect 28354 47631 28410 47640
rect 28368 47025 28396 47631
rect 28460 47258 28488 48214
rect 28540 48204 28592 48210
rect 28540 48146 28592 48152
rect 28552 47462 28580 48146
rect 28540 47456 28592 47462
rect 28540 47398 28592 47404
rect 28448 47252 28500 47258
rect 28448 47194 28500 47200
rect 28552 47190 28580 47398
rect 28540 47184 28592 47190
rect 28540 47126 28592 47132
rect 28354 47016 28410 47025
rect 28644 47002 28672 49710
rect 28736 49298 28764 50866
rect 28920 50182 28948 51206
rect 29000 50720 29052 50726
rect 28998 50688 29000 50697
rect 29052 50688 29054 50697
rect 28998 50623 29054 50632
rect 29104 50538 29132 51478
rect 29288 51241 29316 61095
rect 29274 51232 29330 51241
rect 29274 51167 29330 51176
rect 29012 50510 29132 50538
rect 28908 50176 28960 50182
rect 28908 50118 28960 50124
rect 28814 49600 28870 49609
rect 28814 49535 28870 49544
rect 28828 49298 28856 49535
rect 28724 49292 28776 49298
rect 28724 49234 28776 49240
rect 28816 49292 28868 49298
rect 28816 49234 28868 49240
rect 28736 48890 28764 49234
rect 28724 48884 28776 48890
rect 28724 48826 28776 48832
rect 28816 48544 28868 48550
rect 28816 48486 28868 48492
rect 28724 48340 28776 48346
rect 28724 48282 28776 48288
rect 28354 46951 28410 46960
rect 28460 46974 28672 47002
rect 28354 46064 28410 46073
rect 28354 45999 28356 46008
rect 28408 45999 28410 46008
rect 28356 45970 28408 45976
rect 28460 45286 28488 46974
rect 28632 46640 28684 46646
rect 28632 46582 28684 46588
rect 28644 46170 28672 46582
rect 28632 46164 28684 46170
rect 28632 46106 28684 46112
rect 28540 46096 28592 46102
rect 28540 46038 28592 46044
rect 28448 45280 28500 45286
rect 28448 45222 28500 45228
rect 28356 45076 28408 45082
rect 28356 45018 28408 45024
rect 28368 43858 28396 45018
rect 28356 43852 28408 43858
rect 28356 43794 28408 43800
rect 28368 43450 28396 43794
rect 28356 43444 28408 43450
rect 28356 43386 28408 43392
rect 28276 43302 28396 43330
rect 28184 43166 28304 43194
rect 28078 42392 28134 42401
rect 28078 42327 28080 42336
rect 28132 42327 28134 42336
rect 28080 42298 28132 42304
rect 27988 42288 28040 42294
rect 27988 42230 28040 42236
rect 28092 42158 28120 42298
rect 28080 42152 28132 42158
rect 28000 42100 28080 42106
rect 28000 42094 28132 42100
rect 28000 42078 28120 42094
rect 28172 42084 28224 42090
rect 27896 35080 27948 35086
rect 27896 35022 27948 35028
rect 27908 29850 27936 35022
rect 27896 29844 27948 29850
rect 27896 29786 27948 29792
rect 27896 29708 27948 29714
rect 27896 29650 27948 29656
rect 27908 29238 27936 29650
rect 27896 29232 27948 29238
rect 27896 29174 27948 29180
rect 27802 27432 27858 27441
rect 27802 27367 27858 27376
rect 27804 27328 27856 27334
rect 27802 27296 27804 27305
rect 27856 27296 27858 27305
rect 27802 27231 27858 27240
rect 27448 26540 27568 26568
rect 27344 25492 27396 25498
rect 27344 25434 27396 25440
rect 27448 23089 27476 26540
rect 27528 26444 27580 26450
rect 27528 26386 27580 26392
rect 27540 26194 27568 26386
rect 27620 26376 27672 26382
rect 27618 26344 27620 26353
rect 27672 26344 27674 26353
rect 27618 26279 27674 26288
rect 27540 26166 27660 26194
rect 27632 26042 27660 26166
rect 27620 26036 27672 26042
rect 27620 25978 27672 25984
rect 27434 23080 27490 23089
rect 27434 23015 27490 23024
rect 27158 21448 27214 21457
rect 27158 21383 27214 21392
rect 27066 17912 27122 17921
rect 27066 17847 27122 17856
rect 26882 10568 26938 10577
rect 26882 10503 26938 10512
rect 26514 7848 26570 7857
rect 26514 7783 26570 7792
rect 26698 7576 26754 7585
rect 26698 7511 26754 7520
rect 26146 6896 26202 6905
rect 26146 6831 26202 6840
rect 25962 6352 26018 6361
rect 25962 6287 26018 6296
rect 26160 5681 26188 6831
rect 26146 5672 26202 5681
rect 26146 5607 26202 5616
rect 26160 5522 26188 5607
rect 26160 5494 26280 5522
rect 26252 2938 26280 5494
rect 26160 2910 26280 2938
rect 26160 2446 26188 2910
rect 26148 2440 26200 2446
rect 26148 2382 26200 2388
rect 26712 800 26740 7511
rect 28000 6225 28028 42078
rect 28172 42026 28224 42032
rect 28080 42016 28132 42022
rect 28080 41958 28132 41964
rect 28092 38894 28120 41958
rect 28080 38888 28132 38894
rect 28080 38830 28132 38836
rect 28078 38448 28134 38457
rect 28078 38383 28080 38392
rect 28132 38383 28134 38392
rect 28080 38354 28132 38360
rect 28092 38010 28120 38354
rect 28080 38004 28132 38010
rect 28080 37946 28132 37952
rect 28078 36816 28134 36825
rect 28078 36751 28134 36760
rect 28092 32065 28120 36751
rect 28184 34746 28212 42026
rect 28276 42022 28304 43166
rect 28264 42016 28316 42022
rect 28264 41958 28316 41964
rect 28262 41848 28318 41857
rect 28262 41783 28318 41792
rect 28276 40089 28304 41783
rect 28368 41177 28396 43302
rect 28354 41168 28410 41177
rect 28354 41103 28410 41112
rect 28460 40390 28488 45222
rect 28552 45082 28580 46038
rect 28540 45076 28592 45082
rect 28540 45018 28592 45024
rect 28538 44976 28594 44985
rect 28538 44911 28540 44920
rect 28592 44911 28594 44920
rect 28540 44882 28592 44888
rect 28552 42702 28580 44882
rect 28632 44872 28684 44878
rect 28630 44840 28632 44849
rect 28684 44840 28686 44849
rect 28630 44775 28686 44784
rect 28644 44538 28672 44775
rect 28632 44532 28684 44538
rect 28632 44474 28684 44480
rect 28736 44033 28764 48282
rect 28828 48249 28856 48486
rect 28814 48240 28870 48249
rect 28814 48175 28870 48184
rect 28920 48074 28948 50118
rect 29012 48929 29040 50510
rect 29092 50380 29144 50386
rect 29092 50322 29144 50328
rect 29104 49774 29132 50322
rect 29276 50176 29328 50182
rect 29276 50118 29328 50124
rect 29288 49774 29316 50118
rect 29092 49768 29144 49774
rect 29092 49710 29144 49716
rect 29276 49768 29328 49774
rect 29276 49710 29328 49716
rect 29090 49464 29146 49473
rect 29090 49399 29146 49408
rect 28998 48920 29054 48929
rect 28998 48855 29054 48864
rect 29104 48074 29132 49399
rect 29288 49366 29316 49710
rect 29276 49360 29328 49366
rect 29276 49302 29328 49308
rect 29276 48544 29328 48550
rect 29276 48486 29328 48492
rect 28908 48068 28960 48074
rect 28908 48010 28960 48016
rect 29092 48068 29144 48074
rect 29092 48010 29144 48016
rect 29000 48000 29052 48006
rect 29000 47942 29052 47948
rect 29012 47122 29040 47942
rect 29090 47832 29146 47841
rect 29090 47767 29092 47776
rect 29144 47767 29146 47776
rect 29092 47738 29144 47744
rect 29104 47598 29132 47738
rect 29288 47734 29316 48486
rect 29276 47728 29328 47734
rect 29276 47670 29328 47676
rect 29092 47592 29144 47598
rect 29092 47534 29144 47540
rect 29380 47462 29408 74598
rect 29932 71641 29960 79200
rect 30380 76288 30432 76294
rect 30380 76230 30432 76236
rect 30392 75410 30420 76230
rect 30380 75404 30432 75410
rect 30380 75346 30432 75352
rect 30392 75002 30420 75346
rect 30656 75336 30708 75342
rect 30656 75278 30708 75284
rect 30380 74996 30432 75002
rect 30380 74938 30432 74944
rect 30668 74662 30696 75278
rect 30852 74746 30880 79200
rect 31772 75041 31800 79200
rect 32232 77178 32260 79200
rect 32220 77172 32272 77178
rect 32220 77114 32272 77120
rect 31758 75032 31814 75041
rect 31758 74967 31814 74976
rect 33152 74746 33180 79200
rect 33508 77716 33560 77722
rect 33508 77658 33560 77664
rect 30852 74718 31340 74746
rect 33152 74718 33272 74746
rect 30656 74656 30708 74662
rect 30656 74598 30708 74604
rect 29918 71632 29974 71641
rect 29918 71567 29974 71576
rect 30378 70136 30434 70145
rect 30378 70071 30434 70080
rect 30392 64682 30420 70071
rect 30024 64654 30420 64682
rect 29918 60616 29974 60625
rect 29918 60551 29974 60560
rect 29550 60344 29606 60353
rect 29550 60279 29552 60288
rect 29604 60279 29606 60288
rect 29552 60250 29604 60256
rect 29932 59974 29960 60551
rect 29920 59968 29972 59974
rect 29920 59910 29972 59916
rect 29932 59430 29960 59910
rect 29920 59424 29972 59430
rect 29826 59392 29882 59401
rect 29920 59366 29972 59372
rect 29826 59327 29882 59336
rect 29840 59090 29868 59327
rect 29828 59084 29880 59090
rect 29828 59026 29880 59032
rect 29736 59016 29788 59022
rect 29736 58958 29788 58964
rect 29748 58342 29776 58958
rect 29736 58336 29788 58342
rect 29736 58278 29788 58284
rect 29748 56409 29776 58278
rect 29840 58138 29868 59026
rect 29828 58132 29880 58138
rect 29828 58074 29880 58080
rect 29932 58018 29960 59366
rect 29840 57990 29960 58018
rect 29734 56400 29790 56409
rect 29734 56335 29790 56344
rect 29552 54324 29604 54330
rect 29552 54266 29604 54272
rect 29564 53242 29592 54266
rect 29552 53236 29604 53242
rect 29552 53178 29604 53184
rect 29458 52592 29514 52601
rect 29564 52562 29592 53178
rect 29642 52864 29698 52873
rect 29642 52799 29698 52808
rect 29458 52527 29460 52536
rect 29512 52527 29514 52536
rect 29552 52556 29604 52562
rect 29460 52498 29512 52504
rect 29552 52498 29604 52504
rect 29472 52154 29500 52498
rect 29550 52456 29606 52465
rect 29550 52391 29606 52400
rect 29460 52148 29512 52154
rect 29460 52090 29512 52096
rect 29564 51474 29592 52391
rect 29552 51468 29604 51474
rect 29552 51410 29604 51416
rect 29564 51270 29592 51410
rect 29552 51264 29604 51270
rect 29552 51206 29604 51212
rect 29460 50720 29512 50726
rect 29460 50662 29512 50668
rect 29472 49314 29500 50662
rect 29552 50312 29604 50318
rect 29552 50254 29604 50260
rect 29564 49978 29592 50254
rect 29552 49972 29604 49978
rect 29552 49914 29604 49920
rect 29472 49286 29592 49314
rect 29460 49224 29512 49230
rect 29460 49166 29512 49172
rect 29472 48754 29500 49166
rect 29460 48748 29512 48754
rect 29460 48690 29512 48696
rect 29472 48346 29500 48690
rect 29460 48340 29512 48346
rect 29460 48282 29512 48288
rect 29564 48210 29592 49286
rect 29656 48249 29684 52799
rect 29748 50726 29776 56335
rect 29736 50720 29788 50726
rect 29736 50662 29788 50668
rect 29736 50312 29788 50318
rect 29736 50254 29788 50260
rect 29748 49745 29776 50254
rect 29840 49910 29868 57990
rect 30024 57934 30052 64654
rect 30472 60308 30524 60314
rect 30472 60250 30524 60256
rect 30378 60072 30434 60081
rect 30378 60007 30434 60016
rect 30392 59634 30420 60007
rect 30380 59628 30432 59634
rect 30380 59570 30432 59576
rect 30012 57928 30064 57934
rect 30012 57870 30064 57876
rect 30484 54346 30512 60250
rect 30564 57928 30616 57934
rect 30564 57870 30616 57876
rect 30300 54330 30512 54346
rect 30288 54324 30512 54330
rect 30340 54318 30512 54324
rect 30288 54266 30340 54272
rect 30288 52488 30340 52494
rect 30288 52430 30340 52436
rect 30300 51950 30328 52430
rect 30576 52136 30604 57870
rect 30668 56545 30696 74598
rect 31022 74216 31078 74225
rect 31022 74151 31078 74160
rect 31036 62121 31064 74151
rect 31206 62656 31262 62665
rect 31206 62591 31262 62600
rect 31022 62112 31078 62121
rect 31022 62047 31078 62056
rect 31220 60722 31248 62591
rect 31208 60716 31260 60722
rect 31208 60658 31260 60664
rect 30932 60648 30984 60654
rect 30932 60590 30984 60596
rect 30944 60314 30972 60590
rect 30932 60308 30984 60314
rect 30932 60250 30984 60256
rect 30654 56536 30710 56545
rect 30654 56471 30710 56480
rect 30748 52488 30800 52494
rect 30748 52430 30800 52436
rect 30484 52108 30604 52136
rect 30288 51944 30340 51950
rect 30288 51886 30340 51892
rect 30300 51610 30328 51886
rect 30288 51604 30340 51610
rect 30288 51546 30340 51552
rect 30196 51468 30248 51474
rect 30484 51456 30512 52108
rect 30562 52048 30618 52057
rect 30562 51983 30564 51992
rect 30616 51983 30618 51992
rect 30564 51954 30616 51960
rect 30656 51604 30708 51610
rect 30656 51546 30708 51552
rect 30484 51428 30604 51456
rect 30196 51410 30248 51416
rect 30104 51264 30156 51270
rect 30104 51206 30156 51212
rect 30116 51105 30144 51206
rect 30102 51096 30158 51105
rect 30208 51066 30236 51410
rect 30300 51338 30512 51354
rect 30288 51332 30512 51338
rect 30340 51326 30512 51332
rect 30288 51274 30340 51280
rect 30380 51264 30432 51270
rect 30380 51206 30432 51212
rect 30102 51031 30158 51040
rect 30196 51060 30248 51066
rect 30196 51002 30248 51008
rect 30012 50924 30064 50930
rect 30012 50866 30064 50872
rect 29828 49904 29880 49910
rect 29828 49846 29880 49852
rect 29828 49768 29880 49774
rect 29734 49736 29790 49745
rect 29828 49710 29880 49716
rect 29734 49671 29790 49680
rect 29748 49434 29776 49671
rect 29736 49428 29788 49434
rect 29736 49370 29788 49376
rect 29840 48686 29868 49710
rect 29920 49292 29972 49298
rect 29920 49234 29972 49240
rect 29932 49065 29960 49234
rect 29918 49056 29974 49065
rect 29918 48991 29974 49000
rect 29932 48890 29960 48991
rect 29920 48884 29972 48890
rect 29920 48826 29972 48832
rect 29828 48680 29880 48686
rect 29828 48622 29880 48628
rect 29840 48346 29868 48622
rect 29828 48340 29880 48346
rect 29828 48282 29880 48288
rect 29642 48240 29698 48249
rect 29552 48204 29604 48210
rect 29642 48175 29698 48184
rect 29918 48240 29974 48249
rect 29918 48175 29920 48184
rect 29552 48146 29604 48152
rect 29972 48175 29974 48184
rect 29920 48146 29972 48152
rect 29734 48104 29790 48113
rect 29460 48068 29512 48074
rect 29644 48068 29696 48074
rect 29512 48028 29592 48056
rect 29460 48010 29512 48016
rect 29458 47968 29514 47977
rect 29458 47903 29514 47912
rect 29368 47456 29420 47462
rect 29368 47398 29420 47404
rect 29000 47116 29052 47122
rect 29000 47058 29052 47064
rect 29276 47116 29328 47122
rect 29276 47058 29328 47064
rect 28908 47048 28960 47054
rect 29012 47025 29040 47058
rect 29092 47048 29144 47054
rect 28908 46990 28960 46996
rect 28998 47016 29054 47025
rect 28816 46980 28868 46986
rect 28816 46922 28868 46928
rect 28722 44024 28778 44033
rect 28722 43959 28778 43968
rect 28632 43784 28684 43790
rect 28632 43726 28684 43732
rect 28540 42696 28592 42702
rect 28540 42638 28592 42644
rect 28448 40384 28500 40390
rect 28448 40326 28500 40332
rect 28262 40080 28318 40089
rect 28262 40015 28318 40024
rect 28356 38344 28408 38350
rect 28356 38286 28408 38292
rect 28368 38010 28396 38286
rect 28356 38004 28408 38010
rect 28356 37946 28408 37952
rect 28460 37890 28488 40326
rect 28368 37862 28488 37890
rect 28264 36236 28316 36242
rect 28264 36178 28316 36184
rect 28276 35834 28304 36178
rect 28264 35828 28316 35834
rect 28264 35770 28316 35776
rect 28172 34740 28224 34746
rect 28172 34682 28224 34688
rect 28276 34542 28304 35770
rect 28264 34536 28316 34542
rect 28264 34478 28316 34484
rect 28276 33998 28304 34478
rect 28264 33992 28316 33998
rect 28264 33934 28316 33940
rect 28276 33658 28304 33934
rect 28264 33652 28316 33658
rect 28264 33594 28316 33600
rect 28276 32978 28304 33594
rect 28264 32972 28316 32978
rect 28264 32914 28316 32920
rect 28172 32836 28224 32842
rect 28172 32778 28224 32784
rect 28078 32056 28134 32065
rect 28078 31991 28134 32000
rect 28080 31952 28132 31958
rect 28080 31894 28132 31900
rect 28092 31482 28120 31894
rect 28080 31476 28132 31482
rect 28080 31418 28132 31424
rect 28184 30598 28212 32778
rect 28172 30592 28224 30598
rect 28172 30534 28224 30540
rect 28078 30152 28134 30161
rect 28078 30087 28080 30096
rect 28132 30087 28134 30096
rect 28080 30058 28132 30064
rect 28170 29608 28226 29617
rect 28170 29543 28226 29552
rect 28184 29238 28212 29543
rect 28264 29504 28316 29510
rect 28264 29446 28316 29452
rect 28172 29232 28224 29238
rect 28172 29174 28224 29180
rect 28080 29096 28132 29102
rect 28080 29038 28132 29044
rect 28092 28665 28120 29038
rect 28078 28656 28134 28665
rect 28078 28591 28134 28600
rect 28172 28620 28224 28626
rect 28172 28562 28224 28568
rect 28184 28218 28212 28562
rect 28172 28212 28224 28218
rect 28172 28154 28224 28160
rect 28184 28121 28212 28154
rect 28170 28112 28226 28121
rect 28170 28047 28226 28056
rect 28276 27538 28304 29446
rect 28368 29306 28396 37862
rect 28448 36168 28500 36174
rect 28448 36110 28500 36116
rect 28460 35562 28488 36110
rect 28538 35864 28594 35873
rect 28538 35799 28594 35808
rect 28448 35556 28500 35562
rect 28448 35498 28500 35504
rect 28448 32972 28500 32978
rect 28448 32914 28500 32920
rect 28460 32570 28488 32914
rect 28448 32564 28500 32570
rect 28448 32506 28500 32512
rect 28448 31340 28500 31346
rect 28448 31282 28500 31288
rect 28356 29300 28408 29306
rect 28356 29242 28408 29248
rect 28080 27532 28132 27538
rect 28080 27474 28132 27480
rect 28264 27532 28316 27538
rect 28264 27474 28316 27480
rect 28092 26926 28120 27474
rect 28354 27160 28410 27169
rect 28354 27095 28356 27104
rect 28408 27095 28410 27104
rect 28356 27066 28408 27072
rect 28080 26920 28132 26926
rect 28078 26888 28080 26897
rect 28132 26888 28134 26897
rect 28078 26823 28134 26832
rect 28460 26625 28488 31282
rect 28552 30841 28580 35799
rect 28538 30832 28594 30841
rect 28538 30767 28594 30776
rect 28540 30592 28592 30598
rect 28540 30534 28592 30540
rect 28552 28422 28580 30534
rect 28540 28416 28592 28422
rect 28540 28358 28592 28364
rect 28446 26616 28502 26625
rect 28446 26551 28448 26560
rect 28500 26551 28502 26560
rect 28448 26522 28500 26528
rect 28460 26491 28488 26522
rect 28552 26489 28580 28358
rect 28538 26480 28594 26489
rect 28538 26415 28594 26424
rect 28644 15881 28672 43726
rect 28724 42696 28776 42702
rect 28722 42664 28724 42673
rect 28776 42664 28778 42673
rect 28722 42599 28778 42608
rect 28722 40216 28778 40225
rect 28722 40151 28778 40160
rect 28736 31958 28764 40151
rect 28828 37233 28856 46922
rect 28920 46866 28948 46990
rect 29092 46990 29144 46996
rect 28998 46951 29054 46960
rect 28920 46838 29040 46866
rect 28908 46368 28960 46374
rect 28906 46336 28908 46345
rect 28960 46336 28962 46345
rect 28906 46271 28962 46280
rect 29012 45490 29040 46838
rect 29104 46714 29132 46990
rect 29092 46708 29144 46714
rect 29092 46650 29144 46656
rect 29104 46034 29132 46650
rect 29182 46608 29238 46617
rect 29182 46543 29238 46552
rect 29196 46102 29224 46543
rect 29288 46345 29316 47058
rect 29274 46336 29330 46345
rect 29274 46271 29330 46280
rect 29276 46164 29328 46170
rect 29276 46106 29328 46112
rect 29184 46096 29236 46102
rect 29184 46038 29236 46044
rect 29092 46028 29144 46034
rect 29092 45970 29144 45976
rect 29104 45665 29132 45970
rect 29090 45656 29146 45665
rect 29090 45591 29146 45600
rect 29104 45558 29132 45591
rect 29092 45552 29144 45558
rect 29092 45494 29144 45500
rect 29000 45484 29052 45490
rect 29000 45426 29052 45432
rect 28908 45416 28960 45422
rect 28908 45358 28960 45364
rect 28920 44538 28948 45358
rect 29196 45286 29224 46038
rect 29288 45354 29316 46106
rect 29276 45348 29328 45354
rect 29276 45290 29328 45296
rect 29184 45280 29236 45286
rect 29184 45222 29236 45228
rect 29090 44704 29146 44713
rect 29090 44639 29146 44648
rect 28908 44532 28960 44538
rect 28908 44474 28960 44480
rect 29104 44334 29132 44639
rect 28908 44328 28960 44334
rect 28908 44270 28960 44276
rect 29092 44328 29144 44334
rect 29092 44270 29144 44276
rect 28920 43926 28948 44270
rect 29380 43994 29408 47398
rect 29472 46170 29500 47903
rect 29564 46714 29592 48028
rect 29734 48039 29790 48048
rect 29644 48010 29696 48016
rect 29656 46918 29684 48010
rect 29644 46912 29696 46918
rect 29644 46854 29696 46860
rect 29552 46708 29604 46714
rect 29552 46650 29604 46656
rect 29552 46504 29604 46510
rect 29552 46446 29604 46452
rect 29460 46164 29512 46170
rect 29460 46106 29512 46112
rect 29460 45552 29512 45558
rect 29460 45494 29512 45500
rect 29368 43988 29420 43994
rect 29368 43930 29420 43936
rect 28908 43920 28960 43926
rect 28908 43862 28960 43868
rect 29000 43852 29052 43858
rect 29000 43794 29052 43800
rect 29012 42906 29040 43794
rect 29276 43784 29328 43790
rect 29276 43726 29328 43732
rect 29184 43444 29236 43450
rect 29184 43386 29236 43392
rect 29000 42900 29052 42906
rect 29000 42842 29052 42848
rect 29092 42900 29144 42906
rect 29092 42842 29144 42848
rect 29000 42764 29052 42770
rect 29000 42706 29052 42712
rect 29012 42362 29040 42706
rect 29000 42356 29052 42362
rect 29000 42298 29052 42304
rect 28814 37224 28870 37233
rect 28814 37159 28870 37168
rect 28816 35556 28868 35562
rect 28816 35498 28868 35504
rect 28724 31952 28776 31958
rect 28724 31894 28776 31900
rect 28722 31512 28778 31521
rect 28722 31447 28778 31456
rect 28736 31142 28764 31447
rect 28724 31136 28776 31142
rect 28724 31078 28776 31084
rect 28736 30054 28764 31078
rect 28724 30048 28776 30054
rect 28724 29990 28776 29996
rect 28736 29510 28764 29990
rect 28724 29504 28776 29510
rect 28724 29446 28776 29452
rect 28736 29306 28764 29446
rect 28724 29300 28776 29306
rect 28724 29242 28776 29248
rect 28724 29028 28776 29034
rect 28724 28970 28776 28976
rect 28736 27130 28764 28970
rect 28724 27124 28776 27130
rect 28724 27066 28776 27072
rect 28828 26897 28856 35498
rect 28906 33008 28962 33017
rect 28906 32943 28908 32952
rect 28960 32943 28962 32952
rect 28908 32914 28960 32920
rect 28920 32570 28948 32914
rect 28908 32564 28960 32570
rect 28908 32506 28960 32512
rect 28906 31784 28962 31793
rect 28906 31719 28962 31728
rect 28920 28762 28948 31719
rect 28998 30288 29054 30297
rect 28998 30223 29054 30232
rect 29012 29034 29040 30223
rect 29000 29028 29052 29034
rect 29000 28970 29052 28976
rect 28998 28792 29054 28801
rect 28908 28756 28960 28762
rect 28998 28727 29000 28736
rect 28908 28698 28960 28704
rect 29052 28727 29054 28736
rect 29000 28698 29052 28704
rect 28906 28112 28962 28121
rect 28906 28047 28962 28056
rect 28920 27606 28948 28047
rect 28908 27600 28960 27606
rect 28908 27542 28960 27548
rect 28998 27432 29054 27441
rect 28998 27367 29054 27376
rect 28814 26888 28870 26897
rect 28814 26823 28870 26832
rect 29012 22545 29040 27367
rect 29104 23361 29132 42842
rect 29196 41274 29224 43386
rect 29288 43382 29316 43726
rect 29276 43376 29328 43382
rect 29276 43318 29328 43324
rect 29288 42702 29316 43318
rect 29380 43314 29408 43930
rect 29472 43858 29500 45494
rect 29564 44946 29592 46446
rect 29552 44940 29604 44946
rect 29552 44882 29604 44888
rect 29460 43852 29512 43858
rect 29460 43794 29512 43800
rect 29564 43790 29592 44882
rect 29656 44169 29684 46854
rect 29748 45558 29776 48039
rect 29920 47660 29972 47666
rect 29920 47602 29972 47608
rect 29828 47592 29880 47598
rect 29828 47534 29880 47540
rect 29840 47258 29868 47534
rect 29828 47252 29880 47258
rect 29828 47194 29880 47200
rect 29932 47122 29960 47602
rect 29920 47116 29972 47122
rect 29920 47058 29972 47064
rect 29736 45552 29788 45558
rect 29736 45494 29788 45500
rect 29736 45348 29788 45354
rect 29736 45290 29788 45296
rect 29748 44713 29776 45290
rect 29920 45076 29972 45082
rect 29920 45018 29972 45024
rect 29828 44872 29880 44878
rect 29828 44814 29880 44820
rect 29734 44704 29790 44713
rect 29734 44639 29790 44648
rect 29642 44160 29698 44169
rect 29642 44095 29698 44104
rect 29552 43784 29604 43790
rect 29552 43726 29604 43732
rect 29368 43308 29420 43314
rect 29368 43250 29420 43256
rect 29460 43172 29512 43178
rect 29460 43114 29512 43120
rect 29472 42945 29500 43114
rect 29458 42936 29514 42945
rect 29458 42871 29514 42880
rect 29458 42800 29514 42809
rect 29458 42735 29460 42744
rect 29512 42735 29514 42744
rect 29460 42706 29512 42712
rect 29276 42696 29328 42702
rect 29276 42638 29328 42644
rect 29288 42294 29316 42638
rect 29472 42362 29500 42706
rect 29460 42356 29512 42362
rect 29460 42298 29512 42304
rect 29276 42288 29328 42294
rect 29276 42230 29328 42236
rect 29460 41472 29512 41478
rect 29564 41449 29592 43726
rect 29748 43246 29776 44639
rect 29840 44266 29868 44814
rect 29932 44334 29960 45018
rect 29920 44328 29972 44334
rect 29920 44270 29972 44276
rect 29828 44260 29880 44266
rect 29828 44202 29880 44208
rect 29932 43858 29960 44270
rect 29920 43852 29972 43858
rect 29920 43794 29972 43800
rect 29932 43722 29960 43794
rect 29920 43716 29972 43722
rect 29920 43658 29972 43664
rect 29932 43450 29960 43658
rect 29920 43444 29972 43450
rect 29920 43386 29972 43392
rect 29736 43240 29788 43246
rect 29736 43182 29788 43188
rect 29748 42906 29776 43182
rect 29736 42900 29788 42906
rect 29736 42842 29788 42848
rect 30024 41478 30052 50866
rect 30392 50833 30420 51206
rect 30378 50824 30434 50833
rect 30378 50759 30434 50768
rect 30484 50522 30512 51326
rect 30576 50930 30604 51428
rect 30564 50924 30616 50930
rect 30564 50866 30616 50872
rect 30472 50516 30524 50522
rect 30472 50458 30524 50464
rect 30668 50289 30696 51546
rect 30654 50280 30710 50289
rect 30654 50215 30710 50224
rect 30562 50144 30618 50153
rect 30562 50079 30618 50088
rect 30576 49842 30604 50079
rect 30668 49978 30696 50215
rect 30656 49972 30708 49978
rect 30656 49914 30708 49920
rect 30104 49836 30156 49842
rect 30104 49778 30156 49784
rect 30564 49836 30616 49842
rect 30564 49778 30616 49784
rect 30012 41472 30064 41478
rect 29460 41414 29512 41420
rect 29550 41440 29606 41449
rect 29184 41268 29236 41274
rect 29184 41210 29236 41216
rect 29472 39098 29500 41414
rect 30012 41414 30064 41420
rect 29550 41375 29606 41384
rect 29460 39092 29512 39098
rect 29460 39034 29512 39040
rect 29564 38894 29592 41375
rect 29826 41304 29882 41313
rect 29826 41239 29882 41248
rect 29644 40996 29696 41002
rect 29644 40938 29696 40944
rect 29552 38888 29604 38894
rect 29552 38830 29604 38836
rect 29564 38010 29592 38830
rect 29552 38004 29604 38010
rect 29552 37946 29604 37952
rect 29458 37360 29514 37369
rect 29458 37295 29514 37304
rect 29276 34536 29328 34542
rect 29276 34478 29328 34484
rect 29288 34202 29316 34478
rect 29276 34196 29328 34202
rect 29276 34138 29328 34144
rect 29288 33318 29316 34138
rect 29276 33312 29328 33318
rect 29276 33254 29328 33260
rect 29184 32496 29236 32502
rect 29184 32438 29236 32444
rect 29196 31890 29224 32438
rect 29472 31890 29500 37295
rect 29550 36408 29606 36417
rect 29550 36343 29552 36352
rect 29604 36343 29606 36352
rect 29552 36314 29604 36320
rect 29184 31884 29236 31890
rect 29184 31826 29236 31832
rect 29460 31884 29512 31890
rect 29460 31826 29512 31832
rect 29196 31142 29224 31826
rect 29472 31482 29500 31826
rect 29460 31476 29512 31482
rect 29460 31418 29512 31424
rect 29184 31136 29236 31142
rect 29184 31078 29236 31084
rect 29460 31136 29512 31142
rect 29460 31078 29512 31084
rect 29472 30054 29500 31078
rect 29460 30048 29512 30054
rect 29460 29990 29512 29996
rect 29274 28656 29330 28665
rect 29274 28591 29330 28600
rect 29184 28212 29236 28218
rect 29184 28154 29236 28160
rect 29090 23352 29146 23361
rect 29090 23287 29146 23296
rect 29196 22681 29224 28154
rect 29288 28014 29316 28591
rect 29472 28121 29500 29990
rect 29458 28112 29514 28121
rect 29458 28047 29514 28056
rect 29276 28008 29328 28014
rect 29276 27950 29328 27956
rect 29460 27872 29512 27878
rect 29460 27814 29512 27820
rect 29472 27713 29500 27814
rect 29458 27704 29514 27713
rect 29458 27639 29514 27648
rect 29656 27441 29684 40938
rect 29734 40896 29790 40905
rect 29734 40831 29790 40840
rect 29748 27985 29776 40831
rect 29840 34542 29868 41239
rect 30012 41132 30064 41138
rect 30012 41074 30064 41080
rect 30024 40390 30052 41074
rect 30012 40384 30064 40390
rect 30012 40326 30064 40332
rect 29920 38888 29972 38894
rect 29920 38830 29972 38836
rect 29932 38554 29960 38830
rect 29920 38548 29972 38554
rect 29920 38490 29972 38496
rect 29828 34536 29880 34542
rect 29828 34478 29880 34484
rect 30012 32768 30064 32774
rect 30012 32710 30064 32716
rect 30024 28218 30052 32710
rect 30012 28212 30064 28218
rect 30012 28154 30064 28160
rect 29734 27976 29790 27985
rect 29734 27911 29790 27920
rect 29642 27432 29698 27441
rect 29642 27367 29698 27376
rect 29182 22672 29238 22681
rect 29182 22607 29238 22616
rect 28998 22536 29054 22545
rect 28998 22471 29054 22480
rect 30116 19394 30144 49778
rect 30380 49700 30432 49706
rect 30380 49642 30432 49648
rect 30392 49434 30420 49642
rect 30380 49428 30432 49434
rect 30380 49370 30432 49376
rect 30194 49328 30250 49337
rect 30194 49263 30250 49272
rect 30208 47258 30236 49263
rect 30760 48890 30788 52430
rect 30840 50856 30892 50862
rect 30840 50798 30892 50804
rect 30852 49609 30880 50798
rect 30932 50720 30984 50726
rect 30932 50662 30984 50668
rect 31024 50720 31076 50726
rect 31024 50662 31076 50668
rect 30944 49881 30972 50662
rect 31036 50425 31064 50662
rect 31022 50416 31078 50425
rect 31022 50351 31078 50360
rect 31206 50008 31262 50017
rect 31206 49943 31262 49952
rect 30930 49872 30986 49881
rect 31220 49842 31248 49943
rect 30930 49807 30986 49816
rect 31208 49836 31260 49842
rect 30838 49600 30894 49609
rect 30838 49535 30894 49544
rect 30944 49450 30972 49807
rect 31208 49778 31260 49784
rect 31024 49768 31076 49774
rect 31024 49710 31076 49716
rect 30852 49422 30972 49450
rect 30748 48884 30800 48890
rect 30748 48826 30800 48832
rect 30288 48748 30340 48754
rect 30288 48690 30340 48696
rect 30196 47252 30248 47258
rect 30196 47194 30248 47200
rect 30208 45422 30236 47194
rect 30196 45416 30248 45422
rect 30196 45358 30248 45364
rect 30196 41608 30248 41614
rect 30196 41550 30248 41556
rect 30208 41070 30236 41550
rect 30196 41064 30248 41070
rect 30196 41006 30248 41012
rect 30024 19366 30144 19394
rect 28998 17232 29054 17241
rect 28998 17167 29054 17176
rect 28630 15872 28686 15881
rect 28630 15807 28686 15816
rect 27986 6216 28042 6225
rect 27986 6151 28042 6160
rect 29012 4826 29040 17167
rect 29642 15192 29698 15201
rect 29642 15127 29698 15136
rect 29000 4820 29052 4826
rect 29000 4762 29052 4768
rect 29368 4820 29420 4826
rect 29368 4762 29420 4768
rect 28446 2680 28502 2689
rect 28446 2615 28448 2624
rect 28500 2615 28502 2624
rect 28448 2586 28500 2592
rect 27620 2508 27672 2514
rect 27620 2450 27672 2456
rect 27160 2440 27212 2446
rect 27160 2382 27212 2388
rect 27172 2310 27200 2382
rect 27160 2304 27212 2310
rect 27160 2246 27212 2252
rect 27632 800 27660 2450
rect 28540 2440 28592 2446
rect 28540 2382 28592 2388
rect 28552 800 28580 2382
rect 29380 1986 29408 4762
rect 29656 2009 29684 15127
rect 30024 11121 30052 19366
rect 30104 19304 30156 19310
rect 30104 19246 30156 19252
rect 30116 18630 30144 19246
rect 30104 18624 30156 18630
rect 30102 18592 30104 18601
rect 30156 18592 30158 18601
rect 30102 18527 30158 18536
rect 30300 15065 30328 48690
rect 30656 48544 30708 48550
rect 30656 48486 30708 48492
rect 30668 48385 30696 48486
rect 30654 48376 30710 48385
rect 30654 48311 30710 48320
rect 30380 48204 30432 48210
rect 30380 48146 30432 48152
rect 30392 47530 30420 48146
rect 30746 48104 30802 48113
rect 30746 48039 30802 48048
rect 30380 47524 30432 47530
rect 30380 47466 30432 47472
rect 30656 47456 30708 47462
rect 30654 47424 30656 47433
rect 30708 47424 30710 47433
rect 30654 47359 30710 47368
rect 30760 47190 30788 48039
rect 30852 48006 30880 49422
rect 31036 49201 31064 49710
rect 31022 49192 31078 49201
rect 31022 49127 31078 49136
rect 31208 49088 31260 49094
rect 31208 49030 31260 49036
rect 31220 48890 31248 49030
rect 31208 48884 31260 48890
rect 31208 48826 31260 48832
rect 31206 48784 31262 48793
rect 31206 48719 31262 48728
rect 31220 48686 31248 48719
rect 31208 48680 31260 48686
rect 31208 48622 31260 48628
rect 30840 48000 30892 48006
rect 30840 47942 30892 47948
rect 30852 47598 30880 47942
rect 31116 47796 31168 47802
rect 31116 47738 31168 47744
rect 30840 47592 30892 47598
rect 30840 47534 30892 47540
rect 30932 47592 30984 47598
rect 30932 47534 30984 47540
rect 30748 47184 30800 47190
rect 30748 47126 30800 47132
rect 30564 47116 30616 47122
rect 30564 47058 30616 47064
rect 30380 47048 30432 47054
rect 30380 46990 30432 46996
rect 30392 46170 30420 46990
rect 30576 46617 30604 47058
rect 30562 46608 30618 46617
rect 30562 46543 30618 46552
rect 30576 46170 30604 46543
rect 30380 46164 30432 46170
rect 30380 46106 30432 46112
rect 30564 46164 30616 46170
rect 30564 46106 30616 46112
rect 30472 45824 30524 45830
rect 30472 45766 30524 45772
rect 30484 45082 30512 45766
rect 30852 45082 30880 47534
rect 30944 47297 30972 47534
rect 31024 47524 31076 47530
rect 31024 47466 31076 47472
rect 30930 47288 30986 47297
rect 30930 47223 30986 47232
rect 31036 47122 31064 47466
rect 31128 47161 31156 47738
rect 31114 47152 31170 47161
rect 31024 47116 31076 47122
rect 31114 47087 31170 47096
rect 31024 47058 31076 47064
rect 30932 46164 30984 46170
rect 30932 46106 30984 46112
rect 30944 45354 30972 46106
rect 31036 46034 31064 47058
rect 31116 47048 31168 47054
rect 31116 46990 31168 46996
rect 31128 46073 31156 46990
rect 31208 46368 31260 46374
rect 31208 46310 31260 46316
rect 31114 46064 31170 46073
rect 31024 46028 31076 46034
rect 31114 45999 31170 46008
rect 31024 45970 31076 45976
rect 31036 45626 31064 45970
rect 31024 45620 31076 45626
rect 31024 45562 31076 45568
rect 30932 45348 30984 45354
rect 30932 45290 30984 45296
rect 30472 45076 30524 45082
rect 30472 45018 30524 45024
rect 30840 45076 30892 45082
rect 30840 45018 30892 45024
rect 31220 44985 31248 46310
rect 31206 44976 31262 44985
rect 31206 44911 31262 44920
rect 31114 44840 31170 44849
rect 31114 44775 31170 44784
rect 31128 44538 31156 44775
rect 31116 44532 31168 44538
rect 31116 44474 31168 44480
rect 30840 44396 30892 44402
rect 30840 44338 30892 44344
rect 30748 44328 30800 44334
rect 30746 44296 30748 44305
rect 30800 44296 30802 44305
rect 30746 44231 30802 44240
rect 30380 43648 30432 43654
rect 30380 43590 30432 43596
rect 30392 43382 30420 43590
rect 30380 43376 30432 43382
rect 30380 43318 30432 43324
rect 30852 42401 30880 44338
rect 31116 44260 31168 44266
rect 31116 44202 31168 44208
rect 30838 42392 30894 42401
rect 30838 42327 30894 42336
rect 30472 38752 30524 38758
rect 30472 38694 30524 38700
rect 30484 38049 30512 38694
rect 30470 38040 30526 38049
rect 30470 37975 30526 37984
rect 30656 34604 30708 34610
rect 30656 34546 30708 34552
rect 30668 33697 30696 34546
rect 30654 33688 30710 33697
rect 30654 33623 30710 33632
rect 30564 31816 30616 31822
rect 30562 31784 30564 31793
rect 30616 31784 30618 31793
rect 30562 31719 30618 31728
rect 30470 26888 30526 26897
rect 30470 26823 30526 26832
rect 30286 15056 30342 15065
rect 30286 14991 30342 15000
rect 30484 12646 30512 26823
rect 31128 20369 31156 44202
rect 31312 37369 31340 74718
rect 33140 74656 33192 74662
rect 33140 74598 33192 74604
rect 32312 60512 32364 60518
rect 32312 60454 32364 60460
rect 31390 60344 31446 60353
rect 31390 60279 31446 60288
rect 31404 51474 31432 60279
rect 32324 59634 32352 60454
rect 32312 59628 32364 59634
rect 32312 59570 32364 59576
rect 32954 58984 33010 58993
rect 32954 58919 33010 58928
rect 31758 56536 31814 56545
rect 31758 56471 31814 56480
rect 31574 55312 31630 55321
rect 31574 55247 31576 55256
rect 31628 55247 31630 55256
rect 31576 55218 31628 55224
rect 31772 55214 31800 56471
rect 32680 55616 32732 55622
rect 32680 55558 32732 55564
rect 32692 55214 32720 55558
rect 31760 55208 31812 55214
rect 31760 55150 31812 55156
rect 32680 55208 32732 55214
rect 32680 55150 32732 55156
rect 31772 54534 31800 55150
rect 31944 55140 31996 55146
rect 31944 55082 31996 55088
rect 31760 54528 31812 54534
rect 31760 54470 31812 54476
rect 31772 52465 31800 54470
rect 31956 53961 31984 55082
rect 32586 54088 32642 54097
rect 32586 54023 32642 54032
rect 31942 53952 31998 53961
rect 31942 53887 31998 53896
rect 31758 52456 31814 52465
rect 31758 52391 31814 52400
rect 31760 51808 31812 51814
rect 31760 51750 31812 51756
rect 31392 51468 31444 51474
rect 31392 51410 31444 51416
rect 31404 51066 31432 51410
rect 31484 51264 31536 51270
rect 31484 51206 31536 51212
rect 31392 51060 31444 51066
rect 31392 51002 31444 51008
rect 31496 50697 31524 51206
rect 31482 50688 31538 50697
rect 31482 50623 31538 50632
rect 31496 50386 31524 50623
rect 31484 50380 31536 50386
rect 31484 50322 31536 50328
rect 31772 49722 31800 51750
rect 32218 50280 32274 50289
rect 32218 50215 32274 50224
rect 32232 49978 32260 50215
rect 31944 49972 31996 49978
rect 31944 49914 31996 49920
rect 32220 49972 32272 49978
rect 32220 49914 32272 49920
rect 31680 49694 31800 49722
rect 31680 49434 31708 49694
rect 31668 49428 31720 49434
rect 31668 49370 31720 49376
rect 31390 49328 31446 49337
rect 31390 49263 31446 49272
rect 31404 48890 31432 49263
rect 31392 48884 31444 48890
rect 31392 48826 31444 48832
rect 31392 48136 31444 48142
rect 31392 48078 31444 48084
rect 31404 47258 31432 48078
rect 31392 47252 31444 47258
rect 31392 47194 31444 47200
rect 31852 47184 31904 47190
rect 31852 47126 31904 47132
rect 31864 46646 31892 47126
rect 31852 46640 31904 46646
rect 31852 46582 31904 46588
rect 31956 46578 31984 49914
rect 32404 47728 32456 47734
rect 32402 47696 32404 47705
rect 32456 47696 32458 47705
rect 32402 47631 32458 47640
rect 32034 47152 32090 47161
rect 32034 47087 32090 47096
rect 32128 47116 32180 47122
rect 31944 46572 31996 46578
rect 31944 46514 31996 46520
rect 31760 46368 31812 46374
rect 31760 46310 31812 46316
rect 31772 46170 31800 46310
rect 31760 46164 31812 46170
rect 31760 46106 31812 46112
rect 31392 45824 31444 45830
rect 31392 45766 31444 45772
rect 31404 45354 31432 45766
rect 31484 45416 31536 45422
rect 31484 45358 31536 45364
rect 31392 45348 31444 45354
rect 31392 45290 31444 45296
rect 31404 42809 31432 45290
rect 31496 45082 31524 45358
rect 31576 45348 31628 45354
rect 31576 45290 31628 45296
rect 31484 45076 31536 45082
rect 31484 45018 31536 45024
rect 31588 44577 31616 45290
rect 31852 44736 31904 44742
rect 31850 44704 31852 44713
rect 31904 44704 31906 44713
rect 31850 44639 31906 44648
rect 31574 44568 31630 44577
rect 31574 44503 31630 44512
rect 31390 42800 31446 42809
rect 31390 42735 31446 42744
rect 31298 37360 31354 37369
rect 31298 37295 31354 37304
rect 32048 28626 32076 47087
rect 32128 47058 32180 47064
rect 32140 46714 32168 47058
rect 32128 46708 32180 46714
rect 32128 46650 32180 46656
rect 32126 46336 32182 46345
rect 32126 46271 32182 46280
rect 32140 46034 32168 46271
rect 32218 46200 32274 46209
rect 32218 46135 32274 46144
rect 32232 46034 32260 46135
rect 32128 46028 32180 46034
rect 32128 45970 32180 45976
rect 32220 46028 32272 46034
rect 32220 45970 32272 45976
rect 32140 45626 32168 45970
rect 32232 45626 32260 45970
rect 32402 45928 32458 45937
rect 32402 45863 32458 45872
rect 32416 45830 32444 45863
rect 32404 45824 32456 45830
rect 32404 45766 32456 45772
rect 32128 45620 32180 45626
rect 32128 45562 32180 45568
rect 32220 45620 32272 45626
rect 32220 45562 32272 45568
rect 32220 37324 32272 37330
rect 32220 37266 32272 37272
rect 32232 37210 32260 37266
rect 32140 37182 32260 37210
rect 32496 37256 32548 37262
rect 32496 37198 32548 37204
rect 32140 36582 32168 37182
rect 32508 36922 32536 37198
rect 32496 36916 32548 36922
rect 32496 36858 32548 36864
rect 32128 36576 32180 36582
rect 32128 36518 32180 36524
rect 32036 28620 32088 28626
rect 32036 28562 32088 28568
rect 31482 20632 31538 20641
rect 31482 20567 31538 20576
rect 31114 20360 31170 20369
rect 31114 20295 31170 20304
rect 31496 19514 31524 20567
rect 31484 19508 31536 19514
rect 31484 19450 31536 19456
rect 31668 19304 31720 19310
rect 31720 19252 31800 19258
rect 31668 19246 31800 19252
rect 31680 19230 31800 19246
rect 30288 12640 30340 12646
rect 30288 12582 30340 12588
rect 30472 12640 30524 12646
rect 30472 12582 30524 12588
rect 30010 11112 30066 11121
rect 30010 11047 30066 11056
rect 30300 9761 30328 12582
rect 30286 9752 30342 9761
rect 30286 9687 30342 9696
rect 31298 2272 31354 2281
rect 31298 2207 31354 2216
rect 29642 2000 29698 2009
rect 29380 1958 29500 1986
rect 29472 800 29500 1958
rect 29642 1935 29698 1944
rect 30378 912 30434 921
rect 30378 847 30434 856
rect 30392 800 30420 847
rect 31312 800 31340 2207
rect 31772 800 31800 19230
rect 32140 12481 32168 36518
rect 32402 34096 32458 34105
rect 32402 34031 32404 34040
rect 32456 34031 32458 34040
rect 32404 34002 32456 34008
rect 32416 33658 32444 34002
rect 32508 33998 32536 36858
rect 32600 36825 32628 54023
rect 32678 47016 32734 47025
rect 32678 46951 32734 46960
rect 32586 36816 32642 36825
rect 32586 36751 32642 36760
rect 32496 33992 32548 33998
rect 32496 33934 32548 33940
rect 32508 33658 32536 33934
rect 32404 33652 32456 33658
rect 32404 33594 32456 33600
rect 32496 33652 32548 33658
rect 32496 33594 32548 33600
rect 32508 33318 32536 33594
rect 32496 33312 32548 33318
rect 32496 33254 32548 33260
rect 32692 33017 32720 46951
rect 32968 44985 32996 58919
rect 33152 47161 33180 74598
rect 33244 55978 33272 74718
rect 33244 55950 33364 55978
rect 33232 55820 33284 55826
rect 33232 55762 33284 55768
rect 33244 55418 33272 55762
rect 33232 55412 33284 55418
rect 33232 55354 33284 55360
rect 33336 52873 33364 55950
rect 33322 52864 33378 52873
rect 33322 52799 33378 52808
rect 33138 47152 33194 47161
rect 33138 47087 33194 47096
rect 33046 46200 33102 46209
rect 33046 46135 33102 46144
rect 32954 44976 33010 44985
rect 32954 44911 33010 44920
rect 33060 36689 33088 46135
rect 33520 37466 33548 77658
rect 34072 74662 34100 79200
rect 34992 77466 35020 79200
rect 35346 78296 35402 78305
rect 35346 78231 35402 78240
rect 34808 77438 35020 77466
rect 35360 77450 35388 78231
rect 35348 77444 35400 77450
rect 34808 75585 34836 77438
rect 35348 77386 35400 77392
rect 34940 77276 35236 77296
rect 34996 77274 35020 77276
rect 35076 77274 35100 77276
rect 35156 77274 35180 77276
rect 35018 77222 35020 77274
rect 35082 77222 35094 77274
rect 35156 77222 35158 77274
rect 34996 77220 35020 77222
rect 35076 77220 35100 77222
rect 35156 77220 35180 77222
rect 34940 77200 35236 77220
rect 34940 76188 35236 76208
rect 34996 76186 35020 76188
rect 35076 76186 35100 76188
rect 35156 76186 35180 76188
rect 35018 76134 35020 76186
rect 35082 76134 35094 76186
rect 35156 76134 35158 76186
rect 34996 76132 35020 76134
rect 35076 76132 35100 76134
rect 35156 76132 35180 76134
rect 34940 76112 35236 76132
rect 34794 75576 34850 75585
rect 34794 75511 34850 75520
rect 34940 75100 35236 75120
rect 34996 75098 35020 75100
rect 35076 75098 35100 75100
rect 35156 75098 35180 75100
rect 35018 75046 35020 75098
rect 35082 75046 35094 75098
rect 35156 75046 35158 75098
rect 34996 75044 35020 75046
rect 35076 75044 35100 75046
rect 35156 75044 35180 75046
rect 34940 75024 35236 75044
rect 35452 75018 35480 79591
rect 35898 79200 35954 80000
rect 36818 79200 36874 80000
rect 37738 79200 37794 80000
rect 38658 79200 38714 80000
rect 39578 79200 39634 80000
rect 35806 76936 35862 76945
rect 35806 76871 35862 76880
rect 35622 75576 35678 75585
rect 35622 75511 35678 75520
rect 35360 74990 35480 75018
rect 34060 74656 34112 74662
rect 34060 74598 34112 74604
rect 34940 74012 35236 74032
rect 34996 74010 35020 74012
rect 35076 74010 35100 74012
rect 35156 74010 35180 74012
rect 35018 73958 35020 74010
rect 35082 73958 35094 74010
rect 35156 73958 35158 74010
rect 34996 73956 35020 73958
rect 35076 73956 35100 73958
rect 35156 73956 35180 73958
rect 34940 73936 35236 73956
rect 34940 72924 35236 72944
rect 34996 72922 35020 72924
rect 35076 72922 35100 72924
rect 35156 72922 35180 72924
rect 35018 72870 35020 72922
rect 35082 72870 35094 72922
rect 35156 72870 35158 72922
rect 34996 72868 35020 72870
rect 35076 72868 35100 72870
rect 35156 72868 35180 72870
rect 34940 72848 35236 72868
rect 34940 71836 35236 71856
rect 34996 71834 35020 71836
rect 35076 71834 35100 71836
rect 35156 71834 35180 71836
rect 35018 71782 35020 71834
rect 35082 71782 35094 71834
rect 35156 71782 35158 71834
rect 34996 71780 35020 71782
rect 35076 71780 35100 71782
rect 35156 71780 35180 71782
rect 34940 71760 35236 71780
rect 34518 71496 34574 71505
rect 34518 71431 34574 71440
rect 34532 70009 34560 71431
rect 34940 70748 35236 70768
rect 34996 70746 35020 70748
rect 35076 70746 35100 70748
rect 35156 70746 35180 70748
rect 35018 70694 35020 70746
rect 35082 70694 35094 70746
rect 35156 70694 35158 70746
rect 34996 70692 35020 70694
rect 35076 70692 35100 70694
rect 35156 70692 35180 70694
rect 34940 70672 35236 70692
rect 34518 70000 34574 70009
rect 34518 69935 34574 69944
rect 34940 69660 35236 69680
rect 34996 69658 35020 69660
rect 35076 69658 35100 69660
rect 35156 69658 35180 69660
rect 35018 69606 35020 69658
rect 35082 69606 35094 69658
rect 35156 69606 35158 69658
rect 34996 69604 35020 69606
rect 35076 69604 35100 69606
rect 35156 69604 35180 69606
rect 34940 69584 35236 69604
rect 34940 68572 35236 68592
rect 34996 68570 35020 68572
rect 35076 68570 35100 68572
rect 35156 68570 35180 68572
rect 35018 68518 35020 68570
rect 35082 68518 35094 68570
rect 35156 68518 35158 68570
rect 34996 68516 35020 68518
rect 35076 68516 35100 68518
rect 35156 68516 35180 68518
rect 34940 68496 35236 68516
rect 34940 67484 35236 67504
rect 34996 67482 35020 67484
rect 35076 67482 35100 67484
rect 35156 67482 35180 67484
rect 35018 67430 35020 67482
rect 35082 67430 35094 67482
rect 35156 67430 35158 67482
rect 34996 67428 35020 67430
rect 35076 67428 35100 67430
rect 35156 67428 35180 67430
rect 34940 67408 35236 67428
rect 34940 66396 35236 66416
rect 34996 66394 35020 66396
rect 35076 66394 35100 66396
rect 35156 66394 35180 66396
rect 35018 66342 35020 66394
rect 35082 66342 35094 66394
rect 35156 66342 35158 66394
rect 34996 66340 35020 66342
rect 35076 66340 35100 66342
rect 35156 66340 35180 66342
rect 34940 66320 35236 66340
rect 34940 65308 35236 65328
rect 34996 65306 35020 65308
rect 35076 65306 35100 65308
rect 35156 65306 35180 65308
rect 35018 65254 35020 65306
rect 35082 65254 35094 65306
rect 35156 65254 35158 65306
rect 34996 65252 35020 65254
rect 35076 65252 35100 65254
rect 35156 65252 35180 65254
rect 34940 65232 35236 65252
rect 34940 64220 35236 64240
rect 34996 64218 35020 64220
rect 35076 64218 35100 64220
rect 35156 64218 35180 64220
rect 35018 64166 35020 64218
rect 35082 64166 35094 64218
rect 35156 64166 35158 64218
rect 34996 64164 35020 64166
rect 35076 64164 35100 64166
rect 35156 64164 35180 64166
rect 34940 64144 35236 64164
rect 34940 63132 35236 63152
rect 34996 63130 35020 63132
rect 35076 63130 35100 63132
rect 35156 63130 35180 63132
rect 35018 63078 35020 63130
rect 35082 63078 35094 63130
rect 35156 63078 35158 63130
rect 34996 63076 35020 63078
rect 35076 63076 35100 63078
rect 35156 63076 35180 63078
rect 34940 63056 35236 63076
rect 34940 62044 35236 62064
rect 34996 62042 35020 62044
rect 35076 62042 35100 62044
rect 35156 62042 35180 62044
rect 35018 61990 35020 62042
rect 35082 61990 35094 62042
rect 35156 61990 35158 62042
rect 34996 61988 35020 61990
rect 35076 61988 35100 61990
rect 35156 61988 35180 61990
rect 34940 61968 35236 61988
rect 34940 60956 35236 60976
rect 34996 60954 35020 60956
rect 35076 60954 35100 60956
rect 35156 60954 35180 60956
rect 35018 60902 35020 60954
rect 35082 60902 35094 60954
rect 35156 60902 35158 60954
rect 34996 60900 35020 60902
rect 35076 60900 35100 60902
rect 35156 60900 35180 60902
rect 34940 60880 35236 60900
rect 35360 60058 35388 74990
rect 35438 72856 35494 72865
rect 35438 72791 35494 72800
rect 35452 70961 35480 72791
rect 35438 70952 35494 70961
rect 35438 70887 35494 70896
rect 35530 68776 35586 68785
rect 35530 68711 35586 68720
rect 35438 65376 35494 65385
rect 35438 65311 35494 65320
rect 35452 62257 35480 65311
rect 35544 62801 35572 68711
rect 35530 62792 35586 62801
rect 35530 62727 35586 62736
rect 35438 62248 35494 62257
rect 35438 62183 35494 62192
rect 35636 61441 35664 75511
rect 35622 61432 35678 61441
rect 35622 61367 35678 61376
rect 35438 61296 35494 61305
rect 35438 61231 35494 61240
rect 34716 60030 35388 60058
rect 34518 57216 34574 57225
rect 34518 57151 34574 57160
rect 34532 55842 34560 57151
rect 34612 56704 34664 56710
rect 34612 56646 34664 56652
rect 34440 55826 34560 55842
rect 34428 55820 34560 55826
rect 34480 55814 34560 55820
rect 34428 55762 34480 55768
rect 34624 55758 34652 56646
rect 33600 55752 33652 55758
rect 33600 55694 33652 55700
rect 34612 55752 34664 55758
rect 34612 55694 34664 55700
rect 33612 55282 33640 55694
rect 33600 55276 33652 55282
rect 33600 55218 33652 55224
rect 33612 51270 33640 55218
rect 34716 52601 34744 60030
rect 35256 59968 35308 59974
rect 35256 59910 35308 59916
rect 34940 59868 35236 59888
rect 34996 59866 35020 59868
rect 35076 59866 35100 59868
rect 35156 59866 35180 59868
rect 35018 59814 35020 59866
rect 35082 59814 35094 59866
rect 35156 59814 35158 59866
rect 34996 59812 35020 59814
rect 35076 59812 35100 59814
rect 35156 59812 35180 59814
rect 34940 59792 35236 59812
rect 35268 59090 35296 59910
rect 35452 59090 35480 61231
rect 35820 61169 35848 76871
rect 35912 71641 35940 79200
rect 36832 73273 36860 79200
rect 37752 79098 37780 79200
rect 37476 79070 37780 79098
rect 37372 74792 37424 74798
rect 37372 74734 37424 74740
rect 36818 73264 36874 73273
rect 36818 73199 36874 73208
rect 35898 71632 35954 71641
rect 35898 71567 35954 71576
rect 37384 68241 37412 74734
rect 37370 68232 37426 68241
rect 37370 68167 37426 68176
rect 35806 61160 35862 61169
rect 35806 61095 35862 61104
rect 37476 60722 37504 79070
rect 38672 74798 38700 79200
rect 38660 74792 38712 74798
rect 38660 74734 38712 74740
rect 39592 73817 39620 79200
rect 39578 73808 39634 73817
rect 39578 73743 39634 73752
rect 37464 60716 37516 60722
rect 37464 60658 37516 60664
rect 35808 60648 35860 60654
rect 35808 60590 35860 60596
rect 35820 59974 35848 60590
rect 37372 60512 37424 60518
rect 37372 60454 37424 60460
rect 35808 59968 35860 59974
rect 35808 59910 35860 59916
rect 37384 59401 37412 60454
rect 37370 59392 37426 59401
rect 37370 59327 37426 59336
rect 35256 59084 35308 59090
rect 35256 59026 35308 59032
rect 35440 59084 35492 59090
rect 35440 59026 35492 59032
rect 34940 58780 35236 58800
rect 34996 58778 35020 58780
rect 35076 58778 35100 58780
rect 35156 58778 35180 58780
rect 35018 58726 35020 58778
rect 35082 58726 35094 58778
rect 35156 58726 35158 58778
rect 34996 58724 35020 58726
rect 35076 58724 35100 58726
rect 35156 58724 35180 58726
rect 34940 58704 35236 58724
rect 35268 58342 35296 59026
rect 35452 58682 35480 59026
rect 35808 58880 35860 58886
rect 35808 58822 35860 58828
rect 35440 58676 35492 58682
rect 35440 58618 35492 58624
rect 35346 58576 35402 58585
rect 35346 58511 35402 58520
rect 35256 58336 35308 58342
rect 35256 58278 35308 58284
rect 34940 57692 35236 57712
rect 34996 57690 35020 57692
rect 35076 57690 35100 57692
rect 35156 57690 35180 57692
rect 35018 57638 35020 57690
rect 35082 57638 35094 57690
rect 35156 57638 35158 57690
rect 34996 57636 35020 57638
rect 35076 57636 35100 57638
rect 35156 57636 35180 57638
rect 34940 57616 35236 57636
rect 35268 57390 35296 58278
rect 35256 57384 35308 57390
rect 35256 57326 35308 57332
rect 35268 56710 35296 57326
rect 35256 56704 35308 56710
rect 35256 56646 35308 56652
rect 34940 56604 35236 56624
rect 34996 56602 35020 56604
rect 35076 56602 35100 56604
rect 35156 56602 35180 56604
rect 35018 56550 35020 56602
rect 35082 56550 35094 56602
rect 35156 56550 35158 56602
rect 34996 56548 35020 56550
rect 35076 56548 35100 56550
rect 35156 56548 35180 56550
rect 34940 56528 35236 56548
rect 34940 55516 35236 55536
rect 34996 55514 35020 55516
rect 35076 55514 35100 55516
rect 35156 55514 35180 55516
rect 35018 55462 35020 55514
rect 35082 55462 35094 55514
rect 35156 55462 35158 55514
rect 34996 55460 35020 55462
rect 35076 55460 35100 55462
rect 35156 55460 35180 55462
rect 34940 55440 35236 55460
rect 34940 54428 35236 54448
rect 34996 54426 35020 54428
rect 35076 54426 35100 54428
rect 35156 54426 35180 54428
rect 35018 54374 35020 54426
rect 35082 54374 35094 54426
rect 35156 54374 35158 54426
rect 34996 54372 35020 54374
rect 35076 54372 35100 54374
rect 35156 54372 35180 54374
rect 34940 54352 35236 54372
rect 35254 53952 35310 53961
rect 35254 53887 35310 53896
rect 34940 53340 35236 53360
rect 34996 53338 35020 53340
rect 35076 53338 35100 53340
rect 35156 53338 35180 53340
rect 35018 53286 35020 53338
rect 35082 53286 35094 53338
rect 35156 53286 35158 53338
rect 34996 53284 35020 53286
rect 35076 53284 35100 53286
rect 35156 53284 35180 53286
rect 34940 53264 35236 53284
rect 34702 52592 34758 52601
rect 34702 52527 34758 52536
rect 34704 52488 34756 52494
rect 34610 52456 34666 52465
rect 34704 52430 34756 52436
rect 34610 52391 34666 52400
rect 33692 51468 33744 51474
rect 33692 51410 33744 51416
rect 33600 51264 33652 51270
rect 33600 51206 33652 51212
rect 33704 50862 33732 51410
rect 34152 51264 34204 51270
rect 34152 51206 34204 51212
rect 33692 50856 33744 50862
rect 33692 50798 33744 50804
rect 33704 50697 33732 50798
rect 33690 50688 33746 50697
rect 33690 50623 33746 50632
rect 34164 44334 34192 51206
rect 34624 47025 34652 52391
rect 34610 47016 34666 47025
rect 34610 46951 34666 46960
rect 34152 44328 34204 44334
rect 34152 44270 34204 44276
rect 34164 42770 34192 44270
rect 34518 42936 34574 42945
rect 34518 42871 34574 42880
rect 34152 42764 34204 42770
rect 34152 42706 34204 42712
rect 34060 42696 34112 42702
rect 34060 42638 34112 42644
rect 34072 42022 34100 42638
rect 34164 42362 34192 42706
rect 34152 42356 34204 42362
rect 34152 42298 34204 42304
rect 34060 42016 34112 42022
rect 34060 41958 34112 41964
rect 33508 37460 33560 37466
rect 33508 37402 33560 37408
rect 33046 36680 33102 36689
rect 33046 36615 33102 36624
rect 33508 33856 33560 33862
rect 33508 33798 33560 33804
rect 32678 33008 32734 33017
rect 32678 32943 32734 32952
rect 32496 28620 32548 28626
rect 32496 28562 32548 28568
rect 32508 28218 32536 28562
rect 32772 28552 32824 28558
rect 32772 28494 32824 28500
rect 32784 28218 32812 28494
rect 32496 28212 32548 28218
rect 32496 28154 32548 28160
rect 32772 28212 32824 28218
rect 32772 28154 32824 28160
rect 32784 28121 32812 28154
rect 32770 28112 32826 28121
rect 32770 28047 32826 28056
rect 33520 26353 33548 33798
rect 33784 28416 33836 28422
rect 33784 28358 33836 28364
rect 33506 26344 33562 26353
rect 33506 26279 33562 26288
rect 33796 23633 33824 28358
rect 34072 27577 34100 41958
rect 34532 40905 34560 42871
rect 34612 42356 34664 42362
rect 34612 42298 34664 42304
rect 34518 40896 34574 40905
rect 34518 40831 34574 40840
rect 34624 40526 34652 42298
rect 34716 41274 34744 52430
rect 34940 52252 35236 52272
rect 34996 52250 35020 52252
rect 35076 52250 35100 52252
rect 35156 52250 35180 52252
rect 35018 52198 35020 52250
rect 35082 52198 35094 52250
rect 35156 52198 35158 52250
rect 34996 52196 35020 52198
rect 35076 52196 35100 52198
rect 35156 52196 35180 52198
rect 34940 52176 35236 52196
rect 34940 51164 35236 51184
rect 34996 51162 35020 51164
rect 35076 51162 35100 51164
rect 35156 51162 35180 51164
rect 35018 51110 35020 51162
rect 35082 51110 35094 51162
rect 35156 51110 35158 51162
rect 34996 51108 35020 51110
rect 35076 51108 35100 51110
rect 35156 51108 35180 51110
rect 34940 51088 35236 51108
rect 34796 50720 34848 50726
rect 34796 50662 34848 50668
rect 34808 46209 34836 50662
rect 34940 50076 35236 50096
rect 34996 50074 35020 50076
rect 35076 50074 35100 50076
rect 35156 50074 35180 50076
rect 35018 50022 35020 50074
rect 35082 50022 35094 50074
rect 35156 50022 35158 50074
rect 34996 50020 35020 50022
rect 35076 50020 35100 50022
rect 35156 50020 35180 50022
rect 34940 50000 35236 50020
rect 34940 48988 35236 49008
rect 34996 48986 35020 48988
rect 35076 48986 35100 48988
rect 35156 48986 35180 48988
rect 35018 48934 35020 48986
rect 35082 48934 35094 48986
rect 35156 48934 35158 48986
rect 34996 48932 35020 48934
rect 35076 48932 35100 48934
rect 35156 48932 35180 48934
rect 34940 48912 35236 48932
rect 34940 47900 35236 47920
rect 34996 47898 35020 47900
rect 35076 47898 35100 47900
rect 35156 47898 35180 47900
rect 35018 47846 35020 47898
rect 35082 47846 35094 47898
rect 35156 47846 35158 47898
rect 34996 47844 35020 47846
rect 35076 47844 35100 47846
rect 35156 47844 35180 47846
rect 34940 47824 35236 47844
rect 34940 46812 35236 46832
rect 34996 46810 35020 46812
rect 35076 46810 35100 46812
rect 35156 46810 35180 46812
rect 35018 46758 35020 46810
rect 35082 46758 35094 46810
rect 35156 46758 35158 46810
rect 34996 46756 35020 46758
rect 35076 46756 35100 46758
rect 35156 46756 35180 46758
rect 34940 46736 35236 46756
rect 34794 46200 34850 46209
rect 34794 46135 34850 46144
rect 34940 45724 35236 45744
rect 34996 45722 35020 45724
rect 35076 45722 35100 45724
rect 35156 45722 35180 45724
rect 35018 45670 35020 45722
rect 35082 45670 35094 45722
rect 35156 45670 35158 45722
rect 34996 45668 35020 45670
rect 35076 45668 35100 45670
rect 35156 45668 35180 45670
rect 34940 45648 35236 45668
rect 34940 44636 35236 44656
rect 34996 44634 35020 44636
rect 35076 44634 35100 44636
rect 35156 44634 35180 44636
rect 35018 44582 35020 44634
rect 35082 44582 35094 44634
rect 35156 44582 35158 44634
rect 34996 44580 35020 44582
rect 35076 44580 35100 44582
rect 35156 44580 35180 44582
rect 34940 44560 35236 44580
rect 34940 43548 35236 43568
rect 34996 43546 35020 43548
rect 35076 43546 35100 43548
rect 35156 43546 35180 43548
rect 35018 43494 35020 43546
rect 35082 43494 35094 43546
rect 35156 43494 35158 43546
rect 34996 43492 35020 43494
rect 35076 43492 35100 43494
rect 35156 43492 35180 43494
rect 34940 43472 35236 43492
rect 35162 42800 35218 42809
rect 35162 42735 35218 42744
rect 35176 42702 35204 42735
rect 35164 42696 35216 42702
rect 34794 42664 34850 42673
rect 35164 42638 35216 42644
rect 34794 42599 34850 42608
rect 34704 41268 34756 41274
rect 34704 41210 34756 41216
rect 34612 40520 34664 40526
rect 34612 40462 34664 40468
rect 34808 39545 34836 42599
rect 34940 42460 35236 42480
rect 34996 42458 35020 42460
rect 35076 42458 35100 42460
rect 35156 42458 35180 42460
rect 35018 42406 35020 42458
rect 35082 42406 35094 42458
rect 35156 42406 35158 42458
rect 34996 42404 35020 42406
rect 35076 42404 35100 42406
rect 35156 42404 35180 42406
rect 34940 42384 35236 42404
rect 34940 41372 35236 41392
rect 34996 41370 35020 41372
rect 35076 41370 35100 41372
rect 35156 41370 35180 41372
rect 35018 41318 35020 41370
rect 35082 41318 35094 41370
rect 35156 41318 35158 41370
rect 34996 41316 35020 41318
rect 35076 41316 35100 41318
rect 35156 41316 35180 41318
rect 34940 41296 35236 41316
rect 34888 41200 34940 41206
rect 34888 41142 34940 41148
rect 34900 40594 34928 41142
rect 34888 40588 34940 40594
rect 34888 40530 34940 40536
rect 34940 40284 35236 40304
rect 34996 40282 35020 40284
rect 35076 40282 35100 40284
rect 35156 40282 35180 40284
rect 35018 40230 35020 40282
rect 35082 40230 35094 40282
rect 35156 40230 35158 40282
rect 34996 40228 35020 40230
rect 35076 40228 35100 40230
rect 35156 40228 35180 40230
rect 34940 40208 35236 40228
rect 34794 39536 34850 39545
rect 34794 39471 34850 39480
rect 34704 39432 34756 39438
rect 34704 39374 34756 39380
rect 34716 38321 34744 39374
rect 34940 39196 35236 39216
rect 34996 39194 35020 39196
rect 35076 39194 35100 39196
rect 35156 39194 35180 39196
rect 35018 39142 35020 39194
rect 35082 39142 35094 39194
rect 35156 39142 35158 39194
rect 34996 39140 35020 39142
rect 35076 39140 35100 39142
rect 35156 39140 35180 39142
rect 34940 39120 35236 39140
rect 34702 38312 34758 38321
rect 34702 38247 34758 38256
rect 34940 38108 35236 38128
rect 34996 38106 35020 38108
rect 35076 38106 35100 38108
rect 35156 38106 35180 38108
rect 35018 38054 35020 38106
rect 35082 38054 35094 38106
rect 35156 38054 35158 38106
rect 34996 38052 35020 38054
rect 35076 38052 35100 38054
rect 35156 38052 35180 38054
rect 34940 38032 35236 38052
rect 34940 37020 35236 37040
rect 34996 37018 35020 37020
rect 35076 37018 35100 37020
rect 35156 37018 35180 37020
rect 35018 36966 35020 37018
rect 35082 36966 35094 37018
rect 35156 36966 35158 37018
rect 34996 36964 35020 36966
rect 35076 36964 35100 36966
rect 35156 36964 35180 36966
rect 34940 36944 35236 36964
rect 34940 35932 35236 35952
rect 34996 35930 35020 35932
rect 35076 35930 35100 35932
rect 35156 35930 35180 35932
rect 35018 35878 35020 35930
rect 35082 35878 35094 35930
rect 35156 35878 35158 35930
rect 34996 35876 35020 35878
rect 35076 35876 35100 35878
rect 35156 35876 35180 35878
rect 34940 35856 35236 35876
rect 34940 34844 35236 34864
rect 34996 34842 35020 34844
rect 35076 34842 35100 34844
rect 35156 34842 35180 34844
rect 35018 34790 35020 34842
rect 35082 34790 35094 34842
rect 35156 34790 35158 34842
rect 34996 34788 35020 34790
rect 35076 34788 35100 34790
rect 35156 34788 35180 34790
rect 34940 34768 35236 34788
rect 34940 33756 35236 33776
rect 34996 33754 35020 33756
rect 35076 33754 35100 33756
rect 35156 33754 35180 33756
rect 35018 33702 35020 33754
rect 35082 33702 35094 33754
rect 35156 33702 35158 33754
rect 34996 33700 35020 33702
rect 35076 33700 35100 33702
rect 35156 33700 35180 33702
rect 34940 33680 35236 33700
rect 34940 32668 35236 32688
rect 34996 32666 35020 32668
rect 35076 32666 35100 32668
rect 35156 32666 35180 32668
rect 35018 32614 35020 32666
rect 35082 32614 35094 32666
rect 35156 32614 35158 32666
rect 34996 32612 35020 32614
rect 35076 32612 35100 32614
rect 35156 32612 35180 32614
rect 34940 32592 35236 32612
rect 34940 31580 35236 31600
rect 34996 31578 35020 31580
rect 35076 31578 35100 31580
rect 35156 31578 35180 31580
rect 35018 31526 35020 31578
rect 35082 31526 35094 31578
rect 35156 31526 35158 31578
rect 34996 31524 35020 31526
rect 35076 31524 35100 31526
rect 35156 31524 35180 31526
rect 34940 31504 35236 31524
rect 34940 30492 35236 30512
rect 34996 30490 35020 30492
rect 35076 30490 35100 30492
rect 35156 30490 35180 30492
rect 35018 30438 35020 30490
rect 35082 30438 35094 30490
rect 35156 30438 35158 30490
rect 34996 30436 35020 30438
rect 35076 30436 35100 30438
rect 35156 30436 35180 30438
rect 34940 30416 35236 30436
rect 34940 29404 35236 29424
rect 34996 29402 35020 29404
rect 35076 29402 35100 29404
rect 35156 29402 35180 29404
rect 35018 29350 35020 29402
rect 35082 29350 35094 29402
rect 35156 29350 35158 29402
rect 34996 29348 35020 29350
rect 35076 29348 35100 29350
rect 35156 29348 35180 29350
rect 34940 29328 35236 29348
rect 34940 28316 35236 28336
rect 34996 28314 35020 28316
rect 35076 28314 35100 28316
rect 35156 28314 35180 28316
rect 35018 28262 35020 28314
rect 35082 28262 35094 28314
rect 35156 28262 35158 28314
rect 34996 28260 35020 28262
rect 35076 28260 35100 28262
rect 35156 28260 35180 28262
rect 34940 28240 35236 28260
rect 34058 27568 34114 27577
rect 34058 27503 34114 27512
rect 34702 27568 34758 27577
rect 34702 27503 34758 27512
rect 33782 23624 33838 23633
rect 33782 23559 33838 23568
rect 34518 17912 34574 17921
rect 34518 17847 34574 17856
rect 34532 13705 34560 17847
rect 34518 13696 34574 13705
rect 34518 13631 34574 13640
rect 32126 12472 32182 12481
rect 32126 12407 32182 12416
rect 33138 12472 33194 12481
rect 34716 12442 34744 27503
rect 34940 27228 35236 27248
rect 34996 27226 35020 27228
rect 35076 27226 35100 27228
rect 35156 27226 35180 27228
rect 35018 27174 35020 27226
rect 35082 27174 35094 27226
rect 35156 27174 35158 27226
rect 34996 27172 35020 27174
rect 35076 27172 35100 27174
rect 35156 27172 35180 27174
rect 34940 27152 35236 27172
rect 34940 26140 35236 26160
rect 34996 26138 35020 26140
rect 35076 26138 35100 26140
rect 35156 26138 35180 26140
rect 35018 26086 35020 26138
rect 35082 26086 35094 26138
rect 35156 26086 35158 26138
rect 34996 26084 35020 26086
rect 35076 26084 35100 26086
rect 35156 26084 35180 26086
rect 34940 26064 35236 26084
rect 34940 25052 35236 25072
rect 34996 25050 35020 25052
rect 35076 25050 35100 25052
rect 35156 25050 35180 25052
rect 35018 24998 35020 25050
rect 35082 24998 35094 25050
rect 35156 24998 35158 25050
rect 34996 24996 35020 24998
rect 35076 24996 35100 24998
rect 35156 24996 35180 24998
rect 34940 24976 35236 24996
rect 34940 23964 35236 23984
rect 34996 23962 35020 23964
rect 35076 23962 35100 23964
rect 35156 23962 35180 23964
rect 35018 23910 35020 23962
rect 35082 23910 35094 23962
rect 35156 23910 35158 23962
rect 34996 23908 35020 23910
rect 35076 23908 35100 23910
rect 35156 23908 35180 23910
rect 34940 23888 35236 23908
rect 34940 22876 35236 22896
rect 34996 22874 35020 22876
rect 35076 22874 35100 22876
rect 35156 22874 35180 22876
rect 35018 22822 35020 22874
rect 35082 22822 35094 22874
rect 35156 22822 35158 22874
rect 34996 22820 35020 22822
rect 35076 22820 35100 22822
rect 35156 22820 35180 22822
rect 34940 22800 35236 22820
rect 34940 21788 35236 21808
rect 34996 21786 35020 21788
rect 35076 21786 35100 21788
rect 35156 21786 35180 21788
rect 35018 21734 35020 21786
rect 35082 21734 35094 21786
rect 35156 21734 35158 21786
rect 34996 21732 35020 21734
rect 35076 21732 35100 21734
rect 35156 21732 35180 21734
rect 34940 21712 35236 21732
rect 34940 20700 35236 20720
rect 34996 20698 35020 20700
rect 35076 20698 35100 20700
rect 35156 20698 35180 20700
rect 35018 20646 35020 20698
rect 35082 20646 35094 20698
rect 35156 20646 35158 20698
rect 34996 20644 35020 20646
rect 35076 20644 35100 20646
rect 35156 20644 35180 20646
rect 34940 20624 35236 20644
rect 34940 19612 35236 19632
rect 34996 19610 35020 19612
rect 35076 19610 35100 19612
rect 35156 19610 35180 19612
rect 35018 19558 35020 19610
rect 35082 19558 35094 19610
rect 35156 19558 35158 19610
rect 34996 19556 35020 19558
rect 35076 19556 35100 19558
rect 35156 19556 35180 19558
rect 34940 19536 35236 19556
rect 34940 18524 35236 18544
rect 34996 18522 35020 18524
rect 35076 18522 35100 18524
rect 35156 18522 35180 18524
rect 35018 18470 35020 18522
rect 35082 18470 35094 18522
rect 35156 18470 35158 18522
rect 34996 18468 35020 18470
rect 35076 18468 35100 18470
rect 35156 18468 35180 18470
rect 34940 18448 35236 18468
rect 35268 17785 35296 53887
rect 35360 51898 35388 58511
rect 35820 57390 35848 58822
rect 35808 57384 35860 57390
rect 35808 57326 35860 57332
rect 35900 57248 35952 57254
rect 35900 57190 35952 57196
rect 35438 56808 35494 56817
rect 35438 56743 35494 56752
rect 35452 55185 35480 56743
rect 35530 56536 35586 56545
rect 35530 56471 35586 56480
rect 35438 55176 35494 55185
rect 35438 55111 35494 55120
rect 35438 53816 35494 53825
rect 35438 53751 35494 53760
rect 35452 52057 35480 53751
rect 35438 52048 35494 52057
rect 35438 51983 35494 51992
rect 35360 51870 35480 51898
rect 35452 50726 35480 51870
rect 35440 50720 35492 50726
rect 35440 50662 35492 50668
rect 35438 50552 35494 50561
rect 35438 50487 35494 50496
rect 35452 48385 35480 50487
rect 35438 48376 35494 48385
rect 35438 48311 35494 48320
rect 35346 43616 35402 43625
rect 35346 43551 35402 43560
rect 35360 40633 35388 43551
rect 35544 40769 35572 56471
rect 35912 55264 35940 57190
rect 35820 55236 35940 55264
rect 35820 52494 35848 55236
rect 35808 52488 35860 52494
rect 35808 52430 35860 52436
rect 35622 48648 35678 48657
rect 35622 48583 35678 48592
rect 35636 47025 35664 48583
rect 35622 47016 35678 47025
rect 35622 46951 35678 46960
rect 37646 45520 37702 45529
rect 37646 45455 37702 45464
rect 37660 44538 37688 45455
rect 37648 44532 37700 44538
rect 37648 44474 37700 44480
rect 36084 44328 36136 44334
rect 36084 44270 36136 44276
rect 36360 44328 36412 44334
rect 36360 44270 36412 44276
rect 36096 43994 36124 44270
rect 36084 43988 36136 43994
rect 36084 43930 36136 43936
rect 35622 41168 35678 41177
rect 35622 41103 35678 41112
rect 35530 40760 35586 40769
rect 35530 40695 35586 40704
rect 35346 40624 35402 40633
rect 35346 40559 35402 40568
rect 35532 40588 35584 40594
rect 35532 40530 35584 40536
rect 35440 40520 35492 40526
rect 35440 40462 35492 40468
rect 35452 40186 35480 40462
rect 35440 40180 35492 40186
rect 35440 40122 35492 40128
rect 35544 40118 35572 40530
rect 35532 40112 35584 40118
rect 35532 40054 35584 40060
rect 35636 38185 35664 41103
rect 35716 40384 35768 40390
rect 35716 40326 35768 40332
rect 35728 39506 35756 40326
rect 35716 39500 35768 39506
rect 35716 39442 35768 39448
rect 35728 39098 35756 39442
rect 35716 39092 35768 39098
rect 35716 39034 35768 39040
rect 35622 38176 35678 38185
rect 35622 38111 35678 38120
rect 35530 37224 35586 37233
rect 35530 37159 35586 37168
rect 35438 35456 35494 35465
rect 35438 35391 35494 35400
rect 35452 34241 35480 35391
rect 35438 34232 35494 34241
rect 35438 34167 35494 34176
rect 35544 33425 35572 37159
rect 35530 33416 35586 33425
rect 35530 33351 35586 33360
rect 35346 27432 35402 27441
rect 35346 27367 35402 27376
rect 35254 17776 35310 17785
rect 35254 17711 35310 17720
rect 34940 17436 35236 17456
rect 34996 17434 35020 17436
rect 35076 17434 35100 17436
rect 35156 17434 35180 17436
rect 35018 17382 35020 17434
rect 35082 17382 35094 17434
rect 35156 17382 35158 17434
rect 34996 17380 35020 17382
rect 35076 17380 35100 17382
rect 35156 17380 35180 17382
rect 34940 17360 35236 17380
rect 35360 16425 35388 27367
rect 36372 26353 36400 44270
rect 35806 26344 35862 26353
rect 35806 26279 35862 26288
rect 36358 26344 36414 26353
rect 36358 26279 36414 26288
rect 35622 20496 35678 20505
rect 35622 20431 35678 20440
rect 35438 19952 35494 19961
rect 35438 19887 35494 19896
rect 35346 16416 35402 16425
rect 34940 16348 35236 16368
rect 35346 16351 35402 16360
rect 34996 16346 35020 16348
rect 35076 16346 35100 16348
rect 35156 16346 35180 16348
rect 35018 16294 35020 16346
rect 35082 16294 35094 16346
rect 35156 16294 35158 16346
rect 34996 16292 35020 16294
rect 35076 16292 35100 16294
rect 35156 16292 35180 16294
rect 34940 16272 35236 16292
rect 34940 15260 35236 15280
rect 34996 15258 35020 15260
rect 35076 15258 35100 15260
rect 35156 15258 35180 15260
rect 35018 15206 35020 15258
rect 35082 15206 35094 15258
rect 35156 15206 35158 15258
rect 34996 15204 35020 15206
rect 35076 15204 35100 15206
rect 35156 15204 35180 15206
rect 34940 15184 35236 15204
rect 34940 14172 35236 14192
rect 34996 14170 35020 14172
rect 35076 14170 35100 14172
rect 35156 14170 35180 14172
rect 35018 14118 35020 14170
rect 35082 14118 35094 14170
rect 35156 14118 35158 14170
rect 34996 14116 35020 14118
rect 35076 14116 35100 14118
rect 35156 14116 35180 14118
rect 34940 14096 35236 14116
rect 34940 13084 35236 13104
rect 34996 13082 35020 13084
rect 35076 13082 35100 13084
rect 35156 13082 35180 13084
rect 35018 13030 35020 13082
rect 35082 13030 35094 13082
rect 35156 13030 35158 13082
rect 34996 13028 35020 13030
rect 35076 13028 35100 13030
rect 35156 13028 35180 13030
rect 34940 13008 35236 13028
rect 33138 12407 33194 12416
rect 34704 12436 34756 12442
rect 32678 5264 32734 5273
rect 32678 5199 32734 5208
rect 32692 800 32720 5199
rect 33152 4826 33180 12407
rect 34704 12378 34756 12384
rect 35348 12436 35400 12442
rect 35348 12378 35400 12384
rect 34940 11996 35236 12016
rect 34996 11994 35020 11996
rect 35076 11994 35100 11996
rect 35156 11994 35180 11996
rect 35018 11942 35020 11994
rect 35082 11942 35094 11994
rect 35156 11942 35158 11994
rect 34996 11940 35020 11942
rect 35076 11940 35100 11942
rect 35156 11940 35180 11942
rect 34940 11920 35236 11940
rect 34940 10908 35236 10928
rect 34996 10906 35020 10908
rect 35076 10906 35100 10908
rect 35156 10906 35180 10908
rect 35018 10854 35020 10906
rect 35082 10854 35094 10906
rect 35156 10854 35158 10906
rect 34996 10852 35020 10854
rect 35076 10852 35100 10854
rect 35156 10852 35180 10854
rect 34940 10832 35236 10852
rect 35360 10826 35388 12378
rect 35452 10985 35480 19887
rect 35636 13569 35664 20431
rect 35622 13560 35678 13569
rect 35622 13495 35678 13504
rect 35438 10976 35494 10985
rect 35438 10911 35494 10920
rect 35360 10798 35480 10826
rect 34940 9820 35236 9840
rect 34996 9818 35020 9820
rect 35076 9818 35100 9820
rect 35156 9818 35180 9820
rect 35018 9766 35020 9818
rect 35082 9766 35094 9818
rect 35156 9766 35158 9818
rect 34996 9764 35020 9766
rect 35076 9764 35100 9766
rect 35156 9764 35180 9766
rect 34940 9744 35236 9764
rect 34940 8732 35236 8752
rect 34996 8730 35020 8732
rect 35076 8730 35100 8732
rect 35156 8730 35180 8732
rect 35018 8678 35020 8730
rect 35082 8678 35094 8730
rect 35156 8678 35158 8730
rect 34996 8676 35020 8678
rect 35076 8676 35100 8678
rect 35156 8676 35180 8678
rect 34940 8656 35236 8676
rect 34940 7644 35236 7664
rect 34996 7642 35020 7644
rect 35076 7642 35100 7644
rect 35156 7642 35180 7644
rect 35018 7590 35020 7642
rect 35082 7590 35094 7642
rect 35156 7590 35158 7642
rect 34996 7588 35020 7590
rect 35076 7588 35100 7590
rect 35156 7588 35180 7590
rect 34518 7576 34574 7585
rect 34940 7568 35236 7588
rect 34518 7511 34574 7520
rect 33140 4820 33192 4826
rect 33140 4762 33192 4768
rect 33508 4820 33560 4826
rect 33508 4762 33560 4768
rect 33520 2666 33548 4762
rect 33520 2638 33640 2666
rect 33612 800 33640 2638
rect 34532 800 34560 7511
rect 34940 6556 35236 6576
rect 34996 6554 35020 6556
rect 35076 6554 35100 6556
rect 35156 6554 35180 6556
rect 35018 6502 35020 6554
rect 35082 6502 35094 6554
rect 35156 6502 35158 6554
rect 34996 6500 35020 6502
rect 35076 6500 35100 6502
rect 35156 6500 35180 6502
rect 34940 6480 35236 6500
rect 34940 5468 35236 5488
rect 34996 5466 35020 5468
rect 35076 5466 35100 5468
rect 35156 5466 35180 5468
rect 35018 5414 35020 5466
rect 35082 5414 35094 5466
rect 35156 5414 35158 5466
rect 34996 5412 35020 5414
rect 35076 5412 35100 5414
rect 35156 5412 35180 5414
rect 34940 5392 35236 5412
rect 34940 4380 35236 4400
rect 34996 4378 35020 4380
rect 35076 4378 35100 4380
rect 35156 4378 35180 4380
rect 35018 4326 35020 4378
rect 35082 4326 35094 4378
rect 35156 4326 35158 4378
rect 34996 4324 35020 4326
rect 35076 4324 35100 4326
rect 35156 4324 35180 4326
rect 34940 4304 35236 4324
rect 34940 3292 35236 3312
rect 34996 3290 35020 3292
rect 35076 3290 35100 3292
rect 35156 3290 35180 3292
rect 35018 3238 35020 3290
rect 35082 3238 35094 3290
rect 35156 3238 35158 3290
rect 34996 3236 35020 3238
rect 35076 3236 35100 3238
rect 35156 3236 35180 3238
rect 34940 3216 35236 3236
rect 34940 2204 35236 2224
rect 34996 2202 35020 2204
rect 35076 2202 35100 2204
rect 35156 2202 35180 2204
rect 35018 2150 35020 2202
rect 35082 2150 35094 2202
rect 35156 2150 35158 2202
rect 34996 2148 35020 2150
rect 35076 2148 35100 2150
rect 35156 2148 35180 2150
rect 34940 2128 35236 2148
rect 35452 800 35480 10798
rect 35820 3505 35848 26279
rect 37738 20360 37794 20369
rect 37738 20295 37794 20304
rect 37370 15872 37426 15881
rect 37370 15807 37426 15816
rect 36358 9072 36414 9081
rect 36358 9007 36414 9016
rect 36266 6352 36322 6361
rect 36266 6287 36268 6296
rect 36320 6287 36322 6296
rect 36268 6258 36320 6264
rect 35992 6248 36044 6254
rect 35992 6190 36044 6196
rect 36004 5710 36032 6190
rect 35992 5704 36044 5710
rect 35990 5672 35992 5681
rect 36044 5672 36046 5681
rect 35990 5607 36046 5616
rect 35806 3496 35862 3505
rect 35806 3431 35862 3440
rect 36372 800 36400 9007
rect 37384 6304 37412 15807
rect 37462 15056 37518 15065
rect 37462 14991 37518 15000
rect 37476 7750 37504 14991
rect 37554 13288 37610 13297
rect 37554 13223 37610 13232
rect 37464 7744 37516 7750
rect 37464 7686 37516 7692
rect 37568 7546 37596 13223
rect 37556 7540 37608 7546
rect 37556 7482 37608 7488
rect 37292 6276 37412 6304
rect 37292 800 37320 6276
rect 37370 6216 37426 6225
rect 37370 6151 37426 6160
rect 37384 6118 37412 6151
rect 37372 6112 37424 6118
rect 37372 6054 37424 6060
rect 37752 2802 37780 20295
rect 39580 7744 39632 7750
rect 39580 7686 39632 7692
rect 39120 7540 39172 7546
rect 39120 7482 39172 7488
rect 37752 2774 38056 2802
rect 38028 2530 38056 2774
rect 38028 2502 38240 2530
rect 38212 800 38240 2502
rect 39132 800 39160 7482
rect 39592 800 39620 7686
rect 22742 232 22798 241
rect 22742 167 22798 176
rect 23478 0 23534 800
rect 23938 0 23994 800
rect 24858 0 24914 800
rect 25778 0 25834 800
rect 26698 0 26754 800
rect 27618 0 27674 800
rect 28538 0 28594 800
rect 29458 0 29514 800
rect 30378 0 30434 800
rect 31298 0 31354 800
rect 31758 0 31814 800
rect 32678 0 32734 800
rect 33598 0 33654 800
rect 34518 0 34574 800
rect 35438 0 35494 800
rect 36358 0 36414 800
rect 37278 0 37334 800
rect 38198 0 38254 800
rect 39118 0 39174 800
rect 39578 0 39634 800
<< via2 >>
rect 3974 79600 4030 79656
rect 478 75792 534 75848
rect 1674 75792 1730 75848
rect 110 69808 166 69864
rect 1582 66680 1638 66736
rect 2410 76880 2466 76936
rect 1858 75384 1914 75440
rect 1858 63980 1914 64016
rect 1858 63960 1860 63980
rect 1860 63960 1912 63980
rect 1912 63960 1914 63980
rect 1858 59880 1914 59936
rect 1306 46008 1362 46064
rect 1766 46280 1822 46336
rect 2042 44276 2044 44296
rect 2044 44276 2096 44296
rect 2096 44276 2098 44296
rect 2042 44240 2098 44276
rect 3330 75520 3386 75576
rect 3238 69400 3294 69456
rect 2870 65320 2926 65376
rect 1950 40568 2006 40624
rect 1582 39516 1584 39536
rect 1584 39516 1636 39536
rect 1636 39516 1638 39536
rect 1582 39480 1638 39516
rect 1858 29280 1914 29336
rect 1582 26560 1638 26616
rect 1766 19080 1822 19136
rect 1398 16904 1454 16960
rect 1582 15308 1584 15328
rect 1584 15308 1636 15328
rect 1636 15308 1638 15328
rect 1582 15272 1638 15308
rect 2778 38120 2834 38176
rect 3054 46144 3110 46200
rect 3054 43288 3110 43344
rect 3054 36760 3110 36816
rect 2962 36488 3018 36544
rect 2686 23296 2742 23352
rect 3146 23296 3202 23352
rect 2226 16496 2282 16552
rect 2870 19080 2926 19136
rect 1950 13776 2006 13832
rect 2778 13640 2834 13696
rect 2778 12280 2834 12336
rect 2778 11736 2834 11792
rect 2686 10512 2742 10568
rect 2042 10124 2098 10160
rect 2042 10104 2044 10124
rect 2044 10104 2096 10124
rect 2096 10104 2098 10124
rect 1582 8880 1638 8936
rect 1398 7792 1454 7848
rect 35438 79600 35494 79656
rect 4066 78240 4122 78296
rect 4220 77274 4276 77276
rect 4300 77274 4356 77276
rect 4380 77274 4436 77276
rect 4460 77274 4516 77276
rect 4220 77222 4246 77274
rect 4246 77222 4276 77274
rect 4300 77222 4310 77274
rect 4310 77222 4356 77274
rect 4380 77222 4426 77274
rect 4426 77222 4436 77274
rect 4460 77222 4490 77274
rect 4490 77222 4516 77274
rect 4220 77220 4276 77222
rect 4300 77220 4356 77222
rect 4380 77220 4436 77222
rect 4460 77220 4516 77222
rect 4220 76186 4276 76188
rect 4300 76186 4356 76188
rect 4380 76186 4436 76188
rect 4460 76186 4516 76188
rect 4220 76134 4246 76186
rect 4246 76134 4276 76186
rect 4300 76134 4310 76186
rect 4310 76134 4356 76186
rect 4380 76134 4426 76186
rect 4426 76134 4436 76186
rect 4460 76134 4490 76186
rect 4490 76134 4516 76186
rect 4220 76132 4276 76134
rect 4300 76132 4356 76134
rect 4380 76132 4436 76134
rect 4460 76132 4516 76134
rect 4220 75098 4276 75100
rect 4300 75098 4356 75100
rect 4380 75098 4436 75100
rect 4460 75098 4516 75100
rect 4220 75046 4246 75098
rect 4246 75046 4276 75098
rect 4300 75046 4310 75098
rect 4310 75046 4356 75098
rect 4380 75046 4426 75098
rect 4426 75046 4436 75098
rect 4460 75046 4490 75098
rect 4490 75046 4516 75098
rect 4220 75044 4276 75046
rect 4300 75044 4356 75046
rect 4380 75044 4436 75046
rect 4460 75044 4516 75046
rect 3790 74160 3846 74216
rect 3790 72528 3846 72584
rect 3330 68176 3386 68232
rect 3422 68040 3478 68096
rect 4618 74704 4674 74760
rect 4220 74010 4276 74012
rect 4300 74010 4356 74012
rect 4380 74010 4436 74012
rect 4460 74010 4516 74012
rect 4220 73958 4246 74010
rect 4246 73958 4276 74010
rect 4300 73958 4310 74010
rect 4310 73958 4356 74010
rect 4380 73958 4426 74010
rect 4426 73958 4436 74010
rect 4460 73958 4490 74010
rect 4490 73958 4516 74010
rect 4220 73956 4276 73958
rect 4300 73956 4356 73958
rect 4380 73956 4436 73958
rect 4460 73956 4516 73958
rect 4220 72922 4276 72924
rect 4300 72922 4356 72924
rect 4380 72922 4436 72924
rect 4460 72922 4516 72924
rect 4220 72870 4246 72922
rect 4246 72870 4276 72922
rect 4300 72870 4310 72922
rect 4310 72870 4356 72922
rect 4380 72870 4426 72922
rect 4426 72870 4436 72922
rect 4460 72870 4490 72922
rect 4490 72870 4516 72922
rect 4220 72868 4276 72870
rect 4300 72868 4356 72870
rect 4380 72868 4436 72870
rect 4460 72868 4516 72870
rect 4066 72800 4122 72856
rect 4066 71984 4122 72040
rect 4220 71834 4276 71836
rect 4300 71834 4356 71836
rect 4380 71834 4436 71836
rect 4460 71834 4516 71836
rect 4220 71782 4246 71834
rect 4246 71782 4276 71834
rect 4300 71782 4310 71834
rect 4310 71782 4356 71834
rect 4380 71782 4426 71834
rect 4426 71782 4436 71834
rect 4460 71782 4490 71834
rect 4490 71782 4516 71834
rect 4220 71780 4276 71782
rect 4300 71780 4356 71782
rect 4380 71780 4436 71782
rect 4460 71780 4516 71782
rect 4802 71576 4858 71632
rect 4802 70760 4858 70816
rect 4220 70746 4276 70748
rect 4300 70746 4356 70748
rect 4380 70746 4436 70748
rect 4460 70746 4516 70748
rect 4220 70694 4246 70746
rect 4246 70694 4276 70746
rect 4300 70694 4310 70746
rect 4310 70694 4356 70746
rect 4380 70694 4426 70746
rect 4426 70694 4436 70746
rect 4460 70694 4490 70746
rect 4490 70694 4516 70746
rect 4220 70692 4276 70694
rect 4300 70692 4356 70694
rect 4380 70692 4436 70694
rect 4460 70692 4516 70694
rect 4894 70080 4950 70136
rect 4220 69658 4276 69660
rect 4300 69658 4356 69660
rect 4380 69658 4436 69660
rect 4460 69658 4516 69660
rect 4220 69606 4246 69658
rect 4246 69606 4276 69658
rect 4300 69606 4310 69658
rect 4310 69606 4356 69658
rect 4380 69606 4426 69658
rect 4426 69606 4436 69658
rect 4460 69606 4490 69658
rect 4490 69606 4516 69658
rect 4220 69604 4276 69606
rect 4300 69604 4356 69606
rect 4380 69604 4436 69606
rect 4460 69604 4516 69606
rect 4220 68570 4276 68572
rect 4300 68570 4356 68572
rect 4380 68570 4436 68572
rect 4460 68570 4516 68572
rect 4220 68518 4246 68570
rect 4246 68518 4276 68570
rect 4300 68518 4310 68570
rect 4310 68518 4356 68570
rect 4380 68518 4426 68570
rect 4426 68518 4436 68570
rect 4460 68518 4490 68570
rect 4490 68518 4516 68570
rect 4220 68516 4276 68518
rect 4300 68516 4356 68518
rect 4380 68516 4436 68518
rect 4460 68516 4516 68518
rect 4220 67482 4276 67484
rect 4300 67482 4356 67484
rect 4380 67482 4436 67484
rect 4460 67482 4516 67484
rect 4220 67430 4246 67482
rect 4246 67430 4276 67482
rect 4300 67430 4310 67482
rect 4310 67430 4356 67482
rect 4380 67430 4426 67482
rect 4426 67430 4436 67482
rect 4460 67430 4490 67482
rect 4490 67430 4516 67482
rect 4220 67428 4276 67430
rect 4300 67428 4356 67430
rect 4380 67428 4436 67430
rect 4460 67428 4516 67430
rect 3974 67088 4030 67144
rect 4220 66394 4276 66396
rect 4300 66394 4356 66396
rect 4380 66394 4436 66396
rect 4460 66394 4516 66396
rect 4220 66342 4246 66394
rect 4246 66342 4276 66394
rect 4300 66342 4310 66394
rect 4310 66342 4356 66394
rect 4380 66342 4426 66394
rect 4426 66342 4436 66394
rect 4460 66342 4490 66394
rect 4490 66342 4516 66394
rect 4220 66340 4276 66342
rect 4300 66340 4356 66342
rect 4380 66340 4436 66342
rect 4460 66340 4516 66342
rect 4220 65306 4276 65308
rect 4300 65306 4356 65308
rect 4380 65306 4436 65308
rect 4460 65306 4516 65308
rect 4220 65254 4246 65306
rect 4246 65254 4276 65306
rect 4300 65254 4310 65306
rect 4310 65254 4356 65306
rect 4380 65254 4426 65306
rect 4426 65254 4436 65306
rect 4460 65254 4490 65306
rect 4490 65254 4516 65306
rect 4220 65252 4276 65254
rect 4300 65252 4356 65254
rect 4380 65252 4436 65254
rect 4460 65252 4516 65254
rect 4220 64218 4276 64220
rect 4300 64218 4356 64220
rect 4380 64218 4436 64220
rect 4460 64218 4516 64220
rect 4220 64166 4246 64218
rect 4246 64166 4276 64218
rect 4300 64166 4310 64218
rect 4310 64166 4356 64218
rect 4380 64166 4426 64218
rect 4426 64166 4436 64218
rect 4460 64166 4490 64218
rect 4490 64166 4516 64218
rect 4220 64164 4276 64166
rect 4300 64164 4356 64166
rect 4380 64164 4436 64166
rect 4460 64164 4516 64166
rect 4158 63960 4214 64016
rect 4220 63130 4276 63132
rect 4300 63130 4356 63132
rect 4380 63130 4436 63132
rect 4460 63130 4516 63132
rect 4220 63078 4246 63130
rect 4246 63078 4276 63130
rect 4300 63078 4310 63130
rect 4310 63078 4356 63130
rect 4380 63078 4426 63130
rect 4426 63078 4436 63130
rect 4460 63078 4490 63130
rect 4490 63078 4516 63130
rect 4220 63076 4276 63078
rect 4300 63076 4356 63078
rect 4380 63076 4436 63078
rect 4460 63076 4516 63078
rect 4220 62042 4276 62044
rect 4300 62042 4356 62044
rect 4380 62042 4436 62044
rect 4460 62042 4516 62044
rect 4220 61990 4246 62042
rect 4246 61990 4276 62042
rect 4300 61990 4310 62042
rect 4310 61990 4356 62042
rect 4380 61990 4426 62042
rect 4426 61990 4436 62042
rect 4460 61990 4490 62042
rect 4490 61990 4516 62042
rect 4220 61988 4276 61990
rect 4300 61988 4356 61990
rect 4380 61988 4436 61990
rect 4460 61988 4516 61990
rect 4220 60954 4276 60956
rect 4300 60954 4356 60956
rect 4380 60954 4436 60956
rect 4460 60954 4516 60956
rect 4220 60902 4246 60954
rect 4246 60902 4276 60954
rect 4300 60902 4310 60954
rect 4310 60902 4356 60954
rect 4380 60902 4426 60954
rect 4426 60902 4436 60954
rect 4460 60902 4490 60954
rect 4490 60902 4516 60954
rect 4220 60900 4276 60902
rect 4300 60900 4356 60902
rect 4380 60900 4436 60902
rect 4460 60900 4516 60902
rect 3422 60560 3478 60616
rect 6458 75112 6514 75168
rect 7378 74840 7434 74896
rect 6182 74704 6238 74760
rect 5630 69536 5686 69592
rect 4894 59880 4950 59936
rect 4220 59866 4276 59868
rect 4300 59866 4356 59868
rect 4380 59866 4436 59868
rect 4460 59866 4516 59868
rect 4220 59814 4246 59866
rect 4246 59814 4276 59866
rect 4300 59814 4310 59866
rect 4310 59814 4356 59866
rect 4380 59814 4426 59866
rect 4426 59814 4436 59866
rect 4460 59814 4490 59866
rect 4490 59814 4516 59866
rect 4220 59812 4276 59814
rect 4300 59812 4356 59814
rect 4380 59812 4436 59814
rect 4460 59812 4516 59814
rect 4220 58778 4276 58780
rect 4300 58778 4356 58780
rect 4380 58778 4436 58780
rect 4460 58778 4516 58780
rect 4220 58726 4246 58778
rect 4246 58726 4276 58778
rect 4300 58726 4310 58778
rect 4310 58726 4356 58778
rect 4380 58726 4426 58778
rect 4426 58726 4436 58778
rect 4460 58726 4490 58778
rect 4490 58726 4516 58778
rect 4220 58724 4276 58726
rect 4300 58724 4356 58726
rect 4380 58724 4436 58726
rect 4460 58724 4516 58726
rect 4220 57690 4276 57692
rect 4300 57690 4356 57692
rect 4380 57690 4436 57692
rect 4460 57690 4516 57692
rect 4220 57638 4246 57690
rect 4246 57638 4276 57690
rect 4300 57638 4310 57690
rect 4310 57638 4356 57690
rect 4380 57638 4426 57690
rect 4426 57638 4436 57690
rect 4460 57638 4490 57690
rect 4490 57638 4516 57690
rect 4220 57636 4276 57638
rect 4300 57636 4356 57638
rect 4380 57636 4436 57638
rect 4460 57636 4516 57638
rect 4220 56602 4276 56604
rect 4300 56602 4356 56604
rect 4380 56602 4436 56604
rect 4460 56602 4516 56604
rect 4220 56550 4246 56602
rect 4246 56550 4276 56602
rect 4300 56550 4310 56602
rect 4310 56550 4356 56602
rect 4380 56550 4426 56602
rect 4426 56550 4436 56602
rect 4460 56550 4490 56602
rect 4490 56550 4516 56602
rect 4220 56548 4276 56550
rect 4300 56548 4356 56550
rect 4380 56548 4436 56550
rect 4460 56548 4516 56550
rect 3882 56344 3938 56400
rect 3330 55120 3386 55176
rect 3698 53760 3754 53816
rect 3330 53080 3386 53136
rect 3330 52400 3386 52456
rect 3330 49544 3386 49600
rect 3514 48592 3570 48648
rect 4220 55514 4276 55516
rect 4300 55514 4356 55516
rect 4380 55514 4436 55516
rect 4460 55514 4516 55516
rect 4220 55462 4246 55514
rect 4246 55462 4276 55514
rect 4300 55462 4310 55514
rect 4310 55462 4356 55514
rect 4380 55462 4426 55514
rect 4426 55462 4436 55514
rect 4460 55462 4490 55514
rect 4490 55462 4516 55514
rect 4220 55460 4276 55462
rect 4300 55460 4356 55462
rect 4380 55460 4436 55462
rect 4460 55460 4516 55462
rect 4220 54426 4276 54428
rect 4300 54426 4356 54428
rect 4380 54426 4436 54428
rect 4460 54426 4516 54428
rect 4220 54374 4246 54426
rect 4246 54374 4276 54426
rect 4300 54374 4310 54426
rect 4310 54374 4356 54426
rect 4380 54374 4426 54426
rect 4426 54374 4436 54426
rect 4460 54374 4490 54426
rect 4490 54374 4516 54426
rect 4220 54372 4276 54374
rect 4300 54372 4356 54374
rect 4380 54372 4436 54374
rect 4460 54372 4516 54374
rect 4220 53338 4276 53340
rect 4300 53338 4356 53340
rect 4380 53338 4436 53340
rect 4460 53338 4516 53340
rect 4220 53286 4246 53338
rect 4246 53286 4276 53338
rect 4300 53286 4310 53338
rect 4310 53286 4356 53338
rect 4380 53286 4426 53338
rect 4426 53286 4436 53338
rect 4460 53286 4490 53338
rect 4490 53286 4516 53338
rect 4220 53284 4276 53286
rect 4300 53284 4356 53286
rect 4380 53284 4436 53286
rect 4460 53284 4516 53286
rect 4220 52250 4276 52252
rect 4300 52250 4356 52252
rect 4380 52250 4436 52252
rect 4460 52250 4516 52252
rect 4220 52198 4246 52250
rect 4246 52198 4276 52250
rect 4300 52198 4310 52250
rect 4310 52198 4356 52250
rect 4380 52198 4426 52250
rect 4426 52198 4436 52250
rect 4460 52198 4490 52250
rect 4490 52198 4516 52250
rect 4220 52196 4276 52198
rect 4300 52196 4356 52198
rect 4380 52196 4436 52198
rect 4460 52196 4516 52198
rect 4220 51162 4276 51164
rect 4300 51162 4356 51164
rect 4380 51162 4436 51164
rect 4460 51162 4516 51164
rect 4220 51110 4246 51162
rect 4246 51110 4276 51162
rect 4300 51110 4310 51162
rect 4310 51110 4356 51162
rect 4380 51110 4426 51162
rect 4426 51110 4436 51162
rect 4460 51110 4490 51162
rect 4490 51110 4516 51162
rect 4220 51108 4276 51110
rect 4300 51108 4356 51110
rect 4380 51108 4436 51110
rect 4460 51108 4516 51110
rect 4220 50074 4276 50076
rect 4300 50074 4356 50076
rect 4380 50074 4436 50076
rect 4460 50074 4516 50076
rect 4220 50022 4246 50074
rect 4246 50022 4276 50074
rect 4300 50022 4310 50074
rect 4310 50022 4356 50074
rect 4380 50022 4426 50074
rect 4426 50022 4436 50074
rect 4460 50022 4490 50074
rect 4490 50022 4516 50074
rect 4220 50020 4276 50022
rect 4300 50020 4356 50022
rect 4380 50020 4436 50022
rect 4460 50020 4516 50022
rect 5170 62056 5226 62112
rect 7378 69808 7434 69864
rect 6182 54440 6238 54496
rect 4066 49680 4122 49736
rect 5078 49680 5134 49736
rect 4220 48986 4276 48988
rect 4300 48986 4356 48988
rect 4380 48986 4436 48988
rect 4460 48986 4516 48988
rect 4220 48934 4246 48986
rect 4246 48934 4276 48986
rect 4300 48934 4310 48986
rect 4310 48934 4356 48986
rect 4380 48934 4426 48986
rect 4426 48934 4436 48986
rect 4460 48934 4490 48986
rect 4490 48934 4516 48986
rect 4220 48932 4276 48934
rect 4300 48932 4356 48934
rect 4380 48932 4436 48934
rect 4460 48932 4516 48934
rect 4066 48728 4122 48784
rect 3882 48320 3938 48376
rect 4220 47898 4276 47900
rect 4300 47898 4356 47900
rect 4380 47898 4436 47900
rect 4460 47898 4516 47900
rect 4220 47846 4246 47898
rect 4246 47846 4276 47898
rect 4300 47846 4310 47898
rect 4310 47846 4356 47898
rect 4380 47846 4426 47898
rect 4426 47846 4436 47898
rect 4460 47846 4490 47898
rect 4490 47846 4516 47898
rect 4220 47844 4276 47846
rect 4300 47844 4356 47846
rect 4380 47844 4436 47846
rect 4460 47844 4516 47846
rect 3514 46960 3570 47016
rect 3698 46960 3754 47016
rect 6274 46960 6330 47016
rect 4220 46810 4276 46812
rect 4300 46810 4356 46812
rect 4380 46810 4436 46812
rect 4460 46810 4516 46812
rect 4220 46758 4246 46810
rect 4246 46758 4276 46810
rect 4300 46758 4310 46810
rect 4310 46758 4356 46810
rect 4380 46758 4426 46810
rect 4426 46758 4436 46810
rect 4460 46758 4490 46810
rect 4490 46758 4516 46810
rect 4220 46756 4276 46758
rect 4300 46756 4356 46758
rect 4380 46756 4436 46758
rect 4460 46756 4516 46758
rect 4220 45722 4276 45724
rect 4300 45722 4356 45724
rect 4380 45722 4436 45724
rect 4460 45722 4516 45724
rect 4220 45670 4246 45722
rect 4246 45670 4276 45722
rect 4300 45670 4310 45722
rect 4310 45670 4356 45722
rect 4380 45670 4426 45722
rect 4426 45670 4436 45722
rect 4460 45670 4490 45722
rect 4490 45670 4516 45722
rect 4220 45668 4276 45670
rect 4300 45668 4356 45670
rect 4380 45668 4436 45670
rect 4460 45668 4516 45670
rect 4220 44634 4276 44636
rect 4300 44634 4356 44636
rect 4380 44634 4436 44636
rect 4460 44634 4516 44636
rect 4220 44582 4246 44634
rect 4246 44582 4276 44634
rect 4300 44582 4310 44634
rect 4310 44582 4356 44634
rect 4380 44582 4426 44634
rect 4426 44582 4436 44634
rect 4460 44582 4490 44634
rect 4490 44582 4516 44634
rect 4220 44580 4276 44582
rect 4300 44580 4356 44582
rect 4380 44580 4436 44582
rect 4460 44580 4516 44582
rect 4220 43546 4276 43548
rect 4300 43546 4356 43548
rect 4380 43546 4436 43548
rect 4460 43546 4516 43548
rect 4220 43494 4246 43546
rect 4246 43494 4276 43546
rect 4300 43494 4310 43546
rect 4310 43494 4356 43546
rect 4380 43494 4426 43546
rect 4426 43494 4436 43546
rect 4460 43494 4490 43546
rect 4490 43494 4516 43546
rect 4220 43492 4276 43494
rect 4300 43492 4356 43494
rect 4380 43492 4436 43494
rect 4460 43492 4516 43494
rect 4220 42458 4276 42460
rect 4300 42458 4356 42460
rect 4380 42458 4436 42460
rect 4460 42458 4516 42460
rect 4220 42406 4246 42458
rect 4246 42406 4276 42458
rect 4300 42406 4310 42458
rect 4310 42406 4356 42458
rect 4380 42406 4426 42458
rect 4426 42406 4436 42458
rect 4460 42406 4490 42458
rect 4490 42406 4516 42458
rect 4220 42404 4276 42406
rect 4300 42404 4356 42406
rect 4380 42404 4436 42406
rect 4460 42404 4516 42406
rect 5722 41792 5778 41848
rect 3882 40840 3938 40896
rect 3790 40704 3846 40760
rect 3514 37848 3570 37904
rect 3330 32000 3386 32056
rect 3330 30232 3386 30288
rect 3698 37304 3754 37360
rect 4220 41370 4276 41372
rect 4300 41370 4356 41372
rect 4380 41370 4436 41372
rect 4460 41370 4516 41372
rect 4220 41318 4246 41370
rect 4246 41318 4276 41370
rect 4300 41318 4310 41370
rect 4310 41318 4356 41370
rect 4380 41318 4426 41370
rect 4426 41318 4436 41370
rect 4460 41318 4490 41370
rect 4490 41318 4516 41370
rect 4220 41316 4276 41318
rect 4300 41316 4356 41318
rect 4380 41316 4436 41318
rect 4460 41316 4516 41318
rect 3974 40568 4030 40624
rect 4220 40282 4276 40284
rect 4300 40282 4356 40284
rect 4380 40282 4436 40284
rect 4460 40282 4516 40284
rect 4220 40230 4246 40282
rect 4246 40230 4276 40282
rect 4300 40230 4310 40282
rect 4310 40230 4356 40282
rect 4380 40230 4426 40282
rect 4426 40230 4436 40282
rect 4460 40230 4490 40282
rect 4490 40230 4516 40282
rect 4220 40228 4276 40230
rect 4300 40228 4356 40230
rect 4380 40228 4436 40230
rect 4460 40228 4516 40230
rect 4066 39616 4122 39672
rect 3882 39344 3938 39400
rect 4220 39194 4276 39196
rect 4300 39194 4356 39196
rect 4380 39194 4436 39196
rect 4460 39194 4516 39196
rect 4220 39142 4246 39194
rect 4246 39142 4276 39194
rect 4300 39142 4310 39194
rect 4310 39142 4356 39194
rect 4380 39142 4426 39194
rect 4426 39142 4436 39194
rect 4460 39142 4490 39194
rect 4490 39142 4516 39194
rect 4220 39140 4276 39142
rect 4300 39140 4356 39142
rect 4380 39140 4436 39142
rect 4460 39140 4516 39142
rect 4220 38106 4276 38108
rect 4300 38106 4356 38108
rect 4380 38106 4436 38108
rect 4460 38106 4516 38108
rect 4220 38054 4246 38106
rect 4246 38054 4276 38106
rect 4300 38054 4310 38106
rect 4310 38054 4356 38106
rect 4380 38054 4426 38106
rect 4426 38054 4436 38106
rect 4460 38054 4490 38106
rect 4490 38054 4516 38106
rect 4220 38052 4276 38054
rect 4300 38052 4356 38054
rect 4380 38052 4436 38054
rect 4460 38052 4516 38054
rect 4220 37018 4276 37020
rect 4300 37018 4356 37020
rect 4380 37018 4436 37020
rect 4460 37018 4516 37020
rect 4220 36966 4246 37018
rect 4246 36966 4276 37018
rect 4300 36966 4310 37018
rect 4310 36966 4356 37018
rect 4380 36966 4426 37018
rect 4426 36966 4436 37018
rect 4460 36966 4490 37018
rect 4490 36966 4516 37018
rect 4220 36964 4276 36966
rect 4300 36964 4356 36966
rect 4380 36964 4436 36966
rect 4460 36964 4516 36966
rect 3882 36080 3938 36136
rect 3790 35400 3846 35456
rect 4220 35930 4276 35932
rect 4300 35930 4356 35932
rect 4380 35930 4436 35932
rect 4460 35930 4516 35932
rect 4220 35878 4246 35930
rect 4246 35878 4276 35930
rect 4300 35878 4310 35930
rect 4310 35878 4356 35930
rect 4380 35878 4426 35930
rect 4426 35878 4436 35930
rect 4460 35878 4490 35930
rect 4490 35878 4516 35930
rect 4220 35876 4276 35878
rect 4300 35876 4356 35878
rect 4380 35876 4436 35878
rect 4460 35876 4516 35878
rect 4220 34842 4276 34844
rect 4300 34842 4356 34844
rect 4380 34842 4436 34844
rect 4460 34842 4516 34844
rect 4220 34790 4246 34842
rect 4246 34790 4276 34842
rect 4300 34790 4310 34842
rect 4310 34790 4356 34842
rect 4380 34790 4426 34842
rect 4426 34790 4436 34842
rect 4460 34790 4490 34842
rect 4490 34790 4516 34842
rect 4220 34788 4276 34790
rect 4300 34788 4356 34790
rect 4380 34788 4436 34790
rect 4460 34788 4516 34790
rect 3882 34720 3938 34776
rect 4220 33754 4276 33756
rect 4300 33754 4356 33756
rect 4380 33754 4436 33756
rect 4460 33754 4516 33756
rect 4220 33702 4246 33754
rect 4246 33702 4276 33754
rect 4300 33702 4310 33754
rect 4310 33702 4356 33754
rect 4380 33702 4426 33754
rect 4426 33702 4436 33754
rect 4460 33702 4490 33754
rect 4490 33702 4516 33754
rect 4220 33700 4276 33702
rect 4300 33700 4356 33702
rect 4380 33700 4436 33702
rect 4460 33700 4516 33702
rect 4220 32666 4276 32668
rect 4300 32666 4356 32668
rect 4380 32666 4436 32668
rect 4460 32666 4516 32668
rect 4220 32614 4246 32666
rect 4246 32614 4276 32666
rect 4300 32614 4310 32666
rect 4310 32614 4356 32666
rect 4380 32614 4426 32666
rect 4426 32614 4436 32666
rect 4460 32614 4490 32666
rect 4490 32614 4516 32666
rect 4220 32612 4276 32614
rect 4300 32612 4356 32614
rect 4380 32612 4436 32614
rect 4460 32612 4516 32614
rect 4220 31578 4276 31580
rect 4300 31578 4356 31580
rect 4380 31578 4436 31580
rect 4460 31578 4516 31580
rect 4220 31526 4246 31578
rect 4246 31526 4276 31578
rect 4300 31526 4310 31578
rect 4310 31526 4356 31578
rect 4380 31526 4426 31578
rect 4426 31526 4436 31578
rect 4460 31526 4490 31578
rect 4490 31526 4516 31578
rect 4220 31524 4276 31526
rect 4300 31524 4356 31526
rect 4380 31524 4436 31526
rect 4460 31524 4516 31526
rect 4066 30640 4122 30696
rect 4220 30490 4276 30492
rect 4300 30490 4356 30492
rect 4380 30490 4436 30492
rect 4460 30490 4516 30492
rect 4220 30438 4246 30490
rect 4246 30438 4276 30490
rect 4300 30438 4310 30490
rect 4310 30438 4356 30490
rect 4380 30438 4426 30490
rect 4426 30438 4436 30490
rect 4460 30438 4490 30490
rect 4490 30438 4516 30490
rect 4220 30436 4276 30438
rect 4300 30436 4356 30438
rect 4380 30436 4436 30438
rect 4460 30436 4516 30438
rect 4220 29402 4276 29404
rect 4300 29402 4356 29404
rect 4380 29402 4436 29404
rect 4460 29402 4516 29404
rect 4220 29350 4246 29402
rect 4246 29350 4276 29402
rect 4300 29350 4310 29402
rect 4310 29350 4356 29402
rect 4380 29350 4426 29402
rect 4426 29350 4436 29402
rect 4460 29350 4490 29402
rect 4490 29350 4516 29402
rect 4220 29348 4276 29350
rect 4300 29348 4356 29350
rect 4380 29348 4436 29350
rect 4460 29348 4516 29350
rect 4066 28872 4122 28928
rect 4220 28314 4276 28316
rect 4300 28314 4356 28316
rect 4380 28314 4436 28316
rect 4460 28314 4516 28316
rect 4220 28262 4246 28314
rect 4246 28262 4276 28314
rect 4300 28262 4310 28314
rect 4310 28262 4356 28314
rect 4380 28262 4426 28314
rect 4426 28262 4436 28314
rect 4460 28262 4490 28314
rect 4490 28262 4516 28314
rect 4220 28260 4276 28262
rect 4300 28260 4356 28262
rect 4380 28260 4436 28262
rect 4460 28260 4516 28262
rect 3698 27920 3754 27976
rect 4220 27226 4276 27228
rect 4300 27226 4356 27228
rect 4380 27226 4436 27228
rect 4460 27226 4516 27228
rect 4220 27174 4246 27226
rect 4246 27174 4276 27226
rect 4300 27174 4310 27226
rect 4310 27174 4356 27226
rect 4380 27174 4426 27226
rect 4426 27174 4436 27226
rect 4460 27174 4490 27226
rect 4490 27174 4516 27226
rect 4220 27172 4276 27174
rect 4300 27172 4356 27174
rect 4380 27172 4436 27174
rect 4460 27172 4516 27174
rect 4066 26288 4122 26344
rect 4220 26138 4276 26140
rect 4300 26138 4356 26140
rect 4380 26138 4436 26140
rect 4460 26138 4516 26140
rect 4220 26086 4246 26138
rect 4246 26086 4276 26138
rect 4300 26086 4310 26138
rect 4310 26086 4356 26138
rect 4380 26086 4426 26138
rect 4426 26086 4436 26138
rect 4460 26086 4490 26138
rect 4490 26086 4516 26138
rect 4220 26084 4276 26086
rect 4300 26084 4356 26086
rect 4380 26084 4436 26086
rect 4460 26084 4516 26086
rect 3514 25200 3570 25256
rect 4066 25200 4122 25256
rect 4220 25050 4276 25052
rect 4300 25050 4356 25052
rect 4380 25050 4436 25052
rect 4460 25050 4516 25052
rect 4220 24998 4246 25050
rect 4246 24998 4276 25050
rect 4300 24998 4310 25050
rect 4310 24998 4356 25050
rect 4380 24998 4426 25050
rect 4426 24998 4436 25050
rect 4460 24998 4490 25050
rect 4490 24998 4516 25050
rect 4220 24996 4276 24998
rect 4300 24996 4356 24998
rect 4380 24996 4436 24998
rect 4460 24996 4516 24998
rect 4220 23962 4276 23964
rect 4300 23962 4356 23964
rect 4380 23962 4436 23964
rect 4460 23962 4516 23964
rect 4220 23910 4246 23962
rect 4246 23910 4276 23962
rect 4300 23910 4310 23962
rect 4310 23910 4356 23962
rect 4380 23910 4426 23962
rect 4426 23910 4436 23962
rect 4460 23910 4490 23962
rect 4490 23910 4516 23962
rect 4220 23908 4276 23910
rect 4300 23908 4356 23910
rect 4380 23908 4436 23910
rect 4460 23908 4516 23910
rect 4066 23840 4122 23896
rect 4220 22874 4276 22876
rect 4300 22874 4356 22876
rect 4380 22874 4436 22876
rect 4460 22874 4516 22876
rect 4220 22822 4246 22874
rect 4246 22822 4276 22874
rect 4300 22822 4310 22874
rect 4310 22822 4356 22874
rect 4380 22822 4426 22874
rect 4426 22822 4436 22874
rect 4460 22822 4490 22874
rect 4490 22822 4516 22874
rect 4220 22820 4276 22822
rect 4300 22820 4356 22822
rect 4380 22820 4436 22822
rect 4460 22820 4516 22822
rect 4220 21786 4276 21788
rect 4300 21786 4356 21788
rect 4380 21786 4436 21788
rect 4460 21786 4516 21788
rect 4220 21734 4246 21786
rect 4246 21734 4276 21786
rect 4300 21734 4310 21786
rect 4310 21734 4356 21786
rect 4380 21734 4426 21786
rect 4426 21734 4436 21786
rect 4460 21734 4490 21786
rect 4490 21734 4516 21786
rect 4220 21732 4276 21734
rect 4300 21732 4356 21734
rect 4380 21732 4436 21734
rect 4460 21732 4516 21734
rect 4220 20698 4276 20700
rect 4300 20698 4356 20700
rect 4380 20698 4436 20700
rect 4460 20698 4516 20700
rect 4220 20646 4246 20698
rect 4246 20646 4276 20698
rect 4300 20646 4310 20698
rect 4310 20646 4356 20698
rect 4380 20646 4426 20698
rect 4426 20646 4436 20698
rect 4460 20646 4490 20698
rect 4490 20646 4516 20698
rect 4220 20644 4276 20646
rect 4300 20644 4356 20646
rect 4380 20644 4436 20646
rect 4460 20644 4516 20646
rect 4220 19610 4276 19612
rect 4300 19610 4356 19612
rect 4380 19610 4436 19612
rect 4460 19610 4516 19612
rect 4220 19558 4246 19610
rect 4246 19558 4276 19610
rect 4300 19558 4310 19610
rect 4310 19558 4356 19610
rect 4380 19558 4426 19610
rect 4426 19558 4436 19610
rect 4460 19558 4490 19610
rect 4490 19558 4516 19610
rect 4220 19556 4276 19558
rect 4300 19556 4356 19558
rect 4380 19556 4436 19558
rect 4460 19556 4516 19558
rect 4618 19352 4674 19408
rect 4434 19116 4436 19136
rect 4436 19116 4488 19136
rect 4488 19116 4490 19136
rect 4434 19080 4490 19116
rect 4220 18522 4276 18524
rect 4300 18522 4356 18524
rect 4380 18522 4436 18524
rect 4460 18522 4516 18524
rect 4220 18470 4246 18522
rect 4246 18470 4276 18522
rect 4300 18470 4310 18522
rect 4310 18470 4356 18522
rect 4380 18470 4426 18522
rect 4426 18470 4436 18522
rect 4460 18470 4490 18522
rect 4490 18470 4516 18522
rect 4220 18468 4276 18470
rect 4300 18468 4356 18470
rect 4380 18468 4436 18470
rect 4460 18468 4516 18470
rect 3882 17992 3938 18048
rect 3422 15000 3478 15056
rect 3330 13368 3386 13424
rect 3330 11600 3386 11656
rect 3146 10004 3148 10024
rect 3148 10004 3200 10024
rect 3200 10004 3202 10024
rect 3146 9968 3202 10004
rect 3698 12280 3754 12336
rect 3514 5072 3570 5128
rect 3422 4800 3478 4856
rect 4220 17434 4276 17436
rect 4300 17434 4356 17436
rect 4380 17434 4436 17436
rect 4460 17434 4516 17436
rect 4220 17382 4246 17434
rect 4246 17382 4276 17434
rect 4300 17382 4310 17434
rect 4310 17382 4356 17434
rect 4380 17382 4426 17434
rect 4426 17382 4436 17434
rect 4460 17382 4490 17434
rect 4490 17382 4516 17434
rect 4220 17380 4276 17382
rect 4300 17380 4356 17382
rect 4380 17380 4436 17382
rect 4460 17380 4516 17382
rect 4220 16346 4276 16348
rect 4300 16346 4356 16348
rect 4380 16346 4436 16348
rect 4460 16346 4516 16348
rect 4220 16294 4246 16346
rect 4246 16294 4276 16346
rect 4300 16294 4310 16346
rect 4310 16294 4356 16346
rect 4380 16294 4426 16346
rect 4426 16294 4436 16346
rect 4460 16294 4490 16346
rect 4490 16294 4516 16346
rect 4220 16292 4276 16294
rect 4300 16292 4356 16294
rect 4380 16292 4436 16294
rect 4460 16292 4516 16294
rect 4220 15258 4276 15260
rect 4300 15258 4356 15260
rect 4380 15258 4436 15260
rect 4460 15258 4516 15260
rect 4220 15206 4246 15258
rect 4246 15206 4276 15258
rect 4300 15206 4310 15258
rect 4310 15206 4356 15258
rect 4380 15206 4426 15258
rect 4426 15206 4436 15258
rect 4460 15206 4490 15258
rect 4490 15206 4516 15258
rect 4220 15204 4276 15206
rect 4300 15204 4356 15206
rect 4380 15204 4436 15206
rect 4460 15204 4516 15206
rect 4220 14170 4276 14172
rect 4300 14170 4356 14172
rect 4380 14170 4436 14172
rect 4460 14170 4516 14172
rect 4220 14118 4246 14170
rect 4246 14118 4276 14170
rect 4300 14118 4310 14170
rect 4310 14118 4356 14170
rect 4380 14118 4426 14170
rect 4426 14118 4436 14170
rect 4460 14118 4490 14170
rect 4490 14118 4516 14170
rect 4220 14116 4276 14118
rect 4300 14116 4356 14118
rect 4380 14116 4436 14118
rect 4460 14116 4516 14118
rect 4220 13082 4276 13084
rect 4300 13082 4356 13084
rect 4380 13082 4436 13084
rect 4460 13082 4516 13084
rect 4220 13030 4246 13082
rect 4246 13030 4276 13082
rect 4300 13030 4310 13082
rect 4310 13030 4356 13082
rect 4380 13030 4426 13082
rect 4426 13030 4436 13082
rect 4460 13030 4490 13082
rect 4490 13030 4516 13082
rect 4220 13028 4276 13030
rect 4300 13028 4356 13030
rect 4380 13028 4436 13030
rect 4460 13028 4516 13030
rect 4220 11994 4276 11996
rect 4300 11994 4356 11996
rect 4380 11994 4436 11996
rect 4460 11994 4516 11996
rect 4220 11942 4246 11994
rect 4246 11942 4276 11994
rect 4300 11942 4310 11994
rect 4310 11942 4356 11994
rect 4380 11942 4426 11994
rect 4426 11942 4436 11994
rect 4460 11942 4490 11994
rect 4490 11942 4516 11994
rect 4220 11940 4276 11942
rect 4300 11940 4356 11942
rect 4380 11940 4436 11942
rect 4460 11940 4516 11942
rect 4220 10906 4276 10908
rect 4300 10906 4356 10908
rect 4380 10906 4436 10908
rect 4460 10906 4516 10908
rect 4220 10854 4246 10906
rect 4246 10854 4276 10906
rect 4300 10854 4310 10906
rect 4310 10854 4356 10906
rect 4380 10854 4426 10906
rect 4426 10854 4436 10906
rect 4460 10854 4490 10906
rect 4490 10854 4516 10906
rect 4220 10852 4276 10854
rect 4300 10852 4356 10854
rect 4380 10852 4436 10854
rect 4460 10852 4516 10854
rect 3882 10240 3938 10296
rect 4220 9818 4276 9820
rect 4300 9818 4356 9820
rect 4380 9818 4436 9820
rect 4460 9818 4516 9820
rect 4220 9766 4246 9818
rect 4246 9766 4276 9818
rect 4300 9766 4310 9818
rect 4310 9766 4356 9818
rect 4380 9766 4426 9818
rect 4426 9766 4436 9818
rect 4460 9766 4490 9818
rect 4490 9766 4516 9818
rect 4220 9764 4276 9766
rect 4300 9764 4356 9766
rect 4380 9764 4436 9766
rect 4460 9764 4516 9766
rect 4220 8730 4276 8732
rect 4300 8730 4356 8732
rect 4380 8730 4436 8732
rect 4460 8730 4516 8732
rect 4220 8678 4246 8730
rect 4246 8678 4276 8730
rect 4300 8678 4310 8730
rect 4310 8678 4356 8730
rect 4380 8678 4426 8730
rect 4426 8678 4436 8730
rect 4460 8678 4490 8730
rect 4490 8678 4516 8730
rect 4220 8676 4276 8678
rect 4300 8676 4356 8678
rect 4380 8676 4436 8678
rect 4460 8676 4516 8678
rect 4220 7642 4276 7644
rect 4300 7642 4356 7644
rect 4380 7642 4436 7644
rect 4460 7642 4516 7644
rect 4220 7590 4246 7642
rect 4246 7590 4276 7642
rect 4300 7590 4310 7642
rect 4310 7590 4356 7642
rect 4380 7590 4426 7642
rect 4426 7590 4436 7642
rect 4460 7590 4490 7642
rect 4490 7590 4516 7642
rect 4220 7588 4276 7590
rect 4300 7588 4356 7590
rect 4380 7588 4436 7590
rect 4460 7588 4516 7590
rect 6734 33768 6790 33824
rect 9402 74840 9458 74896
rect 8758 74704 8814 74760
rect 8942 72800 8998 72856
rect 8390 67632 8446 67688
rect 7378 62192 7434 62248
rect 8758 49680 8814 49736
rect 8850 46164 8906 46200
rect 8850 46144 8852 46164
rect 8852 46144 8904 46164
rect 8904 46144 8906 46164
rect 8114 44920 8170 44976
rect 8298 44276 8300 44296
rect 8300 44276 8352 44296
rect 8352 44276 8354 44296
rect 8298 44240 8354 44276
rect 8850 42336 8906 42392
rect 8666 36488 8722 36544
rect 8482 34448 8538 34504
rect 8574 33904 8630 33960
rect 8482 33804 8484 33824
rect 8484 33804 8536 33824
rect 8536 33804 8538 33824
rect 7746 32680 7802 32736
rect 7010 31184 7066 31240
rect 7562 31864 7618 31920
rect 7654 31764 7656 31784
rect 7656 31764 7708 31784
rect 7708 31764 7710 31784
rect 7654 31728 7710 31764
rect 7470 31084 7472 31104
rect 7472 31084 7524 31104
rect 7524 31084 7526 31104
rect 7470 31048 7526 31084
rect 7746 30776 7802 30832
rect 7654 30252 7710 30288
rect 7654 30232 7656 30252
rect 7656 30232 7708 30252
rect 7708 30232 7710 30252
rect 7562 29960 7618 30016
rect 7562 28872 7618 28928
rect 7102 26732 7104 26752
rect 7104 26732 7156 26752
rect 7156 26732 7158 26752
rect 7102 26696 7158 26732
rect 8482 33768 8538 33804
rect 8114 32816 8170 32872
rect 8022 31048 8078 31104
rect 8574 32680 8630 32736
rect 8206 29280 8262 29336
rect 8206 29144 8262 29200
rect 8390 29144 8446 29200
rect 8114 28872 8170 28928
rect 8114 28736 8170 28792
rect 8758 33108 8814 33144
rect 8758 33088 8760 33108
rect 8760 33088 8812 33108
rect 8812 33088 8814 33108
rect 8758 32680 8814 32736
rect 8298 28872 8354 28928
rect 8482 28872 8538 28928
rect 8206 28600 8262 28656
rect 8022 27820 8024 27840
rect 8024 27820 8076 27840
rect 8076 27820 8078 27840
rect 8022 27784 8078 27820
rect 7838 23704 7894 23760
rect 6274 21800 6330 21856
rect 6090 19352 6146 19408
rect 4894 17720 4950 17776
rect 4894 16904 4950 16960
rect 8114 23976 8170 24032
rect 7930 16224 7986 16280
rect 8482 26424 8538 26480
rect 8390 17720 8446 17776
rect 4710 13776 4766 13832
rect 4066 6840 4122 6896
rect 4220 6554 4276 6556
rect 4300 6554 4356 6556
rect 4380 6554 4436 6556
rect 4460 6554 4516 6556
rect 4220 6502 4246 6554
rect 4246 6502 4276 6554
rect 4300 6502 4310 6554
rect 4310 6502 4356 6554
rect 4380 6502 4426 6554
rect 4426 6502 4436 6554
rect 4460 6502 4490 6554
rect 4490 6502 4516 6554
rect 4220 6500 4276 6502
rect 4300 6500 4356 6502
rect 4380 6500 4436 6502
rect 4460 6500 4516 6502
rect 4066 6160 4122 6216
rect 4220 5466 4276 5468
rect 4300 5466 4356 5468
rect 4380 5466 4436 5468
rect 4460 5466 4516 5468
rect 4220 5414 4246 5466
rect 4246 5414 4276 5466
rect 4300 5414 4310 5466
rect 4310 5414 4356 5466
rect 4380 5414 4426 5466
rect 4426 5414 4436 5466
rect 4460 5414 4490 5466
rect 4490 5414 4516 5466
rect 4220 5412 4276 5414
rect 4300 5412 4356 5414
rect 4380 5412 4436 5414
rect 4460 5412 4516 5414
rect 4220 4378 4276 4380
rect 4300 4378 4356 4380
rect 4380 4378 4436 4380
rect 4460 4378 4516 4380
rect 4220 4326 4246 4378
rect 4246 4326 4276 4378
rect 4300 4326 4310 4378
rect 4310 4326 4356 4378
rect 4380 4326 4426 4378
rect 4426 4326 4436 4378
rect 4460 4326 4490 4378
rect 4490 4326 4516 4378
rect 4220 4324 4276 4326
rect 4300 4324 4356 4326
rect 4380 4324 4436 4326
rect 4460 4324 4516 4326
rect 3698 3440 3754 3496
rect 4220 3290 4276 3292
rect 4300 3290 4356 3292
rect 4380 3290 4436 3292
rect 4460 3290 4516 3292
rect 4220 3238 4246 3290
rect 4246 3238 4276 3290
rect 4300 3238 4310 3290
rect 4310 3238 4356 3290
rect 4380 3238 4426 3290
rect 4426 3238 4436 3290
rect 4460 3238 4490 3290
rect 4490 3238 4516 3290
rect 4220 3236 4276 3238
rect 4300 3236 4356 3238
rect 4380 3236 4436 3238
rect 4460 3236 4516 3238
rect 4220 2202 4276 2204
rect 4300 2202 4356 2204
rect 4380 2202 4436 2204
rect 4460 2202 4516 2204
rect 4220 2150 4246 2202
rect 4246 2150 4276 2202
rect 4300 2150 4310 2202
rect 4310 2150 4356 2202
rect 4380 2150 4426 2202
rect 4426 2150 4436 2202
rect 4460 2150 4490 2202
rect 4490 2150 4516 2202
rect 4220 2148 4276 2150
rect 4300 2148 4356 2150
rect 4380 2148 4436 2150
rect 4460 2148 4516 2150
rect 7102 10124 7158 10160
rect 7102 10104 7104 10124
rect 7104 10104 7156 10124
rect 7156 10104 7158 10124
rect 7194 8336 7250 8392
rect 5998 7520 6054 7576
rect 4802 6160 4858 6216
rect 7838 6296 7894 6352
rect 10598 75248 10654 75304
rect 10414 74704 10470 74760
rect 9218 60560 9274 60616
rect 9126 43696 9182 43752
rect 8942 41792 8998 41848
rect 9034 36896 9090 36952
rect 8942 35128 8998 35184
rect 9954 53080 10010 53136
rect 9862 45328 9918 45384
rect 9402 39344 9458 39400
rect 9310 36352 9366 36408
rect 9218 32564 9274 32600
rect 9218 32544 9220 32564
rect 9220 32544 9272 32564
rect 9272 32544 9274 32564
rect 9402 33768 9458 33824
rect 10230 39888 10286 39944
rect 10138 34856 10194 34912
rect 10046 34720 10102 34776
rect 8942 28620 8998 28656
rect 8942 28600 8944 28620
rect 8944 28600 8996 28620
rect 8996 28600 8998 28620
rect 8942 27956 8944 27976
rect 8944 27956 8996 27976
rect 8996 27956 8998 27976
rect 8942 27920 8998 27956
rect 8942 23704 8998 23760
rect 8850 21936 8906 21992
rect 9126 29708 9182 29744
rect 9126 29688 9128 29708
rect 9128 29688 9180 29708
rect 9180 29688 9182 29708
rect 9126 28192 9182 28248
rect 9126 26968 9182 27024
rect 9310 25472 9366 25528
rect 9034 19896 9090 19952
rect 8298 9016 8354 9072
rect 9586 33496 9642 33552
rect 9862 32952 9918 33008
rect 9586 32544 9642 32600
rect 9678 32136 9734 32192
rect 9494 31456 9550 31512
rect 9494 30640 9550 30696
rect 9586 30504 9642 30560
rect 9862 31864 9918 31920
rect 9586 29280 9642 29336
rect 9678 28736 9734 28792
rect 9494 28328 9550 28384
rect 9954 29416 10010 29472
rect 9862 27648 9918 27704
rect 9862 26288 9918 26344
rect 9678 25236 9680 25256
rect 9680 25236 9732 25256
rect 9732 25236 9734 25256
rect 9678 25200 9734 25236
rect 10322 28464 10378 28520
rect 10230 27784 10286 27840
rect 10138 27412 10140 27432
rect 10140 27412 10192 27432
rect 10192 27412 10194 27432
rect 10138 27376 10194 27412
rect 9678 23296 9734 23352
rect 10046 22208 10102 22264
rect 10690 69672 10746 69728
rect 10506 59880 10562 59936
rect 10598 34040 10654 34096
rect 10506 33632 10562 33688
rect 10598 31592 10654 31648
rect 10598 28872 10654 28928
rect 10506 28600 10562 28656
rect 10506 27548 10508 27568
rect 10508 27548 10560 27568
rect 10560 27548 10562 27568
rect 10506 27512 10562 27548
rect 9678 17856 9734 17912
rect 10230 16224 10286 16280
rect 10598 15000 10654 15056
rect 9586 4256 9642 4312
rect 12346 75384 12402 75440
rect 11518 70488 11574 70544
rect 12346 68312 12402 68368
rect 11242 67632 11298 67688
rect 10874 67224 10930 67280
rect 10782 62056 10838 62112
rect 10966 61512 11022 61568
rect 10782 57568 10838 57624
rect 10966 36624 11022 36680
rect 10782 35828 10838 35864
rect 10782 35808 10784 35828
rect 10784 35808 10836 35828
rect 10836 35808 10838 35828
rect 10966 35692 11022 35728
rect 10966 35672 10968 35692
rect 10968 35672 11020 35692
rect 11020 35672 11022 35692
rect 11150 35128 11206 35184
rect 10966 33904 11022 33960
rect 10874 32544 10930 32600
rect 11150 32952 11206 33008
rect 11058 32816 11114 32872
rect 10966 32428 11022 32464
rect 10966 32408 10968 32428
rect 10968 32408 11020 32428
rect 11020 32408 11022 32428
rect 10874 32292 10930 32328
rect 10874 32272 10876 32292
rect 10876 32272 10928 32292
rect 10928 32272 10930 32292
rect 10782 31184 10838 31240
rect 10966 31084 10968 31104
rect 10968 31084 11020 31104
rect 11020 31084 11022 31104
rect 10966 31048 11022 31084
rect 10966 30368 11022 30424
rect 10874 30096 10930 30152
rect 10966 29824 11022 29880
rect 10966 29572 11022 29608
rect 10966 29552 10968 29572
rect 10968 29552 11020 29572
rect 11020 29552 11022 29572
rect 10874 29144 10930 29200
rect 10874 29044 10876 29064
rect 10876 29044 10928 29064
rect 10928 29044 10930 29064
rect 10874 29008 10930 29044
rect 13358 75792 13414 75848
rect 16394 75792 16450 75848
rect 14278 73888 14334 73944
rect 15382 73752 15438 73808
rect 14094 71848 14150 71904
rect 12622 67768 12678 67824
rect 12254 55412 12310 55448
rect 12254 55392 12256 55412
rect 12256 55392 12308 55412
rect 12308 55392 12310 55412
rect 11886 50496 11942 50552
rect 11610 49544 11666 49600
rect 11426 46316 11428 46336
rect 11428 46316 11480 46336
rect 11480 46316 11482 46336
rect 11426 46280 11482 46316
rect 11334 37304 11390 37360
rect 11334 36216 11390 36272
rect 12254 40840 12310 40896
rect 11702 35536 11758 35592
rect 11518 33768 11574 33824
rect 11426 32952 11482 33008
rect 11334 31728 11390 31784
rect 11242 30776 11298 30832
rect 10966 28600 11022 28656
rect 10782 27920 10838 27976
rect 10874 26832 10930 26888
rect 11334 29280 11390 29336
rect 11702 32816 11758 32872
rect 11702 32544 11758 32600
rect 11886 34992 11942 35048
rect 12254 35944 12310 36000
rect 11886 33940 11888 33960
rect 11888 33940 11940 33960
rect 11940 33940 11942 33960
rect 11886 33904 11942 33940
rect 11886 33360 11942 33416
rect 12162 32972 12218 33008
rect 12162 32952 12164 32972
rect 12164 32952 12216 32972
rect 12216 32952 12218 32972
rect 12070 32716 12072 32736
rect 12072 32716 12124 32736
rect 12124 32716 12126 32736
rect 12070 32680 12126 32716
rect 11610 32136 11666 32192
rect 11334 26560 11390 26616
rect 11242 26424 11298 26480
rect 11334 25492 11390 25528
rect 11334 25472 11336 25492
rect 11336 25472 11388 25492
rect 11388 25472 11390 25492
rect 10966 21412 11022 21448
rect 10966 21392 10968 21412
rect 10968 21392 11020 21412
rect 11020 21392 11022 21412
rect 11886 32136 11942 32192
rect 11978 31220 11980 31240
rect 11980 31220 12032 31240
rect 12032 31220 12034 31240
rect 11978 31184 12034 31220
rect 11886 30776 11942 30832
rect 11794 30640 11850 30696
rect 12254 32000 12310 32056
rect 12254 31456 12310 31512
rect 12162 31184 12218 31240
rect 11886 29960 11942 30016
rect 11886 29300 11942 29336
rect 11886 29280 11888 29300
rect 11888 29280 11940 29300
rect 11940 29280 11942 29300
rect 11518 26424 11574 26480
rect 11518 25916 11520 25936
rect 11520 25916 11572 25936
rect 11572 25916 11574 25936
rect 11518 25880 11574 25916
rect 12070 29688 12126 29744
rect 12254 31084 12256 31104
rect 12256 31084 12308 31104
rect 12308 31084 12310 31104
rect 12254 31048 12310 31084
rect 15198 70760 15254 70816
rect 15198 69808 15254 69864
rect 14094 65456 14150 65512
rect 13174 61548 13176 61568
rect 13176 61548 13228 61568
rect 13228 61548 13230 61568
rect 13174 61512 13230 61548
rect 13818 61512 13874 61568
rect 13358 57976 13414 58032
rect 13266 56616 13322 56672
rect 13450 55120 13506 55176
rect 13266 54440 13322 54496
rect 13542 54440 13598 54496
rect 13358 54032 13414 54088
rect 12806 46824 12862 46880
rect 12714 42628 12770 42664
rect 12714 42608 12716 42628
rect 12716 42608 12768 42628
rect 12768 42608 12770 42628
rect 12622 40296 12678 40352
rect 12530 33516 12586 33552
rect 12530 33496 12532 33516
rect 12532 33496 12584 33516
rect 12584 33496 12586 33516
rect 12806 34604 12862 34640
rect 12806 34584 12808 34604
rect 12808 34584 12860 34604
rect 12860 34584 12862 34604
rect 12806 33632 12862 33688
rect 12714 32836 12770 32872
rect 12714 32816 12716 32836
rect 12716 32816 12768 32836
rect 12768 32816 12770 32836
rect 13634 46280 13690 46336
rect 13174 40296 13230 40352
rect 13082 39924 13084 39944
rect 13084 39924 13136 39944
rect 13136 39924 13138 39944
rect 13082 39888 13138 39924
rect 12990 36760 13046 36816
rect 13082 32816 13138 32872
rect 12898 31592 12954 31648
rect 12530 30912 12586 30968
rect 12438 29552 12494 29608
rect 12714 30640 12770 30696
rect 12898 30676 12900 30696
rect 12900 30676 12952 30696
rect 12952 30676 12954 30696
rect 12898 30640 12954 30676
rect 12622 30232 12678 30288
rect 12622 29416 12678 29472
rect 12162 25744 12218 25800
rect 11978 25336 12034 25392
rect 11794 23296 11850 23352
rect 12162 22752 12218 22808
rect 11610 21800 11666 21856
rect 11426 18128 11482 18184
rect 11886 20304 11942 20360
rect 13082 30504 13138 30560
rect 12806 28500 12808 28520
rect 12808 28500 12860 28520
rect 12860 28500 12862 28520
rect 12806 28464 12862 28500
rect 12990 27548 12992 27568
rect 12992 27548 13044 27568
rect 13044 27548 13046 27568
rect 12990 27512 13046 27548
rect 13266 31592 13322 31648
rect 13542 38256 13598 38312
rect 14554 63824 14610 63880
rect 14278 57588 14334 57624
rect 14278 57568 14280 57588
rect 14280 57568 14332 57588
rect 14332 57568 14334 57588
rect 14186 56364 14242 56400
rect 14186 56344 14188 56364
rect 14188 56344 14240 56364
rect 14240 56344 14242 56364
rect 14370 56752 14426 56808
rect 14278 55256 14334 55312
rect 14370 54596 14426 54632
rect 14370 54576 14372 54596
rect 14372 54576 14424 54596
rect 14424 54576 14426 54596
rect 15014 57316 15070 57352
rect 15014 57296 15016 57316
rect 15016 57296 15068 57316
rect 15068 57296 15070 57316
rect 14646 55936 14702 55992
rect 14738 53932 14740 53952
rect 14740 53932 14792 53952
rect 14792 53932 14794 53952
rect 14738 53896 14794 53932
rect 14922 53896 14978 53952
rect 15106 53760 15162 53816
rect 14738 52692 14794 52728
rect 14738 52672 14740 52692
rect 14740 52672 14792 52692
rect 14792 52672 14794 52692
rect 14738 51212 14740 51232
rect 14740 51212 14792 51232
rect 14792 51212 14794 51232
rect 14738 51176 14794 51212
rect 15198 53352 15254 53408
rect 15290 52536 15346 52592
rect 15106 52128 15162 52184
rect 14830 50496 14886 50552
rect 14462 45464 14518 45520
rect 14002 40332 14004 40352
rect 14004 40332 14056 40352
rect 14056 40332 14058 40352
rect 14002 40296 14058 40332
rect 14370 41792 14426 41848
rect 13726 37324 13782 37360
rect 13726 37304 13728 37324
rect 13728 37304 13780 37324
rect 13780 37304 13782 37324
rect 14094 37032 14150 37088
rect 14002 36896 14058 36952
rect 13542 36488 13598 36544
rect 13542 34040 13598 34096
rect 13542 33632 13598 33688
rect 13266 29144 13322 29200
rect 12622 25608 12678 25664
rect 12346 23740 12348 23760
rect 12348 23740 12400 23760
rect 12400 23740 12402 23760
rect 12346 23704 12402 23740
rect 12530 22924 12532 22944
rect 12532 22924 12584 22944
rect 12584 22924 12586 22944
rect 12530 22888 12586 22924
rect 12438 22344 12494 22400
rect 11886 17992 11942 18048
rect 11978 16088 12034 16144
rect 11702 14456 11758 14512
rect 12346 7284 12348 7304
rect 12348 7284 12400 7304
rect 12400 7284 12402 7304
rect 12346 7248 12402 7284
rect 12898 26288 12954 26344
rect 12806 24792 12862 24848
rect 13358 28872 13414 28928
rect 13542 30504 13598 30560
rect 13450 28192 13506 28248
rect 13450 27820 13452 27840
rect 13452 27820 13504 27840
rect 13504 27820 13506 27840
rect 13450 27784 13506 27820
rect 13082 26424 13138 26480
rect 13542 26968 13598 27024
rect 14370 38412 14426 38448
rect 14370 38392 14372 38412
rect 14372 38392 14424 38412
rect 14424 38392 14426 38412
rect 14186 36488 14242 36544
rect 13910 34584 13966 34640
rect 14370 35572 14372 35592
rect 14372 35572 14424 35592
rect 14424 35572 14426 35592
rect 14370 35536 14426 35572
rect 13910 33088 13966 33144
rect 13818 32000 13874 32056
rect 13818 29144 13874 29200
rect 14370 33632 14426 33688
rect 14278 33360 14334 33416
rect 14370 31884 14426 31920
rect 14370 31864 14372 31884
rect 14372 31864 14424 31884
rect 14424 31864 14426 31884
rect 14278 31592 14334 31648
rect 13910 28872 13966 28928
rect 14186 29552 14242 29608
rect 14094 29144 14150 29200
rect 13174 26288 13230 26344
rect 13082 24112 13138 24168
rect 13174 22616 13230 22672
rect 13082 21392 13138 21448
rect 12990 19352 13046 19408
rect 13174 12316 13176 12336
rect 13176 12316 13228 12336
rect 13228 12316 13230 12336
rect 13174 12280 13230 12316
rect 14186 28192 14242 28248
rect 14002 27376 14058 27432
rect 14094 27240 14150 27296
rect 14002 26152 14058 26208
rect 13634 24520 13690 24576
rect 13910 24404 13966 24440
rect 13910 24384 13912 24404
rect 13912 24384 13964 24404
rect 13964 24384 13966 24404
rect 14094 24384 14150 24440
rect 14002 23296 14058 23352
rect 14370 27784 14426 27840
rect 14462 27412 14464 27432
rect 14464 27412 14516 27432
rect 14516 27412 14518 27432
rect 14462 27376 14518 27412
rect 16394 72800 16450 72856
rect 15842 71984 15898 72040
rect 15566 71576 15622 71632
rect 15474 55700 15476 55720
rect 15476 55700 15528 55720
rect 15528 55700 15530 55720
rect 15474 55664 15530 55700
rect 15474 53624 15530 53680
rect 15106 48864 15162 48920
rect 15382 48764 15384 48784
rect 15384 48764 15436 48784
rect 15436 48764 15438 48784
rect 15382 48728 15438 48764
rect 15750 70896 15806 70952
rect 15934 70488 15990 70544
rect 15842 64096 15898 64152
rect 15934 63416 15990 63472
rect 16486 59336 16542 59392
rect 16670 56208 16726 56264
rect 16302 55528 16358 55584
rect 16118 54168 16174 54224
rect 16854 55820 16910 55856
rect 16854 55800 16856 55820
rect 16856 55800 16908 55820
rect 16908 55800 16910 55820
rect 16578 55120 16634 55176
rect 16210 52944 16266 53000
rect 15658 51040 15714 51096
rect 15658 46824 15714 46880
rect 15566 45464 15622 45520
rect 16118 52012 16174 52048
rect 16118 51992 16120 52012
rect 16120 51992 16172 52012
rect 16172 51992 16174 52012
rect 16854 54324 16910 54360
rect 16854 54304 16856 54324
rect 16856 54304 16908 54324
rect 16908 54304 16910 54324
rect 16854 54032 16910 54088
rect 16946 52672 17002 52728
rect 16578 52400 16634 52456
rect 16486 51856 16542 51912
rect 16670 52128 16726 52184
rect 16670 49272 16726 49328
rect 16854 46824 16910 46880
rect 17498 77152 17554 77208
rect 19580 77818 19636 77820
rect 19660 77818 19716 77820
rect 19740 77818 19796 77820
rect 19820 77818 19876 77820
rect 19580 77766 19606 77818
rect 19606 77766 19636 77818
rect 19660 77766 19670 77818
rect 19670 77766 19716 77818
rect 19740 77766 19786 77818
rect 19786 77766 19796 77818
rect 19820 77766 19850 77818
rect 19850 77766 19876 77818
rect 19580 77764 19636 77766
rect 19660 77764 19716 77766
rect 19740 77764 19796 77766
rect 19820 77764 19876 77766
rect 17130 57740 17132 57760
rect 17132 57740 17184 57760
rect 17184 57740 17186 57760
rect 17130 57704 17186 57740
rect 17222 55700 17224 55720
rect 17224 55700 17276 55720
rect 17276 55700 17278 55720
rect 17222 55664 17278 55700
rect 17222 55392 17278 55448
rect 17498 54712 17554 54768
rect 17498 53760 17554 53816
rect 17038 46416 17094 46472
rect 17222 50924 17278 50960
rect 17222 50904 17224 50924
rect 17224 50904 17276 50924
rect 17276 50904 17278 50924
rect 17222 49972 17278 50008
rect 17590 51176 17646 51232
rect 17590 50768 17646 50824
rect 17406 50260 17408 50280
rect 17408 50260 17460 50280
rect 17460 50260 17462 50280
rect 17406 50224 17462 50260
rect 17222 49952 17224 49972
rect 17224 49952 17276 49972
rect 17276 49952 17278 49972
rect 17406 48884 17462 48920
rect 17406 48864 17408 48884
rect 17408 48864 17460 48884
rect 17460 48864 17462 48884
rect 14830 39752 14886 39808
rect 15106 38528 15162 38584
rect 14830 37848 14886 37904
rect 15014 37848 15070 37904
rect 15106 37440 15162 37496
rect 14738 37068 14740 37088
rect 14740 37068 14792 37088
rect 14792 37068 14794 37088
rect 14738 37032 14794 37068
rect 14646 35400 14702 35456
rect 14646 35128 14702 35184
rect 14646 33396 14648 33416
rect 14648 33396 14700 33416
rect 14700 33396 14702 33416
rect 14646 33360 14702 33396
rect 14922 36660 14924 36680
rect 14924 36660 14976 36680
rect 14976 36660 14978 36680
rect 14922 36624 14978 36660
rect 14922 34720 14978 34776
rect 15198 36488 15254 36544
rect 15198 36352 15254 36408
rect 15474 37712 15530 37768
rect 15290 36216 15346 36272
rect 15198 35128 15254 35184
rect 14830 34584 14886 34640
rect 14830 33904 14886 33960
rect 14830 33632 14886 33688
rect 14830 32000 14886 32056
rect 14922 31728 14978 31784
rect 15106 31728 15162 31784
rect 15106 31456 15162 31512
rect 14830 30796 14886 30832
rect 14830 30776 14832 30796
rect 14832 30776 14884 30796
rect 14884 30776 14886 30796
rect 14922 30640 14978 30696
rect 14830 29552 14886 29608
rect 14646 26580 14702 26616
rect 14646 26560 14648 26580
rect 14648 26560 14700 26580
rect 14700 26560 14702 26580
rect 14462 25200 14518 25256
rect 14646 25064 14702 25120
rect 14554 24928 14610 24984
rect 14738 24656 14794 24712
rect 14554 23704 14610 23760
rect 15290 32680 15346 32736
rect 15106 29552 15162 29608
rect 15106 29280 15162 29336
rect 15474 31340 15530 31376
rect 15474 31320 15476 31340
rect 15476 31320 15528 31340
rect 15528 31320 15530 31340
rect 16486 40024 16542 40080
rect 15934 36624 15990 36680
rect 15934 35808 15990 35864
rect 15934 34040 15990 34096
rect 15842 33904 15898 33960
rect 15842 32292 15898 32328
rect 15842 32272 15844 32292
rect 15844 32272 15896 32292
rect 15896 32272 15898 32292
rect 15842 31728 15898 31784
rect 15750 30776 15806 30832
rect 15474 29844 15530 29880
rect 15474 29824 15476 29844
rect 15476 29824 15528 29844
rect 15528 29824 15530 29844
rect 15842 29960 15898 30016
rect 15566 29008 15622 29064
rect 15106 28600 15162 28656
rect 14646 22752 14702 22808
rect 14830 22752 14886 22808
rect 14738 22344 14794 22400
rect 14278 20576 14334 20632
rect 13634 19488 13690 19544
rect 13910 20476 13912 20496
rect 13912 20476 13964 20496
rect 13964 20476 13966 20496
rect 13910 20440 13966 20476
rect 13726 18808 13782 18864
rect 13266 8472 13322 8528
rect 13450 7284 13452 7304
rect 13452 7284 13504 7304
rect 13504 7284 13506 7304
rect 13450 7248 13506 7284
rect 13818 15020 13874 15056
rect 13818 15000 13820 15020
rect 13820 15000 13872 15020
rect 13872 15000 13874 15020
rect 13634 5480 13690 5536
rect 14002 4820 14058 4856
rect 14002 4800 14004 4820
rect 14004 4800 14056 4820
rect 14056 4800 14058 4820
rect 14462 19488 14518 19544
rect 14462 18420 14518 18456
rect 14462 18400 14464 18420
rect 14464 18400 14516 18420
rect 14516 18400 14518 18420
rect 14830 17992 14886 18048
rect 14738 5480 14794 5536
rect 14278 3984 14334 4040
rect 15106 24828 15108 24848
rect 15108 24828 15160 24848
rect 15160 24828 15162 24848
rect 15106 24792 15162 24828
rect 15658 28328 15714 28384
rect 16026 32564 16082 32600
rect 16026 32544 16028 32564
rect 16028 32544 16080 32564
rect 16080 32544 16082 32564
rect 16210 36760 16266 36816
rect 16302 35672 16358 35728
rect 16486 38256 16542 38312
rect 16670 38800 16726 38856
rect 16578 37848 16634 37904
rect 16486 35944 16542 36000
rect 16210 34992 16266 35048
rect 16394 34856 16450 34912
rect 16302 34720 16358 34776
rect 16394 34620 16396 34640
rect 16396 34620 16448 34640
rect 16448 34620 16450 34640
rect 16394 34584 16450 34620
rect 16302 33360 16358 33416
rect 16026 31728 16082 31784
rect 16026 31592 16082 31648
rect 15934 27920 15990 27976
rect 15658 25472 15714 25528
rect 15106 24012 15108 24032
rect 15108 24012 15160 24032
rect 15160 24012 15162 24032
rect 15106 23976 15162 24012
rect 15106 23860 15162 23896
rect 15106 23840 15108 23860
rect 15108 23840 15160 23860
rect 15160 23840 15162 23860
rect 15290 23296 15346 23352
rect 15198 22108 15200 22128
rect 15200 22108 15252 22128
rect 15252 22108 15254 22128
rect 15198 22072 15254 22108
rect 15566 21836 15568 21856
rect 15568 21836 15620 21856
rect 15620 21836 15622 21856
rect 15566 21800 15622 21836
rect 15566 20596 15622 20632
rect 15566 20576 15568 20596
rect 15568 20576 15620 20596
rect 15620 20576 15622 20596
rect 15842 24384 15898 24440
rect 15934 22616 15990 22672
rect 16394 31048 16450 31104
rect 16302 26016 16358 26072
rect 16210 25780 16212 25800
rect 16212 25780 16264 25800
rect 16264 25780 16266 25800
rect 16210 25744 16266 25780
rect 15658 20304 15714 20360
rect 15566 17992 15622 18048
rect 15382 15680 15438 15736
rect 15290 14456 15346 14512
rect 16854 38528 16910 38584
rect 16762 38392 16818 38448
rect 16946 37748 16948 37768
rect 16948 37748 17000 37768
rect 17000 37748 17002 37768
rect 16946 37712 17002 37748
rect 16946 37440 17002 37496
rect 16854 37204 16856 37224
rect 16856 37204 16908 37224
rect 16908 37204 16910 37224
rect 16854 37168 16910 37204
rect 16670 36236 16726 36272
rect 16670 36216 16672 36236
rect 16672 36216 16724 36236
rect 16724 36216 16726 36236
rect 17314 40840 17370 40896
rect 17314 40160 17370 40216
rect 17406 38004 17462 38040
rect 17406 37984 17408 38004
rect 17408 37984 17460 38004
rect 17460 37984 17462 38004
rect 17314 37440 17370 37496
rect 17130 36352 17186 36408
rect 16670 35828 16726 35864
rect 16670 35808 16672 35828
rect 16672 35808 16724 35828
rect 16724 35808 16726 35828
rect 16762 35672 16818 35728
rect 16578 35536 16634 35592
rect 16578 35128 16634 35184
rect 16762 34448 16818 34504
rect 16854 33768 16910 33824
rect 16578 32172 16580 32192
rect 16580 32172 16632 32192
rect 16632 32172 16634 32192
rect 16578 32136 16634 32172
rect 16762 31592 16818 31648
rect 16854 31456 16910 31512
rect 16762 29960 16818 30016
rect 16578 29416 16634 29472
rect 16670 28872 16726 28928
rect 16578 26988 16634 27024
rect 16578 26968 16580 26988
rect 16580 26968 16632 26988
rect 16632 26968 16634 26988
rect 17130 35400 17186 35456
rect 17222 30368 17278 30424
rect 17130 29028 17186 29064
rect 17130 29008 17132 29028
rect 17132 29008 17184 29028
rect 17184 29008 17186 29028
rect 17038 28872 17094 28928
rect 16946 26968 17002 27024
rect 16762 26152 16818 26208
rect 16486 25100 16488 25120
rect 16488 25100 16540 25120
rect 16540 25100 16542 25120
rect 16486 25064 16542 25100
rect 16762 24792 16818 24848
rect 16670 24520 16726 24576
rect 17038 24792 17094 24848
rect 17314 25880 17370 25936
rect 17222 25200 17278 25256
rect 17774 74976 17830 75032
rect 19580 76730 19636 76732
rect 19660 76730 19716 76732
rect 19740 76730 19796 76732
rect 19820 76730 19876 76732
rect 19580 76678 19606 76730
rect 19606 76678 19636 76730
rect 19660 76678 19670 76730
rect 19670 76678 19716 76730
rect 19740 76678 19786 76730
rect 19786 76678 19796 76730
rect 19820 76678 19850 76730
rect 19850 76678 19876 76730
rect 19580 76676 19636 76678
rect 19660 76676 19716 76678
rect 19740 76676 19796 76678
rect 19820 76676 19876 76678
rect 19580 75642 19636 75644
rect 19660 75642 19716 75644
rect 19740 75642 19796 75644
rect 19820 75642 19876 75644
rect 19580 75590 19606 75642
rect 19606 75590 19636 75642
rect 19660 75590 19670 75642
rect 19670 75590 19716 75642
rect 19740 75590 19786 75642
rect 19786 75590 19796 75642
rect 19820 75590 19850 75642
rect 19850 75590 19876 75642
rect 19580 75588 19636 75590
rect 19660 75588 19716 75590
rect 19740 75588 19796 75590
rect 19820 75588 19876 75590
rect 19982 75112 20038 75168
rect 19580 74554 19636 74556
rect 19660 74554 19716 74556
rect 19740 74554 19796 74556
rect 19820 74554 19876 74556
rect 19580 74502 19606 74554
rect 19606 74502 19636 74554
rect 19660 74502 19670 74554
rect 19670 74502 19716 74554
rect 19740 74502 19786 74554
rect 19786 74502 19796 74554
rect 19820 74502 19850 74554
rect 19850 74502 19876 74554
rect 19580 74500 19636 74502
rect 19660 74500 19716 74502
rect 19740 74500 19796 74502
rect 19820 74500 19876 74502
rect 19580 73466 19636 73468
rect 19660 73466 19716 73468
rect 19740 73466 19796 73468
rect 19820 73466 19876 73468
rect 19580 73414 19606 73466
rect 19606 73414 19636 73466
rect 19660 73414 19670 73466
rect 19670 73414 19716 73466
rect 19740 73414 19786 73466
rect 19786 73414 19796 73466
rect 19820 73414 19850 73466
rect 19850 73414 19876 73466
rect 19580 73412 19636 73414
rect 19660 73412 19716 73414
rect 19740 73412 19796 73414
rect 19820 73412 19876 73414
rect 19338 72972 19340 72992
rect 19340 72972 19392 72992
rect 19392 72972 19394 72992
rect 19338 72936 19394 72972
rect 19338 72548 19394 72584
rect 19338 72528 19340 72548
rect 19340 72528 19392 72548
rect 19392 72528 19394 72548
rect 19580 72378 19636 72380
rect 19660 72378 19716 72380
rect 19740 72378 19796 72380
rect 19820 72378 19876 72380
rect 19580 72326 19606 72378
rect 19606 72326 19636 72378
rect 19660 72326 19670 72378
rect 19670 72326 19716 72378
rect 19740 72326 19786 72378
rect 19786 72326 19796 72378
rect 19820 72326 19850 72378
rect 19850 72326 19876 72378
rect 19580 72324 19636 72326
rect 19660 72324 19716 72326
rect 19740 72324 19796 72326
rect 19820 72324 19876 72326
rect 19522 71884 19524 71904
rect 19524 71884 19576 71904
rect 19576 71884 19578 71904
rect 19522 71848 19578 71884
rect 18234 71440 18290 71496
rect 17866 59764 17922 59800
rect 17866 59744 17868 59764
rect 17868 59744 17920 59764
rect 17920 59744 17922 59764
rect 17958 59336 18014 59392
rect 17866 56788 17868 56808
rect 17868 56788 17920 56808
rect 17920 56788 17922 56808
rect 17866 56752 17922 56788
rect 17866 56500 17922 56536
rect 17866 56480 17868 56500
rect 17868 56480 17920 56500
rect 17920 56480 17922 56500
rect 17774 56344 17830 56400
rect 17866 53488 17922 53544
rect 18142 56772 18198 56808
rect 18142 56752 18144 56772
rect 18144 56752 18196 56772
rect 18196 56752 18198 56772
rect 19580 71290 19636 71292
rect 19660 71290 19716 71292
rect 19740 71290 19796 71292
rect 19820 71290 19876 71292
rect 19580 71238 19606 71290
rect 19606 71238 19636 71290
rect 19660 71238 19670 71290
rect 19670 71238 19716 71290
rect 19740 71238 19786 71290
rect 19786 71238 19796 71290
rect 19820 71238 19850 71290
rect 19850 71238 19876 71290
rect 19580 71236 19636 71238
rect 19660 71236 19716 71238
rect 19740 71236 19796 71238
rect 19820 71236 19876 71238
rect 19580 70202 19636 70204
rect 19660 70202 19716 70204
rect 19740 70202 19796 70204
rect 19820 70202 19876 70204
rect 19580 70150 19606 70202
rect 19606 70150 19636 70202
rect 19660 70150 19670 70202
rect 19670 70150 19716 70202
rect 19740 70150 19786 70202
rect 19786 70150 19796 70202
rect 19820 70150 19850 70202
rect 19850 70150 19876 70202
rect 19580 70148 19636 70150
rect 19660 70148 19716 70150
rect 19740 70148 19796 70150
rect 19820 70148 19876 70150
rect 19580 69114 19636 69116
rect 19660 69114 19716 69116
rect 19740 69114 19796 69116
rect 19820 69114 19876 69116
rect 19580 69062 19606 69114
rect 19606 69062 19636 69114
rect 19660 69062 19670 69114
rect 19670 69062 19716 69114
rect 19740 69062 19786 69114
rect 19786 69062 19796 69114
rect 19820 69062 19850 69114
rect 19850 69062 19876 69114
rect 19580 69060 19636 69062
rect 19660 69060 19716 69062
rect 19740 69060 19796 69062
rect 19820 69060 19876 69062
rect 19580 68026 19636 68028
rect 19660 68026 19716 68028
rect 19740 68026 19796 68028
rect 19820 68026 19876 68028
rect 19580 67974 19606 68026
rect 19606 67974 19636 68026
rect 19660 67974 19670 68026
rect 19670 67974 19716 68026
rect 19740 67974 19786 68026
rect 19786 67974 19796 68026
rect 19820 67974 19850 68026
rect 19850 67974 19876 68026
rect 19580 67972 19636 67974
rect 19660 67972 19716 67974
rect 19740 67972 19796 67974
rect 19820 67972 19876 67974
rect 19338 67768 19394 67824
rect 19580 66938 19636 66940
rect 19660 66938 19716 66940
rect 19740 66938 19796 66940
rect 19820 66938 19876 66940
rect 19580 66886 19606 66938
rect 19606 66886 19636 66938
rect 19660 66886 19670 66938
rect 19670 66886 19716 66938
rect 19740 66886 19786 66938
rect 19786 66886 19796 66938
rect 19820 66886 19850 66938
rect 19850 66886 19876 66938
rect 19580 66884 19636 66886
rect 19660 66884 19716 66886
rect 19740 66884 19796 66886
rect 19820 66884 19876 66886
rect 19580 65850 19636 65852
rect 19660 65850 19716 65852
rect 19740 65850 19796 65852
rect 19820 65850 19876 65852
rect 19580 65798 19606 65850
rect 19606 65798 19636 65850
rect 19660 65798 19670 65850
rect 19670 65798 19716 65850
rect 19740 65798 19786 65850
rect 19786 65798 19796 65850
rect 19820 65798 19850 65850
rect 19850 65798 19876 65850
rect 19580 65796 19636 65798
rect 19660 65796 19716 65798
rect 19740 65796 19796 65798
rect 19820 65796 19876 65798
rect 19580 64762 19636 64764
rect 19660 64762 19716 64764
rect 19740 64762 19796 64764
rect 19820 64762 19876 64764
rect 19580 64710 19606 64762
rect 19606 64710 19636 64762
rect 19660 64710 19670 64762
rect 19670 64710 19716 64762
rect 19740 64710 19786 64762
rect 19786 64710 19796 64762
rect 19820 64710 19850 64762
rect 19850 64710 19876 64762
rect 19580 64708 19636 64710
rect 19660 64708 19716 64710
rect 19740 64708 19796 64710
rect 19820 64708 19876 64710
rect 19580 63674 19636 63676
rect 19660 63674 19716 63676
rect 19740 63674 19796 63676
rect 19820 63674 19876 63676
rect 19580 63622 19606 63674
rect 19606 63622 19636 63674
rect 19660 63622 19670 63674
rect 19670 63622 19716 63674
rect 19740 63622 19786 63674
rect 19786 63622 19796 63674
rect 19820 63622 19850 63674
rect 19850 63622 19876 63674
rect 19580 63620 19636 63622
rect 19660 63620 19716 63622
rect 19740 63620 19796 63622
rect 19820 63620 19876 63622
rect 19580 62586 19636 62588
rect 19660 62586 19716 62588
rect 19740 62586 19796 62588
rect 19820 62586 19876 62588
rect 19580 62534 19606 62586
rect 19606 62534 19636 62586
rect 19660 62534 19670 62586
rect 19670 62534 19716 62586
rect 19740 62534 19786 62586
rect 19786 62534 19796 62586
rect 19820 62534 19850 62586
rect 19850 62534 19876 62586
rect 19580 62532 19636 62534
rect 19660 62532 19716 62534
rect 19740 62532 19796 62534
rect 19820 62532 19876 62534
rect 18418 62056 18474 62112
rect 20258 74432 20314 74488
rect 20718 68312 20774 68368
rect 19062 62212 19118 62248
rect 19062 62192 19064 62212
rect 19064 62192 19116 62212
rect 19116 62192 19118 62212
rect 19982 62192 20038 62248
rect 18326 57976 18382 58032
rect 18418 55936 18474 55992
rect 18602 59508 18604 59528
rect 18604 59508 18656 59528
rect 18656 59508 18658 59528
rect 18602 59472 18658 59508
rect 18326 53896 18382 53952
rect 18602 53388 18604 53408
rect 18604 53388 18656 53408
rect 18656 53388 18658 53408
rect 18602 53352 18658 53388
rect 17774 51484 17776 51504
rect 17776 51484 17828 51504
rect 17828 51484 17830 51504
rect 17774 51448 17830 51484
rect 18418 51176 18474 51232
rect 18418 50768 18474 50824
rect 18050 46008 18106 46064
rect 17774 44376 17830 44432
rect 17866 40588 17922 40624
rect 17866 40568 17868 40588
rect 17868 40568 17920 40588
rect 17920 40568 17922 40588
rect 17866 39924 17868 39944
rect 17868 39924 17920 39944
rect 17920 39924 17922 39944
rect 17866 39888 17922 39924
rect 17866 36236 17922 36272
rect 17866 36216 17868 36236
rect 17868 36216 17920 36236
rect 17920 36216 17922 36236
rect 18050 36080 18106 36136
rect 17774 34448 17830 34504
rect 17958 34312 18014 34368
rect 17958 34076 17960 34096
rect 17960 34076 18012 34096
rect 18012 34076 18014 34096
rect 17958 34040 18014 34076
rect 17682 32952 17738 33008
rect 17682 30504 17738 30560
rect 17590 30368 17646 30424
rect 17590 28464 17646 28520
rect 17590 27648 17646 27704
rect 17590 27240 17646 27296
rect 16670 20848 16726 20904
rect 17038 23160 17094 23216
rect 17314 23976 17370 24032
rect 16302 18828 16358 18864
rect 16302 18808 16304 18828
rect 16304 18808 16356 18828
rect 16356 18808 16358 18828
rect 17314 19352 17370 19408
rect 17958 32972 18014 33008
rect 17958 32952 17960 32972
rect 17960 32952 18012 32972
rect 18012 32952 18014 32972
rect 18050 32816 18106 32872
rect 18050 30368 18106 30424
rect 17774 28464 17830 28520
rect 18050 27412 18052 27432
rect 18052 27412 18104 27432
rect 18104 27412 18106 27432
rect 18050 27376 18106 27412
rect 17590 25200 17646 25256
rect 17682 24656 17738 24712
rect 17590 24268 17646 24304
rect 17590 24248 17592 24268
rect 17592 24248 17644 24268
rect 17644 24248 17646 24268
rect 17498 22616 17554 22672
rect 17774 24112 17830 24168
rect 17774 23976 17830 24032
rect 18234 48884 18290 48920
rect 18234 48864 18236 48884
rect 18236 48864 18288 48884
rect 18288 48864 18290 48884
rect 18694 52400 18750 52456
rect 19580 61498 19636 61500
rect 19660 61498 19716 61500
rect 19740 61498 19796 61500
rect 19820 61498 19876 61500
rect 19580 61446 19606 61498
rect 19606 61446 19636 61498
rect 19660 61446 19670 61498
rect 19670 61446 19716 61498
rect 19740 61446 19786 61498
rect 19786 61446 19796 61498
rect 19820 61446 19850 61498
rect 19850 61446 19876 61498
rect 19580 61444 19636 61446
rect 19660 61444 19716 61446
rect 19740 61444 19796 61446
rect 19820 61444 19876 61446
rect 20626 62328 20682 62384
rect 19246 59100 19248 59120
rect 19248 59100 19300 59120
rect 19300 59100 19302 59120
rect 19246 59064 19302 59100
rect 19580 60410 19636 60412
rect 19660 60410 19716 60412
rect 19740 60410 19796 60412
rect 19820 60410 19876 60412
rect 19580 60358 19606 60410
rect 19606 60358 19636 60410
rect 19660 60358 19670 60410
rect 19670 60358 19716 60410
rect 19740 60358 19786 60410
rect 19786 60358 19796 60410
rect 19820 60358 19850 60410
rect 19850 60358 19876 60410
rect 19580 60356 19636 60358
rect 19660 60356 19716 60358
rect 19740 60356 19796 60358
rect 19820 60356 19876 60358
rect 19580 59322 19636 59324
rect 19660 59322 19716 59324
rect 19740 59322 19796 59324
rect 19820 59322 19876 59324
rect 19580 59270 19606 59322
rect 19606 59270 19636 59322
rect 19660 59270 19670 59322
rect 19670 59270 19716 59322
rect 19740 59270 19786 59322
rect 19786 59270 19796 59322
rect 19820 59270 19850 59322
rect 19850 59270 19876 59322
rect 19580 59268 19636 59270
rect 19660 59268 19716 59270
rect 19740 59268 19796 59270
rect 19820 59268 19876 59270
rect 19580 58234 19636 58236
rect 19660 58234 19716 58236
rect 19740 58234 19796 58236
rect 19820 58234 19876 58236
rect 19580 58182 19606 58234
rect 19606 58182 19636 58234
rect 19660 58182 19670 58234
rect 19670 58182 19716 58234
rect 19740 58182 19786 58234
rect 19786 58182 19796 58234
rect 19820 58182 19850 58234
rect 19850 58182 19876 58234
rect 19580 58180 19636 58182
rect 19660 58180 19716 58182
rect 19740 58180 19796 58182
rect 19820 58180 19876 58182
rect 19614 57704 19670 57760
rect 19580 57146 19636 57148
rect 19660 57146 19716 57148
rect 19740 57146 19796 57148
rect 19820 57146 19876 57148
rect 19580 57094 19606 57146
rect 19606 57094 19636 57146
rect 19660 57094 19670 57146
rect 19670 57094 19716 57146
rect 19740 57094 19786 57146
rect 19786 57094 19796 57146
rect 19820 57094 19850 57146
rect 19850 57094 19876 57146
rect 19580 57092 19636 57094
rect 19660 57092 19716 57094
rect 19740 57092 19796 57094
rect 19820 57092 19876 57094
rect 19522 56652 19524 56672
rect 19524 56652 19576 56672
rect 19576 56652 19578 56672
rect 19522 56616 19578 56652
rect 18970 55392 19026 55448
rect 19614 56380 19616 56400
rect 19616 56380 19668 56400
rect 19668 56380 19670 56400
rect 19614 56344 19670 56380
rect 19890 56344 19946 56400
rect 20166 59608 20222 59664
rect 20626 59744 20682 59800
rect 19580 56058 19636 56060
rect 19660 56058 19716 56060
rect 19740 56058 19796 56060
rect 19820 56058 19876 56060
rect 19580 56006 19606 56058
rect 19606 56006 19636 56058
rect 19660 56006 19670 56058
rect 19670 56006 19716 56058
rect 19740 56006 19786 56058
rect 19786 56006 19796 56058
rect 19820 56006 19850 56058
rect 19850 56006 19876 56058
rect 19580 56004 19636 56006
rect 19660 56004 19716 56006
rect 19740 56004 19796 56006
rect 19820 56004 19876 56006
rect 19430 55256 19486 55312
rect 19614 55156 19616 55176
rect 19616 55156 19668 55176
rect 19668 55156 19670 55176
rect 19614 55120 19670 55156
rect 19580 54970 19636 54972
rect 19660 54970 19716 54972
rect 19740 54970 19796 54972
rect 19820 54970 19876 54972
rect 19580 54918 19606 54970
rect 19606 54918 19636 54970
rect 19660 54918 19670 54970
rect 19670 54918 19716 54970
rect 19740 54918 19786 54970
rect 19786 54918 19796 54970
rect 19820 54918 19850 54970
rect 19850 54918 19876 54970
rect 19580 54916 19636 54918
rect 19660 54916 19716 54918
rect 19740 54916 19796 54918
rect 19820 54916 19876 54918
rect 19246 54576 19302 54632
rect 19338 54324 19394 54360
rect 19338 54304 19340 54324
rect 19340 54304 19392 54324
rect 19392 54304 19394 54324
rect 19430 53896 19486 53952
rect 19580 53882 19636 53884
rect 19660 53882 19716 53884
rect 19740 53882 19796 53884
rect 19820 53882 19876 53884
rect 19580 53830 19606 53882
rect 19606 53830 19636 53882
rect 19660 53830 19670 53882
rect 19670 53830 19716 53882
rect 19740 53830 19786 53882
rect 19786 53830 19796 53882
rect 19820 53830 19850 53882
rect 19850 53830 19876 53882
rect 19580 53828 19636 53830
rect 19660 53828 19716 53830
rect 19740 53828 19796 53830
rect 19820 53828 19876 53830
rect 18878 51992 18934 52048
rect 19062 51992 19118 52048
rect 19614 53660 19616 53680
rect 19616 53660 19668 53680
rect 19668 53660 19670 53680
rect 19614 53624 19670 53660
rect 19522 53236 19578 53272
rect 19522 53216 19524 53236
rect 19524 53216 19576 53236
rect 19576 53216 19578 53236
rect 19580 52794 19636 52796
rect 19660 52794 19716 52796
rect 19740 52794 19796 52796
rect 19820 52794 19876 52796
rect 19580 52742 19606 52794
rect 19606 52742 19636 52794
rect 19660 52742 19670 52794
rect 19670 52742 19716 52794
rect 19740 52742 19786 52794
rect 19786 52742 19796 52794
rect 19820 52742 19850 52794
rect 19850 52742 19876 52794
rect 19580 52740 19636 52742
rect 19660 52740 19716 52742
rect 19740 52740 19796 52742
rect 19820 52740 19876 52742
rect 19982 56072 20038 56128
rect 19982 55392 20038 55448
rect 20258 55392 20314 55448
rect 18234 40024 18290 40080
rect 18602 39788 18604 39808
rect 18604 39788 18656 39808
rect 18656 39788 18658 39808
rect 18602 39752 18658 39788
rect 18326 37848 18382 37904
rect 19246 49000 19302 49056
rect 19062 48204 19118 48240
rect 19062 48184 19064 48204
rect 19064 48184 19116 48204
rect 19116 48184 19118 48204
rect 19580 51706 19636 51708
rect 19660 51706 19716 51708
rect 19740 51706 19796 51708
rect 19820 51706 19876 51708
rect 19580 51654 19606 51706
rect 19606 51654 19636 51706
rect 19660 51654 19670 51706
rect 19670 51654 19716 51706
rect 19740 51654 19786 51706
rect 19786 51654 19796 51706
rect 19820 51654 19850 51706
rect 19850 51654 19876 51706
rect 19580 51652 19636 51654
rect 19660 51652 19716 51654
rect 19740 51652 19796 51654
rect 19820 51652 19876 51654
rect 19522 50768 19578 50824
rect 19580 50618 19636 50620
rect 19660 50618 19716 50620
rect 19740 50618 19796 50620
rect 19820 50618 19876 50620
rect 19580 50566 19606 50618
rect 19606 50566 19636 50618
rect 19660 50566 19670 50618
rect 19670 50566 19716 50618
rect 19740 50566 19786 50618
rect 19786 50566 19796 50618
rect 19820 50566 19850 50618
rect 19850 50566 19876 50618
rect 19580 50564 19636 50566
rect 19660 50564 19716 50566
rect 19740 50564 19796 50566
rect 19820 50564 19876 50566
rect 19982 51720 20038 51776
rect 19982 51448 20038 51504
rect 20442 55020 20444 55040
rect 20444 55020 20496 55040
rect 20496 55020 20498 55040
rect 20442 54984 20498 55020
rect 20442 54848 20498 54904
rect 20718 55564 20720 55584
rect 20720 55564 20772 55584
rect 20772 55564 20774 55584
rect 20718 55528 20774 55564
rect 20718 53100 20774 53136
rect 20718 53080 20720 53100
rect 20720 53080 20772 53100
rect 20772 53080 20774 53100
rect 20626 52808 20682 52864
rect 20350 51856 20406 51912
rect 20166 50904 20222 50960
rect 20074 50632 20130 50688
rect 19890 49952 19946 50008
rect 19580 49530 19636 49532
rect 19660 49530 19716 49532
rect 19740 49530 19796 49532
rect 19820 49530 19876 49532
rect 19580 49478 19606 49530
rect 19606 49478 19636 49530
rect 19660 49478 19670 49530
rect 19670 49478 19716 49530
rect 19740 49478 19786 49530
rect 19786 49478 19796 49530
rect 19820 49478 19850 49530
rect 19850 49478 19876 49530
rect 19580 49476 19636 49478
rect 19660 49476 19716 49478
rect 19740 49476 19796 49478
rect 19820 49476 19876 49478
rect 19982 48728 20038 48784
rect 19522 48592 19578 48648
rect 19580 48442 19636 48444
rect 19660 48442 19716 48444
rect 19740 48442 19796 48444
rect 19820 48442 19876 48444
rect 19580 48390 19606 48442
rect 19606 48390 19636 48442
rect 19660 48390 19670 48442
rect 19670 48390 19716 48442
rect 19740 48390 19786 48442
rect 19786 48390 19796 48442
rect 19820 48390 19850 48442
rect 19850 48390 19876 48442
rect 19580 48388 19636 48390
rect 19660 48388 19716 48390
rect 19740 48388 19796 48390
rect 19820 48388 19876 48390
rect 19580 47354 19636 47356
rect 19660 47354 19716 47356
rect 19740 47354 19796 47356
rect 19820 47354 19876 47356
rect 19580 47302 19606 47354
rect 19606 47302 19636 47354
rect 19660 47302 19670 47354
rect 19670 47302 19716 47354
rect 19740 47302 19786 47354
rect 19786 47302 19796 47354
rect 19820 47302 19850 47354
rect 19850 47302 19876 47354
rect 19580 47300 19636 47302
rect 19660 47300 19716 47302
rect 19740 47300 19796 47302
rect 19820 47300 19876 47302
rect 19982 46960 20038 47016
rect 20074 46824 20130 46880
rect 19580 46266 19636 46268
rect 19660 46266 19716 46268
rect 19740 46266 19796 46268
rect 19820 46266 19876 46268
rect 19580 46214 19606 46266
rect 19606 46214 19636 46266
rect 19660 46214 19670 46266
rect 19670 46214 19716 46266
rect 19740 46214 19786 46266
rect 19786 46214 19796 46266
rect 19820 46214 19850 46266
rect 19850 46214 19876 46266
rect 19580 46212 19636 46214
rect 19660 46212 19716 46214
rect 19740 46212 19796 46214
rect 19820 46212 19876 46214
rect 19338 46144 19394 46200
rect 19580 45178 19636 45180
rect 19660 45178 19716 45180
rect 19740 45178 19796 45180
rect 19820 45178 19876 45180
rect 19580 45126 19606 45178
rect 19606 45126 19636 45178
rect 19660 45126 19670 45178
rect 19670 45126 19716 45178
rect 19740 45126 19786 45178
rect 19786 45126 19796 45178
rect 19820 45126 19850 45178
rect 19850 45126 19876 45178
rect 19580 45124 19636 45126
rect 19660 45124 19716 45126
rect 19740 45124 19796 45126
rect 19820 45124 19876 45126
rect 19580 44090 19636 44092
rect 19660 44090 19716 44092
rect 19740 44090 19796 44092
rect 19820 44090 19876 44092
rect 19580 44038 19606 44090
rect 19606 44038 19636 44090
rect 19660 44038 19670 44090
rect 19670 44038 19716 44090
rect 19740 44038 19786 44090
rect 19786 44038 19796 44090
rect 19820 44038 19850 44090
rect 19850 44038 19876 44090
rect 19580 44036 19636 44038
rect 19660 44036 19716 44038
rect 19740 44036 19796 44038
rect 19820 44036 19876 44038
rect 19246 43152 19302 43208
rect 18878 42336 18934 42392
rect 19580 43002 19636 43004
rect 19660 43002 19716 43004
rect 19740 43002 19796 43004
rect 19820 43002 19876 43004
rect 19580 42950 19606 43002
rect 19606 42950 19636 43002
rect 19660 42950 19670 43002
rect 19670 42950 19716 43002
rect 19740 42950 19786 43002
rect 19786 42950 19796 43002
rect 19820 42950 19850 43002
rect 19850 42950 19876 43002
rect 19580 42948 19636 42950
rect 19660 42948 19716 42950
rect 19740 42948 19796 42950
rect 19820 42948 19876 42950
rect 19580 41914 19636 41916
rect 19660 41914 19716 41916
rect 19740 41914 19796 41916
rect 19820 41914 19876 41916
rect 19580 41862 19606 41914
rect 19606 41862 19636 41914
rect 19660 41862 19670 41914
rect 19670 41862 19716 41914
rect 19740 41862 19786 41914
rect 19786 41862 19796 41914
rect 19820 41862 19850 41914
rect 19850 41862 19876 41914
rect 19580 41860 19636 41862
rect 19660 41860 19716 41862
rect 19740 41860 19796 41862
rect 19820 41860 19876 41862
rect 19246 40704 19302 40760
rect 19580 40826 19636 40828
rect 19660 40826 19716 40828
rect 19740 40826 19796 40828
rect 19820 40826 19876 40828
rect 19580 40774 19606 40826
rect 19606 40774 19636 40826
rect 19660 40774 19670 40826
rect 19670 40774 19716 40826
rect 19740 40774 19786 40826
rect 19786 40774 19796 40826
rect 19820 40774 19850 40826
rect 19850 40774 19876 40826
rect 19580 40772 19636 40774
rect 19660 40772 19716 40774
rect 19740 40772 19796 40774
rect 19820 40772 19876 40774
rect 19062 39636 19118 39672
rect 19062 39616 19064 39636
rect 19064 39616 19116 39636
rect 19116 39616 19118 39636
rect 19706 39888 19762 39944
rect 19580 39738 19636 39740
rect 19660 39738 19716 39740
rect 19740 39738 19796 39740
rect 19820 39738 19876 39740
rect 19580 39686 19606 39738
rect 19606 39686 19636 39738
rect 19660 39686 19670 39738
rect 19670 39686 19716 39738
rect 19740 39686 19786 39738
rect 19786 39686 19796 39738
rect 19820 39686 19850 39738
rect 19850 39686 19876 39738
rect 19580 39684 19636 39686
rect 19660 39684 19716 39686
rect 19740 39684 19796 39686
rect 19820 39684 19876 39686
rect 18694 38664 18750 38720
rect 19580 38650 19636 38652
rect 19660 38650 19716 38652
rect 19740 38650 19796 38652
rect 19820 38650 19876 38652
rect 19580 38598 19606 38650
rect 19606 38598 19636 38650
rect 19660 38598 19670 38650
rect 19670 38598 19716 38650
rect 19740 38598 19786 38650
rect 19786 38598 19796 38650
rect 19820 38598 19850 38650
rect 19850 38598 19876 38650
rect 19580 38596 19636 38598
rect 19660 38596 19716 38598
rect 19740 38596 19796 38598
rect 19820 38596 19876 38598
rect 18786 38256 18842 38312
rect 18602 37848 18658 37904
rect 18418 37304 18474 37360
rect 18326 34584 18382 34640
rect 18326 33496 18382 33552
rect 18326 32408 18382 32464
rect 18786 37032 18842 37088
rect 18326 31884 18382 31920
rect 18326 31864 18328 31884
rect 18328 31864 18380 31884
rect 18380 31864 18382 31884
rect 18234 31728 18290 31784
rect 18418 31728 18474 31784
rect 18602 36216 18658 36272
rect 18970 37712 19026 37768
rect 19798 38004 19854 38040
rect 19798 37984 19800 38004
rect 19800 37984 19852 38004
rect 19852 37984 19854 38004
rect 19580 37562 19636 37564
rect 19660 37562 19716 37564
rect 19740 37562 19796 37564
rect 19820 37562 19876 37564
rect 19580 37510 19606 37562
rect 19606 37510 19636 37562
rect 19660 37510 19670 37562
rect 19670 37510 19716 37562
rect 19740 37510 19786 37562
rect 19786 37510 19796 37562
rect 19820 37510 19850 37562
rect 19850 37510 19876 37562
rect 19580 37508 19636 37510
rect 19660 37508 19716 37510
rect 19740 37508 19796 37510
rect 19820 37508 19876 37510
rect 20074 37576 20130 37632
rect 18694 33632 18750 33688
rect 18694 32952 18750 33008
rect 18234 30232 18290 30288
rect 18510 31456 18566 31512
rect 18418 30504 18474 30560
rect 18418 28736 18474 28792
rect 18234 24112 18290 24168
rect 18786 32836 18842 32872
rect 18786 32816 18788 32836
rect 18788 32816 18840 32836
rect 18840 32816 18842 32836
rect 18786 32544 18842 32600
rect 18786 32000 18842 32056
rect 19580 36474 19636 36476
rect 19660 36474 19716 36476
rect 19740 36474 19796 36476
rect 19820 36474 19876 36476
rect 19580 36422 19606 36474
rect 19606 36422 19636 36474
rect 19660 36422 19670 36474
rect 19670 36422 19716 36474
rect 19740 36422 19786 36474
rect 19786 36422 19796 36474
rect 19820 36422 19850 36474
rect 19850 36422 19876 36474
rect 19580 36420 19636 36422
rect 19660 36420 19716 36422
rect 19740 36420 19796 36422
rect 19820 36420 19876 36422
rect 19338 36352 19394 36408
rect 19154 35808 19210 35864
rect 19338 35944 19394 36000
rect 19580 35386 19636 35388
rect 19660 35386 19716 35388
rect 19740 35386 19796 35388
rect 19820 35386 19876 35388
rect 19580 35334 19606 35386
rect 19606 35334 19636 35386
rect 19660 35334 19670 35386
rect 19670 35334 19716 35386
rect 19740 35334 19786 35386
rect 19786 35334 19796 35386
rect 19820 35334 19850 35386
rect 19850 35334 19876 35386
rect 19580 35332 19636 35334
rect 19660 35332 19716 35334
rect 19740 35332 19796 35334
rect 19820 35332 19876 35334
rect 19338 35148 19394 35184
rect 19338 35128 19340 35148
rect 19340 35128 19392 35148
rect 19392 35128 19394 35148
rect 19614 34720 19670 34776
rect 19338 34176 19394 34232
rect 19154 33224 19210 33280
rect 19580 34298 19636 34300
rect 19660 34298 19716 34300
rect 19740 34298 19796 34300
rect 19820 34298 19876 34300
rect 19580 34246 19606 34298
rect 19606 34246 19636 34298
rect 19660 34246 19670 34298
rect 19670 34246 19716 34298
rect 19740 34246 19786 34298
rect 19786 34246 19796 34298
rect 19820 34246 19850 34298
rect 19850 34246 19876 34298
rect 19580 34244 19636 34246
rect 19660 34244 19716 34246
rect 19740 34244 19796 34246
rect 19820 34244 19876 34246
rect 19430 33904 19486 33960
rect 19614 33904 19670 33960
rect 18878 31320 18934 31376
rect 18602 30640 18658 30696
rect 19062 30640 19118 30696
rect 18786 30116 18842 30152
rect 18786 30096 18788 30116
rect 18788 30096 18840 30116
rect 18840 30096 18842 30116
rect 18970 29416 19026 29472
rect 18878 28620 18934 28656
rect 18878 28600 18880 28620
rect 18880 28600 18932 28620
rect 18932 28600 18934 28620
rect 18878 28328 18934 28384
rect 18786 28056 18842 28112
rect 18694 27240 18750 27296
rect 18970 27376 19026 27432
rect 18326 23860 18382 23896
rect 18326 23840 18328 23860
rect 18328 23840 18380 23860
rect 18380 23840 18382 23860
rect 18694 25780 18696 25800
rect 18696 25780 18748 25800
rect 18748 25780 18750 25800
rect 18694 25744 18750 25780
rect 18786 25608 18842 25664
rect 18694 24928 18750 24984
rect 18326 22500 18382 22536
rect 18326 22480 18328 22500
rect 18328 22480 18380 22500
rect 18380 22480 18382 22500
rect 18510 22344 18566 22400
rect 18602 22072 18658 22128
rect 18418 21936 18474 21992
rect 18142 19760 18198 19816
rect 17958 18400 18014 18456
rect 15566 8472 15622 8528
rect 16486 13368 16542 13424
rect 18050 15680 18106 15736
rect 18326 15156 18382 15192
rect 18326 15136 18328 15156
rect 18328 15136 18380 15156
rect 18380 15136 18382 15156
rect 18326 14356 18328 14376
rect 18328 14356 18380 14376
rect 18380 14356 18382 14376
rect 18326 14320 18382 14356
rect 16118 9696 16174 9752
rect 17038 9696 17094 9752
rect 16026 5208 16082 5264
rect 15842 3984 15898 4040
rect 17038 3984 17094 4040
rect 18970 26460 18972 26480
rect 18972 26460 19024 26480
rect 19024 26460 19026 26480
rect 18970 26424 19026 26460
rect 19580 33210 19636 33212
rect 19660 33210 19716 33212
rect 19740 33210 19796 33212
rect 19820 33210 19876 33212
rect 19580 33158 19606 33210
rect 19606 33158 19636 33210
rect 19660 33158 19670 33210
rect 19670 33158 19716 33210
rect 19740 33158 19786 33210
rect 19786 33158 19796 33210
rect 19820 33158 19850 33210
rect 19850 33158 19876 33210
rect 19580 33156 19636 33158
rect 19660 33156 19716 33158
rect 19740 33156 19796 33158
rect 19820 33156 19876 33158
rect 20074 35012 20130 35048
rect 20074 34992 20076 35012
rect 20076 34992 20128 35012
rect 20128 34992 20130 35012
rect 20074 34856 20130 34912
rect 19982 34312 20038 34368
rect 19580 32122 19636 32124
rect 19660 32122 19716 32124
rect 19740 32122 19796 32124
rect 19820 32122 19876 32124
rect 19580 32070 19606 32122
rect 19606 32070 19636 32122
rect 19660 32070 19670 32122
rect 19670 32070 19716 32122
rect 19740 32070 19786 32122
rect 19786 32070 19796 32122
rect 19820 32070 19850 32122
rect 19850 32070 19876 32122
rect 19580 32068 19636 32070
rect 19660 32068 19716 32070
rect 19740 32068 19796 32070
rect 19820 32068 19876 32070
rect 19890 31456 19946 31512
rect 19614 31184 19670 31240
rect 19890 31184 19946 31240
rect 19580 31034 19636 31036
rect 19660 31034 19716 31036
rect 19740 31034 19796 31036
rect 19820 31034 19876 31036
rect 19580 30982 19606 31034
rect 19606 30982 19636 31034
rect 19660 30982 19670 31034
rect 19670 30982 19716 31034
rect 19740 30982 19786 31034
rect 19786 30982 19796 31034
rect 19820 30982 19850 31034
rect 19850 30982 19876 31034
rect 19580 30980 19636 30982
rect 19660 30980 19716 30982
rect 19740 30980 19796 30982
rect 19820 30980 19876 30982
rect 19246 30232 19302 30288
rect 19154 29164 19210 29200
rect 19154 29144 19156 29164
rect 19156 29144 19208 29164
rect 19208 29144 19210 29164
rect 19246 28872 19302 28928
rect 19580 29946 19636 29948
rect 19660 29946 19716 29948
rect 19740 29946 19796 29948
rect 19820 29946 19876 29948
rect 19580 29894 19606 29946
rect 19606 29894 19636 29946
rect 19660 29894 19670 29946
rect 19670 29894 19716 29946
rect 19740 29894 19786 29946
rect 19786 29894 19796 29946
rect 19820 29894 19850 29946
rect 19850 29894 19876 29946
rect 19580 29892 19636 29894
rect 19660 29892 19716 29894
rect 19740 29892 19796 29894
rect 19820 29892 19876 29894
rect 19982 30776 20038 30832
rect 20074 29960 20130 30016
rect 19982 29280 20038 29336
rect 19522 29144 19578 29200
rect 19580 28858 19636 28860
rect 19660 28858 19716 28860
rect 19740 28858 19796 28860
rect 19820 28858 19876 28860
rect 19580 28806 19606 28858
rect 19606 28806 19636 28858
rect 19660 28806 19670 28858
rect 19670 28806 19716 28858
rect 19740 28806 19786 28858
rect 19786 28806 19796 28858
rect 19820 28806 19850 28858
rect 19850 28806 19876 28858
rect 19580 28804 19636 28806
rect 19660 28804 19716 28806
rect 19740 28804 19796 28806
rect 19820 28804 19876 28806
rect 19890 28328 19946 28384
rect 19580 27770 19636 27772
rect 19660 27770 19716 27772
rect 19740 27770 19796 27772
rect 19820 27770 19876 27772
rect 19580 27718 19606 27770
rect 19606 27718 19636 27770
rect 19660 27718 19670 27770
rect 19670 27718 19716 27770
rect 19740 27718 19786 27770
rect 19786 27718 19796 27770
rect 19820 27718 19850 27770
rect 19850 27718 19876 27770
rect 19580 27716 19636 27718
rect 19660 27716 19716 27718
rect 19740 27716 19796 27718
rect 19820 27716 19876 27718
rect 19430 27648 19486 27704
rect 19430 27104 19486 27160
rect 19430 26868 19432 26888
rect 19432 26868 19484 26888
rect 19484 26868 19486 26888
rect 19430 26832 19486 26868
rect 19580 26682 19636 26684
rect 19660 26682 19716 26684
rect 19740 26682 19796 26684
rect 19820 26682 19876 26684
rect 19580 26630 19606 26682
rect 19606 26630 19636 26682
rect 19660 26630 19670 26682
rect 19670 26630 19716 26682
rect 19740 26630 19786 26682
rect 19786 26630 19796 26682
rect 19820 26630 19850 26682
rect 19850 26630 19876 26682
rect 19580 26628 19636 26630
rect 19660 26628 19716 26630
rect 19740 26628 19796 26630
rect 19820 26628 19876 26630
rect 19154 25880 19210 25936
rect 19614 26152 19670 26208
rect 19580 25594 19636 25596
rect 19660 25594 19716 25596
rect 19740 25594 19796 25596
rect 19820 25594 19876 25596
rect 19580 25542 19606 25594
rect 19606 25542 19636 25594
rect 19660 25542 19670 25594
rect 19670 25542 19716 25594
rect 19740 25542 19786 25594
rect 19786 25542 19796 25594
rect 19820 25542 19850 25594
rect 19850 25542 19876 25594
rect 19580 25540 19636 25542
rect 19660 25540 19716 25542
rect 19740 25540 19796 25542
rect 19820 25540 19876 25542
rect 19798 25200 19854 25256
rect 19580 24506 19636 24508
rect 19660 24506 19716 24508
rect 19740 24506 19796 24508
rect 19820 24506 19876 24508
rect 19580 24454 19606 24506
rect 19606 24454 19636 24506
rect 19660 24454 19670 24506
rect 19670 24454 19716 24506
rect 19740 24454 19786 24506
rect 19786 24454 19796 24506
rect 19820 24454 19850 24506
rect 19850 24454 19876 24506
rect 19580 24452 19636 24454
rect 19660 24452 19716 24454
rect 19740 24452 19796 24454
rect 19820 24452 19876 24454
rect 18786 22208 18842 22264
rect 19430 24248 19486 24304
rect 19246 23840 19302 23896
rect 19154 23024 19210 23080
rect 18786 21664 18842 21720
rect 19580 23418 19636 23420
rect 19660 23418 19716 23420
rect 19740 23418 19796 23420
rect 19820 23418 19876 23420
rect 19580 23366 19606 23418
rect 19606 23366 19636 23418
rect 19660 23366 19670 23418
rect 19670 23366 19716 23418
rect 19740 23366 19786 23418
rect 19786 23366 19796 23418
rect 19820 23366 19850 23418
rect 19850 23366 19876 23418
rect 19580 23364 19636 23366
rect 19660 23364 19716 23366
rect 19740 23364 19796 23366
rect 19820 23364 19876 23366
rect 20074 23976 20130 24032
rect 19154 21528 19210 21584
rect 18786 20984 18842 21040
rect 18970 20848 19026 20904
rect 19580 22330 19636 22332
rect 19660 22330 19716 22332
rect 19740 22330 19796 22332
rect 19820 22330 19876 22332
rect 19580 22278 19606 22330
rect 19606 22278 19636 22330
rect 19660 22278 19670 22330
rect 19670 22278 19716 22330
rect 19740 22278 19786 22330
rect 19786 22278 19796 22330
rect 19820 22278 19850 22330
rect 19850 22278 19876 22330
rect 19580 22276 19636 22278
rect 19660 22276 19716 22278
rect 19740 22276 19796 22278
rect 19820 22276 19876 22278
rect 20074 23024 20130 23080
rect 19890 21936 19946 21992
rect 19614 21548 19670 21584
rect 19614 21528 19616 21548
rect 19616 21528 19668 21548
rect 19668 21528 19670 21548
rect 19580 21242 19636 21244
rect 19660 21242 19716 21244
rect 19740 21242 19796 21244
rect 19820 21242 19876 21244
rect 19580 21190 19606 21242
rect 19606 21190 19636 21242
rect 19660 21190 19670 21242
rect 19670 21190 19716 21242
rect 19740 21190 19786 21242
rect 19786 21190 19796 21242
rect 19820 21190 19850 21242
rect 19850 21190 19876 21242
rect 19580 21188 19636 21190
rect 19660 21188 19716 21190
rect 19740 21188 19796 21190
rect 19820 21188 19876 21190
rect 19522 20440 19578 20496
rect 19580 20154 19636 20156
rect 19660 20154 19716 20156
rect 19740 20154 19796 20156
rect 19820 20154 19876 20156
rect 19580 20102 19606 20154
rect 19606 20102 19636 20154
rect 19660 20102 19670 20154
rect 19670 20102 19716 20154
rect 19740 20102 19786 20154
rect 19786 20102 19796 20154
rect 19820 20102 19850 20154
rect 19850 20102 19876 20154
rect 19580 20100 19636 20102
rect 19660 20100 19716 20102
rect 19740 20100 19796 20102
rect 19820 20100 19876 20102
rect 19154 19252 19156 19272
rect 19156 19252 19208 19272
rect 19208 19252 19210 19272
rect 19154 19216 19210 19252
rect 19580 19066 19636 19068
rect 19660 19066 19716 19068
rect 19740 19066 19796 19068
rect 19820 19066 19876 19068
rect 19580 19014 19606 19066
rect 19606 19014 19636 19066
rect 19660 19014 19670 19066
rect 19670 19014 19716 19066
rect 19740 19014 19786 19066
rect 19786 19014 19796 19066
rect 19820 19014 19850 19066
rect 19850 19014 19876 19066
rect 19580 19012 19636 19014
rect 19660 19012 19716 19014
rect 19740 19012 19796 19014
rect 19820 19012 19876 19014
rect 19580 17978 19636 17980
rect 19660 17978 19716 17980
rect 19740 17978 19796 17980
rect 19820 17978 19876 17980
rect 19580 17926 19606 17978
rect 19606 17926 19636 17978
rect 19660 17926 19670 17978
rect 19670 17926 19716 17978
rect 19740 17926 19786 17978
rect 19786 17926 19796 17978
rect 19820 17926 19850 17978
rect 19850 17926 19876 17978
rect 19580 17924 19636 17926
rect 19660 17924 19716 17926
rect 19740 17924 19796 17926
rect 19820 17924 19876 17926
rect 20074 17856 20130 17912
rect 19580 16890 19636 16892
rect 19660 16890 19716 16892
rect 19740 16890 19796 16892
rect 19820 16890 19876 16892
rect 19580 16838 19606 16890
rect 19606 16838 19636 16890
rect 19660 16838 19670 16890
rect 19670 16838 19716 16890
rect 19740 16838 19786 16890
rect 19786 16838 19796 16890
rect 19820 16838 19850 16890
rect 19850 16838 19876 16890
rect 19580 16836 19636 16838
rect 19660 16836 19716 16838
rect 19740 16836 19796 16838
rect 19820 16836 19876 16838
rect 19154 16496 19210 16552
rect 18970 14456 19026 14512
rect 18510 9016 18566 9072
rect 18878 9016 18934 9072
rect 18234 3304 18290 3360
rect 19580 15802 19636 15804
rect 19660 15802 19716 15804
rect 19740 15802 19796 15804
rect 19820 15802 19876 15804
rect 19580 15750 19606 15802
rect 19606 15750 19636 15802
rect 19660 15750 19670 15802
rect 19670 15750 19716 15802
rect 19740 15750 19786 15802
rect 19786 15750 19796 15802
rect 19820 15750 19850 15802
rect 19850 15750 19876 15802
rect 19580 15748 19636 15750
rect 19660 15748 19716 15750
rect 19740 15748 19796 15750
rect 19820 15748 19876 15750
rect 20350 48864 20406 48920
rect 20258 48320 20314 48376
rect 20718 51584 20774 51640
rect 20626 49136 20682 49192
rect 20718 40568 20774 40624
rect 20258 37168 20314 37224
rect 20350 34176 20406 34232
rect 21178 76356 21234 76392
rect 21178 76336 21180 76356
rect 21180 76336 21232 76356
rect 21232 76336 21234 76356
rect 21362 75248 21418 75304
rect 21270 74432 21326 74488
rect 21086 71848 21142 71904
rect 20902 69672 20958 69728
rect 20902 67924 20958 67960
rect 20902 67904 20904 67924
rect 20904 67904 20956 67924
rect 20956 67904 20958 67924
rect 20902 59084 20958 59120
rect 20902 59064 20904 59084
rect 20904 59064 20956 59084
rect 20956 59064 20958 59084
rect 20902 56228 20958 56264
rect 20902 56208 20904 56228
rect 20904 56208 20956 56228
rect 20956 56208 20958 56228
rect 20902 54168 20958 54224
rect 20994 52400 21050 52456
rect 20902 51856 20958 51912
rect 20902 50768 20958 50824
rect 21086 49716 21088 49736
rect 21088 49716 21140 49736
rect 21140 49716 21142 49736
rect 21086 49680 21142 49716
rect 21178 48864 21234 48920
rect 20994 47232 21050 47288
rect 21178 47096 21234 47152
rect 20810 37460 20866 37496
rect 20810 37440 20812 37460
rect 20812 37440 20864 37460
rect 20864 37440 20866 37460
rect 21086 38292 21088 38312
rect 21088 38292 21140 38312
rect 21140 38292 21142 38312
rect 21086 38256 21142 38292
rect 20994 37848 21050 37904
rect 20902 37168 20958 37224
rect 20902 36216 20958 36272
rect 21086 35672 21142 35728
rect 20994 35536 21050 35592
rect 20534 34448 20590 34504
rect 20902 34856 20958 34912
rect 20810 34620 20812 34640
rect 20812 34620 20864 34640
rect 20864 34620 20866 34640
rect 20810 34584 20866 34620
rect 20902 34448 20958 34504
rect 20534 33224 20590 33280
rect 20718 33632 20774 33688
rect 20994 33360 21050 33416
rect 20718 33088 20774 33144
rect 20626 32136 20682 32192
rect 20810 32680 20866 32736
rect 21822 73208 21878 73264
rect 21362 67496 21418 67552
rect 21730 63416 21786 63472
rect 21546 59472 21602 59528
rect 21454 58248 21510 58304
rect 21638 57840 21694 57896
rect 21362 56752 21418 56808
rect 21454 56616 21510 56672
rect 21546 56480 21602 56536
rect 21454 55664 21510 55720
rect 21362 55120 21418 55176
rect 21546 54576 21602 54632
rect 21362 54032 21418 54088
rect 21638 53896 21694 53952
rect 21546 51892 21548 51912
rect 21548 51892 21600 51912
rect 21600 51892 21602 51912
rect 21546 51856 21602 51892
rect 21546 51584 21602 51640
rect 22834 69808 22890 69864
rect 22190 67496 22246 67552
rect 22006 62092 22008 62112
rect 22008 62092 22060 62112
rect 22060 62092 22062 62112
rect 22006 62056 22062 62092
rect 22006 60288 22062 60344
rect 22282 66680 22338 66736
rect 22466 62192 22522 62248
rect 22374 59744 22430 59800
rect 22098 59608 22154 59664
rect 22558 59744 22614 59800
rect 21914 56616 21970 56672
rect 24398 77172 24454 77208
rect 24398 77152 24400 77172
rect 24400 77152 24452 77172
rect 24452 77152 24454 77172
rect 24122 76336 24178 76392
rect 24674 76064 24730 76120
rect 25870 76064 25926 76120
rect 24766 74432 24822 74488
rect 23938 73208 23994 73264
rect 23018 70896 23074 70952
rect 24306 70932 24308 70952
rect 24308 70932 24360 70952
rect 24360 70932 24362 70952
rect 24306 70896 24362 70932
rect 22650 57976 22706 58032
rect 22098 55936 22154 55992
rect 22466 55700 22468 55720
rect 22468 55700 22520 55720
rect 22520 55700 22522 55720
rect 22466 55664 22522 55700
rect 22466 54440 22522 54496
rect 22282 52980 22284 53000
rect 22284 52980 22336 53000
rect 22336 52980 22338 53000
rect 22282 52944 22338 52980
rect 22374 52536 22430 52592
rect 21822 51992 21878 52048
rect 22282 52128 22338 52184
rect 21730 51040 21786 51096
rect 22006 50924 22062 50960
rect 22006 50904 22008 50924
rect 22008 50904 22060 50924
rect 22060 50904 22062 50924
rect 21822 50768 21878 50824
rect 21362 47776 21418 47832
rect 21362 41012 21364 41032
rect 21364 41012 21416 41032
rect 21416 41012 21418 41032
rect 21362 40976 21418 41012
rect 21638 38800 21694 38856
rect 21638 37984 21694 38040
rect 21546 37868 21602 37904
rect 21546 37848 21548 37868
rect 21548 37848 21600 37868
rect 21600 37848 21602 37868
rect 21638 37304 21694 37360
rect 21362 34584 21418 34640
rect 21178 32680 21234 32736
rect 20350 31048 20406 31104
rect 20258 27920 20314 27976
rect 20258 27668 20314 27704
rect 20258 27648 20260 27668
rect 20260 27648 20312 27668
rect 20312 27648 20314 27668
rect 20442 24928 20498 24984
rect 20442 24656 20498 24712
rect 20442 22208 20498 22264
rect 20350 22072 20406 22128
rect 20718 30368 20774 30424
rect 20810 29824 20866 29880
rect 20718 28464 20774 28520
rect 20626 26852 20682 26888
rect 20626 26832 20628 26852
rect 20628 26832 20680 26852
rect 20680 26832 20682 26852
rect 20994 32136 21050 32192
rect 20994 31728 21050 31784
rect 21454 33088 21510 33144
rect 21730 33768 21786 33824
rect 21638 33632 21694 33688
rect 21546 32272 21602 32328
rect 21454 31320 21510 31376
rect 21362 30640 21418 30696
rect 21270 30368 21326 30424
rect 21454 30504 21510 30560
rect 21178 29688 21234 29744
rect 20810 27956 20812 27976
rect 20812 27956 20864 27976
rect 20864 27956 20866 27976
rect 20810 27920 20866 27956
rect 20994 28464 21050 28520
rect 20902 26424 20958 26480
rect 20902 26016 20958 26072
rect 21730 32544 21786 32600
rect 21270 28600 21326 28656
rect 21178 27648 21234 27704
rect 21270 27512 21326 27568
rect 21086 26016 21142 26072
rect 20810 25608 20866 25664
rect 20810 24792 20866 24848
rect 20994 25744 21050 25800
rect 21546 29552 21602 29608
rect 21454 27784 21510 27840
rect 21730 28076 21786 28112
rect 21730 28056 21732 28076
rect 21732 28056 21784 28076
rect 21784 28056 21786 28076
rect 21454 26696 21510 26752
rect 21454 26444 21510 26480
rect 21454 26424 21456 26444
rect 21456 26424 21508 26444
rect 21508 26424 21510 26444
rect 21270 25472 21326 25528
rect 21086 24692 21088 24712
rect 21088 24692 21140 24712
rect 21140 24692 21142 24712
rect 21086 24656 21142 24692
rect 20442 21428 20444 21448
rect 20444 21428 20496 21448
rect 20496 21428 20498 21448
rect 20442 21392 20498 21428
rect 21178 23160 21234 23216
rect 21178 22480 21234 22536
rect 21178 22344 21234 22400
rect 21086 20984 21142 21040
rect 21730 27240 21786 27296
rect 21454 24112 21510 24168
rect 21546 23976 21602 24032
rect 21546 23604 21548 23624
rect 21548 23604 21600 23624
rect 21600 23604 21602 23624
rect 21546 23568 21602 23604
rect 21638 23024 21694 23080
rect 21546 22888 21602 22944
rect 21454 22616 21510 22672
rect 21362 21664 21418 21720
rect 21086 19780 21142 19816
rect 21086 19760 21088 19780
rect 21088 19760 21140 19780
rect 21140 19760 21142 19780
rect 21178 15564 21234 15600
rect 21178 15544 21180 15564
rect 21180 15544 21232 15564
rect 21232 15544 21234 15564
rect 20166 15408 20222 15464
rect 19580 14714 19636 14716
rect 19660 14714 19716 14716
rect 19740 14714 19796 14716
rect 19820 14714 19876 14716
rect 19580 14662 19606 14714
rect 19606 14662 19636 14714
rect 19660 14662 19670 14714
rect 19670 14662 19716 14714
rect 19740 14662 19786 14714
rect 19786 14662 19796 14714
rect 19820 14662 19850 14714
rect 19850 14662 19876 14714
rect 19580 14660 19636 14662
rect 19660 14660 19716 14662
rect 19740 14660 19796 14662
rect 19820 14660 19876 14662
rect 21270 14320 21326 14376
rect 19580 13626 19636 13628
rect 19660 13626 19716 13628
rect 19740 13626 19796 13628
rect 19820 13626 19876 13628
rect 19580 13574 19606 13626
rect 19606 13574 19636 13626
rect 19660 13574 19670 13626
rect 19670 13574 19716 13626
rect 19740 13574 19786 13626
rect 19786 13574 19796 13626
rect 19820 13574 19850 13626
rect 19850 13574 19876 13626
rect 19580 13572 19636 13574
rect 19660 13572 19716 13574
rect 19740 13572 19796 13574
rect 19820 13572 19876 13574
rect 19580 12538 19636 12540
rect 19660 12538 19716 12540
rect 19740 12538 19796 12540
rect 19820 12538 19876 12540
rect 19580 12486 19606 12538
rect 19606 12486 19636 12538
rect 19660 12486 19670 12538
rect 19670 12486 19716 12538
rect 19740 12486 19786 12538
rect 19786 12486 19796 12538
rect 19820 12486 19850 12538
rect 19850 12486 19876 12538
rect 19580 12484 19636 12486
rect 19660 12484 19716 12486
rect 19740 12484 19796 12486
rect 19820 12484 19876 12486
rect 21638 19488 21694 19544
rect 19580 11450 19636 11452
rect 19660 11450 19716 11452
rect 19740 11450 19796 11452
rect 19820 11450 19876 11452
rect 19580 11398 19606 11450
rect 19606 11398 19636 11450
rect 19660 11398 19670 11450
rect 19670 11398 19716 11450
rect 19740 11398 19786 11450
rect 19786 11398 19796 11450
rect 19820 11398 19850 11450
rect 19850 11398 19876 11450
rect 19580 11396 19636 11398
rect 19660 11396 19716 11398
rect 19740 11396 19796 11398
rect 19820 11396 19876 11398
rect 19580 10362 19636 10364
rect 19660 10362 19716 10364
rect 19740 10362 19796 10364
rect 19820 10362 19876 10364
rect 19580 10310 19606 10362
rect 19606 10310 19636 10362
rect 19660 10310 19670 10362
rect 19670 10310 19716 10362
rect 19740 10310 19786 10362
rect 19786 10310 19796 10362
rect 19820 10310 19850 10362
rect 19850 10310 19876 10362
rect 19580 10308 19636 10310
rect 19660 10308 19716 10310
rect 19740 10308 19796 10310
rect 19820 10308 19876 10310
rect 19982 10240 20038 10296
rect 19430 9424 19486 9480
rect 19580 9274 19636 9276
rect 19660 9274 19716 9276
rect 19740 9274 19796 9276
rect 19820 9274 19876 9276
rect 19580 9222 19606 9274
rect 19606 9222 19636 9274
rect 19660 9222 19670 9274
rect 19670 9222 19716 9274
rect 19740 9222 19786 9274
rect 19786 9222 19796 9274
rect 19820 9222 19850 9274
rect 19850 9222 19876 9274
rect 19580 9220 19636 9222
rect 19660 9220 19716 9222
rect 19740 9220 19796 9222
rect 19820 9220 19876 9222
rect 19580 8186 19636 8188
rect 19660 8186 19716 8188
rect 19740 8186 19796 8188
rect 19820 8186 19876 8188
rect 19580 8134 19606 8186
rect 19606 8134 19636 8186
rect 19660 8134 19670 8186
rect 19670 8134 19716 8186
rect 19740 8134 19786 8186
rect 19786 8134 19796 8186
rect 19820 8134 19850 8186
rect 19850 8134 19876 8186
rect 19580 8132 19636 8134
rect 19660 8132 19716 8134
rect 19740 8132 19796 8134
rect 19820 8132 19876 8134
rect 19580 7098 19636 7100
rect 19660 7098 19716 7100
rect 19740 7098 19796 7100
rect 19820 7098 19876 7100
rect 19580 7046 19606 7098
rect 19606 7046 19636 7098
rect 19660 7046 19670 7098
rect 19670 7046 19716 7098
rect 19740 7046 19786 7098
rect 19786 7046 19796 7098
rect 19820 7046 19850 7098
rect 19850 7046 19876 7098
rect 19580 7044 19636 7046
rect 19660 7044 19716 7046
rect 19740 7044 19796 7046
rect 19820 7044 19876 7046
rect 19430 6840 19486 6896
rect 19580 6010 19636 6012
rect 19660 6010 19716 6012
rect 19740 6010 19796 6012
rect 19820 6010 19876 6012
rect 19580 5958 19606 6010
rect 19606 5958 19636 6010
rect 19660 5958 19670 6010
rect 19670 5958 19716 6010
rect 19740 5958 19786 6010
rect 19786 5958 19796 6010
rect 19820 5958 19850 6010
rect 19850 5958 19876 6010
rect 19580 5956 19636 5958
rect 19660 5956 19716 5958
rect 19740 5956 19796 5958
rect 19820 5956 19876 5958
rect 19580 4922 19636 4924
rect 19660 4922 19716 4924
rect 19740 4922 19796 4924
rect 19820 4922 19876 4924
rect 19580 4870 19606 4922
rect 19606 4870 19636 4922
rect 19660 4870 19670 4922
rect 19670 4870 19716 4922
rect 19740 4870 19786 4922
rect 19786 4870 19796 4922
rect 19820 4870 19850 4922
rect 19850 4870 19876 4922
rect 19580 4868 19636 4870
rect 19660 4868 19716 4870
rect 19740 4868 19796 4870
rect 19820 4868 19876 4870
rect 19246 4256 19302 4312
rect 19430 4256 19486 4312
rect 19580 3834 19636 3836
rect 19660 3834 19716 3836
rect 19740 3834 19796 3836
rect 19820 3834 19876 3836
rect 19580 3782 19606 3834
rect 19606 3782 19636 3834
rect 19660 3782 19670 3834
rect 19670 3782 19716 3834
rect 19740 3782 19786 3834
rect 19786 3782 19796 3834
rect 19820 3782 19850 3834
rect 19850 3782 19876 3834
rect 19580 3780 19636 3782
rect 19660 3780 19716 3782
rect 19740 3780 19796 3782
rect 19820 3780 19876 3782
rect 19430 3340 19432 3360
rect 19432 3340 19484 3360
rect 19484 3340 19486 3360
rect 19430 3304 19486 3340
rect 19580 2746 19636 2748
rect 19660 2746 19716 2748
rect 19740 2746 19796 2748
rect 19820 2746 19876 2748
rect 19580 2694 19606 2746
rect 19606 2694 19636 2746
rect 19660 2694 19670 2746
rect 19670 2694 19716 2746
rect 19740 2694 19786 2746
rect 19786 2694 19796 2746
rect 19820 2694 19850 2746
rect 19850 2694 19876 2746
rect 19580 2692 19636 2694
rect 19660 2692 19716 2694
rect 19740 2692 19796 2694
rect 19820 2692 19876 2694
rect 18970 2216 19026 2272
rect 22190 49272 22246 49328
rect 22834 58112 22890 58168
rect 23018 55936 23074 55992
rect 22742 54576 22798 54632
rect 22466 49000 22522 49056
rect 22374 48220 22376 48240
rect 22376 48220 22428 48240
rect 22428 48220 22430 48240
rect 22374 48184 22430 48220
rect 22742 48628 22744 48648
rect 22744 48628 22796 48648
rect 22796 48628 22798 48648
rect 22742 48592 22798 48628
rect 21914 46980 21970 47016
rect 21914 46960 21916 46980
rect 21916 46960 21968 46980
rect 21968 46960 21970 46980
rect 22466 46824 22522 46880
rect 22282 37168 22338 37224
rect 22374 36080 22430 36136
rect 22098 34348 22100 34368
rect 22100 34348 22152 34368
rect 22152 34348 22154 34368
rect 22098 34312 22154 34348
rect 22006 33360 22062 33416
rect 22006 30676 22008 30696
rect 22008 30676 22060 30696
rect 22060 30676 22062 30696
rect 22006 30640 22062 30676
rect 22742 37712 22798 37768
rect 22650 35808 22706 35864
rect 22098 29960 22154 30016
rect 22098 28464 22154 28520
rect 22282 29008 22338 29064
rect 22190 27512 22246 27568
rect 22006 24384 22062 24440
rect 22006 23024 22062 23080
rect 22006 22652 22008 22672
rect 22008 22652 22060 22672
rect 22060 22652 22062 22672
rect 22006 22616 22062 22652
rect 21914 21800 21970 21856
rect 22282 27104 22338 27160
rect 22190 25336 22246 25392
rect 22190 25064 22246 25120
rect 22190 20576 22246 20632
rect 22190 17856 22246 17912
rect 22006 13912 22062 13968
rect 22098 13504 22154 13560
rect 22098 9968 22154 10024
rect 22466 33496 22522 33552
rect 22558 30388 22614 30424
rect 22558 30368 22560 30388
rect 22560 30368 22612 30388
rect 22612 30368 22614 30388
rect 22558 29996 22560 30016
rect 22560 29996 22612 30016
rect 22612 29996 22614 30016
rect 22558 29960 22614 29996
rect 22466 29044 22468 29064
rect 22468 29044 22520 29064
rect 22520 29044 22522 29064
rect 22466 29008 22522 29044
rect 22558 26288 22614 26344
rect 22926 51720 22982 51776
rect 23110 53352 23166 53408
rect 23018 48456 23074 48512
rect 23110 38664 23166 38720
rect 22834 36760 22890 36816
rect 22926 32172 22928 32192
rect 22928 32172 22980 32192
rect 22980 32172 22982 32192
rect 22926 32136 22982 32172
rect 22926 32000 22982 32056
rect 22834 31900 22836 31920
rect 22836 31900 22888 31920
rect 22888 31900 22890 31920
rect 22834 31864 22890 31900
rect 22926 31592 22982 31648
rect 22834 28328 22890 28384
rect 22742 26968 22798 27024
rect 22834 26324 22836 26344
rect 22836 26324 22888 26344
rect 22888 26324 22890 26344
rect 22834 26288 22890 26324
rect 22834 25744 22890 25800
rect 22926 25336 22982 25392
rect 22834 23568 22890 23624
rect 22834 23044 22890 23080
rect 22834 23024 22836 23044
rect 22836 23024 22888 23044
rect 22888 23024 22890 23044
rect 22926 22208 22982 22264
rect 22466 19896 22522 19952
rect 22742 19080 22798 19136
rect 22650 16360 22706 16416
rect 22466 13776 22522 13832
rect 22650 11192 22706 11248
rect 23110 33260 23112 33280
rect 23112 33260 23164 33280
rect 23164 33260 23166 33280
rect 23110 33224 23166 33260
rect 23110 31184 23166 31240
rect 23110 29300 23166 29336
rect 23110 29280 23112 29300
rect 23112 29280 23164 29300
rect 23164 29280 23166 29300
rect 23110 28756 23166 28792
rect 23110 28736 23112 28756
rect 23112 28736 23164 28756
rect 23164 28736 23166 28756
rect 23110 28092 23112 28112
rect 23112 28092 23164 28112
rect 23164 28092 23166 28112
rect 23110 28056 23166 28092
rect 23110 22516 23112 22536
rect 23112 22516 23164 22536
rect 23164 22516 23166 22536
rect 23110 22480 23166 22516
rect 24214 69944 24270 70000
rect 23386 61376 23442 61432
rect 23846 60288 23902 60344
rect 24306 68176 24362 68232
rect 23938 59336 23994 59392
rect 23386 58948 23442 58984
rect 23386 58928 23388 58948
rect 23388 58928 23440 58948
rect 23440 58928 23442 58948
rect 23294 51604 23350 51640
rect 23294 51584 23296 51604
rect 23296 51584 23348 51604
rect 23348 51584 23350 51604
rect 23662 56344 23718 56400
rect 23478 53896 23534 53952
rect 23754 53488 23810 53544
rect 23662 53352 23718 53408
rect 23938 52844 23940 52864
rect 23940 52844 23992 52864
rect 23992 52844 23994 52864
rect 23938 52808 23994 52844
rect 23662 48728 23718 48784
rect 23570 47096 23626 47152
rect 24490 58248 24546 58304
rect 24306 57860 24362 57896
rect 24306 57840 24308 57860
rect 24308 57840 24360 57860
rect 24360 57840 24362 57860
rect 24122 53488 24178 53544
rect 24398 56788 24400 56808
rect 24400 56788 24452 56808
rect 24452 56788 24454 56808
rect 24398 56752 24454 56788
rect 24490 56108 24492 56128
rect 24492 56108 24544 56128
rect 24544 56108 24546 56128
rect 24490 56072 24546 56108
rect 24490 54168 24546 54224
rect 24490 53896 24546 53952
rect 24214 50496 24270 50552
rect 24030 49000 24086 49056
rect 24214 48864 24270 48920
rect 23754 46960 23810 47016
rect 24214 47232 24270 47288
rect 23938 45600 23994 45656
rect 23570 44376 23626 44432
rect 24030 44276 24032 44296
rect 24032 44276 24084 44296
rect 24084 44276 24086 44296
rect 24030 44240 24086 44276
rect 23386 41384 23442 41440
rect 23754 41556 23756 41576
rect 23756 41556 23808 41576
rect 23808 41556 23810 41576
rect 23754 41520 23810 41556
rect 23846 41384 23902 41440
rect 23478 40976 23534 41032
rect 23754 37576 23810 37632
rect 23386 36236 23442 36272
rect 23386 36216 23388 36236
rect 23388 36216 23440 36236
rect 23440 36216 23442 36236
rect 23294 32020 23350 32056
rect 23294 32000 23296 32020
rect 23296 32000 23348 32020
rect 23348 32000 23350 32020
rect 23846 34892 23848 34912
rect 23848 34892 23900 34912
rect 23900 34892 23902 34912
rect 23846 34856 23902 34892
rect 23662 32852 23664 32872
rect 23664 32852 23716 32872
rect 23716 32852 23718 32872
rect 23662 32816 23718 32852
rect 23662 32136 23718 32192
rect 23570 31592 23626 31648
rect 23478 30232 23534 30288
rect 23386 27920 23442 27976
rect 23294 27512 23350 27568
rect 23294 27104 23350 27160
rect 23386 26288 23442 26344
rect 23294 25608 23350 25664
rect 23754 31456 23810 31512
rect 23938 32308 23940 32328
rect 23940 32308 23992 32328
rect 23992 32308 23994 32328
rect 23938 32272 23994 32308
rect 24214 32272 24270 32328
rect 24030 30232 24086 30288
rect 23938 29824 23994 29880
rect 23846 29688 23902 29744
rect 23662 29552 23718 29608
rect 23754 28736 23810 28792
rect 23938 28212 23994 28248
rect 23938 28192 23940 28212
rect 23940 28192 23992 28212
rect 23992 28192 23994 28212
rect 24122 28328 24178 28384
rect 23938 26288 23994 26344
rect 24214 26288 24270 26344
rect 23846 25200 23902 25256
rect 23754 24520 23810 24576
rect 23846 24384 23902 24440
rect 23754 24248 23810 24304
rect 23662 23840 23718 23896
rect 23662 23704 23718 23760
rect 23294 23024 23350 23080
rect 24030 22752 24086 22808
rect 23846 22616 23902 22672
rect 23386 21972 23388 21992
rect 23388 21972 23440 21992
rect 23440 21972 23442 21992
rect 23386 21936 23442 21972
rect 23846 19216 23902 19272
rect 24306 22344 24362 22400
rect 24122 17176 24178 17232
rect 23202 14184 23258 14240
rect 23110 13912 23166 13968
rect 23478 13368 23534 13424
rect 23478 7384 23534 7440
rect 23938 11056 23994 11112
rect 23846 7248 23902 7304
rect 23018 5072 23074 5128
rect 3422 720 3478 776
rect 23754 2372 23810 2408
rect 23754 2352 23756 2372
rect 23756 2352 23808 2372
rect 23808 2352 23810 2372
rect 24490 50224 24546 50280
rect 24490 48204 24546 48240
rect 24490 48184 24492 48204
rect 24492 48184 24544 48204
rect 24544 48184 24546 48204
rect 24490 46960 24546 47016
rect 24490 37304 24546 37360
rect 24490 26560 24546 26616
rect 24490 23044 24546 23080
rect 24490 23024 24492 23044
rect 24492 23024 24544 23044
rect 24544 23024 24546 23044
rect 24490 21836 24492 21856
rect 24492 21836 24544 21856
rect 24544 21836 24546 21856
rect 24490 21800 24546 21836
rect 24398 7656 24454 7712
rect 25686 73888 25742 73944
rect 25318 68176 25374 68232
rect 24950 61240 25006 61296
rect 25042 59336 25098 59392
rect 25318 60560 25374 60616
rect 24674 55664 24730 55720
rect 25042 52944 25098 53000
rect 24858 51856 24914 51912
rect 25502 56652 25504 56672
rect 25504 56652 25556 56672
rect 25556 56652 25558 56672
rect 25502 56616 25558 56652
rect 25318 56480 25374 56536
rect 25226 52128 25282 52184
rect 24858 51312 24914 51368
rect 24950 51176 25006 51232
rect 24674 50768 24730 50824
rect 24674 49680 24730 49736
rect 24674 48320 24730 48376
rect 24674 43968 24730 44024
rect 24674 43172 24730 43208
rect 24674 43152 24676 43172
rect 24676 43152 24728 43172
rect 24728 43152 24730 43172
rect 25410 52128 25466 52184
rect 25226 50088 25282 50144
rect 25502 51040 25558 51096
rect 25594 50904 25650 50960
rect 25226 48320 25282 48376
rect 24858 47776 24914 47832
rect 24858 41420 24860 41440
rect 24860 41420 24912 41440
rect 24912 41420 24914 41440
rect 24858 41384 24914 41420
rect 24766 40840 24822 40896
rect 24766 40704 24822 40760
rect 24674 34740 24730 34776
rect 24674 34720 24676 34740
rect 24676 34720 24728 34740
rect 24728 34720 24730 34740
rect 25318 47368 25374 47424
rect 25226 47232 25282 47288
rect 25042 34584 25098 34640
rect 25042 33360 25098 33416
rect 24858 32408 24914 32464
rect 25042 31320 25098 31376
rect 24858 31048 24914 31104
rect 24674 29996 24676 30016
rect 24676 29996 24728 30016
rect 24728 29996 24730 30016
rect 24674 29960 24730 29996
rect 24766 29824 24822 29880
rect 24950 30232 25006 30288
rect 24766 26732 24768 26752
rect 24768 26732 24820 26752
rect 24820 26732 24822 26752
rect 24766 26696 24822 26732
rect 24674 26560 24730 26616
rect 24858 25880 24914 25936
rect 25042 26968 25098 27024
rect 25042 26152 25098 26208
rect 24674 24812 24730 24848
rect 24674 24792 24676 24812
rect 24676 24792 24728 24812
rect 24728 24792 24730 24812
rect 25410 45772 25412 45792
rect 25412 45772 25464 45792
rect 25464 45772 25466 45792
rect 25410 45736 25466 45772
rect 25594 46960 25650 47016
rect 25502 44104 25558 44160
rect 25410 40024 25466 40080
rect 26146 69536 26202 69592
rect 25778 64096 25834 64152
rect 25778 54032 25834 54088
rect 25778 53080 25834 53136
rect 25778 52556 25834 52592
rect 25778 52536 25780 52556
rect 25780 52536 25832 52556
rect 25832 52536 25834 52556
rect 25778 49952 25834 50008
rect 25778 46316 25780 46336
rect 25780 46316 25832 46336
rect 25832 46316 25834 46336
rect 25778 46280 25834 46316
rect 25778 38836 25780 38856
rect 25780 38836 25832 38856
rect 25832 38836 25834 38856
rect 25778 38800 25834 38836
rect 25686 36660 25688 36680
rect 25688 36660 25740 36680
rect 25740 36660 25742 36680
rect 25686 36624 25742 36660
rect 26054 56364 26110 56400
rect 26054 56344 26056 56364
rect 26056 56344 26108 56364
rect 26108 56344 26110 56364
rect 25962 48728 26018 48784
rect 25962 44684 25964 44704
rect 25964 44684 26016 44704
rect 26016 44684 26018 44704
rect 25962 44648 26018 44684
rect 25962 44240 26018 44296
rect 26330 65456 26386 65512
rect 26238 60596 26240 60616
rect 26240 60596 26292 60616
rect 26292 60596 26294 60616
rect 26238 60560 26294 60596
rect 26514 55800 26570 55856
rect 27434 72800 27490 72856
rect 27250 67224 27306 67280
rect 27158 63960 27214 64016
rect 27066 60288 27122 60344
rect 26330 55256 26386 55312
rect 26238 54576 26294 54632
rect 26422 47912 26478 47968
rect 26238 45872 26294 45928
rect 26790 54848 26846 54904
rect 26698 53216 26754 53272
rect 26882 50668 26884 50688
rect 26884 50668 26936 50688
rect 26936 50668 26938 50688
rect 26882 50632 26938 50668
rect 26790 49952 26846 50008
rect 26606 47776 26662 47832
rect 27986 74432 28042 74488
rect 27526 68992 27582 69048
rect 27710 58384 27766 58440
rect 28814 76064 28870 76120
rect 28814 72972 28816 72992
rect 28816 72972 28868 72992
rect 28868 72972 28870 72992
rect 28814 72936 28870 72972
rect 29826 75520 29882 75576
rect 28078 57568 28134 57624
rect 27986 55392 28042 55448
rect 27894 54984 27950 55040
rect 27618 53488 27674 53544
rect 27158 49000 27214 49056
rect 27618 49680 27674 49736
rect 29090 62056 29146 62112
rect 28446 51176 28502 51232
rect 27894 49816 27950 49872
rect 27342 48048 27398 48104
rect 27158 47116 27214 47152
rect 27158 47096 27160 47116
rect 27160 47096 27212 47116
rect 27212 47096 27214 47116
rect 28078 50360 28134 50416
rect 27986 49272 28042 49328
rect 27986 48492 27988 48512
rect 27988 48492 28040 48512
rect 28040 48492 28042 48512
rect 27986 48456 28042 48492
rect 27250 46824 27306 46880
rect 26882 46280 26938 46336
rect 26422 44276 26424 44296
rect 26424 44276 26476 44296
rect 26476 44276 26478 44296
rect 26422 44240 26478 44276
rect 26330 43988 26386 44024
rect 26330 43968 26332 43988
rect 26332 43968 26384 43988
rect 26384 43968 26386 43988
rect 27526 46960 27582 47016
rect 27434 46008 27490 46064
rect 27526 45872 27582 45928
rect 26606 43696 26662 43752
rect 27158 43288 27214 43344
rect 26146 38664 26202 38720
rect 25870 34720 25926 34776
rect 25318 33904 25374 33960
rect 25594 33652 25650 33688
rect 25594 33632 25596 33652
rect 25596 33632 25648 33652
rect 25648 33632 25650 33652
rect 25318 31048 25374 31104
rect 25594 32952 25650 33008
rect 25594 31900 25596 31920
rect 25596 31900 25648 31920
rect 25648 31900 25650 31920
rect 25594 31864 25650 31900
rect 25410 30640 25466 30696
rect 25686 30096 25742 30152
rect 25410 26968 25466 27024
rect 25502 26424 25558 26480
rect 25318 26036 25374 26072
rect 25318 26016 25320 26036
rect 25320 26016 25372 26036
rect 25372 26016 25374 26036
rect 25318 25492 25374 25528
rect 25318 25472 25320 25492
rect 25320 25472 25372 25492
rect 25372 25472 25374 25492
rect 25870 30116 25926 30152
rect 25870 30096 25872 30116
rect 25872 30096 25924 30116
rect 25924 30096 25926 30116
rect 25778 26832 25834 26888
rect 25778 26560 25834 26616
rect 25870 25780 25872 25800
rect 25872 25780 25924 25800
rect 25924 25780 25926 25800
rect 25870 25744 25926 25780
rect 25226 24656 25282 24712
rect 24674 23180 24730 23216
rect 24674 23160 24676 23180
rect 24676 23160 24728 23180
rect 24728 23160 24730 23180
rect 24950 18536 25006 18592
rect 24858 15408 24914 15464
rect 24674 7792 24730 7848
rect 25410 24012 25412 24032
rect 25412 24012 25464 24032
rect 25464 24012 25466 24032
rect 25410 23976 25466 24012
rect 25134 13912 25190 13968
rect 25778 7656 25834 7712
rect 25042 7520 25098 7576
rect 24950 6840 25006 6896
rect 26054 33632 26110 33688
rect 26974 38800 27030 38856
rect 26790 37440 26846 37496
rect 26330 32000 26386 32056
rect 26422 31728 26478 31784
rect 26054 27376 26110 27432
rect 26238 30232 26294 30288
rect 26238 29824 26294 29880
rect 26514 31320 26570 31376
rect 26422 29688 26478 29744
rect 26606 30776 26662 30832
rect 26514 29008 26570 29064
rect 26238 24792 26294 24848
rect 26146 24112 26202 24168
rect 26422 28464 26478 28520
rect 26422 23704 26478 23760
rect 26422 23296 26478 23352
rect 26330 14456 26386 14512
rect 26790 32272 26846 32328
rect 26790 28328 26846 28384
rect 26790 26288 26846 26344
rect 26606 22616 26662 22672
rect 27802 45328 27858 45384
rect 28170 48184 28226 48240
rect 28078 45872 28134 45928
rect 27250 41384 27306 41440
rect 27526 41656 27582 41712
rect 27710 41384 27766 41440
rect 27434 36352 27490 36408
rect 27066 35808 27122 35864
rect 26974 32272 27030 32328
rect 26974 29452 26976 29472
rect 26976 29452 27028 29472
rect 27028 29452 27030 29472
rect 26974 29416 27030 29452
rect 27618 34176 27674 34232
rect 27434 33768 27490 33824
rect 27158 31592 27214 31648
rect 27250 31320 27306 31376
rect 27526 31592 27582 31648
rect 27250 29960 27306 30016
rect 27894 44512 27950 44568
rect 29274 61104 29330 61160
rect 28998 57588 29054 57624
rect 28998 57568 29000 57588
rect 29000 57568 29052 57588
rect 29052 57568 29054 57588
rect 28906 54032 28962 54088
rect 28998 53352 29054 53408
rect 29182 52672 29238 52728
rect 28538 50360 28594 50416
rect 28354 47640 28410 47696
rect 28354 46960 28410 47016
rect 28998 50668 29000 50688
rect 29000 50668 29052 50688
rect 29052 50668 29054 50688
rect 28998 50632 29054 50668
rect 29274 51176 29330 51232
rect 28814 49544 28870 49600
rect 28354 46028 28410 46064
rect 28354 46008 28356 46028
rect 28356 46008 28408 46028
rect 28408 46008 28410 46028
rect 28078 42356 28134 42392
rect 28078 42336 28080 42356
rect 28080 42336 28132 42356
rect 28132 42336 28134 42356
rect 27802 27376 27858 27432
rect 27802 27276 27804 27296
rect 27804 27276 27856 27296
rect 27856 27276 27858 27296
rect 27802 27240 27858 27276
rect 27618 26324 27620 26344
rect 27620 26324 27672 26344
rect 27672 26324 27674 26344
rect 27618 26288 27674 26324
rect 27434 23024 27490 23080
rect 27158 21392 27214 21448
rect 27066 17856 27122 17912
rect 26882 10512 26938 10568
rect 26514 7792 26570 7848
rect 26698 7520 26754 7576
rect 26146 6840 26202 6896
rect 25962 6296 26018 6352
rect 26146 5616 26202 5672
rect 28078 38412 28134 38448
rect 28078 38392 28080 38412
rect 28080 38392 28132 38412
rect 28132 38392 28134 38412
rect 28078 36760 28134 36816
rect 28262 41792 28318 41848
rect 28354 41112 28410 41168
rect 28538 44940 28594 44976
rect 28538 44920 28540 44940
rect 28540 44920 28592 44940
rect 28592 44920 28594 44940
rect 28630 44820 28632 44840
rect 28632 44820 28684 44840
rect 28684 44820 28686 44840
rect 28630 44784 28686 44820
rect 28814 48184 28870 48240
rect 29090 49408 29146 49464
rect 28998 48864 29054 48920
rect 29090 47796 29146 47832
rect 29090 47776 29092 47796
rect 29092 47776 29144 47796
rect 29144 47776 29146 47796
rect 31758 74976 31814 75032
rect 29918 71576 29974 71632
rect 30378 70080 30434 70136
rect 29918 60560 29974 60616
rect 29550 60308 29606 60344
rect 29550 60288 29552 60308
rect 29552 60288 29604 60308
rect 29604 60288 29606 60308
rect 29826 59336 29882 59392
rect 29734 56344 29790 56400
rect 29458 52556 29514 52592
rect 29642 52808 29698 52864
rect 29458 52536 29460 52556
rect 29460 52536 29512 52556
rect 29512 52536 29514 52556
rect 29550 52400 29606 52456
rect 30378 60016 30434 60072
rect 31022 74160 31078 74216
rect 31206 62600 31262 62656
rect 31022 62056 31078 62112
rect 30654 56480 30710 56536
rect 30562 52012 30618 52048
rect 30562 51992 30564 52012
rect 30564 51992 30616 52012
rect 30616 51992 30618 52012
rect 30102 51040 30158 51096
rect 29734 49680 29790 49736
rect 29918 49000 29974 49056
rect 29642 48184 29698 48240
rect 29918 48204 29974 48240
rect 29918 48184 29920 48204
rect 29920 48184 29972 48204
rect 29972 48184 29974 48204
rect 29458 47912 29514 47968
rect 28722 43968 28778 44024
rect 28262 40024 28318 40080
rect 28078 32000 28134 32056
rect 28078 30116 28134 30152
rect 28078 30096 28080 30116
rect 28080 30096 28132 30116
rect 28132 30096 28134 30116
rect 28170 29552 28226 29608
rect 28078 28600 28134 28656
rect 28170 28056 28226 28112
rect 28538 35808 28594 35864
rect 28354 27124 28410 27160
rect 28354 27104 28356 27124
rect 28356 27104 28408 27124
rect 28408 27104 28410 27124
rect 28078 26868 28080 26888
rect 28080 26868 28132 26888
rect 28132 26868 28134 26888
rect 28078 26832 28134 26868
rect 28538 30776 28594 30832
rect 28446 26580 28502 26616
rect 28446 26560 28448 26580
rect 28448 26560 28500 26580
rect 28500 26560 28502 26580
rect 28538 26424 28594 26480
rect 28722 42644 28724 42664
rect 28724 42644 28776 42664
rect 28776 42644 28778 42664
rect 28722 42608 28778 42644
rect 28722 40160 28778 40216
rect 28998 46960 29054 47016
rect 28906 46316 28908 46336
rect 28908 46316 28960 46336
rect 28960 46316 28962 46336
rect 28906 46280 28962 46316
rect 29182 46552 29238 46608
rect 29274 46280 29330 46336
rect 29090 45600 29146 45656
rect 29090 44648 29146 44704
rect 29734 48048 29790 48104
rect 28814 37168 28870 37224
rect 28722 31456 28778 31512
rect 28906 32972 28962 33008
rect 28906 32952 28908 32972
rect 28908 32952 28960 32972
rect 28960 32952 28962 32972
rect 28906 31728 28962 31784
rect 28998 30232 29054 30288
rect 28998 28756 29054 28792
rect 28998 28736 29000 28756
rect 29000 28736 29052 28756
rect 29052 28736 29054 28756
rect 28906 28056 28962 28112
rect 28998 27376 29054 27432
rect 28814 26832 28870 26888
rect 29734 44648 29790 44704
rect 29642 44104 29698 44160
rect 29458 42880 29514 42936
rect 29458 42764 29514 42800
rect 29458 42744 29460 42764
rect 29460 42744 29512 42764
rect 29512 42744 29514 42764
rect 30378 50768 30434 50824
rect 30654 50224 30710 50280
rect 30562 50088 30618 50144
rect 29550 41384 29606 41440
rect 29826 41248 29882 41304
rect 29458 37304 29514 37360
rect 29550 36372 29606 36408
rect 29550 36352 29552 36372
rect 29552 36352 29604 36372
rect 29604 36352 29606 36372
rect 29274 28600 29330 28656
rect 29090 23296 29146 23352
rect 29458 28056 29514 28112
rect 29458 27648 29514 27704
rect 29734 40840 29790 40896
rect 29734 27920 29790 27976
rect 29642 27376 29698 27432
rect 29182 22616 29238 22672
rect 28998 22480 29054 22536
rect 30194 49272 30250 49328
rect 31022 50360 31078 50416
rect 31206 49952 31262 50008
rect 30930 49816 30986 49872
rect 30838 49544 30894 49600
rect 28998 17176 29054 17232
rect 28630 15816 28686 15872
rect 27986 6160 28042 6216
rect 29642 15136 29698 15192
rect 28446 2644 28502 2680
rect 28446 2624 28448 2644
rect 28448 2624 28500 2644
rect 28500 2624 28502 2644
rect 30102 18572 30104 18592
rect 30104 18572 30156 18592
rect 30156 18572 30158 18592
rect 30102 18536 30158 18572
rect 30654 48320 30710 48376
rect 30746 48048 30802 48104
rect 30654 47404 30656 47424
rect 30656 47404 30708 47424
rect 30708 47404 30710 47424
rect 30654 47368 30710 47404
rect 31022 49136 31078 49192
rect 31206 48728 31262 48784
rect 30562 46552 30618 46608
rect 30930 47232 30986 47288
rect 31114 47096 31170 47152
rect 31114 46008 31170 46064
rect 31206 44920 31262 44976
rect 31114 44784 31170 44840
rect 30746 44276 30748 44296
rect 30748 44276 30800 44296
rect 30800 44276 30802 44296
rect 30746 44240 30802 44276
rect 30838 42336 30894 42392
rect 30470 37984 30526 38040
rect 30654 33632 30710 33688
rect 30562 31764 30564 31784
rect 30564 31764 30616 31784
rect 30616 31764 30618 31784
rect 30562 31728 30618 31764
rect 30470 26832 30526 26888
rect 30286 15000 30342 15056
rect 31390 60288 31446 60344
rect 32954 58928 33010 58984
rect 31758 56480 31814 56536
rect 31574 55276 31630 55312
rect 31574 55256 31576 55276
rect 31576 55256 31628 55276
rect 31628 55256 31630 55276
rect 32586 54032 32642 54088
rect 31942 53896 31998 53952
rect 31758 52400 31814 52456
rect 31482 50632 31538 50688
rect 32218 50224 32274 50280
rect 31390 49272 31446 49328
rect 32402 47676 32404 47696
rect 32404 47676 32456 47696
rect 32456 47676 32458 47696
rect 32402 47640 32458 47676
rect 32034 47096 32090 47152
rect 31850 44684 31852 44704
rect 31852 44684 31904 44704
rect 31904 44684 31906 44704
rect 31850 44648 31906 44684
rect 31574 44512 31630 44568
rect 31390 42744 31446 42800
rect 31298 37304 31354 37360
rect 32126 46280 32182 46336
rect 32218 46144 32274 46200
rect 32402 45872 32458 45928
rect 31482 20576 31538 20632
rect 31114 20304 31170 20360
rect 30010 11056 30066 11112
rect 30286 9696 30342 9752
rect 31298 2216 31354 2272
rect 29642 1944 29698 2000
rect 30378 856 30434 912
rect 32402 34060 32458 34096
rect 32402 34040 32404 34060
rect 32404 34040 32456 34060
rect 32456 34040 32458 34060
rect 32678 46960 32734 47016
rect 32586 36760 32642 36816
rect 33322 52808 33378 52864
rect 33138 47096 33194 47152
rect 33046 46144 33102 46200
rect 32954 44920 33010 44976
rect 35346 78240 35402 78296
rect 34940 77274 34996 77276
rect 35020 77274 35076 77276
rect 35100 77274 35156 77276
rect 35180 77274 35236 77276
rect 34940 77222 34966 77274
rect 34966 77222 34996 77274
rect 35020 77222 35030 77274
rect 35030 77222 35076 77274
rect 35100 77222 35146 77274
rect 35146 77222 35156 77274
rect 35180 77222 35210 77274
rect 35210 77222 35236 77274
rect 34940 77220 34996 77222
rect 35020 77220 35076 77222
rect 35100 77220 35156 77222
rect 35180 77220 35236 77222
rect 34940 76186 34996 76188
rect 35020 76186 35076 76188
rect 35100 76186 35156 76188
rect 35180 76186 35236 76188
rect 34940 76134 34966 76186
rect 34966 76134 34996 76186
rect 35020 76134 35030 76186
rect 35030 76134 35076 76186
rect 35100 76134 35146 76186
rect 35146 76134 35156 76186
rect 35180 76134 35210 76186
rect 35210 76134 35236 76186
rect 34940 76132 34996 76134
rect 35020 76132 35076 76134
rect 35100 76132 35156 76134
rect 35180 76132 35236 76134
rect 34794 75520 34850 75576
rect 34940 75098 34996 75100
rect 35020 75098 35076 75100
rect 35100 75098 35156 75100
rect 35180 75098 35236 75100
rect 34940 75046 34966 75098
rect 34966 75046 34996 75098
rect 35020 75046 35030 75098
rect 35030 75046 35076 75098
rect 35100 75046 35146 75098
rect 35146 75046 35156 75098
rect 35180 75046 35210 75098
rect 35210 75046 35236 75098
rect 34940 75044 34996 75046
rect 35020 75044 35076 75046
rect 35100 75044 35156 75046
rect 35180 75044 35236 75046
rect 35806 76880 35862 76936
rect 35622 75520 35678 75576
rect 34940 74010 34996 74012
rect 35020 74010 35076 74012
rect 35100 74010 35156 74012
rect 35180 74010 35236 74012
rect 34940 73958 34966 74010
rect 34966 73958 34996 74010
rect 35020 73958 35030 74010
rect 35030 73958 35076 74010
rect 35100 73958 35146 74010
rect 35146 73958 35156 74010
rect 35180 73958 35210 74010
rect 35210 73958 35236 74010
rect 34940 73956 34996 73958
rect 35020 73956 35076 73958
rect 35100 73956 35156 73958
rect 35180 73956 35236 73958
rect 34940 72922 34996 72924
rect 35020 72922 35076 72924
rect 35100 72922 35156 72924
rect 35180 72922 35236 72924
rect 34940 72870 34966 72922
rect 34966 72870 34996 72922
rect 35020 72870 35030 72922
rect 35030 72870 35076 72922
rect 35100 72870 35146 72922
rect 35146 72870 35156 72922
rect 35180 72870 35210 72922
rect 35210 72870 35236 72922
rect 34940 72868 34996 72870
rect 35020 72868 35076 72870
rect 35100 72868 35156 72870
rect 35180 72868 35236 72870
rect 34940 71834 34996 71836
rect 35020 71834 35076 71836
rect 35100 71834 35156 71836
rect 35180 71834 35236 71836
rect 34940 71782 34966 71834
rect 34966 71782 34996 71834
rect 35020 71782 35030 71834
rect 35030 71782 35076 71834
rect 35100 71782 35146 71834
rect 35146 71782 35156 71834
rect 35180 71782 35210 71834
rect 35210 71782 35236 71834
rect 34940 71780 34996 71782
rect 35020 71780 35076 71782
rect 35100 71780 35156 71782
rect 35180 71780 35236 71782
rect 34518 71440 34574 71496
rect 34940 70746 34996 70748
rect 35020 70746 35076 70748
rect 35100 70746 35156 70748
rect 35180 70746 35236 70748
rect 34940 70694 34966 70746
rect 34966 70694 34996 70746
rect 35020 70694 35030 70746
rect 35030 70694 35076 70746
rect 35100 70694 35146 70746
rect 35146 70694 35156 70746
rect 35180 70694 35210 70746
rect 35210 70694 35236 70746
rect 34940 70692 34996 70694
rect 35020 70692 35076 70694
rect 35100 70692 35156 70694
rect 35180 70692 35236 70694
rect 34518 69944 34574 70000
rect 34940 69658 34996 69660
rect 35020 69658 35076 69660
rect 35100 69658 35156 69660
rect 35180 69658 35236 69660
rect 34940 69606 34966 69658
rect 34966 69606 34996 69658
rect 35020 69606 35030 69658
rect 35030 69606 35076 69658
rect 35100 69606 35146 69658
rect 35146 69606 35156 69658
rect 35180 69606 35210 69658
rect 35210 69606 35236 69658
rect 34940 69604 34996 69606
rect 35020 69604 35076 69606
rect 35100 69604 35156 69606
rect 35180 69604 35236 69606
rect 34940 68570 34996 68572
rect 35020 68570 35076 68572
rect 35100 68570 35156 68572
rect 35180 68570 35236 68572
rect 34940 68518 34966 68570
rect 34966 68518 34996 68570
rect 35020 68518 35030 68570
rect 35030 68518 35076 68570
rect 35100 68518 35146 68570
rect 35146 68518 35156 68570
rect 35180 68518 35210 68570
rect 35210 68518 35236 68570
rect 34940 68516 34996 68518
rect 35020 68516 35076 68518
rect 35100 68516 35156 68518
rect 35180 68516 35236 68518
rect 34940 67482 34996 67484
rect 35020 67482 35076 67484
rect 35100 67482 35156 67484
rect 35180 67482 35236 67484
rect 34940 67430 34966 67482
rect 34966 67430 34996 67482
rect 35020 67430 35030 67482
rect 35030 67430 35076 67482
rect 35100 67430 35146 67482
rect 35146 67430 35156 67482
rect 35180 67430 35210 67482
rect 35210 67430 35236 67482
rect 34940 67428 34996 67430
rect 35020 67428 35076 67430
rect 35100 67428 35156 67430
rect 35180 67428 35236 67430
rect 34940 66394 34996 66396
rect 35020 66394 35076 66396
rect 35100 66394 35156 66396
rect 35180 66394 35236 66396
rect 34940 66342 34966 66394
rect 34966 66342 34996 66394
rect 35020 66342 35030 66394
rect 35030 66342 35076 66394
rect 35100 66342 35146 66394
rect 35146 66342 35156 66394
rect 35180 66342 35210 66394
rect 35210 66342 35236 66394
rect 34940 66340 34996 66342
rect 35020 66340 35076 66342
rect 35100 66340 35156 66342
rect 35180 66340 35236 66342
rect 34940 65306 34996 65308
rect 35020 65306 35076 65308
rect 35100 65306 35156 65308
rect 35180 65306 35236 65308
rect 34940 65254 34966 65306
rect 34966 65254 34996 65306
rect 35020 65254 35030 65306
rect 35030 65254 35076 65306
rect 35100 65254 35146 65306
rect 35146 65254 35156 65306
rect 35180 65254 35210 65306
rect 35210 65254 35236 65306
rect 34940 65252 34996 65254
rect 35020 65252 35076 65254
rect 35100 65252 35156 65254
rect 35180 65252 35236 65254
rect 34940 64218 34996 64220
rect 35020 64218 35076 64220
rect 35100 64218 35156 64220
rect 35180 64218 35236 64220
rect 34940 64166 34966 64218
rect 34966 64166 34996 64218
rect 35020 64166 35030 64218
rect 35030 64166 35076 64218
rect 35100 64166 35146 64218
rect 35146 64166 35156 64218
rect 35180 64166 35210 64218
rect 35210 64166 35236 64218
rect 34940 64164 34996 64166
rect 35020 64164 35076 64166
rect 35100 64164 35156 64166
rect 35180 64164 35236 64166
rect 34940 63130 34996 63132
rect 35020 63130 35076 63132
rect 35100 63130 35156 63132
rect 35180 63130 35236 63132
rect 34940 63078 34966 63130
rect 34966 63078 34996 63130
rect 35020 63078 35030 63130
rect 35030 63078 35076 63130
rect 35100 63078 35146 63130
rect 35146 63078 35156 63130
rect 35180 63078 35210 63130
rect 35210 63078 35236 63130
rect 34940 63076 34996 63078
rect 35020 63076 35076 63078
rect 35100 63076 35156 63078
rect 35180 63076 35236 63078
rect 34940 62042 34996 62044
rect 35020 62042 35076 62044
rect 35100 62042 35156 62044
rect 35180 62042 35236 62044
rect 34940 61990 34966 62042
rect 34966 61990 34996 62042
rect 35020 61990 35030 62042
rect 35030 61990 35076 62042
rect 35100 61990 35146 62042
rect 35146 61990 35156 62042
rect 35180 61990 35210 62042
rect 35210 61990 35236 62042
rect 34940 61988 34996 61990
rect 35020 61988 35076 61990
rect 35100 61988 35156 61990
rect 35180 61988 35236 61990
rect 34940 60954 34996 60956
rect 35020 60954 35076 60956
rect 35100 60954 35156 60956
rect 35180 60954 35236 60956
rect 34940 60902 34966 60954
rect 34966 60902 34996 60954
rect 35020 60902 35030 60954
rect 35030 60902 35076 60954
rect 35100 60902 35146 60954
rect 35146 60902 35156 60954
rect 35180 60902 35210 60954
rect 35210 60902 35236 60954
rect 34940 60900 34996 60902
rect 35020 60900 35076 60902
rect 35100 60900 35156 60902
rect 35180 60900 35236 60902
rect 35438 72800 35494 72856
rect 35438 70896 35494 70952
rect 35530 68720 35586 68776
rect 35438 65320 35494 65376
rect 35530 62736 35586 62792
rect 35438 62192 35494 62248
rect 35622 61376 35678 61432
rect 35438 61240 35494 61296
rect 34518 57160 34574 57216
rect 34940 59866 34996 59868
rect 35020 59866 35076 59868
rect 35100 59866 35156 59868
rect 35180 59866 35236 59868
rect 34940 59814 34966 59866
rect 34966 59814 34996 59866
rect 35020 59814 35030 59866
rect 35030 59814 35076 59866
rect 35100 59814 35146 59866
rect 35146 59814 35156 59866
rect 35180 59814 35210 59866
rect 35210 59814 35236 59866
rect 34940 59812 34996 59814
rect 35020 59812 35076 59814
rect 35100 59812 35156 59814
rect 35180 59812 35236 59814
rect 36818 73208 36874 73264
rect 35898 71576 35954 71632
rect 37370 68176 37426 68232
rect 35806 61104 35862 61160
rect 39578 73752 39634 73808
rect 37370 59336 37426 59392
rect 34940 58778 34996 58780
rect 35020 58778 35076 58780
rect 35100 58778 35156 58780
rect 35180 58778 35236 58780
rect 34940 58726 34966 58778
rect 34966 58726 34996 58778
rect 35020 58726 35030 58778
rect 35030 58726 35076 58778
rect 35100 58726 35146 58778
rect 35146 58726 35156 58778
rect 35180 58726 35210 58778
rect 35210 58726 35236 58778
rect 34940 58724 34996 58726
rect 35020 58724 35076 58726
rect 35100 58724 35156 58726
rect 35180 58724 35236 58726
rect 35346 58520 35402 58576
rect 34940 57690 34996 57692
rect 35020 57690 35076 57692
rect 35100 57690 35156 57692
rect 35180 57690 35236 57692
rect 34940 57638 34966 57690
rect 34966 57638 34996 57690
rect 35020 57638 35030 57690
rect 35030 57638 35076 57690
rect 35100 57638 35146 57690
rect 35146 57638 35156 57690
rect 35180 57638 35210 57690
rect 35210 57638 35236 57690
rect 34940 57636 34996 57638
rect 35020 57636 35076 57638
rect 35100 57636 35156 57638
rect 35180 57636 35236 57638
rect 34940 56602 34996 56604
rect 35020 56602 35076 56604
rect 35100 56602 35156 56604
rect 35180 56602 35236 56604
rect 34940 56550 34966 56602
rect 34966 56550 34996 56602
rect 35020 56550 35030 56602
rect 35030 56550 35076 56602
rect 35100 56550 35146 56602
rect 35146 56550 35156 56602
rect 35180 56550 35210 56602
rect 35210 56550 35236 56602
rect 34940 56548 34996 56550
rect 35020 56548 35076 56550
rect 35100 56548 35156 56550
rect 35180 56548 35236 56550
rect 34940 55514 34996 55516
rect 35020 55514 35076 55516
rect 35100 55514 35156 55516
rect 35180 55514 35236 55516
rect 34940 55462 34966 55514
rect 34966 55462 34996 55514
rect 35020 55462 35030 55514
rect 35030 55462 35076 55514
rect 35100 55462 35146 55514
rect 35146 55462 35156 55514
rect 35180 55462 35210 55514
rect 35210 55462 35236 55514
rect 34940 55460 34996 55462
rect 35020 55460 35076 55462
rect 35100 55460 35156 55462
rect 35180 55460 35236 55462
rect 34940 54426 34996 54428
rect 35020 54426 35076 54428
rect 35100 54426 35156 54428
rect 35180 54426 35236 54428
rect 34940 54374 34966 54426
rect 34966 54374 34996 54426
rect 35020 54374 35030 54426
rect 35030 54374 35076 54426
rect 35100 54374 35146 54426
rect 35146 54374 35156 54426
rect 35180 54374 35210 54426
rect 35210 54374 35236 54426
rect 34940 54372 34996 54374
rect 35020 54372 35076 54374
rect 35100 54372 35156 54374
rect 35180 54372 35236 54374
rect 35254 53896 35310 53952
rect 34940 53338 34996 53340
rect 35020 53338 35076 53340
rect 35100 53338 35156 53340
rect 35180 53338 35236 53340
rect 34940 53286 34966 53338
rect 34966 53286 34996 53338
rect 35020 53286 35030 53338
rect 35030 53286 35076 53338
rect 35100 53286 35146 53338
rect 35146 53286 35156 53338
rect 35180 53286 35210 53338
rect 35210 53286 35236 53338
rect 34940 53284 34996 53286
rect 35020 53284 35076 53286
rect 35100 53284 35156 53286
rect 35180 53284 35236 53286
rect 34702 52536 34758 52592
rect 34610 52400 34666 52456
rect 33690 50632 33746 50688
rect 34610 46960 34666 47016
rect 34518 42880 34574 42936
rect 33046 36624 33102 36680
rect 32678 32952 32734 33008
rect 32770 28056 32826 28112
rect 33506 26288 33562 26344
rect 34518 40840 34574 40896
rect 34940 52250 34996 52252
rect 35020 52250 35076 52252
rect 35100 52250 35156 52252
rect 35180 52250 35236 52252
rect 34940 52198 34966 52250
rect 34966 52198 34996 52250
rect 35020 52198 35030 52250
rect 35030 52198 35076 52250
rect 35100 52198 35146 52250
rect 35146 52198 35156 52250
rect 35180 52198 35210 52250
rect 35210 52198 35236 52250
rect 34940 52196 34996 52198
rect 35020 52196 35076 52198
rect 35100 52196 35156 52198
rect 35180 52196 35236 52198
rect 34940 51162 34996 51164
rect 35020 51162 35076 51164
rect 35100 51162 35156 51164
rect 35180 51162 35236 51164
rect 34940 51110 34966 51162
rect 34966 51110 34996 51162
rect 35020 51110 35030 51162
rect 35030 51110 35076 51162
rect 35100 51110 35146 51162
rect 35146 51110 35156 51162
rect 35180 51110 35210 51162
rect 35210 51110 35236 51162
rect 34940 51108 34996 51110
rect 35020 51108 35076 51110
rect 35100 51108 35156 51110
rect 35180 51108 35236 51110
rect 34940 50074 34996 50076
rect 35020 50074 35076 50076
rect 35100 50074 35156 50076
rect 35180 50074 35236 50076
rect 34940 50022 34966 50074
rect 34966 50022 34996 50074
rect 35020 50022 35030 50074
rect 35030 50022 35076 50074
rect 35100 50022 35146 50074
rect 35146 50022 35156 50074
rect 35180 50022 35210 50074
rect 35210 50022 35236 50074
rect 34940 50020 34996 50022
rect 35020 50020 35076 50022
rect 35100 50020 35156 50022
rect 35180 50020 35236 50022
rect 34940 48986 34996 48988
rect 35020 48986 35076 48988
rect 35100 48986 35156 48988
rect 35180 48986 35236 48988
rect 34940 48934 34966 48986
rect 34966 48934 34996 48986
rect 35020 48934 35030 48986
rect 35030 48934 35076 48986
rect 35100 48934 35146 48986
rect 35146 48934 35156 48986
rect 35180 48934 35210 48986
rect 35210 48934 35236 48986
rect 34940 48932 34996 48934
rect 35020 48932 35076 48934
rect 35100 48932 35156 48934
rect 35180 48932 35236 48934
rect 34940 47898 34996 47900
rect 35020 47898 35076 47900
rect 35100 47898 35156 47900
rect 35180 47898 35236 47900
rect 34940 47846 34966 47898
rect 34966 47846 34996 47898
rect 35020 47846 35030 47898
rect 35030 47846 35076 47898
rect 35100 47846 35146 47898
rect 35146 47846 35156 47898
rect 35180 47846 35210 47898
rect 35210 47846 35236 47898
rect 34940 47844 34996 47846
rect 35020 47844 35076 47846
rect 35100 47844 35156 47846
rect 35180 47844 35236 47846
rect 34940 46810 34996 46812
rect 35020 46810 35076 46812
rect 35100 46810 35156 46812
rect 35180 46810 35236 46812
rect 34940 46758 34966 46810
rect 34966 46758 34996 46810
rect 35020 46758 35030 46810
rect 35030 46758 35076 46810
rect 35100 46758 35146 46810
rect 35146 46758 35156 46810
rect 35180 46758 35210 46810
rect 35210 46758 35236 46810
rect 34940 46756 34996 46758
rect 35020 46756 35076 46758
rect 35100 46756 35156 46758
rect 35180 46756 35236 46758
rect 34794 46144 34850 46200
rect 34940 45722 34996 45724
rect 35020 45722 35076 45724
rect 35100 45722 35156 45724
rect 35180 45722 35236 45724
rect 34940 45670 34966 45722
rect 34966 45670 34996 45722
rect 35020 45670 35030 45722
rect 35030 45670 35076 45722
rect 35100 45670 35146 45722
rect 35146 45670 35156 45722
rect 35180 45670 35210 45722
rect 35210 45670 35236 45722
rect 34940 45668 34996 45670
rect 35020 45668 35076 45670
rect 35100 45668 35156 45670
rect 35180 45668 35236 45670
rect 34940 44634 34996 44636
rect 35020 44634 35076 44636
rect 35100 44634 35156 44636
rect 35180 44634 35236 44636
rect 34940 44582 34966 44634
rect 34966 44582 34996 44634
rect 35020 44582 35030 44634
rect 35030 44582 35076 44634
rect 35100 44582 35146 44634
rect 35146 44582 35156 44634
rect 35180 44582 35210 44634
rect 35210 44582 35236 44634
rect 34940 44580 34996 44582
rect 35020 44580 35076 44582
rect 35100 44580 35156 44582
rect 35180 44580 35236 44582
rect 34940 43546 34996 43548
rect 35020 43546 35076 43548
rect 35100 43546 35156 43548
rect 35180 43546 35236 43548
rect 34940 43494 34966 43546
rect 34966 43494 34996 43546
rect 35020 43494 35030 43546
rect 35030 43494 35076 43546
rect 35100 43494 35146 43546
rect 35146 43494 35156 43546
rect 35180 43494 35210 43546
rect 35210 43494 35236 43546
rect 34940 43492 34996 43494
rect 35020 43492 35076 43494
rect 35100 43492 35156 43494
rect 35180 43492 35236 43494
rect 35162 42744 35218 42800
rect 34794 42608 34850 42664
rect 34940 42458 34996 42460
rect 35020 42458 35076 42460
rect 35100 42458 35156 42460
rect 35180 42458 35236 42460
rect 34940 42406 34966 42458
rect 34966 42406 34996 42458
rect 35020 42406 35030 42458
rect 35030 42406 35076 42458
rect 35100 42406 35146 42458
rect 35146 42406 35156 42458
rect 35180 42406 35210 42458
rect 35210 42406 35236 42458
rect 34940 42404 34996 42406
rect 35020 42404 35076 42406
rect 35100 42404 35156 42406
rect 35180 42404 35236 42406
rect 34940 41370 34996 41372
rect 35020 41370 35076 41372
rect 35100 41370 35156 41372
rect 35180 41370 35236 41372
rect 34940 41318 34966 41370
rect 34966 41318 34996 41370
rect 35020 41318 35030 41370
rect 35030 41318 35076 41370
rect 35100 41318 35146 41370
rect 35146 41318 35156 41370
rect 35180 41318 35210 41370
rect 35210 41318 35236 41370
rect 34940 41316 34996 41318
rect 35020 41316 35076 41318
rect 35100 41316 35156 41318
rect 35180 41316 35236 41318
rect 34940 40282 34996 40284
rect 35020 40282 35076 40284
rect 35100 40282 35156 40284
rect 35180 40282 35236 40284
rect 34940 40230 34966 40282
rect 34966 40230 34996 40282
rect 35020 40230 35030 40282
rect 35030 40230 35076 40282
rect 35100 40230 35146 40282
rect 35146 40230 35156 40282
rect 35180 40230 35210 40282
rect 35210 40230 35236 40282
rect 34940 40228 34996 40230
rect 35020 40228 35076 40230
rect 35100 40228 35156 40230
rect 35180 40228 35236 40230
rect 34794 39480 34850 39536
rect 34940 39194 34996 39196
rect 35020 39194 35076 39196
rect 35100 39194 35156 39196
rect 35180 39194 35236 39196
rect 34940 39142 34966 39194
rect 34966 39142 34996 39194
rect 35020 39142 35030 39194
rect 35030 39142 35076 39194
rect 35100 39142 35146 39194
rect 35146 39142 35156 39194
rect 35180 39142 35210 39194
rect 35210 39142 35236 39194
rect 34940 39140 34996 39142
rect 35020 39140 35076 39142
rect 35100 39140 35156 39142
rect 35180 39140 35236 39142
rect 34702 38256 34758 38312
rect 34940 38106 34996 38108
rect 35020 38106 35076 38108
rect 35100 38106 35156 38108
rect 35180 38106 35236 38108
rect 34940 38054 34966 38106
rect 34966 38054 34996 38106
rect 35020 38054 35030 38106
rect 35030 38054 35076 38106
rect 35100 38054 35146 38106
rect 35146 38054 35156 38106
rect 35180 38054 35210 38106
rect 35210 38054 35236 38106
rect 34940 38052 34996 38054
rect 35020 38052 35076 38054
rect 35100 38052 35156 38054
rect 35180 38052 35236 38054
rect 34940 37018 34996 37020
rect 35020 37018 35076 37020
rect 35100 37018 35156 37020
rect 35180 37018 35236 37020
rect 34940 36966 34966 37018
rect 34966 36966 34996 37018
rect 35020 36966 35030 37018
rect 35030 36966 35076 37018
rect 35100 36966 35146 37018
rect 35146 36966 35156 37018
rect 35180 36966 35210 37018
rect 35210 36966 35236 37018
rect 34940 36964 34996 36966
rect 35020 36964 35076 36966
rect 35100 36964 35156 36966
rect 35180 36964 35236 36966
rect 34940 35930 34996 35932
rect 35020 35930 35076 35932
rect 35100 35930 35156 35932
rect 35180 35930 35236 35932
rect 34940 35878 34966 35930
rect 34966 35878 34996 35930
rect 35020 35878 35030 35930
rect 35030 35878 35076 35930
rect 35100 35878 35146 35930
rect 35146 35878 35156 35930
rect 35180 35878 35210 35930
rect 35210 35878 35236 35930
rect 34940 35876 34996 35878
rect 35020 35876 35076 35878
rect 35100 35876 35156 35878
rect 35180 35876 35236 35878
rect 34940 34842 34996 34844
rect 35020 34842 35076 34844
rect 35100 34842 35156 34844
rect 35180 34842 35236 34844
rect 34940 34790 34966 34842
rect 34966 34790 34996 34842
rect 35020 34790 35030 34842
rect 35030 34790 35076 34842
rect 35100 34790 35146 34842
rect 35146 34790 35156 34842
rect 35180 34790 35210 34842
rect 35210 34790 35236 34842
rect 34940 34788 34996 34790
rect 35020 34788 35076 34790
rect 35100 34788 35156 34790
rect 35180 34788 35236 34790
rect 34940 33754 34996 33756
rect 35020 33754 35076 33756
rect 35100 33754 35156 33756
rect 35180 33754 35236 33756
rect 34940 33702 34966 33754
rect 34966 33702 34996 33754
rect 35020 33702 35030 33754
rect 35030 33702 35076 33754
rect 35100 33702 35146 33754
rect 35146 33702 35156 33754
rect 35180 33702 35210 33754
rect 35210 33702 35236 33754
rect 34940 33700 34996 33702
rect 35020 33700 35076 33702
rect 35100 33700 35156 33702
rect 35180 33700 35236 33702
rect 34940 32666 34996 32668
rect 35020 32666 35076 32668
rect 35100 32666 35156 32668
rect 35180 32666 35236 32668
rect 34940 32614 34966 32666
rect 34966 32614 34996 32666
rect 35020 32614 35030 32666
rect 35030 32614 35076 32666
rect 35100 32614 35146 32666
rect 35146 32614 35156 32666
rect 35180 32614 35210 32666
rect 35210 32614 35236 32666
rect 34940 32612 34996 32614
rect 35020 32612 35076 32614
rect 35100 32612 35156 32614
rect 35180 32612 35236 32614
rect 34940 31578 34996 31580
rect 35020 31578 35076 31580
rect 35100 31578 35156 31580
rect 35180 31578 35236 31580
rect 34940 31526 34966 31578
rect 34966 31526 34996 31578
rect 35020 31526 35030 31578
rect 35030 31526 35076 31578
rect 35100 31526 35146 31578
rect 35146 31526 35156 31578
rect 35180 31526 35210 31578
rect 35210 31526 35236 31578
rect 34940 31524 34996 31526
rect 35020 31524 35076 31526
rect 35100 31524 35156 31526
rect 35180 31524 35236 31526
rect 34940 30490 34996 30492
rect 35020 30490 35076 30492
rect 35100 30490 35156 30492
rect 35180 30490 35236 30492
rect 34940 30438 34966 30490
rect 34966 30438 34996 30490
rect 35020 30438 35030 30490
rect 35030 30438 35076 30490
rect 35100 30438 35146 30490
rect 35146 30438 35156 30490
rect 35180 30438 35210 30490
rect 35210 30438 35236 30490
rect 34940 30436 34996 30438
rect 35020 30436 35076 30438
rect 35100 30436 35156 30438
rect 35180 30436 35236 30438
rect 34940 29402 34996 29404
rect 35020 29402 35076 29404
rect 35100 29402 35156 29404
rect 35180 29402 35236 29404
rect 34940 29350 34966 29402
rect 34966 29350 34996 29402
rect 35020 29350 35030 29402
rect 35030 29350 35076 29402
rect 35100 29350 35146 29402
rect 35146 29350 35156 29402
rect 35180 29350 35210 29402
rect 35210 29350 35236 29402
rect 34940 29348 34996 29350
rect 35020 29348 35076 29350
rect 35100 29348 35156 29350
rect 35180 29348 35236 29350
rect 34940 28314 34996 28316
rect 35020 28314 35076 28316
rect 35100 28314 35156 28316
rect 35180 28314 35236 28316
rect 34940 28262 34966 28314
rect 34966 28262 34996 28314
rect 35020 28262 35030 28314
rect 35030 28262 35076 28314
rect 35100 28262 35146 28314
rect 35146 28262 35156 28314
rect 35180 28262 35210 28314
rect 35210 28262 35236 28314
rect 34940 28260 34996 28262
rect 35020 28260 35076 28262
rect 35100 28260 35156 28262
rect 35180 28260 35236 28262
rect 34058 27512 34114 27568
rect 34702 27512 34758 27568
rect 33782 23568 33838 23624
rect 34518 17856 34574 17912
rect 34518 13640 34574 13696
rect 32126 12416 32182 12472
rect 33138 12416 33194 12472
rect 34940 27226 34996 27228
rect 35020 27226 35076 27228
rect 35100 27226 35156 27228
rect 35180 27226 35236 27228
rect 34940 27174 34966 27226
rect 34966 27174 34996 27226
rect 35020 27174 35030 27226
rect 35030 27174 35076 27226
rect 35100 27174 35146 27226
rect 35146 27174 35156 27226
rect 35180 27174 35210 27226
rect 35210 27174 35236 27226
rect 34940 27172 34996 27174
rect 35020 27172 35076 27174
rect 35100 27172 35156 27174
rect 35180 27172 35236 27174
rect 34940 26138 34996 26140
rect 35020 26138 35076 26140
rect 35100 26138 35156 26140
rect 35180 26138 35236 26140
rect 34940 26086 34966 26138
rect 34966 26086 34996 26138
rect 35020 26086 35030 26138
rect 35030 26086 35076 26138
rect 35100 26086 35146 26138
rect 35146 26086 35156 26138
rect 35180 26086 35210 26138
rect 35210 26086 35236 26138
rect 34940 26084 34996 26086
rect 35020 26084 35076 26086
rect 35100 26084 35156 26086
rect 35180 26084 35236 26086
rect 34940 25050 34996 25052
rect 35020 25050 35076 25052
rect 35100 25050 35156 25052
rect 35180 25050 35236 25052
rect 34940 24998 34966 25050
rect 34966 24998 34996 25050
rect 35020 24998 35030 25050
rect 35030 24998 35076 25050
rect 35100 24998 35146 25050
rect 35146 24998 35156 25050
rect 35180 24998 35210 25050
rect 35210 24998 35236 25050
rect 34940 24996 34996 24998
rect 35020 24996 35076 24998
rect 35100 24996 35156 24998
rect 35180 24996 35236 24998
rect 34940 23962 34996 23964
rect 35020 23962 35076 23964
rect 35100 23962 35156 23964
rect 35180 23962 35236 23964
rect 34940 23910 34966 23962
rect 34966 23910 34996 23962
rect 35020 23910 35030 23962
rect 35030 23910 35076 23962
rect 35100 23910 35146 23962
rect 35146 23910 35156 23962
rect 35180 23910 35210 23962
rect 35210 23910 35236 23962
rect 34940 23908 34996 23910
rect 35020 23908 35076 23910
rect 35100 23908 35156 23910
rect 35180 23908 35236 23910
rect 34940 22874 34996 22876
rect 35020 22874 35076 22876
rect 35100 22874 35156 22876
rect 35180 22874 35236 22876
rect 34940 22822 34966 22874
rect 34966 22822 34996 22874
rect 35020 22822 35030 22874
rect 35030 22822 35076 22874
rect 35100 22822 35146 22874
rect 35146 22822 35156 22874
rect 35180 22822 35210 22874
rect 35210 22822 35236 22874
rect 34940 22820 34996 22822
rect 35020 22820 35076 22822
rect 35100 22820 35156 22822
rect 35180 22820 35236 22822
rect 34940 21786 34996 21788
rect 35020 21786 35076 21788
rect 35100 21786 35156 21788
rect 35180 21786 35236 21788
rect 34940 21734 34966 21786
rect 34966 21734 34996 21786
rect 35020 21734 35030 21786
rect 35030 21734 35076 21786
rect 35100 21734 35146 21786
rect 35146 21734 35156 21786
rect 35180 21734 35210 21786
rect 35210 21734 35236 21786
rect 34940 21732 34996 21734
rect 35020 21732 35076 21734
rect 35100 21732 35156 21734
rect 35180 21732 35236 21734
rect 34940 20698 34996 20700
rect 35020 20698 35076 20700
rect 35100 20698 35156 20700
rect 35180 20698 35236 20700
rect 34940 20646 34966 20698
rect 34966 20646 34996 20698
rect 35020 20646 35030 20698
rect 35030 20646 35076 20698
rect 35100 20646 35146 20698
rect 35146 20646 35156 20698
rect 35180 20646 35210 20698
rect 35210 20646 35236 20698
rect 34940 20644 34996 20646
rect 35020 20644 35076 20646
rect 35100 20644 35156 20646
rect 35180 20644 35236 20646
rect 34940 19610 34996 19612
rect 35020 19610 35076 19612
rect 35100 19610 35156 19612
rect 35180 19610 35236 19612
rect 34940 19558 34966 19610
rect 34966 19558 34996 19610
rect 35020 19558 35030 19610
rect 35030 19558 35076 19610
rect 35100 19558 35146 19610
rect 35146 19558 35156 19610
rect 35180 19558 35210 19610
rect 35210 19558 35236 19610
rect 34940 19556 34996 19558
rect 35020 19556 35076 19558
rect 35100 19556 35156 19558
rect 35180 19556 35236 19558
rect 34940 18522 34996 18524
rect 35020 18522 35076 18524
rect 35100 18522 35156 18524
rect 35180 18522 35236 18524
rect 34940 18470 34966 18522
rect 34966 18470 34996 18522
rect 35020 18470 35030 18522
rect 35030 18470 35076 18522
rect 35100 18470 35146 18522
rect 35146 18470 35156 18522
rect 35180 18470 35210 18522
rect 35210 18470 35236 18522
rect 34940 18468 34996 18470
rect 35020 18468 35076 18470
rect 35100 18468 35156 18470
rect 35180 18468 35236 18470
rect 35438 56752 35494 56808
rect 35530 56480 35586 56536
rect 35438 55120 35494 55176
rect 35438 53760 35494 53816
rect 35438 51992 35494 52048
rect 35438 50496 35494 50552
rect 35438 48320 35494 48376
rect 35346 43560 35402 43616
rect 35622 48592 35678 48648
rect 35622 46960 35678 47016
rect 37646 45464 37702 45520
rect 35622 41112 35678 41168
rect 35530 40704 35586 40760
rect 35346 40568 35402 40624
rect 35622 38120 35678 38176
rect 35530 37168 35586 37224
rect 35438 35400 35494 35456
rect 35438 34176 35494 34232
rect 35530 33360 35586 33416
rect 35346 27376 35402 27432
rect 35254 17720 35310 17776
rect 34940 17434 34996 17436
rect 35020 17434 35076 17436
rect 35100 17434 35156 17436
rect 35180 17434 35236 17436
rect 34940 17382 34966 17434
rect 34966 17382 34996 17434
rect 35020 17382 35030 17434
rect 35030 17382 35076 17434
rect 35100 17382 35146 17434
rect 35146 17382 35156 17434
rect 35180 17382 35210 17434
rect 35210 17382 35236 17434
rect 34940 17380 34996 17382
rect 35020 17380 35076 17382
rect 35100 17380 35156 17382
rect 35180 17380 35236 17382
rect 35806 26288 35862 26344
rect 36358 26288 36414 26344
rect 35622 20440 35678 20496
rect 35438 19896 35494 19952
rect 35346 16360 35402 16416
rect 34940 16346 34996 16348
rect 35020 16346 35076 16348
rect 35100 16346 35156 16348
rect 35180 16346 35236 16348
rect 34940 16294 34966 16346
rect 34966 16294 34996 16346
rect 35020 16294 35030 16346
rect 35030 16294 35076 16346
rect 35100 16294 35146 16346
rect 35146 16294 35156 16346
rect 35180 16294 35210 16346
rect 35210 16294 35236 16346
rect 34940 16292 34996 16294
rect 35020 16292 35076 16294
rect 35100 16292 35156 16294
rect 35180 16292 35236 16294
rect 34940 15258 34996 15260
rect 35020 15258 35076 15260
rect 35100 15258 35156 15260
rect 35180 15258 35236 15260
rect 34940 15206 34966 15258
rect 34966 15206 34996 15258
rect 35020 15206 35030 15258
rect 35030 15206 35076 15258
rect 35100 15206 35146 15258
rect 35146 15206 35156 15258
rect 35180 15206 35210 15258
rect 35210 15206 35236 15258
rect 34940 15204 34996 15206
rect 35020 15204 35076 15206
rect 35100 15204 35156 15206
rect 35180 15204 35236 15206
rect 34940 14170 34996 14172
rect 35020 14170 35076 14172
rect 35100 14170 35156 14172
rect 35180 14170 35236 14172
rect 34940 14118 34966 14170
rect 34966 14118 34996 14170
rect 35020 14118 35030 14170
rect 35030 14118 35076 14170
rect 35100 14118 35146 14170
rect 35146 14118 35156 14170
rect 35180 14118 35210 14170
rect 35210 14118 35236 14170
rect 34940 14116 34996 14118
rect 35020 14116 35076 14118
rect 35100 14116 35156 14118
rect 35180 14116 35236 14118
rect 34940 13082 34996 13084
rect 35020 13082 35076 13084
rect 35100 13082 35156 13084
rect 35180 13082 35236 13084
rect 34940 13030 34966 13082
rect 34966 13030 34996 13082
rect 35020 13030 35030 13082
rect 35030 13030 35076 13082
rect 35100 13030 35146 13082
rect 35146 13030 35156 13082
rect 35180 13030 35210 13082
rect 35210 13030 35236 13082
rect 34940 13028 34996 13030
rect 35020 13028 35076 13030
rect 35100 13028 35156 13030
rect 35180 13028 35236 13030
rect 32678 5208 32734 5264
rect 34940 11994 34996 11996
rect 35020 11994 35076 11996
rect 35100 11994 35156 11996
rect 35180 11994 35236 11996
rect 34940 11942 34966 11994
rect 34966 11942 34996 11994
rect 35020 11942 35030 11994
rect 35030 11942 35076 11994
rect 35100 11942 35146 11994
rect 35146 11942 35156 11994
rect 35180 11942 35210 11994
rect 35210 11942 35236 11994
rect 34940 11940 34996 11942
rect 35020 11940 35076 11942
rect 35100 11940 35156 11942
rect 35180 11940 35236 11942
rect 34940 10906 34996 10908
rect 35020 10906 35076 10908
rect 35100 10906 35156 10908
rect 35180 10906 35236 10908
rect 34940 10854 34966 10906
rect 34966 10854 34996 10906
rect 35020 10854 35030 10906
rect 35030 10854 35076 10906
rect 35100 10854 35146 10906
rect 35146 10854 35156 10906
rect 35180 10854 35210 10906
rect 35210 10854 35236 10906
rect 34940 10852 34996 10854
rect 35020 10852 35076 10854
rect 35100 10852 35156 10854
rect 35180 10852 35236 10854
rect 35622 13504 35678 13560
rect 35438 10920 35494 10976
rect 34940 9818 34996 9820
rect 35020 9818 35076 9820
rect 35100 9818 35156 9820
rect 35180 9818 35236 9820
rect 34940 9766 34966 9818
rect 34966 9766 34996 9818
rect 35020 9766 35030 9818
rect 35030 9766 35076 9818
rect 35100 9766 35146 9818
rect 35146 9766 35156 9818
rect 35180 9766 35210 9818
rect 35210 9766 35236 9818
rect 34940 9764 34996 9766
rect 35020 9764 35076 9766
rect 35100 9764 35156 9766
rect 35180 9764 35236 9766
rect 34940 8730 34996 8732
rect 35020 8730 35076 8732
rect 35100 8730 35156 8732
rect 35180 8730 35236 8732
rect 34940 8678 34966 8730
rect 34966 8678 34996 8730
rect 35020 8678 35030 8730
rect 35030 8678 35076 8730
rect 35100 8678 35146 8730
rect 35146 8678 35156 8730
rect 35180 8678 35210 8730
rect 35210 8678 35236 8730
rect 34940 8676 34996 8678
rect 35020 8676 35076 8678
rect 35100 8676 35156 8678
rect 35180 8676 35236 8678
rect 34940 7642 34996 7644
rect 35020 7642 35076 7644
rect 35100 7642 35156 7644
rect 35180 7642 35236 7644
rect 34940 7590 34966 7642
rect 34966 7590 34996 7642
rect 35020 7590 35030 7642
rect 35030 7590 35076 7642
rect 35100 7590 35146 7642
rect 35146 7590 35156 7642
rect 35180 7590 35210 7642
rect 35210 7590 35236 7642
rect 34940 7588 34996 7590
rect 35020 7588 35076 7590
rect 35100 7588 35156 7590
rect 35180 7588 35236 7590
rect 34518 7520 34574 7576
rect 34940 6554 34996 6556
rect 35020 6554 35076 6556
rect 35100 6554 35156 6556
rect 35180 6554 35236 6556
rect 34940 6502 34966 6554
rect 34966 6502 34996 6554
rect 35020 6502 35030 6554
rect 35030 6502 35076 6554
rect 35100 6502 35146 6554
rect 35146 6502 35156 6554
rect 35180 6502 35210 6554
rect 35210 6502 35236 6554
rect 34940 6500 34996 6502
rect 35020 6500 35076 6502
rect 35100 6500 35156 6502
rect 35180 6500 35236 6502
rect 34940 5466 34996 5468
rect 35020 5466 35076 5468
rect 35100 5466 35156 5468
rect 35180 5466 35236 5468
rect 34940 5414 34966 5466
rect 34966 5414 34996 5466
rect 35020 5414 35030 5466
rect 35030 5414 35076 5466
rect 35100 5414 35146 5466
rect 35146 5414 35156 5466
rect 35180 5414 35210 5466
rect 35210 5414 35236 5466
rect 34940 5412 34996 5414
rect 35020 5412 35076 5414
rect 35100 5412 35156 5414
rect 35180 5412 35236 5414
rect 34940 4378 34996 4380
rect 35020 4378 35076 4380
rect 35100 4378 35156 4380
rect 35180 4378 35236 4380
rect 34940 4326 34966 4378
rect 34966 4326 34996 4378
rect 35020 4326 35030 4378
rect 35030 4326 35076 4378
rect 35100 4326 35146 4378
rect 35146 4326 35156 4378
rect 35180 4326 35210 4378
rect 35210 4326 35236 4378
rect 34940 4324 34996 4326
rect 35020 4324 35076 4326
rect 35100 4324 35156 4326
rect 35180 4324 35236 4326
rect 34940 3290 34996 3292
rect 35020 3290 35076 3292
rect 35100 3290 35156 3292
rect 35180 3290 35236 3292
rect 34940 3238 34966 3290
rect 34966 3238 34996 3290
rect 35020 3238 35030 3290
rect 35030 3238 35076 3290
rect 35100 3238 35146 3290
rect 35146 3238 35156 3290
rect 35180 3238 35210 3290
rect 35210 3238 35236 3290
rect 34940 3236 34996 3238
rect 35020 3236 35076 3238
rect 35100 3236 35156 3238
rect 35180 3236 35236 3238
rect 34940 2202 34996 2204
rect 35020 2202 35076 2204
rect 35100 2202 35156 2204
rect 35180 2202 35236 2204
rect 34940 2150 34966 2202
rect 34966 2150 34996 2202
rect 35020 2150 35030 2202
rect 35030 2150 35076 2202
rect 35100 2150 35146 2202
rect 35146 2150 35156 2202
rect 35180 2150 35210 2202
rect 35210 2150 35236 2202
rect 34940 2148 34996 2150
rect 35020 2148 35076 2150
rect 35100 2148 35156 2150
rect 35180 2148 35236 2150
rect 37738 20304 37794 20360
rect 37370 15816 37426 15872
rect 36358 9016 36414 9072
rect 36266 6316 36322 6352
rect 36266 6296 36268 6316
rect 36268 6296 36320 6316
rect 36320 6296 36322 6316
rect 35990 5652 35992 5672
rect 35992 5652 36044 5672
rect 36044 5652 36046 5672
rect 35990 5616 36046 5652
rect 35806 3440 35862 3496
rect 37462 15000 37518 15056
rect 37554 13232 37610 13288
rect 37370 6160 37426 6216
rect 22742 176 22798 232
<< metal3 >>
rect 0 79658 800 79688
rect 3969 79658 4035 79661
rect 0 79656 4035 79658
rect 0 79600 3974 79656
rect 4030 79600 4035 79656
rect 0 79598 4035 79600
rect 0 79568 800 79598
rect 3969 79595 4035 79598
rect 35433 79658 35499 79661
rect 39200 79658 40000 79688
rect 35433 79656 40000 79658
rect 35433 79600 35438 79656
rect 35494 79600 40000 79656
rect 35433 79598 40000 79600
rect 35433 79595 35499 79598
rect 39200 79568 40000 79598
rect 0 78298 800 78328
rect 4061 78298 4127 78301
rect 0 78296 4127 78298
rect 0 78240 4066 78296
rect 4122 78240 4127 78296
rect 0 78238 4127 78240
rect 0 78208 800 78238
rect 4061 78235 4127 78238
rect 35341 78298 35407 78301
rect 39200 78298 40000 78328
rect 35341 78296 40000 78298
rect 35341 78240 35346 78296
rect 35402 78240 40000 78296
rect 35341 78238 40000 78240
rect 35341 78235 35407 78238
rect 39200 78208 40000 78238
rect 19568 77824 19888 77825
rect 19568 77760 19576 77824
rect 19640 77760 19656 77824
rect 19720 77760 19736 77824
rect 19800 77760 19816 77824
rect 19880 77760 19888 77824
rect 19568 77759 19888 77760
rect 4208 77280 4528 77281
rect 4208 77216 4216 77280
rect 4280 77216 4296 77280
rect 4360 77216 4376 77280
rect 4440 77216 4456 77280
rect 4520 77216 4528 77280
rect 4208 77215 4528 77216
rect 34928 77280 35248 77281
rect 34928 77216 34936 77280
rect 35000 77216 35016 77280
rect 35080 77216 35096 77280
rect 35160 77216 35176 77280
rect 35240 77216 35248 77280
rect 34928 77215 35248 77216
rect 17493 77210 17559 77213
rect 24393 77210 24459 77213
rect 17493 77208 24459 77210
rect 17493 77152 17498 77208
rect 17554 77152 24398 77208
rect 24454 77152 24459 77208
rect 17493 77150 24459 77152
rect 17493 77147 17559 77150
rect 24393 77147 24459 77150
rect 0 76938 800 76968
rect 2405 76938 2471 76941
rect 0 76936 2471 76938
rect 0 76880 2410 76936
rect 2466 76880 2471 76936
rect 0 76878 2471 76880
rect 0 76848 800 76878
rect 2405 76875 2471 76878
rect 35801 76938 35867 76941
rect 39200 76938 40000 76968
rect 35801 76936 40000 76938
rect 35801 76880 35806 76936
rect 35862 76880 40000 76936
rect 35801 76878 40000 76880
rect 35801 76875 35867 76878
rect 39200 76848 40000 76878
rect 19568 76736 19888 76737
rect 19568 76672 19576 76736
rect 19640 76672 19656 76736
rect 19720 76672 19736 76736
rect 19800 76672 19816 76736
rect 19880 76672 19888 76736
rect 19568 76671 19888 76672
rect 21173 76394 21239 76397
rect 24117 76394 24183 76397
rect 21173 76392 24183 76394
rect 21173 76336 21178 76392
rect 21234 76336 24122 76392
rect 24178 76336 24183 76392
rect 21173 76334 24183 76336
rect 21173 76331 21239 76334
rect 24117 76331 24183 76334
rect 4208 76192 4528 76193
rect 4208 76128 4216 76192
rect 4280 76128 4296 76192
rect 4360 76128 4376 76192
rect 4440 76128 4456 76192
rect 4520 76128 4528 76192
rect 4208 76127 4528 76128
rect 34928 76192 35248 76193
rect 34928 76128 34936 76192
rect 35000 76128 35016 76192
rect 35080 76128 35096 76192
rect 35160 76128 35176 76192
rect 35240 76128 35248 76192
rect 34928 76127 35248 76128
rect 24669 76122 24735 76125
rect 25865 76122 25931 76125
rect 28809 76122 28875 76125
rect 24669 76120 28875 76122
rect 24669 76064 24674 76120
rect 24730 76064 25870 76120
rect 25926 76064 28814 76120
rect 28870 76064 28875 76120
rect 24669 76062 28875 76064
rect 24669 76059 24735 76062
rect 25865 76059 25931 76062
rect 28809 76059 28875 76062
rect 473 75850 539 75853
rect 1669 75850 1735 75853
rect 473 75848 1735 75850
rect 473 75792 478 75848
rect 534 75792 1674 75848
rect 1730 75792 1735 75848
rect 473 75790 1735 75792
rect 473 75787 539 75790
rect 1669 75787 1735 75790
rect 13353 75850 13419 75853
rect 16389 75850 16455 75853
rect 13353 75848 16455 75850
rect 13353 75792 13358 75848
rect 13414 75792 16394 75848
rect 16450 75792 16455 75848
rect 13353 75790 16455 75792
rect 13353 75787 13419 75790
rect 16389 75787 16455 75790
rect 19568 75648 19888 75649
rect 0 75578 800 75608
rect 19568 75584 19576 75648
rect 19640 75584 19656 75648
rect 19720 75584 19736 75648
rect 19800 75584 19816 75648
rect 19880 75584 19888 75648
rect 19568 75583 19888 75584
rect 3325 75578 3391 75581
rect 0 75576 3391 75578
rect 0 75520 3330 75576
rect 3386 75520 3391 75576
rect 0 75518 3391 75520
rect 0 75488 800 75518
rect 3325 75515 3391 75518
rect 29821 75578 29887 75581
rect 34789 75578 34855 75581
rect 29821 75576 34855 75578
rect 29821 75520 29826 75576
rect 29882 75520 34794 75576
rect 34850 75520 34855 75576
rect 29821 75518 34855 75520
rect 29821 75515 29887 75518
rect 34789 75515 34855 75518
rect 35617 75578 35683 75581
rect 39200 75578 40000 75608
rect 35617 75576 40000 75578
rect 35617 75520 35622 75576
rect 35678 75520 40000 75576
rect 35617 75518 40000 75520
rect 35617 75515 35683 75518
rect 39200 75488 40000 75518
rect 1853 75442 1919 75445
rect 12341 75442 12407 75445
rect 1853 75440 12407 75442
rect 1853 75384 1858 75440
rect 1914 75384 12346 75440
rect 12402 75384 12407 75440
rect 1853 75382 12407 75384
rect 1853 75379 1919 75382
rect 12341 75379 12407 75382
rect 10593 75306 10659 75309
rect 21357 75306 21423 75309
rect 10593 75304 21423 75306
rect 10593 75248 10598 75304
rect 10654 75248 21362 75304
rect 21418 75248 21423 75304
rect 10593 75246 21423 75248
rect 10593 75243 10659 75246
rect 21357 75243 21423 75246
rect 6453 75170 6519 75173
rect 19977 75170 20043 75173
rect 6453 75168 20043 75170
rect 6453 75112 6458 75168
rect 6514 75112 19982 75168
rect 20038 75112 20043 75168
rect 6453 75110 20043 75112
rect 6453 75107 6519 75110
rect 19977 75107 20043 75110
rect 4208 75104 4528 75105
rect 4208 75040 4216 75104
rect 4280 75040 4296 75104
rect 4360 75040 4376 75104
rect 4440 75040 4456 75104
rect 4520 75040 4528 75104
rect 4208 75039 4528 75040
rect 34928 75104 35248 75105
rect 34928 75040 34936 75104
rect 35000 75040 35016 75104
rect 35080 75040 35096 75104
rect 35160 75040 35176 75104
rect 35240 75040 35248 75104
rect 34928 75039 35248 75040
rect 17769 75034 17835 75037
rect 31753 75034 31819 75037
rect 17769 75032 31819 75034
rect 17769 74976 17774 75032
rect 17830 74976 31758 75032
rect 31814 74976 31819 75032
rect 17769 74974 31819 74976
rect 17769 74971 17835 74974
rect 31753 74971 31819 74974
rect 7373 74898 7439 74901
rect 9397 74898 9463 74901
rect 7373 74896 9463 74898
rect 7373 74840 7378 74896
rect 7434 74840 9402 74896
rect 9458 74840 9463 74896
rect 7373 74838 9463 74840
rect 7373 74835 7439 74838
rect 9397 74835 9463 74838
rect 4613 74762 4679 74765
rect 6177 74762 6243 74765
rect 4613 74760 6243 74762
rect 4613 74704 4618 74760
rect 4674 74704 6182 74760
rect 6238 74704 6243 74760
rect 4613 74702 6243 74704
rect 4613 74699 4679 74702
rect 6177 74699 6243 74702
rect 8753 74762 8819 74765
rect 10409 74762 10475 74765
rect 8753 74760 10475 74762
rect 8753 74704 8758 74760
rect 8814 74704 10414 74760
rect 10470 74704 10475 74760
rect 8753 74702 10475 74704
rect 8753 74699 8819 74702
rect 10409 74699 10475 74702
rect 19568 74560 19888 74561
rect 19568 74496 19576 74560
rect 19640 74496 19656 74560
rect 19720 74496 19736 74560
rect 19800 74496 19816 74560
rect 19880 74496 19888 74560
rect 19568 74495 19888 74496
rect 20253 74490 20319 74493
rect 21265 74490 21331 74493
rect 20253 74488 21331 74490
rect 20253 74432 20258 74488
rect 20314 74432 21270 74488
rect 21326 74432 21331 74488
rect 20253 74430 21331 74432
rect 20253 74427 20319 74430
rect 21265 74427 21331 74430
rect 24761 74490 24827 74493
rect 27981 74490 28047 74493
rect 24761 74488 28047 74490
rect 24761 74432 24766 74488
rect 24822 74432 27986 74488
rect 28042 74432 28047 74488
rect 24761 74430 28047 74432
rect 24761 74427 24827 74430
rect 27981 74427 28047 74430
rect 0 74218 800 74248
rect 3785 74218 3851 74221
rect 0 74216 3851 74218
rect 0 74160 3790 74216
rect 3846 74160 3851 74216
rect 0 74158 3851 74160
rect 0 74128 800 74158
rect 3785 74155 3851 74158
rect 31017 74218 31083 74221
rect 39200 74218 40000 74248
rect 31017 74216 40000 74218
rect 31017 74160 31022 74216
rect 31078 74160 40000 74216
rect 31017 74158 40000 74160
rect 31017 74155 31083 74158
rect 39200 74128 40000 74158
rect 4208 74016 4528 74017
rect 4208 73952 4216 74016
rect 4280 73952 4296 74016
rect 4360 73952 4376 74016
rect 4440 73952 4456 74016
rect 4520 73952 4528 74016
rect 4208 73951 4528 73952
rect 34928 74016 35248 74017
rect 34928 73952 34936 74016
rect 35000 73952 35016 74016
rect 35080 73952 35096 74016
rect 35160 73952 35176 74016
rect 35240 73952 35248 74016
rect 34928 73951 35248 73952
rect 14273 73946 14339 73949
rect 25681 73946 25747 73949
rect 14273 73944 25747 73946
rect 14273 73888 14278 73944
rect 14334 73888 25686 73944
rect 25742 73888 25747 73944
rect 14273 73886 25747 73888
rect 14273 73883 14339 73886
rect 25681 73883 25747 73886
rect 15377 73810 15443 73813
rect 39573 73810 39639 73813
rect 15377 73808 39639 73810
rect 15377 73752 15382 73808
rect 15438 73752 39578 73808
rect 39634 73752 39639 73808
rect 15377 73750 39639 73752
rect 15377 73747 15443 73750
rect 39573 73747 39639 73750
rect 19568 73472 19888 73473
rect 19568 73408 19576 73472
rect 19640 73408 19656 73472
rect 19720 73408 19736 73472
rect 19800 73408 19816 73472
rect 19880 73408 19888 73472
rect 19568 73407 19888 73408
rect 21817 73266 21883 73269
rect 23933 73266 23999 73269
rect 21817 73264 23999 73266
rect 21817 73208 21822 73264
rect 21878 73208 23938 73264
rect 23994 73208 23999 73264
rect 21817 73206 23999 73208
rect 21817 73203 21883 73206
rect 23933 73203 23999 73206
rect 28942 73204 28948 73268
rect 29012 73266 29018 73268
rect 36813 73266 36879 73269
rect 29012 73264 36879 73266
rect 29012 73208 36818 73264
rect 36874 73208 36879 73264
rect 29012 73206 36879 73208
rect 29012 73204 29018 73206
rect 36813 73203 36879 73206
rect 19333 72994 19399 72997
rect 16254 72992 19399 72994
rect 16254 72936 19338 72992
rect 19394 72936 19399 72992
rect 16254 72934 19399 72936
rect 4208 72928 4528 72929
rect 0 72858 800 72888
rect 4208 72864 4216 72928
rect 4280 72864 4296 72928
rect 4360 72864 4376 72928
rect 4440 72864 4456 72928
rect 4520 72864 4528 72928
rect 4208 72863 4528 72864
rect 4061 72858 4127 72861
rect 0 72856 4127 72858
rect 0 72800 4066 72856
rect 4122 72800 4127 72856
rect 0 72798 4127 72800
rect 0 72768 800 72798
rect 4061 72795 4127 72798
rect 8937 72858 9003 72861
rect 16254 72858 16314 72934
rect 19333 72931 19399 72934
rect 28809 72994 28875 72997
rect 28942 72994 28948 72996
rect 28809 72992 28948 72994
rect 28809 72936 28814 72992
rect 28870 72936 28948 72992
rect 28809 72934 28948 72936
rect 28809 72931 28875 72934
rect 28942 72932 28948 72934
rect 29012 72932 29018 72996
rect 34928 72928 35248 72929
rect 34928 72864 34936 72928
rect 35000 72864 35016 72928
rect 35080 72864 35096 72928
rect 35160 72864 35176 72928
rect 35240 72864 35248 72928
rect 34928 72863 35248 72864
rect 8937 72856 16314 72858
rect 8937 72800 8942 72856
rect 8998 72800 16314 72856
rect 8937 72798 16314 72800
rect 16389 72858 16455 72861
rect 27429 72858 27495 72861
rect 16389 72856 27495 72858
rect 16389 72800 16394 72856
rect 16450 72800 27434 72856
rect 27490 72800 27495 72856
rect 16389 72798 27495 72800
rect 8937 72795 9003 72798
rect 16389 72795 16455 72798
rect 27429 72795 27495 72798
rect 35433 72858 35499 72861
rect 39200 72858 40000 72888
rect 35433 72856 40000 72858
rect 35433 72800 35438 72856
rect 35494 72800 40000 72856
rect 35433 72798 40000 72800
rect 35433 72795 35499 72798
rect 39200 72768 40000 72798
rect 3785 72586 3851 72589
rect 19333 72586 19399 72589
rect 3785 72584 19399 72586
rect 3785 72528 3790 72584
rect 3846 72528 19338 72584
rect 19394 72528 19399 72584
rect 3785 72526 19399 72528
rect 3785 72523 3851 72526
rect 19333 72523 19399 72526
rect 19568 72384 19888 72385
rect 19568 72320 19576 72384
rect 19640 72320 19656 72384
rect 19720 72320 19736 72384
rect 19800 72320 19816 72384
rect 19880 72320 19888 72384
rect 19568 72319 19888 72320
rect 4061 72042 4127 72045
rect 15837 72042 15903 72045
rect 4061 72040 15903 72042
rect 4061 71984 4066 72040
rect 4122 71984 15842 72040
rect 15898 71984 15903 72040
rect 4061 71982 15903 71984
rect 4061 71979 4127 71982
rect 15837 71979 15903 71982
rect 14089 71906 14155 71909
rect 19517 71906 19583 71909
rect 21081 71908 21147 71909
rect 21030 71906 21036 71908
rect 14089 71904 19583 71906
rect 14089 71848 14094 71904
rect 14150 71848 19522 71904
rect 19578 71848 19583 71904
rect 14089 71846 19583 71848
rect 20990 71846 21036 71906
rect 21100 71904 21147 71908
rect 21142 71848 21147 71904
rect 14089 71843 14155 71846
rect 19517 71843 19583 71846
rect 21030 71844 21036 71846
rect 21100 71844 21147 71848
rect 21081 71843 21147 71844
rect 4208 71840 4528 71841
rect 4208 71776 4216 71840
rect 4280 71776 4296 71840
rect 4360 71776 4376 71840
rect 4440 71776 4456 71840
rect 4520 71776 4528 71840
rect 4208 71775 4528 71776
rect 34928 71840 35248 71841
rect 34928 71776 34936 71840
rect 35000 71776 35016 71840
rect 35080 71776 35096 71840
rect 35160 71776 35176 71840
rect 35240 71776 35248 71840
rect 34928 71775 35248 71776
rect 4797 71634 4863 71637
rect 798 71632 4863 71634
rect 798 71576 4802 71632
rect 4858 71576 4863 71632
rect 798 71574 4863 71576
rect 798 71528 858 71574
rect 4797 71571 4863 71574
rect 15561 71634 15627 71637
rect 29913 71634 29979 71637
rect 35893 71634 35959 71637
rect 15561 71632 29979 71634
rect 15561 71576 15566 71632
rect 15622 71576 29918 71632
rect 29974 71576 29979 71632
rect 15561 71574 29979 71576
rect 15561 71571 15627 71574
rect 29913 71571 29979 71574
rect 30054 71632 35959 71634
rect 30054 71576 35898 71632
rect 35954 71576 35959 71632
rect 30054 71574 35959 71576
rect 0 71438 858 71528
rect 18229 71498 18295 71501
rect 18229 71496 20730 71498
rect 18229 71440 18234 71496
rect 18290 71440 20730 71496
rect 18229 71438 20730 71440
rect 0 71408 800 71438
rect 18229 71435 18295 71438
rect 19568 71296 19888 71297
rect 19568 71232 19576 71296
rect 19640 71232 19656 71296
rect 19720 71232 19736 71296
rect 19800 71232 19816 71296
rect 19880 71232 19888 71296
rect 19568 71231 19888 71232
rect 20670 71226 20730 71438
rect 30054 71362 30114 71574
rect 35893 71571 35959 71574
rect 34513 71498 34579 71501
rect 39200 71498 40000 71528
rect 34513 71496 40000 71498
rect 34513 71440 34518 71496
rect 34574 71440 40000 71496
rect 34513 71438 40000 71440
rect 34513 71435 34579 71438
rect 39200 71408 40000 71438
rect 22188 71302 30114 71362
rect 22188 71226 22248 71302
rect 20670 71166 22248 71226
rect 15745 70954 15811 70957
rect 23013 70954 23079 70957
rect 15745 70952 23079 70954
rect 15745 70896 15750 70952
rect 15806 70896 23018 70952
rect 23074 70896 23079 70952
rect 15745 70894 23079 70896
rect 15745 70891 15811 70894
rect 23013 70891 23079 70894
rect 24301 70954 24367 70957
rect 35433 70954 35499 70957
rect 24301 70952 35499 70954
rect 24301 70896 24306 70952
rect 24362 70896 35438 70952
rect 35494 70896 35499 70952
rect 24301 70894 35499 70896
rect 24301 70891 24367 70894
rect 35433 70891 35499 70894
rect 4797 70818 4863 70821
rect 15193 70818 15259 70821
rect 4797 70816 15259 70818
rect 4797 70760 4802 70816
rect 4858 70760 15198 70816
rect 15254 70760 15259 70816
rect 4797 70758 15259 70760
rect 4797 70755 4863 70758
rect 15193 70755 15259 70758
rect 4208 70752 4528 70753
rect 4208 70688 4216 70752
rect 4280 70688 4296 70752
rect 4360 70688 4376 70752
rect 4440 70688 4456 70752
rect 4520 70688 4528 70752
rect 4208 70687 4528 70688
rect 34928 70752 35248 70753
rect 34928 70688 34936 70752
rect 35000 70688 35016 70752
rect 35080 70688 35096 70752
rect 35160 70688 35176 70752
rect 35240 70688 35248 70752
rect 34928 70687 35248 70688
rect 11513 70546 11579 70549
rect 15929 70546 15995 70549
rect 11513 70544 15995 70546
rect 11513 70488 11518 70544
rect 11574 70488 15934 70544
rect 15990 70488 15995 70544
rect 11513 70486 15995 70488
rect 11513 70483 11579 70486
rect 15929 70483 15995 70486
rect 19568 70208 19888 70209
rect 0 70138 800 70168
rect 19568 70144 19576 70208
rect 19640 70144 19656 70208
rect 19720 70144 19736 70208
rect 19800 70144 19816 70208
rect 19880 70144 19888 70208
rect 19568 70143 19888 70144
rect 4889 70138 4955 70141
rect 0 70136 4955 70138
rect 0 70080 4894 70136
rect 4950 70080 4955 70136
rect 0 70078 4955 70080
rect 0 70048 800 70078
rect 4889 70075 4955 70078
rect 30373 70138 30439 70141
rect 39200 70138 40000 70168
rect 30373 70136 40000 70138
rect 30373 70080 30378 70136
rect 30434 70080 40000 70136
rect 30373 70078 40000 70080
rect 30373 70075 30439 70078
rect 39200 70048 40000 70078
rect 24209 70002 24275 70005
rect 34513 70002 34579 70005
rect 24209 70000 34579 70002
rect 24209 69944 24214 70000
rect 24270 69944 34518 70000
rect 34574 69944 34579 70000
rect 24209 69942 34579 69944
rect 24209 69939 24275 69942
rect 34513 69939 34579 69942
rect 105 69866 171 69869
rect 7373 69866 7439 69869
rect 105 69864 7439 69866
rect 105 69808 110 69864
rect 166 69808 7378 69864
rect 7434 69808 7439 69864
rect 105 69806 7439 69808
rect 105 69803 171 69806
rect 7373 69803 7439 69806
rect 15193 69866 15259 69869
rect 22829 69866 22895 69869
rect 15193 69864 22895 69866
rect 15193 69808 15198 69864
rect 15254 69808 22834 69864
rect 22890 69808 22895 69864
rect 15193 69806 22895 69808
rect 15193 69803 15259 69806
rect 22829 69803 22895 69806
rect 10685 69730 10751 69733
rect 20897 69730 20963 69733
rect 10685 69728 20963 69730
rect 10685 69672 10690 69728
rect 10746 69672 20902 69728
rect 20958 69672 20963 69728
rect 10685 69670 20963 69672
rect 10685 69667 10751 69670
rect 20897 69667 20963 69670
rect 4208 69664 4528 69665
rect 4208 69600 4216 69664
rect 4280 69600 4296 69664
rect 4360 69600 4376 69664
rect 4440 69600 4456 69664
rect 4520 69600 4528 69664
rect 4208 69599 4528 69600
rect 34928 69664 35248 69665
rect 34928 69600 34936 69664
rect 35000 69600 35016 69664
rect 35080 69600 35096 69664
rect 35160 69600 35176 69664
rect 35240 69600 35248 69664
rect 34928 69599 35248 69600
rect 5625 69594 5691 69597
rect 26141 69594 26207 69597
rect 5625 69592 26207 69594
rect 5625 69536 5630 69592
rect 5686 69536 26146 69592
rect 26202 69536 26207 69592
rect 5625 69534 26207 69536
rect 5625 69531 5691 69534
rect 26141 69531 26207 69534
rect 0 69458 800 69488
rect 3233 69458 3299 69461
rect 0 69456 3299 69458
rect 0 69400 3238 69456
rect 3294 69400 3299 69456
rect 0 69398 3299 69400
rect 0 69368 800 69398
rect 3233 69395 3299 69398
rect 19568 69120 19888 69121
rect 19568 69056 19576 69120
rect 19640 69056 19656 69120
rect 19720 69056 19736 69120
rect 19800 69056 19816 69120
rect 19880 69056 19888 69120
rect 19568 69055 19888 69056
rect 27521 69050 27587 69053
rect 30046 69050 30052 69052
rect 27521 69048 30052 69050
rect 27521 68992 27526 69048
rect 27582 68992 30052 69048
rect 27521 68990 30052 68992
rect 27521 68987 27587 68990
rect 30046 68988 30052 68990
rect 30116 68988 30122 69052
rect 35525 68778 35591 68781
rect 39200 68778 40000 68808
rect 35525 68776 40000 68778
rect 35525 68720 35530 68776
rect 35586 68720 40000 68776
rect 35525 68718 40000 68720
rect 35525 68715 35591 68718
rect 39200 68688 40000 68718
rect 4208 68576 4528 68577
rect 4208 68512 4216 68576
rect 4280 68512 4296 68576
rect 4360 68512 4376 68576
rect 4440 68512 4456 68576
rect 4520 68512 4528 68576
rect 4208 68511 4528 68512
rect 34928 68576 35248 68577
rect 34928 68512 34936 68576
rect 35000 68512 35016 68576
rect 35080 68512 35096 68576
rect 35160 68512 35176 68576
rect 35240 68512 35248 68576
rect 34928 68511 35248 68512
rect 12341 68370 12407 68373
rect 20713 68370 20779 68373
rect 12341 68368 20779 68370
rect 12341 68312 12346 68368
rect 12402 68312 20718 68368
rect 20774 68312 20779 68368
rect 12341 68310 20779 68312
rect 12341 68307 12407 68310
rect 20713 68307 20779 68310
rect 28942 68308 28948 68372
rect 29012 68370 29018 68372
rect 29012 68310 39130 68370
rect 29012 68308 29018 68310
rect 3325 68234 3391 68237
rect 24301 68234 24367 68237
rect 3325 68232 24367 68234
rect 3325 68176 3330 68232
rect 3386 68176 24306 68232
rect 24362 68176 24367 68232
rect 3325 68174 24367 68176
rect 3325 68171 3391 68174
rect 24301 68171 24367 68174
rect 25313 68234 25379 68237
rect 37365 68234 37431 68237
rect 25313 68232 37431 68234
rect 25313 68176 25318 68232
rect 25374 68176 37370 68232
rect 37426 68176 37431 68232
rect 25313 68174 37431 68176
rect 25313 68171 25379 68174
rect 37365 68171 37431 68174
rect 0 68098 800 68128
rect 3417 68098 3483 68101
rect 0 68096 3483 68098
rect 0 68040 3422 68096
rect 3478 68040 3483 68096
rect 0 68038 3483 68040
rect 39070 68098 39130 68310
rect 39200 68098 40000 68128
rect 39070 68038 40000 68098
rect 0 68008 800 68038
rect 3417 68035 3483 68038
rect 19568 68032 19888 68033
rect 19568 67968 19576 68032
rect 19640 67968 19656 68032
rect 19720 67968 19736 68032
rect 19800 67968 19816 68032
rect 19880 67968 19888 68032
rect 39200 68008 40000 68038
rect 19568 67967 19888 67968
rect 20897 67962 20963 67965
rect 28942 67962 28948 67964
rect 20897 67960 28948 67962
rect 20897 67904 20902 67960
rect 20958 67904 28948 67960
rect 20897 67902 28948 67904
rect 20897 67899 20963 67902
rect 28942 67900 28948 67902
rect 29012 67900 29018 67964
rect 12617 67826 12683 67829
rect 19333 67826 19399 67829
rect 12617 67824 19399 67826
rect 12617 67768 12622 67824
rect 12678 67768 19338 67824
rect 19394 67768 19399 67824
rect 12617 67766 19399 67768
rect 12617 67763 12683 67766
rect 19333 67763 19399 67766
rect 8385 67690 8451 67693
rect 11237 67690 11303 67693
rect 8385 67688 11303 67690
rect 8385 67632 8390 67688
rect 8446 67632 11242 67688
rect 11298 67632 11303 67688
rect 8385 67630 11303 67632
rect 8385 67627 8451 67630
rect 11237 67627 11303 67630
rect 21357 67554 21423 67557
rect 22185 67554 22251 67557
rect 21357 67552 22251 67554
rect 21357 67496 21362 67552
rect 21418 67496 22190 67552
rect 22246 67496 22251 67552
rect 21357 67494 22251 67496
rect 21357 67491 21423 67494
rect 22185 67491 22251 67494
rect 4208 67488 4528 67489
rect 4208 67424 4216 67488
rect 4280 67424 4296 67488
rect 4360 67424 4376 67488
rect 4440 67424 4456 67488
rect 4520 67424 4528 67488
rect 4208 67423 4528 67424
rect 34928 67488 35248 67489
rect 34928 67424 34936 67488
rect 35000 67424 35016 67488
rect 35080 67424 35096 67488
rect 35160 67424 35176 67488
rect 35240 67424 35248 67488
rect 34928 67423 35248 67424
rect 10869 67282 10935 67285
rect 27245 67282 27311 67285
rect 10869 67280 27311 67282
rect 10869 67224 10874 67280
rect 10930 67224 27250 67280
rect 27306 67224 27311 67280
rect 10869 67222 27311 67224
rect 10869 67219 10935 67222
rect 27245 67219 27311 67222
rect 3969 67146 4035 67149
rect 28390 67146 28396 67148
rect 3969 67144 28396 67146
rect 3969 67088 3974 67144
rect 4030 67088 28396 67144
rect 3969 67086 28396 67088
rect 3969 67083 4035 67086
rect 28390 67084 28396 67086
rect 28460 67084 28466 67148
rect 19568 66944 19888 66945
rect 19568 66880 19576 66944
rect 19640 66880 19656 66944
rect 19720 66880 19736 66944
rect 19800 66880 19816 66944
rect 19880 66880 19888 66944
rect 19568 66879 19888 66880
rect 0 66738 800 66768
rect 1577 66738 1643 66741
rect 0 66736 1643 66738
rect 0 66680 1582 66736
rect 1638 66680 1643 66736
rect 0 66678 1643 66680
rect 0 66648 800 66678
rect 1577 66675 1643 66678
rect 22277 66738 22343 66741
rect 39200 66738 40000 66768
rect 22277 66736 40000 66738
rect 22277 66680 22282 66736
rect 22338 66680 40000 66736
rect 22277 66678 40000 66680
rect 22277 66675 22343 66678
rect 39200 66648 40000 66678
rect 4208 66400 4528 66401
rect 4208 66336 4216 66400
rect 4280 66336 4296 66400
rect 4360 66336 4376 66400
rect 4440 66336 4456 66400
rect 4520 66336 4528 66400
rect 4208 66335 4528 66336
rect 34928 66400 35248 66401
rect 34928 66336 34936 66400
rect 35000 66336 35016 66400
rect 35080 66336 35096 66400
rect 35160 66336 35176 66400
rect 35240 66336 35248 66400
rect 34928 66335 35248 66336
rect 19568 65856 19888 65857
rect 19568 65792 19576 65856
rect 19640 65792 19656 65856
rect 19720 65792 19736 65856
rect 19800 65792 19816 65856
rect 19880 65792 19888 65856
rect 19568 65791 19888 65792
rect 14089 65514 14155 65517
rect 26325 65514 26391 65517
rect 14089 65512 26391 65514
rect 14089 65456 14094 65512
rect 14150 65456 26330 65512
rect 26386 65456 26391 65512
rect 14089 65454 26391 65456
rect 14089 65451 14155 65454
rect 26325 65451 26391 65454
rect 0 65378 800 65408
rect 2865 65378 2931 65381
rect 0 65376 2931 65378
rect 0 65320 2870 65376
rect 2926 65320 2931 65376
rect 0 65318 2931 65320
rect 0 65288 800 65318
rect 2865 65315 2931 65318
rect 35433 65378 35499 65381
rect 39200 65378 40000 65408
rect 35433 65376 40000 65378
rect 35433 65320 35438 65376
rect 35494 65320 40000 65376
rect 35433 65318 40000 65320
rect 35433 65315 35499 65318
rect 4208 65312 4528 65313
rect 4208 65248 4216 65312
rect 4280 65248 4296 65312
rect 4360 65248 4376 65312
rect 4440 65248 4456 65312
rect 4520 65248 4528 65312
rect 4208 65247 4528 65248
rect 34928 65312 35248 65313
rect 34928 65248 34936 65312
rect 35000 65248 35016 65312
rect 35080 65248 35096 65312
rect 35160 65248 35176 65312
rect 35240 65248 35248 65312
rect 39200 65288 40000 65318
rect 34928 65247 35248 65248
rect 19568 64768 19888 64769
rect 19568 64704 19576 64768
rect 19640 64704 19656 64768
rect 19720 64704 19736 64768
rect 19800 64704 19816 64768
rect 19880 64704 19888 64768
rect 19568 64703 19888 64704
rect 4208 64224 4528 64225
rect 4208 64160 4216 64224
rect 4280 64160 4296 64224
rect 4360 64160 4376 64224
rect 4440 64160 4456 64224
rect 4520 64160 4528 64224
rect 4208 64159 4528 64160
rect 34928 64224 35248 64225
rect 34928 64160 34936 64224
rect 35000 64160 35016 64224
rect 35080 64160 35096 64224
rect 35160 64160 35176 64224
rect 35240 64160 35248 64224
rect 34928 64159 35248 64160
rect 15837 64154 15903 64157
rect 25773 64154 25839 64157
rect 15837 64152 25839 64154
rect 15837 64096 15842 64152
rect 15898 64096 25778 64152
rect 25834 64096 25839 64152
rect 15837 64094 25839 64096
rect 15837 64091 15903 64094
rect 25773 64091 25839 64094
rect 0 64018 800 64048
rect 1853 64018 1919 64021
rect 0 64016 1919 64018
rect 0 63960 1858 64016
rect 1914 63960 1919 64016
rect 0 63958 1919 63960
rect 0 63928 800 63958
rect 1853 63955 1919 63958
rect 4153 64018 4219 64021
rect 27153 64018 27219 64021
rect 39200 64018 40000 64048
rect 4153 64016 27219 64018
rect 4153 63960 4158 64016
rect 4214 63960 27158 64016
rect 27214 63960 27219 64016
rect 4153 63958 27219 63960
rect 4153 63955 4219 63958
rect 27153 63955 27219 63958
rect 39070 63958 40000 64018
rect 14549 63882 14615 63885
rect 39070 63882 39130 63958
rect 39200 63928 40000 63958
rect 14549 63880 39130 63882
rect 14549 63824 14554 63880
rect 14610 63824 39130 63880
rect 14549 63822 39130 63824
rect 14549 63819 14615 63822
rect 19568 63680 19888 63681
rect 19568 63616 19576 63680
rect 19640 63616 19656 63680
rect 19720 63616 19736 63680
rect 19800 63616 19816 63680
rect 19880 63616 19888 63680
rect 19568 63615 19888 63616
rect 15929 63474 15995 63477
rect 21725 63474 21791 63477
rect 15929 63472 21791 63474
rect 15929 63416 15934 63472
rect 15990 63416 21730 63472
rect 21786 63416 21791 63472
rect 15929 63414 21791 63416
rect 15929 63411 15995 63414
rect 21725 63411 21791 63414
rect 4208 63136 4528 63137
rect 4208 63072 4216 63136
rect 4280 63072 4296 63136
rect 4360 63072 4376 63136
rect 4440 63072 4456 63136
rect 4520 63072 4528 63136
rect 4208 63071 4528 63072
rect 34928 63136 35248 63137
rect 34928 63072 34936 63136
rect 35000 63072 35016 63136
rect 35080 63072 35096 63136
rect 35160 63072 35176 63136
rect 35240 63072 35248 63136
rect 34928 63071 35248 63072
rect 22502 62732 22508 62796
rect 22572 62794 22578 62796
rect 35525 62794 35591 62797
rect 22572 62792 35591 62794
rect 22572 62736 35530 62792
rect 35586 62736 35591 62792
rect 22572 62734 35591 62736
rect 22572 62732 22578 62734
rect 35525 62731 35591 62734
rect 0 62658 800 62688
rect 31201 62658 31267 62661
rect 39200 62658 40000 62688
rect 0 62568 858 62658
rect 31201 62656 40000 62658
rect 31201 62600 31206 62656
rect 31262 62600 40000 62656
rect 31201 62598 40000 62600
rect 31201 62595 31267 62598
rect 798 62386 858 62568
rect 19568 62592 19888 62593
rect 19568 62528 19576 62592
rect 19640 62528 19656 62592
rect 19720 62528 19736 62592
rect 19800 62528 19816 62592
rect 19880 62528 19888 62592
rect 39200 62568 40000 62598
rect 19568 62527 19888 62528
rect 20621 62386 20687 62389
rect 798 62384 20687 62386
rect 798 62328 20626 62384
rect 20682 62328 20687 62384
rect 798 62326 20687 62328
rect 20621 62323 20687 62326
rect 7373 62250 7439 62253
rect 19057 62250 19123 62253
rect 7373 62248 19123 62250
rect 7373 62192 7378 62248
rect 7434 62192 19062 62248
rect 19118 62192 19123 62248
rect 7373 62190 19123 62192
rect 7373 62187 7439 62190
rect 19057 62187 19123 62190
rect 19977 62250 20043 62253
rect 22461 62250 22527 62253
rect 19977 62248 22527 62250
rect 19977 62192 19982 62248
rect 20038 62192 22466 62248
rect 22522 62192 22527 62248
rect 19977 62190 22527 62192
rect 19977 62187 20043 62190
rect 22461 62187 22527 62190
rect 28022 62188 28028 62252
rect 28092 62250 28098 62252
rect 35433 62250 35499 62253
rect 28092 62248 35499 62250
rect 28092 62192 35438 62248
rect 35494 62192 35499 62248
rect 28092 62190 35499 62192
rect 28092 62188 28098 62190
rect 35433 62187 35499 62190
rect 5165 62114 5231 62117
rect 10777 62114 10843 62117
rect 5165 62112 10843 62114
rect 5165 62056 5170 62112
rect 5226 62056 10782 62112
rect 10838 62056 10843 62112
rect 5165 62054 10843 62056
rect 5165 62051 5231 62054
rect 10777 62051 10843 62054
rect 18413 62114 18479 62117
rect 22001 62114 22067 62117
rect 18413 62112 22067 62114
rect 18413 62056 18418 62112
rect 18474 62056 22006 62112
rect 22062 62056 22067 62112
rect 18413 62054 22067 62056
rect 18413 62051 18479 62054
rect 22001 62051 22067 62054
rect 29085 62114 29151 62117
rect 31017 62114 31083 62117
rect 29085 62112 31083 62114
rect 29085 62056 29090 62112
rect 29146 62056 31022 62112
rect 31078 62056 31083 62112
rect 29085 62054 31083 62056
rect 29085 62051 29151 62054
rect 31017 62051 31083 62054
rect 4208 62048 4528 62049
rect 4208 61984 4216 62048
rect 4280 61984 4296 62048
rect 4360 61984 4376 62048
rect 4440 61984 4456 62048
rect 4520 61984 4528 62048
rect 4208 61983 4528 61984
rect 34928 62048 35248 62049
rect 34928 61984 34936 62048
rect 35000 61984 35016 62048
rect 35080 61984 35096 62048
rect 35160 61984 35176 62048
rect 35240 61984 35248 62048
rect 34928 61983 35248 61984
rect 10961 61570 11027 61573
rect 13169 61570 13235 61573
rect 13813 61570 13879 61573
rect 10961 61568 13879 61570
rect 10961 61512 10966 61568
rect 11022 61512 13174 61568
rect 13230 61512 13818 61568
rect 13874 61512 13879 61568
rect 10961 61510 13879 61512
rect 10961 61507 11027 61510
rect 13169 61507 13235 61510
rect 13813 61507 13879 61510
rect 19568 61504 19888 61505
rect 19568 61440 19576 61504
rect 19640 61440 19656 61504
rect 19720 61440 19736 61504
rect 19800 61440 19816 61504
rect 19880 61440 19888 61504
rect 19568 61439 19888 61440
rect 23381 61434 23447 61437
rect 35617 61434 35683 61437
rect 23381 61432 35683 61434
rect 23381 61376 23386 61432
rect 23442 61376 35622 61432
rect 35678 61376 35683 61432
rect 23381 61374 35683 61376
rect 23381 61371 23447 61374
rect 35617 61371 35683 61374
rect 0 61298 800 61328
rect 24945 61298 25011 61301
rect 0 61296 25011 61298
rect 0 61240 24950 61296
rect 25006 61240 25011 61296
rect 0 61238 25011 61240
rect 0 61208 800 61238
rect 24945 61235 25011 61238
rect 35433 61298 35499 61301
rect 39200 61298 40000 61328
rect 35433 61296 40000 61298
rect 35433 61240 35438 61296
rect 35494 61240 40000 61296
rect 35433 61238 40000 61240
rect 35433 61235 35499 61238
rect 39200 61208 40000 61238
rect 29269 61162 29335 61165
rect 35801 61162 35867 61165
rect 29269 61160 35867 61162
rect 29269 61104 29274 61160
rect 29330 61104 35806 61160
rect 35862 61104 35867 61160
rect 29269 61102 35867 61104
rect 29269 61099 29335 61102
rect 35801 61099 35867 61102
rect 4208 60960 4528 60961
rect 4208 60896 4216 60960
rect 4280 60896 4296 60960
rect 4360 60896 4376 60960
rect 4440 60896 4456 60960
rect 4520 60896 4528 60960
rect 4208 60895 4528 60896
rect 34928 60960 35248 60961
rect 34928 60896 34936 60960
rect 35000 60896 35016 60960
rect 35080 60896 35096 60960
rect 35160 60896 35176 60960
rect 35240 60896 35248 60960
rect 34928 60895 35248 60896
rect 3417 60618 3483 60621
rect 9213 60618 9279 60621
rect 3417 60616 9279 60618
rect 3417 60560 3422 60616
rect 3478 60560 9218 60616
rect 9274 60560 9279 60616
rect 3417 60558 9279 60560
rect 3417 60555 3483 60558
rect 9213 60555 9279 60558
rect 25313 60618 25379 60621
rect 26233 60618 26299 60621
rect 29913 60618 29979 60621
rect 25313 60616 29979 60618
rect 25313 60560 25318 60616
rect 25374 60560 26238 60616
rect 26294 60560 29918 60616
rect 29974 60560 29979 60616
rect 25313 60558 29979 60560
rect 25313 60555 25379 60558
rect 26233 60555 26299 60558
rect 29913 60555 29979 60558
rect 19568 60416 19888 60417
rect 19568 60352 19576 60416
rect 19640 60352 19656 60416
rect 19720 60352 19736 60416
rect 19800 60352 19816 60416
rect 19880 60352 19888 60416
rect 19568 60351 19888 60352
rect 22001 60346 22067 60349
rect 23841 60346 23907 60349
rect 22001 60344 23907 60346
rect 22001 60288 22006 60344
rect 22062 60288 23846 60344
rect 23902 60288 23907 60344
rect 22001 60286 23907 60288
rect 22001 60283 22067 60286
rect 23841 60283 23907 60286
rect 27061 60346 27127 60349
rect 29545 60346 29611 60349
rect 31385 60346 31451 60349
rect 27061 60344 31451 60346
rect 27061 60288 27066 60344
rect 27122 60288 29550 60344
rect 29606 60288 31390 60344
rect 31446 60288 31451 60344
rect 27061 60286 31451 60288
rect 27061 60283 27127 60286
rect 29545 60283 29611 60286
rect 31385 60283 31451 60286
rect 30373 60074 30439 60077
rect 30373 60072 35588 60074
rect 30373 60016 30378 60072
rect 30434 60016 35588 60072
rect 30373 60014 35588 60016
rect 30373 60011 30439 60014
rect 0 59938 800 59968
rect 1853 59938 1919 59941
rect 0 59936 1919 59938
rect 0 59880 1858 59936
rect 1914 59880 1919 59936
rect 0 59878 1919 59880
rect 0 59848 800 59878
rect 1853 59875 1919 59878
rect 4889 59938 4955 59941
rect 10501 59938 10567 59941
rect 4889 59936 10567 59938
rect 4889 59880 4894 59936
rect 4950 59880 10506 59936
rect 10562 59880 10567 59936
rect 4889 59878 10567 59880
rect 35528 59938 35588 60014
rect 39200 59938 40000 59968
rect 35528 59878 40000 59938
rect 4889 59875 4955 59878
rect 10501 59875 10567 59878
rect 4208 59872 4528 59873
rect 4208 59808 4216 59872
rect 4280 59808 4296 59872
rect 4360 59808 4376 59872
rect 4440 59808 4456 59872
rect 4520 59808 4528 59872
rect 4208 59807 4528 59808
rect 34928 59872 35248 59873
rect 34928 59808 34936 59872
rect 35000 59808 35016 59872
rect 35080 59808 35096 59872
rect 35160 59808 35176 59872
rect 35240 59808 35248 59872
rect 39200 59848 40000 59878
rect 34928 59807 35248 59808
rect 17861 59802 17927 59805
rect 20621 59802 20687 59805
rect 22369 59802 22435 59805
rect 22553 59802 22619 59805
rect 17861 59800 22619 59802
rect 17861 59744 17866 59800
rect 17922 59744 20626 59800
rect 20682 59744 22374 59800
rect 22430 59744 22558 59800
rect 22614 59744 22619 59800
rect 17861 59742 22619 59744
rect 17861 59739 17927 59742
rect 20621 59739 20687 59742
rect 22369 59739 22435 59742
rect 22553 59739 22619 59742
rect 20161 59666 20227 59669
rect 22093 59666 22159 59669
rect 20161 59664 22159 59666
rect 20161 59608 20166 59664
rect 20222 59608 22098 59664
rect 22154 59608 22159 59664
rect 20161 59606 22159 59608
rect 20161 59603 20227 59606
rect 22093 59603 22159 59606
rect 18597 59530 18663 59533
rect 21541 59530 21607 59533
rect 18597 59528 21607 59530
rect 18597 59472 18602 59528
rect 18658 59472 21546 59528
rect 21602 59472 21607 59528
rect 18597 59470 21607 59472
rect 18597 59467 18663 59470
rect 21541 59467 21607 59470
rect 16481 59394 16547 59397
rect 17953 59394 18019 59397
rect 16481 59392 18019 59394
rect 16481 59336 16486 59392
rect 16542 59336 17958 59392
rect 18014 59336 18019 59392
rect 16481 59334 18019 59336
rect 16481 59331 16547 59334
rect 17953 59331 18019 59334
rect 23933 59394 23999 59397
rect 25037 59394 25103 59397
rect 23933 59392 25103 59394
rect 23933 59336 23938 59392
rect 23994 59336 25042 59392
rect 25098 59336 25103 59392
rect 23933 59334 25103 59336
rect 23933 59331 23999 59334
rect 25037 59331 25103 59334
rect 29821 59394 29887 59397
rect 37365 59394 37431 59397
rect 29821 59392 37431 59394
rect 29821 59336 29826 59392
rect 29882 59336 37370 59392
rect 37426 59336 37431 59392
rect 29821 59334 37431 59336
rect 29821 59331 29887 59334
rect 37365 59331 37431 59334
rect 19568 59328 19888 59329
rect 19568 59264 19576 59328
rect 19640 59264 19656 59328
rect 19720 59264 19736 59328
rect 19800 59264 19816 59328
rect 19880 59264 19888 59328
rect 19568 59263 19888 59264
rect 19241 59122 19307 59125
rect 20897 59122 20963 59125
rect 19241 59120 20963 59122
rect 19241 59064 19246 59120
rect 19302 59064 20902 59120
rect 20958 59064 20963 59120
rect 19241 59062 20963 59064
rect 19241 59059 19307 59062
rect 20897 59059 20963 59062
rect 23381 58986 23447 58989
rect 32949 58986 33015 58989
rect 23381 58984 33015 58986
rect 23381 58928 23386 58984
rect 23442 58928 32954 58984
rect 33010 58928 33015 58984
rect 23381 58926 33015 58928
rect 23381 58923 23447 58926
rect 32949 58923 33015 58926
rect 4208 58784 4528 58785
rect 4208 58720 4216 58784
rect 4280 58720 4296 58784
rect 4360 58720 4376 58784
rect 4440 58720 4456 58784
rect 4520 58720 4528 58784
rect 4208 58719 4528 58720
rect 34928 58784 35248 58785
rect 34928 58720 34936 58784
rect 35000 58720 35016 58784
rect 35080 58720 35096 58784
rect 35160 58720 35176 58784
rect 35240 58720 35248 58784
rect 34928 58719 35248 58720
rect 0 58578 800 58608
rect 35341 58578 35407 58581
rect 39200 58578 40000 58608
rect 0 58488 858 58578
rect 35341 58576 40000 58578
rect 35341 58520 35346 58576
rect 35402 58520 40000 58576
rect 35341 58518 40000 58520
rect 35341 58515 35407 58518
rect 39200 58488 40000 58518
rect 798 58442 858 58488
rect 27705 58442 27771 58445
rect 798 58440 27771 58442
rect 798 58384 27710 58440
rect 27766 58384 27771 58440
rect 798 58382 27771 58384
rect 27705 58379 27771 58382
rect 21449 58306 21515 58309
rect 24485 58306 24551 58309
rect 21449 58304 24551 58306
rect 21449 58248 21454 58304
rect 21510 58248 24490 58304
rect 24546 58248 24551 58304
rect 21449 58246 24551 58248
rect 21449 58243 21515 58246
rect 24485 58243 24551 58246
rect 19568 58240 19888 58241
rect 19568 58176 19576 58240
rect 19640 58176 19656 58240
rect 19720 58176 19736 58240
rect 19800 58176 19816 58240
rect 19880 58176 19888 58240
rect 19568 58175 19888 58176
rect 22829 58170 22895 58173
rect 22694 58168 22895 58170
rect 22694 58112 22834 58168
rect 22890 58112 22895 58168
rect 22694 58110 22895 58112
rect 22694 58037 22754 58110
rect 22829 58107 22895 58110
rect 13353 58034 13419 58037
rect 18321 58034 18387 58037
rect 13353 58032 18387 58034
rect 13353 57976 13358 58032
rect 13414 57976 18326 58032
rect 18382 57976 18387 58032
rect 13353 57974 18387 57976
rect 13353 57971 13419 57974
rect 18321 57971 18387 57974
rect 22645 58032 22754 58037
rect 22645 57976 22650 58032
rect 22706 57976 22754 58032
rect 22645 57974 22754 57976
rect 22645 57971 22711 57974
rect 0 57898 800 57928
rect 21633 57898 21699 57901
rect 24301 57898 24367 57901
rect 0 57808 858 57898
rect 21633 57896 24367 57898
rect 21633 57840 21638 57896
rect 21694 57840 24306 57896
rect 24362 57840 24367 57896
rect 21633 57838 24367 57840
rect 21633 57835 21699 57838
rect 24301 57835 24367 57838
rect 798 57354 858 57808
rect 17125 57762 17191 57765
rect 19609 57762 19675 57765
rect 17125 57760 19675 57762
rect 17125 57704 17130 57760
rect 17186 57704 19614 57760
rect 19670 57704 19675 57760
rect 17125 57702 19675 57704
rect 17125 57699 17191 57702
rect 19609 57699 19675 57702
rect 4208 57696 4528 57697
rect 4208 57632 4216 57696
rect 4280 57632 4296 57696
rect 4360 57632 4376 57696
rect 4440 57632 4456 57696
rect 4520 57632 4528 57696
rect 4208 57631 4528 57632
rect 34928 57696 35248 57697
rect 34928 57632 34936 57696
rect 35000 57632 35016 57696
rect 35080 57632 35096 57696
rect 35160 57632 35176 57696
rect 35240 57632 35248 57696
rect 34928 57631 35248 57632
rect 10777 57626 10843 57629
rect 14273 57626 14339 57629
rect 10777 57624 14339 57626
rect 10777 57568 10782 57624
rect 10838 57568 14278 57624
rect 14334 57568 14339 57624
rect 10777 57566 14339 57568
rect 10777 57563 10843 57566
rect 14273 57563 14339 57566
rect 28073 57626 28139 57629
rect 28993 57626 29059 57629
rect 28073 57624 29059 57626
rect 28073 57568 28078 57624
rect 28134 57568 28998 57624
rect 29054 57568 29059 57624
rect 28073 57566 29059 57568
rect 28073 57563 28139 57566
rect 28993 57563 29059 57566
rect 15009 57354 15075 57357
rect 798 57352 15075 57354
rect 798 57296 15014 57352
rect 15070 57296 15075 57352
rect 798 57294 15075 57296
rect 15009 57291 15075 57294
rect 34513 57218 34579 57221
rect 39200 57218 40000 57248
rect 34513 57216 40000 57218
rect 34513 57160 34518 57216
rect 34574 57160 40000 57216
rect 34513 57158 40000 57160
rect 34513 57155 34579 57158
rect 19568 57152 19888 57153
rect 19568 57088 19576 57152
rect 19640 57088 19656 57152
rect 19720 57088 19736 57152
rect 19800 57088 19816 57152
rect 19880 57088 19888 57152
rect 39200 57128 40000 57158
rect 19568 57087 19888 57088
rect 14365 56810 14431 56813
rect 17861 56810 17927 56813
rect 14365 56808 17927 56810
rect 14365 56752 14370 56808
rect 14426 56752 17866 56808
rect 17922 56752 17927 56808
rect 14365 56750 17927 56752
rect 14365 56747 14431 56750
rect 17861 56747 17927 56750
rect 18137 56810 18203 56813
rect 21357 56810 21423 56813
rect 18137 56808 21423 56810
rect 18137 56752 18142 56808
rect 18198 56752 21362 56808
rect 21418 56752 21423 56808
rect 18137 56750 21423 56752
rect 18137 56747 18203 56750
rect 21357 56747 21423 56750
rect 24393 56810 24459 56813
rect 35433 56810 35499 56813
rect 24393 56808 35499 56810
rect 24393 56752 24398 56808
rect 24454 56752 35438 56808
rect 35494 56752 35499 56808
rect 24393 56750 35499 56752
rect 24393 56747 24459 56750
rect 35433 56747 35499 56750
rect 13261 56674 13327 56677
rect 19517 56674 19583 56677
rect 13261 56672 19583 56674
rect 13261 56616 13266 56672
rect 13322 56616 19522 56672
rect 19578 56616 19583 56672
rect 13261 56614 19583 56616
rect 13261 56611 13327 56614
rect 19517 56611 19583 56614
rect 21449 56674 21515 56677
rect 21909 56674 21975 56677
rect 25497 56674 25563 56677
rect 21449 56672 21834 56674
rect 21449 56616 21454 56672
rect 21510 56616 21834 56672
rect 21449 56614 21834 56616
rect 21449 56611 21515 56614
rect 4208 56608 4528 56609
rect 0 56538 800 56568
rect 4208 56544 4216 56608
rect 4280 56544 4296 56608
rect 4360 56544 4376 56608
rect 4440 56544 4456 56608
rect 4520 56544 4528 56608
rect 4208 56543 4528 56544
rect 17861 56538 17927 56541
rect 21541 56538 21607 56541
rect 0 56478 3250 56538
rect 0 56448 800 56478
rect 3190 55722 3250 56478
rect 17861 56536 21607 56538
rect 17861 56480 17866 56536
rect 17922 56480 21546 56536
rect 21602 56480 21607 56536
rect 17861 56478 21607 56480
rect 21774 56538 21834 56614
rect 21909 56672 25563 56674
rect 21909 56616 21914 56672
rect 21970 56616 25502 56672
rect 25558 56616 25563 56672
rect 21909 56614 25563 56616
rect 21909 56611 21975 56614
rect 25497 56611 25563 56614
rect 34928 56608 35248 56609
rect 34928 56544 34936 56608
rect 35000 56544 35016 56608
rect 35080 56544 35096 56608
rect 35160 56544 35176 56608
rect 35240 56544 35248 56608
rect 34928 56543 35248 56544
rect 25313 56538 25379 56541
rect 21774 56536 25379 56538
rect 21774 56480 25318 56536
rect 25374 56480 25379 56536
rect 21774 56478 25379 56480
rect 17861 56475 17927 56478
rect 21541 56475 21607 56478
rect 25313 56475 25379 56478
rect 30649 56538 30715 56541
rect 31753 56538 31819 56541
rect 30649 56536 31819 56538
rect 30649 56480 30654 56536
rect 30710 56480 31758 56536
rect 31814 56480 31819 56536
rect 30649 56478 31819 56480
rect 30649 56475 30715 56478
rect 31753 56475 31819 56478
rect 35525 56538 35591 56541
rect 39200 56538 40000 56568
rect 35525 56536 40000 56538
rect 35525 56480 35530 56536
rect 35586 56480 40000 56536
rect 35525 56478 40000 56480
rect 35525 56475 35591 56478
rect 39200 56448 40000 56478
rect 3877 56402 3943 56405
rect 14181 56402 14247 56405
rect 3877 56400 14247 56402
rect 3877 56344 3882 56400
rect 3938 56344 14186 56400
rect 14242 56344 14247 56400
rect 3877 56342 14247 56344
rect 3877 56339 3943 56342
rect 14181 56339 14247 56342
rect 17769 56402 17835 56405
rect 19609 56402 19675 56405
rect 17769 56400 19675 56402
rect 17769 56344 17774 56400
rect 17830 56344 19614 56400
rect 19670 56344 19675 56400
rect 17769 56342 19675 56344
rect 17769 56339 17835 56342
rect 19609 56339 19675 56342
rect 19885 56402 19951 56405
rect 23657 56402 23723 56405
rect 19885 56400 23723 56402
rect 19885 56344 19890 56400
rect 19946 56344 23662 56400
rect 23718 56344 23723 56400
rect 19885 56342 23723 56344
rect 19885 56339 19951 56342
rect 23657 56339 23723 56342
rect 26049 56402 26115 56405
rect 29729 56402 29795 56405
rect 26049 56400 29795 56402
rect 26049 56344 26054 56400
rect 26110 56344 29734 56400
rect 29790 56344 29795 56400
rect 26049 56342 29795 56344
rect 26049 56339 26115 56342
rect 29729 56339 29795 56342
rect 16665 56266 16731 56269
rect 20897 56266 20963 56269
rect 16665 56264 20963 56266
rect 16665 56208 16670 56264
rect 16726 56208 20902 56264
rect 20958 56208 20963 56264
rect 16665 56206 20963 56208
rect 16665 56203 16731 56206
rect 20897 56203 20963 56206
rect 19977 56130 20043 56133
rect 24485 56130 24551 56133
rect 19977 56128 24551 56130
rect 19977 56072 19982 56128
rect 20038 56072 24490 56128
rect 24546 56072 24551 56128
rect 19977 56070 24551 56072
rect 19977 56067 20043 56070
rect 24485 56067 24551 56070
rect 19568 56064 19888 56065
rect 19568 56000 19576 56064
rect 19640 56000 19656 56064
rect 19720 56000 19736 56064
rect 19800 56000 19816 56064
rect 19880 56000 19888 56064
rect 19568 55999 19888 56000
rect 14641 55994 14707 55997
rect 18413 55994 18479 55997
rect 14641 55992 18479 55994
rect 14641 55936 14646 55992
rect 14702 55936 18418 55992
rect 18474 55936 18479 55992
rect 14641 55934 18479 55936
rect 14641 55931 14707 55934
rect 18413 55931 18479 55934
rect 22093 55994 22159 55997
rect 23013 55994 23079 55997
rect 22093 55992 23079 55994
rect 22093 55936 22098 55992
rect 22154 55936 23018 55992
rect 23074 55936 23079 55992
rect 22093 55934 23079 55936
rect 22093 55931 22159 55934
rect 23013 55931 23079 55934
rect 16849 55858 16915 55861
rect 26509 55858 26575 55861
rect 16849 55856 26575 55858
rect 16849 55800 16854 55856
rect 16910 55800 26514 55856
rect 26570 55800 26575 55856
rect 16849 55798 26575 55800
rect 16849 55795 16915 55798
rect 26509 55795 26575 55798
rect 15469 55722 15535 55725
rect 3190 55720 15535 55722
rect 3190 55664 15474 55720
rect 15530 55664 15535 55720
rect 3190 55662 15535 55664
rect 15469 55659 15535 55662
rect 17217 55722 17283 55725
rect 21449 55722 21515 55725
rect 17217 55720 21515 55722
rect 17217 55664 17222 55720
rect 17278 55664 21454 55720
rect 21510 55664 21515 55720
rect 17217 55662 21515 55664
rect 17217 55659 17283 55662
rect 21449 55659 21515 55662
rect 22461 55722 22527 55725
rect 24669 55722 24735 55725
rect 22461 55720 24735 55722
rect 22461 55664 22466 55720
rect 22522 55664 24674 55720
rect 24730 55664 24735 55720
rect 22461 55662 24735 55664
rect 22461 55659 22527 55662
rect 24669 55659 24735 55662
rect 16297 55586 16363 55589
rect 20713 55586 20779 55589
rect 16297 55584 20779 55586
rect 16297 55528 16302 55584
rect 16358 55528 20718 55584
rect 20774 55528 20779 55584
rect 16297 55526 20779 55528
rect 16297 55523 16363 55526
rect 20713 55523 20779 55526
rect 4208 55520 4528 55521
rect 4208 55456 4216 55520
rect 4280 55456 4296 55520
rect 4360 55456 4376 55520
rect 4440 55456 4456 55520
rect 4520 55456 4528 55520
rect 4208 55455 4528 55456
rect 34928 55520 35248 55521
rect 34928 55456 34936 55520
rect 35000 55456 35016 55520
rect 35080 55456 35096 55520
rect 35160 55456 35176 55520
rect 35240 55456 35248 55520
rect 34928 55455 35248 55456
rect 12249 55450 12315 55453
rect 17217 55450 17283 55453
rect 12249 55448 17283 55450
rect 12249 55392 12254 55448
rect 12310 55392 17222 55448
rect 17278 55392 17283 55448
rect 12249 55390 17283 55392
rect 12249 55387 12315 55390
rect 17217 55387 17283 55390
rect 18965 55450 19031 55453
rect 19977 55450 20043 55453
rect 18965 55448 20043 55450
rect 18965 55392 18970 55448
rect 19026 55392 19982 55448
rect 20038 55392 20043 55448
rect 18965 55390 20043 55392
rect 18965 55387 19031 55390
rect 19977 55387 20043 55390
rect 20253 55450 20319 55453
rect 27981 55450 28047 55453
rect 20253 55448 28047 55450
rect 20253 55392 20258 55448
rect 20314 55392 27986 55448
rect 28042 55392 28047 55448
rect 20253 55390 28047 55392
rect 20253 55387 20319 55390
rect 27981 55387 28047 55390
rect 14273 55314 14339 55317
rect 19425 55314 19491 55317
rect 14273 55312 19491 55314
rect 14273 55256 14278 55312
rect 14334 55256 19430 55312
rect 19486 55256 19491 55312
rect 14273 55254 19491 55256
rect 14273 55251 14339 55254
rect 19425 55251 19491 55254
rect 26325 55314 26391 55317
rect 31569 55314 31635 55317
rect 26325 55312 31635 55314
rect 26325 55256 26330 55312
rect 26386 55256 31574 55312
rect 31630 55256 31635 55312
rect 26325 55254 31635 55256
rect 26325 55251 26391 55254
rect 31569 55251 31635 55254
rect 0 55178 800 55208
rect 3325 55178 3391 55181
rect 0 55176 3391 55178
rect 0 55120 3330 55176
rect 3386 55120 3391 55176
rect 0 55118 3391 55120
rect 0 55088 800 55118
rect 3325 55115 3391 55118
rect 13445 55178 13511 55181
rect 16573 55178 16639 55181
rect 13445 55176 16639 55178
rect 13445 55120 13450 55176
rect 13506 55120 16578 55176
rect 16634 55120 16639 55176
rect 13445 55118 16639 55120
rect 13445 55115 13511 55118
rect 16573 55115 16639 55118
rect 19609 55178 19675 55181
rect 21357 55178 21423 55181
rect 19609 55176 21423 55178
rect 19609 55120 19614 55176
rect 19670 55120 21362 55176
rect 21418 55120 21423 55176
rect 19609 55118 21423 55120
rect 19609 55115 19675 55118
rect 21357 55115 21423 55118
rect 35433 55178 35499 55181
rect 39200 55178 40000 55208
rect 35433 55176 40000 55178
rect 35433 55120 35438 55176
rect 35494 55120 40000 55176
rect 35433 55118 40000 55120
rect 35433 55115 35499 55118
rect 39200 55088 40000 55118
rect 20437 55042 20503 55045
rect 27889 55042 27955 55045
rect 20437 55040 27955 55042
rect 20437 54984 20442 55040
rect 20498 54984 27894 55040
rect 27950 54984 27955 55040
rect 20437 54982 27955 54984
rect 20437 54979 20503 54982
rect 27889 54979 27955 54982
rect 19568 54976 19888 54977
rect 19568 54912 19576 54976
rect 19640 54912 19656 54976
rect 19720 54912 19736 54976
rect 19800 54912 19816 54976
rect 19880 54912 19888 54976
rect 19568 54911 19888 54912
rect 20437 54906 20503 54909
rect 26785 54906 26851 54909
rect 20118 54904 26851 54906
rect 20118 54848 20442 54904
rect 20498 54848 26790 54904
rect 26846 54848 26851 54904
rect 20118 54846 26851 54848
rect 17493 54770 17559 54773
rect 20118 54770 20178 54846
rect 20437 54843 20503 54846
rect 26785 54843 26851 54846
rect 17493 54768 20178 54770
rect 17493 54712 17498 54768
rect 17554 54712 20178 54768
rect 17493 54710 20178 54712
rect 17493 54707 17559 54710
rect 14365 54634 14431 54637
rect 19241 54634 19307 54637
rect 14365 54632 19307 54634
rect 14365 54576 14370 54632
rect 14426 54576 19246 54632
rect 19302 54576 19307 54632
rect 14365 54574 19307 54576
rect 14365 54571 14431 54574
rect 19241 54571 19307 54574
rect 21541 54634 21607 54637
rect 22737 54634 22803 54637
rect 26233 54634 26299 54637
rect 21541 54632 26299 54634
rect 21541 54576 21546 54632
rect 21602 54576 22742 54632
rect 22798 54576 26238 54632
rect 26294 54576 26299 54632
rect 21541 54574 26299 54576
rect 21541 54571 21607 54574
rect 22737 54571 22803 54574
rect 26233 54571 26299 54574
rect 6177 54498 6243 54501
rect 13261 54498 13327 54501
rect 6177 54496 13327 54498
rect 6177 54440 6182 54496
rect 6238 54440 13266 54496
rect 13322 54440 13327 54496
rect 6177 54438 13327 54440
rect 6177 54435 6243 54438
rect 13261 54435 13327 54438
rect 13537 54498 13603 54501
rect 22461 54498 22527 54501
rect 13537 54496 22527 54498
rect 13537 54440 13542 54496
rect 13598 54440 22466 54496
rect 22522 54440 22527 54496
rect 13537 54438 22527 54440
rect 13537 54435 13603 54438
rect 22461 54435 22527 54438
rect 4208 54432 4528 54433
rect 4208 54368 4216 54432
rect 4280 54368 4296 54432
rect 4360 54368 4376 54432
rect 4440 54368 4456 54432
rect 4520 54368 4528 54432
rect 4208 54367 4528 54368
rect 34928 54432 35248 54433
rect 34928 54368 34936 54432
rect 35000 54368 35016 54432
rect 35080 54368 35096 54432
rect 35160 54368 35176 54432
rect 35240 54368 35248 54432
rect 34928 54367 35248 54368
rect 16849 54362 16915 54365
rect 19333 54362 19399 54365
rect 16849 54360 19399 54362
rect 16849 54304 16854 54360
rect 16910 54304 19338 54360
rect 19394 54304 19399 54360
rect 16849 54302 19399 54304
rect 16849 54299 16915 54302
rect 19333 54299 19399 54302
rect 16113 54226 16179 54229
rect 20897 54226 20963 54229
rect 16113 54224 20963 54226
rect 16113 54168 16118 54224
rect 16174 54168 20902 54224
rect 20958 54168 20963 54224
rect 16113 54166 20963 54168
rect 16113 54163 16179 54166
rect 20897 54163 20963 54166
rect 24485 54226 24551 54229
rect 24710 54226 24716 54228
rect 24485 54224 24716 54226
rect 24485 54168 24490 54224
rect 24546 54168 24716 54224
rect 24485 54166 24716 54168
rect 24485 54163 24551 54166
rect 24710 54164 24716 54166
rect 24780 54164 24786 54228
rect 13353 54090 13419 54093
rect 16849 54090 16915 54093
rect 13353 54088 16915 54090
rect 13353 54032 13358 54088
rect 13414 54032 16854 54088
rect 16910 54032 16915 54088
rect 13353 54030 16915 54032
rect 13353 54027 13419 54030
rect 16849 54027 16915 54030
rect 21357 54090 21423 54093
rect 21766 54090 21772 54092
rect 21357 54088 21772 54090
rect 21357 54032 21362 54088
rect 21418 54032 21772 54088
rect 21357 54030 21772 54032
rect 21357 54027 21423 54030
rect 21766 54028 21772 54030
rect 21836 54090 21842 54092
rect 25773 54090 25839 54093
rect 21836 54088 25839 54090
rect 21836 54032 25778 54088
rect 25834 54032 25839 54088
rect 21836 54030 25839 54032
rect 21836 54028 21842 54030
rect 25773 54027 25839 54030
rect 28901 54090 28967 54093
rect 32581 54090 32647 54093
rect 28901 54088 32647 54090
rect 28901 54032 28906 54088
rect 28962 54032 32586 54088
rect 32642 54032 32647 54088
rect 28901 54030 32647 54032
rect 28901 54027 28967 54030
rect 32581 54027 32647 54030
rect 14733 53956 14799 53957
rect 14733 53954 14780 53956
rect 14688 53952 14780 53954
rect 14688 53896 14738 53952
rect 14688 53894 14780 53896
rect 14733 53892 14780 53894
rect 14844 53892 14850 53956
rect 14917 53954 14983 53957
rect 18321 53954 18387 53957
rect 19425 53954 19491 53957
rect 14917 53952 19491 53954
rect 14917 53896 14922 53952
rect 14978 53896 18326 53952
rect 18382 53896 19430 53952
rect 19486 53896 19491 53952
rect 14917 53894 19491 53896
rect 14733 53891 14799 53892
rect 14917 53891 14983 53894
rect 18321 53891 18387 53894
rect 19425 53891 19491 53894
rect 21633 53954 21699 53957
rect 23473 53954 23539 53957
rect 21633 53952 23539 53954
rect 21633 53896 21638 53952
rect 21694 53896 23478 53952
rect 23534 53896 23539 53952
rect 21633 53894 23539 53896
rect 21633 53891 21699 53894
rect 23473 53891 23539 53894
rect 24485 53956 24551 53957
rect 24485 53952 24532 53956
rect 24596 53954 24602 53956
rect 31937 53954 32003 53957
rect 35249 53954 35315 53957
rect 24485 53896 24490 53952
rect 24485 53892 24532 53896
rect 24596 53894 24642 53954
rect 31937 53952 35315 53954
rect 31937 53896 31942 53952
rect 31998 53896 35254 53952
rect 35310 53896 35315 53952
rect 31937 53894 35315 53896
rect 24596 53892 24602 53894
rect 24485 53891 24551 53892
rect 31937 53891 32003 53894
rect 35249 53891 35315 53894
rect 19568 53888 19888 53889
rect 0 53818 800 53848
rect 19568 53824 19576 53888
rect 19640 53824 19656 53888
rect 19720 53824 19736 53888
rect 19800 53824 19816 53888
rect 19880 53824 19888 53888
rect 19568 53823 19888 53824
rect 3693 53818 3759 53821
rect 0 53816 3759 53818
rect 0 53760 3698 53816
rect 3754 53760 3759 53816
rect 0 53758 3759 53760
rect 0 53728 800 53758
rect 3693 53755 3759 53758
rect 15101 53818 15167 53821
rect 17493 53818 17559 53821
rect 15101 53816 17559 53818
rect 15101 53760 15106 53816
rect 15162 53760 17498 53816
rect 17554 53760 17559 53816
rect 15101 53758 17559 53760
rect 15101 53755 15167 53758
rect 17493 53755 17559 53758
rect 35433 53818 35499 53821
rect 39200 53818 40000 53848
rect 35433 53816 40000 53818
rect 35433 53760 35438 53816
rect 35494 53760 40000 53816
rect 35433 53758 40000 53760
rect 35433 53755 35499 53758
rect 39200 53728 40000 53758
rect 15469 53682 15535 53685
rect 19609 53682 19675 53685
rect 15469 53680 19675 53682
rect 15469 53624 15474 53680
rect 15530 53624 19614 53680
rect 19670 53624 19675 53680
rect 15469 53622 19675 53624
rect 15469 53619 15535 53622
rect 19609 53619 19675 53622
rect 17861 53546 17927 53549
rect 23749 53546 23815 53549
rect 17861 53544 23815 53546
rect 17861 53488 17866 53544
rect 17922 53488 23754 53544
rect 23810 53488 23815 53544
rect 17861 53486 23815 53488
rect 17861 53483 17927 53486
rect 23749 53483 23815 53486
rect 24117 53546 24183 53549
rect 27613 53546 27679 53549
rect 24117 53544 27679 53546
rect 24117 53488 24122 53544
rect 24178 53488 27618 53544
rect 27674 53488 27679 53544
rect 24117 53486 27679 53488
rect 24117 53483 24183 53486
rect 27613 53483 27679 53486
rect 15193 53410 15259 53413
rect 18597 53410 18663 53413
rect 15193 53408 18663 53410
rect 15193 53352 15198 53408
rect 15254 53352 18602 53408
rect 18658 53352 18663 53408
rect 15193 53350 18663 53352
rect 15193 53347 15259 53350
rect 18597 53347 18663 53350
rect 23105 53410 23171 53413
rect 23657 53410 23723 53413
rect 28993 53410 29059 53413
rect 23105 53408 29059 53410
rect 23105 53352 23110 53408
rect 23166 53352 23662 53408
rect 23718 53352 28998 53408
rect 29054 53352 29059 53408
rect 23105 53350 29059 53352
rect 23105 53347 23171 53350
rect 23657 53347 23723 53350
rect 28993 53347 29059 53350
rect 4208 53344 4528 53345
rect 4208 53280 4216 53344
rect 4280 53280 4296 53344
rect 4360 53280 4376 53344
rect 4440 53280 4456 53344
rect 4520 53280 4528 53344
rect 4208 53279 4528 53280
rect 34928 53344 35248 53345
rect 34928 53280 34936 53344
rect 35000 53280 35016 53344
rect 35080 53280 35096 53344
rect 35160 53280 35176 53344
rect 35240 53280 35248 53344
rect 34928 53279 35248 53280
rect 19517 53274 19583 53277
rect 26693 53274 26759 53277
rect 19517 53272 26759 53274
rect 19517 53216 19522 53272
rect 19578 53216 26698 53272
rect 26754 53216 26759 53272
rect 19517 53214 26759 53216
rect 19517 53211 19583 53214
rect 26693 53211 26759 53214
rect 3325 53138 3391 53141
rect 9949 53138 10015 53141
rect 3325 53136 10015 53138
rect 3325 53080 3330 53136
rect 3386 53080 9954 53136
rect 10010 53080 10015 53136
rect 3325 53078 10015 53080
rect 3325 53075 3391 53078
rect 9949 53075 10015 53078
rect 20713 53138 20779 53141
rect 25773 53138 25839 53141
rect 20713 53136 25839 53138
rect 20713 53080 20718 53136
rect 20774 53080 25778 53136
rect 25834 53080 25839 53136
rect 20713 53078 25839 53080
rect 20713 53075 20779 53078
rect 25773 53075 25839 53078
rect 16205 53002 16271 53005
rect 22277 53002 22343 53005
rect 25037 53002 25103 53005
rect 16205 53000 25103 53002
rect 16205 52944 16210 53000
rect 16266 52944 22282 53000
rect 22338 52944 25042 53000
rect 25098 52944 25103 53000
rect 16205 52942 25103 52944
rect 16205 52939 16271 52942
rect 22277 52939 22343 52942
rect 25037 52939 25103 52942
rect 20621 52866 20687 52869
rect 23933 52866 23999 52869
rect 20621 52864 23999 52866
rect 20621 52808 20626 52864
rect 20682 52808 23938 52864
rect 23994 52808 23999 52864
rect 20621 52806 23999 52808
rect 20621 52803 20687 52806
rect 23933 52803 23999 52806
rect 29637 52866 29703 52869
rect 33317 52866 33383 52869
rect 29637 52864 33383 52866
rect 29637 52808 29642 52864
rect 29698 52808 33322 52864
rect 33378 52808 33383 52864
rect 29637 52806 33383 52808
rect 29637 52803 29703 52806
rect 33317 52803 33383 52806
rect 19568 52800 19888 52801
rect 19568 52736 19576 52800
rect 19640 52736 19656 52800
rect 19720 52736 19736 52800
rect 19800 52736 19816 52800
rect 19880 52736 19888 52800
rect 19568 52735 19888 52736
rect 14733 52730 14799 52733
rect 16941 52730 17007 52733
rect 29177 52730 29243 52733
rect 14733 52728 17007 52730
rect 14733 52672 14738 52728
rect 14794 52672 16946 52728
rect 17002 52672 17007 52728
rect 14733 52670 17007 52672
rect 14733 52667 14799 52670
rect 16941 52667 17007 52670
rect 22188 52728 29243 52730
rect 22188 52672 29182 52728
rect 29238 52672 29243 52728
rect 22188 52670 29243 52672
rect 15285 52594 15351 52597
rect 22188 52594 22248 52670
rect 29177 52667 29243 52670
rect 15285 52592 22248 52594
rect 15285 52536 15290 52592
rect 15346 52536 22248 52592
rect 15285 52534 22248 52536
rect 22369 52594 22435 52597
rect 25773 52594 25839 52597
rect 22369 52592 25839 52594
rect 22369 52536 22374 52592
rect 22430 52536 25778 52592
rect 25834 52536 25839 52592
rect 22369 52534 25839 52536
rect 15285 52531 15351 52534
rect 0 52458 800 52488
rect 20992 52461 21052 52534
rect 22369 52531 22435 52534
rect 25773 52531 25839 52534
rect 29453 52594 29519 52597
rect 34697 52594 34763 52597
rect 29453 52592 34763 52594
rect 29453 52536 29458 52592
rect 29514 52536 34702 52592
rect 34758 52536 34763 52592
rect 29453 52534 34763 52536
rect 29453 52531 29519 52534
rect 34697 52531 34763 52534
rect 3325 52458 3391 52461
rect 0 52456 3391 52458
rect 0 52400 3330 52456
rect 3386 52400 3391 52456
rect 0 52398 3391 52400
rect 0 52368 800 52398
rect 3325 52395 3391 52398
rect 16573 52458 16639 52461
rect 18689 52458 18755 52461
rect 16573 52456 18755 52458
rect 16573 52400 16578 52456
rect 16634 52400 18694 52456
rect 18750 52400 18755 52456
rect 16573 52398 18755 52400
rect 16573 52395 16639 52398
rect 18689 52395 18755 52398
rect 20989 52456 21055 52461
rect 20989 52400 20994 52456
rect 21050 52400 21055 52456
rect 20989 52395 21055 52400
rect 29545 52458 29611 52461
rect 31753 52458 31819 52461
rect 29545 52456 31819 52458
rect 29545 52400 29550 52456
rect 29606 52400 31758 52456
rect 31814 52400 31819 52456
rect 29545 52398 31819 52400
rect 29545 52395 29611 52398
rect 31753 52395 31819 52398
rect 34605 52458 34671 52461
rect 39200 52458 40000 52488
rect 34605 52456 40000 52458
rect 34605 52400 34610 52456
rect 34666 52400 40000 52456
rect 34605 52398 40000 52400
rect 34605 52395 34671 52398
rect 39200 52368 40000 52398
rect 4208 52256 4528 52257
rect 4208 52192 4216 52256
rect 4280 52192 4296 52256
rect 4360 52192 4376 52256
rect 4440 52192 4456 52256
rect 4520 52192 4528 52256
rect 4208 52191 4528 52192
rect 34928 52256 35248 52257
rect 34928 52192 34936 52256
rect 35000 52192 35016 52256
rect 35080 52192 35096 52256
rect 35160 52192 35176 52256
rect 35240 52192 35248 52256
rect 34928 52191 35248 52192
rect 15101 52186 15167 52189
rect 16665 52186 16731 52189
rect 22277 52186 22343 52189
rect 15101 52184 22343 52186
rect 15101 52128 15106 52184
rect 15162 52128 16670 52184
rect 16726 52128 22282 52184
rect 22338 52128 22343 52184
rect 15101 52126 22343 52128
rect 15101 52123 15167 52126
rect 16665 52123 16731 52126
rect 22277 52123 22343 52126
rect 25221 52186 25287 52189
rect 25405 52186 25471 52189
rect 25221 52184 25471 52186
rect 25221 52128 25226 52184
rect 25282 52128 25410 52184
rect 25466 52128 25471 52184
rect 25221 52126 25471 52128
rect 25221 52123 25287 52126
rect 25405 52123 25471 52126
rect 16113 52050 16179 52053
rect 18873 52050 18939 52053
rect 16113 52048 18939 52050
rect 16113 51992 16118 52048
rect 16174 51992 18878 52048
rect 18934 51992 18939 52048
rect 16113 51990 18939 51992
rect 16113 51987 16179 51990
rect 18873 51987 18939 51990
rect 19057 52050 19123 52053
rect 21817 52050 21883 52053
rect 19057 52048 21883 52050
rect 19057 51992 19062 52048
rect 19118 51992 21822 52048
rect 21878 51992 21883 52048
rect 19057 51990 21883 51992
rect 19057 51987 19123 51990
rect 21817 51987 21883 51990
rect 30557 52050 30623 52053
rect 35433 52050 35499 52053
rect 30557 52048 35499 52050
rect 30557 51992 30562 52048
rect 30618 51992 35438 52048
rect 35494 51992 35499 52048
rect 30557 51990 35499 51992
rect 30557 51987 30623 51990
rect 35433 51987 35499 51990
rect 16481 51914 16547 51917
rect 20345 51914 20411 51917
rect 20897 51914 20963 51917
rect 16481 51912 20963 51914
rect 16481 51856 16486 51912
rect 16542 51856 20350 51912
rect 20406 51856 20902 51912
rect 20958 51856 20963 51912
rect 16481 51854 20963 51856
rect 16481 51851 16547 51854
rect 20345 51851 20411 51854
rect 20897 51851 20963 51854
rect 21541 51914 21607 51917
rect 24853 51914 24919 51917
rect 21541 51912 24919 51914
rect 21541 51856 21546 51912
rect 21602 51856 24858 51912
rect 24914 51856 24919 51912
rect 21541 51854 24919 51856
rect 21541 51851 21607 51854
rect 24853 51851 24919 51854
rect 19977 51778 20043 51781
rect 22921 51778 22987 51781
rect 19977 51776 22987 51778
rect 19977 51720 19982 51776
rect 20038 51720 22926 51776
rect 22982 51720 22987 51776
rect 19977 51718 22987 51720
rect 19977 51715 20043 51718
rect 22921 51715 22987 51718
rect 19568 51712 19888 51713
rect 19568 51648 19576 51712
rect 19640 51648 19656 51712
rect 19720 51648 19736 51712
rect 19800 51648 19816 51712
rect 19880 51648 19888 51712
rect 19568 51647 19888 51648
rect 20713 51642 20779 51645
rect 21541 51642 21607 51645
rect 23289 51642 23355 51645
rect 20713 51640 23355 51642
rect 20713 51584 20718 51640
rect 20774 51584 21546 51640
rect 21602 51584 23294 51640
rect 23350 51584 23355 51640
rect 20713 51582 23355 51584
rect 20713 51579 20779 51582
rect 21541 51579 21607 51582
rect 23289 51579 23355 51582
rect 17769 51506 17835 51509
rect 19977 51506 20043 51509
rect 17769 51504 20043 51506
rect 17769 51448 17774 51504
rect 17830 51448 19982 51504
rect 20038 51448 20043 51504
rect 17769 51446 20043 51448
rect 17769 51443 17835 51446
rect 19977 51443 20043 51446
rect 24853 51370 24919 51373
rect 3374 51368 24919 51370
rect 3374 51312 24858 51368
rect 24914 51312 24919 51368
rect 3374 51310 24919 51312
rect 0 51098 800 51128
rect 3374 51098 3434 51310
rect 24853 51307 24919 51310
rect 27838 51308 27844 51372
rect 27908 51370 27914 51372
rect 27908 51310 35588 51370
rect 27908 51308 27914 51310
rect 14733 51234 14799 51237
rect 17585 51234 17651 51237
rect 14733 51232 17651 51234
rect 14733 51176 14738 51232
rect 14794 51176 17590 51232
rect 17646 51176 17651 51232
rect 14733 51174 17651 51176
rect 14733 51171 14799 51174
rect 17585 51171 17651 51174
rect 18413 51234 18479 51237
rect 24945 51234 25011 51237
rect 18413 51232 25011 51234
rect 18413 51176 18418 51232
rect 18474 51176 24950 51232
rect 25006 51176 25011 51232
rect 18413 51174 25011 51176
rect 18413 51171 18479 51174
rect 24945 51171 25011 51174
rect 28441 51234 28507 51237
rect 28574 51234 28580 51236
rect 28441 51232 28580 51234
rect 28441 51176 28446 51232
rect 28502 51176 28580 51232
rect 28441 51174 28580 51176
rect 28441 51171 28507 51174
rect 28574 51172 28580 51174
rect 28644 51172 28650 51236
rect 29126 51172 29132 51236
rect 29196 51234 29202 51236
rect 29269 51234 29335 51237
rect 29196 51232 29335 51234
rect 29196 51176 29274 51232
rect 29330 51176 29335 51232
rect 29196 51174 29335 51176
rect 29196 51172 29202 51174
rect 29269 51171 29335 51174
rect 4208 51168 4528 51169
rect 4208 51104 4216 51168
rect 4280 51104 4296 51168
rect 4360 51104 4376 51168
rect 4440 51104 4456 51168
rect 4520 51104 4528 51168
rect 4208 51103 4528 51104
rect 34928 51168 35248 51169
rect 34928 51104 34936 51168
rect 35000 51104 35016 51168
rect 35080 51104 35096 51168
rect 35160 51104 35176 51168
rect 35240 51104 35248 51168
rect 34928 51103 35248 51104
rect 0 51038 3434 51098
rect 15653 51098 15719 51101
rect 21725 51098 21791 51101
rect 15653 51096 21791 51098
rect 15653 51040 15658 51096
rect 15714 51040 21730 51096
rect 21786 51040 21791 51096
rect 15653 51038 21791 51040
rect 0 51008 800 51038
rect 15653 51035 15719 51038
rect 21725 51035 21791 51038
rect 25497 51098 25563 51101
rect 30097 51098 30163 51101
rect 25497 51096 30163 51098
rect 25497 51040 25502 51096
rect 25558 51040 30102 51096
rect 30158 51040 30163 51096
rect 25497 51038 30163 51040
rect 35528 51098 35588 51310
rect 39200 51098 40000 51128
rect 35528 51038 40000 51098
rect 25497 51035 25563 51038
rect 30097 51035 30163 51038
rect 39200 51008 40000 51038
rect 17217 50962 17283 50965
rect 20161 50962 20227 50965
rect 17217 50960 20227 50962
rect 17217 50904 17222 50960
rect 17278 50904 20166 50960
rect 20222 50904 20227 50960
rect 17217 50902 20227 50904
rect 17217 50899 17283 50902
rect 20161 50899 20227 50902
rect 22001 50962 22067 50965
rect 25589 50962 25655 50965
rect 22001 50960 25655 50962
rect 22001 50904 22006 50960
rect 22062 50904 25594 50960
rect 25650 50904 25655 50960
rect 22001 50902 25655 50904
rect 22001 50899 22067 50902
rect 25589 50899 25655 50902
rect 17585 50826 17651 50829
rect 18413 50826 18479 50829
rect 19517 50826 19583 50829
rect 20897 50826 20963 50829
rect 21817 50828 21883 50829
rect 21766 50826 21772 50828
rect 17585 50824 20963 50826
rect 17585 50768 17590 50824
rect 17646 50768 18418 50824
rect 18474 50768 19522 50824
rect 19578 50768 20902 50824
rect 20958 50768 20963 50824
rect 17585 50766 20963 50768
rect 21726 50766 21772 50826
rect 21836 50824 21883 50828
rect 21878 50768 21883 50824
rect 17585 50763 17651 50766
rect 18413 50763 18479 50766
rect 19517 50763 19583 50766
rect 20897 50763 20963 50766
rect 21766 50764 21772 50766
rect 21836 50764 21883 50768
rect 21817 50763 21883 50764
rect 24669 50826 24735 50829
rect 30373 50826 30439 50829
rect 24669 50824 30439 50826
rect 24669 50768 24674 50824
rect 24730 50768 30378 50824
rect 30434 50768 30439 50824
rect 24669 50766 30439 50768
rect 24669 50763 24735 50766
rect 30373 50763 30439 50766
rect 20069 50690 20135 50693
rect 24672 50690 24732 50763
rect 20069 50688 24732 50690
rect 20069 50632 20074 50688
rect 20130 50632 24732 50688
rect 20069 50630 24732 50632
rect 26877 50690 26943 50693
rect 28993 50690 29059 50693
rect 26877 50688 29059 50690
rect 26877 50632 26882 50688
rect 26938 50632 28998 50688
rect 29054 50632 29059 50688
rect 26877 50630 29059 50632
rect 20069 50627 20135 50630
rect 26877 50627 26943 50630
rect 28993 50627 29059 50630
rect 31477 50690 31543 50693
rect 33685 50690 33751 50693
rect 31477 50688 33751 50690
rect 31477 50632 31482 50688
rect 31538 50632 33690 50688
rect 33746 50632 33751 50688
rect 31477 50630 33751 50632
rect 31477 50627 31543 50630
rect 33685 50627 33751 50630
rect 19568 50624 19888 50625
rect 19568 50560 19576 50624
rect 19640 50560 19656 50624
rect 19720 50560 19736 50624
rect 19800 50560 19816 50624
rect 19880 50560 19888 50624
rect 19568 50559 19888 50560
rect 11881 50554 11947 50557
rect 14825 50554 14891 50557
rect 11881 50552 14891 50554
rect 11881 50496 11886 50552
rect 11942 50496 14830 50552
rect 14886 50496 14891 50552
rect 11881 50494 14891 50496
rect 11881 50491 11947 50494
rect 14825 50491 14891 50494
rect 24209 50554 24275 50557
rect 35433 50554 35499 50557
rect 24209 50552 35499 50554
rect 24209 50496 24214 50552
rect 24270 50496 35438 50552
rect 35494 50496 35499 50552
rect 24209 50494 35499 50496
rect 24209 50491 24275 50494
rect 35433 50491 35499 50494
rect 28073 50418 28139 50421
rect 28533 50418 28599 50421
rect 31017 50418 31083 50421
rect 28073 50416 31083 50418
rect 28073 50360 28078 50416
rect 28134 50360 28538 50416
rect 28594 50360 31022 50416
rect 31078 50360 31083 50416
rect 28073 50358 31083 50360
rect 28073 50355 28139 50358
rect 28533 50355 28599 50358
rect 31017 50355 31083 50358
rect 17401 50282 17467 50285
rect 24485 50282 24551 50285
rect 17401 50280 24551 50282
rect 17401 50224 17406 50280
rect 17462 50224 24490 50280
rect 24546 50224 24551 50280
rect 17401 50222 24551 50224
rect 17401 50219 17467 50222
rect 24485 50219 24551 50222
rect 30649 50282 30715 50285
rect 32213 50282 32279 50285
rect 30649 50280 32279 50282
rect 30649 50224 30654 50280
rect 30710 50224 32218 50280
rect 32274 50224 32279 50280
rect 30649 50222 32279 50224
rect 30649 50219 30715 50222
rect 32213 50219 32279 50222
rect 25221 50146 25287 50149
rect 30557 50146 30623 50149
rect 25221 50144 30623 50146
rect 25221 50088 25226 50144
rect 25282 50088 30562 50144
rect 30618 50088 30623 50144
rect 25221 50086 30623 50088
rect 25221 50083 25287 50086
rect 30557 50083 30623 50086
rect 4208 50080 4528 50081
rect 4208 50016 4216 50080
rect 4280 50016 4296 50080
rect 4360 50016 4376 50080
rect 4440 50016 4456 50080
rect 4520 50016 4528 50080
rect 4208 50015 4528 50016
rect 34928 50080 35248 50081
rect 34928 50016 34936 50080
rect 35000 50016 35016 50080
rect 35080 50016 35096 50080
rect 35160 50016 35176 50080
rect 35240 50016 35248 50080
rect 34928 50015 35248 50016
rect 17217 50010 17283 50013
rect 19885 50010 19951 50013
rect 17217 50008 19951 50010
rect 17217 49952 17222 50008
rect 17278 49952 19890 50008
rect 19946 49952 19951 50008
rect 17217 49950 19951 49952
rect 17217 49947 17283 49950
rect 19885 49947 19951 49950
rect 25773 50010 25839 50013
rect 26785 50010 26851 50013
rect 31201 50010 31267 50013
rect 25773 50008 31267 50010
rect 25773 49952 25778 50008
rect 25834 49952 26790 50008
rect 26846 49952 31206 50008
rect 31262 49952 31267 50008
rect 25773 49950 31267 49952
rect 25773 49947 25839 49950
rect 26785 49947 26851 49950
rect 31201 49947 31267 49950
rect 27889 49874 27955 49877
rect 30925 49874 30991 49877
rect 27889 49872 30991 49874
rect 27889 49816 27894 49872
rect 27950 49816 30930 49872
rect 30986 49816 30991 49872
rect 27889 49814 30991 49816
rect 27889 49811 27955 49814
rect 30925 49811 30991 49814
rect 0 49738 800 49768
rect 4061 49738 4127 49741
rect 0 49736 4127 49738
rect 0 49680 4066 49736
rect 4122 49680 4127 49736
rect 0 49678 4127 49680
rect 0 49648 800 49678
rect 4061 49675 4127 49678
rect 5073 49738 5139 49741
rect 8753 49738 8819 49741
rect 5073 49736 8819 49738
rect 5073 49680 5078 49736
rect 5134 49680 8758 49736
rect 8814 49680 8819 49736
rect 5073 49678 8819 49680
rect 5073 49675 5139 49678
rect 8753 49675 8819 49678
rect 21081 49738 21147 49741
rect 21214 49738 21220 49740
rect 21081 49736 21220 49738
rect 21081 49680 21086 49736
rect 21142 49680 21220 49736
rect 21081 49678 21220 49680
rect 21081 49675 21147 49678
rect 21214 49676 21220 49678
rect 21284 49676 21290 49740
rect 24669 49738 24735 49741
rect 27613 49738 27679 49741
rect 24669 49736 27679 49738
rect 24669 49680 24674 49736
rect 24730 49680 27618 49736
rect 27674 49680 27679 49736
rect 24669 49678 27679 49680
rect 24669 49675 24735 49678
rect 27613 49675 27679 49678
rect 29729 49738 29795 49741
rect 39200 49738 40000 49768
rect 29729 49736 40000 49738
rect 29729 49680 29734 49736
rect 29790 49680 40000 49736
rect 29729 49678 40000 49680
rect 29729 49675 29795 49678
rect 39200 49648 40000 49678
rect 3325 49602 3391 49605
rect 11605 49602 11671 49605
rect 3325 49600 11671 49602
rect 3325 49544 3330 49600
rect 3386 49544 11610 49600
rect 11666 49544 11671 49600
rect 3325 49542 11671 49544
rect 3325 49539 3391 49542
rect 11605 49539 11671 49542
rect 28809 49602 28875 49605
rect 30833 49602 30899 49605
rect 28809 49600 30899 49602
rect 28809 49544 28814 49600
rect 28870 49544 30838 49600
rect 30894 49544 30899 49600
rect 28809 49542 30899 49544
rect 28809 49539 28875 49542
rect 30833 49539 30899 49542
rect 19568 49536 19888 49537
rect 19568 49472 19576 49536
rect 19640 49472 19656 49536
rect 19720 49472 19736 49536
rect 19800 49472 19816 49536
rect 19880 49472 19888 49536
rect 19568 49471 19888 49472
rect 29085 49468 29151 49469
rect 29085 49466 29132 49468
rect 29040 49464 29132 49466
rect 29040 49408 29090 49464
rect 29040 49406 29132 49408
rect 29085 49404 29132 49406
rect 29196 49404 29202 49468
rect 29085 49403 29151 49404
rect 16665 49330 16731 49333
rect 22185 49330 22251 49333
rect 16665 49328 22251 49330
rect 16665 49272 16670 49328
rect 16726 49272 22190 49328
rect 22246 49272 22251 49328
rect 16665 49270 22251 49272
rect 16665 49267 16731 49270
rect 22185 49267 22251 49270
rect 27981 49330 28047 49333
rect 30189 49330 30255 49333
rect 31385 49330 31451 49333
rect 27981 49328 31451 49330
rect 27981 49272 27986 49328
rect 28042 49272 30194 49328
rect 30250 49272 31390 49328
rect 31446 49272 31451 49328
rect 27981 49270 31451 49272
rect 27981 49267 28047 49270
rect 30189 49267 30255 49270
rect 31385 49267 31451 49270
rect 20621 49194 20687 49197
rect 31017 49194 31083 49197
rect 20621 49192 31083 49194
rect 20621 49136 20626 49192
rect 20682 49136 31022 49192
rect 31078 49136 31083 49192
rect 20621 49134 31083 49136
rect 20621 49131 20687 49134
rect 31017 49131 31083 49134
rect 19241 49058 19307 49061
rect 22461 49058 22527 49061
rect 24025 49058 24091 49061
rect 19241 49056 24091 49058
rect 19241 49000 19246 49056
rect 19302 49000 22466 49056
rect 22522 49000 24030 49056
rect 24086 49000 24091 49056
rect 19241 48998 24091 49000
rect 19241 48995 19307 48998
rect 22461 48995 22527 48998
rect 24025 48995 24091 48998
rect 27153 49058 27219 49061
rect 29913 49058 29979 49061
rect 27153 49056 29979 49058
rect 27153 49000 27158 49056
rect 27214 49000 29918 49056
rect 29974 49000 29979 49056
rect 27153 48998 29979 49000
rect 27153 48995 27219 48998
rect 29913 48995 29979 48998
rect 4208 48992 4528 48993
rect 4208 48928 4216 48992
rect 4280 48928 4296 48992
rect 4360 48928 4376 48992
rect 4440 48928 4456 48992
rect 4520 48928 4528 48992
rect 4208 48927 4528 48928
rect 34928 48992 35248 48993
rect 34928 48928 34936 48992
rect 35000 48928 35016 48992
rect 35080 48928 35096 48992
rect 35160 48928 35176 48992
rect 35240 48928 35248 48992
rect 34928 48927 35248 48928
rect 15101 48922 15167 48925
rect 17401 48922 17467 48925
rect 15101 48920 17467 48922
rect 15101 48864 15106 48920
rect 15162 48864 17406 48920
rect 17462 48864 17467 48920
rect 15101 48862 17467 48864
rect 15101 48859 15167 48862
rect 17401 48859 17467 48862
rect 18229 48922 18295 48925
rect 20345 48922 20411 48925
rect 21173 48922 21239 48925
rect 18229 48920 21239 48922
rect 18229 48864 18234 48920
rect 18290 48864 20350 48920
rect 20406 48864 21178 48920
rect 21234 48864 21239 48920
rect 18229 48862 21239 48864
rect 18229 48859 18295 48862
rect 20345 48859 20411 48862
rect 21173 48859 21239 48862
rect 24209 48922 24275 48925
rect 28993 48922 29059 48925
rect 24209 48920 29059 48922
rect 24209 48864 24214 48920
rect 24270 48864 28998 48920
rect 29054 48864 29059 48920
rect 24209 48862 29059 48864
rect 24209 48859 24275 48862
rect 28993 48859 29059 48862
rect 4061 48786 4127 48789
rect 15377 48786 15443 48789
rect 4061 48784 15443 48786
rect 4061 48728 4066 48784
rect 4122 48728 15382 48784
rect 15438 48728 15443 48784
rect 4061 48726 15443 48728
rect 4061 48723 4127 48726
rect 15377 48723 15443 48726
rect 19977 48786 20043 48789
rect 23657 48786 23723 48789
rect 19977 48784 23723 48786
rect 19977 48728 19982 48784
rect 20038 48728 23662 48784
rect 23718 48728 23723 48784
rect 19977 48726 23723 48728
rect 19977 48723 20043 48726
rect 23657 48723 23723 48726
rect 25957 48786 26023 48789
rect 31201 48786 31267 48789
rect 25957 48784 31267 48786
rect 25957 48728 25962 48784
rect 26018 48728 31206 48784
rect 31262 48728 31267 48784
rect 25957 48726 31267 48728
rect 25957 48723 26023 48726
rect 31201 48723 31267 48726
rect 3509 48650 3575 48653
rect 19517 48650 19583 48653
rect 3509 48648 19583 48650
rect 3509 48592 3514 48648
rect 3570 48592 19522 48648
rect 19578 48592 19583 48648
rect 3509 48590 19583 48592
rect 3509 48587 3575 48590
rect 19517 48587 19583 48590
rect 22737 48650 22803 48653
rect 35617 48650 35683 48653
rect 22737 48648 35683 48650
rect 22737 48592 22742 48648
rect 22798 48592 35622 48648
rect 35678 48592 35683 48648
rect 22737 48590 35683 48592
rect 22737 48587 22803 48590
rect 35617 48587 35683 48590
rect 23013 48514 23079 48517
rect 27981 48514 28047 48517
rect 23013 48512 28047 48514
rect 23013 48456 23018 48512
rect 23074 48456 27986 48512
rect 28042 48456 28047 48512
rect 23013 48454 28047 48456
rect 23013 48451 23079 48454
rect 27981 48451 28047 48454
rect 19568 48448 19888 48449
rect 0 48378 800 48408
rect 19568 48384 19576 48448
rect 19640 48384 19656 48448
rect 19720 48384 19736 48448
rect 19800 48384 19816 48448
rect 19880 48384 19888 48448
rect 19568 48383 19888 48384
rect 3877 48378 3943 48381
rect 0 48376 3943 48378
rect 0 48320 3882 48376
rect 3938 48320 3943 48376
rect 0 48318 3943 48320
rect 0 48288 800 48318
rect 3877 48315 3943 48318
rect 20253 48378 20319 48381
rect 24669 48378 24735 48381
rect 20253 48376 24735 48378
rect 20253 48320 20258 48376
rect 20314 48320 24674 48376
rect 24730 48320 24735 48376
rect 20253 48318 24735 48320
rect 20253 48315 20319 48318
rect 24669 48315 24735 48318
rect 25221 48378 25287 48381
rect 30649 48378 30715 48381
rect 25221 48376 30715 48378
rect 25221 48320 25226 48376
rect 25282 48320 30654 48376
rect 30710 48320 30715 48376
rect 25221 48318 30715 48320
rect 25221 48315 25287 48318
rect 30649 48315 30715 48318
rect 35433 48378 35499 48381
rect 39200 48378 40000 48408
rect 35433 48376 40000 48378
rect 35433 48320 35438 48376
rect 35494 48320 40000 48376
rect 35433 48318 40000 48320
rect 35433 48315 35499 48318
rect 39200 48288 40000 48318
rect 19057 48242 19123 48245
rect 22369 48242 22435 48245
rect 19057 48240 22435 48242
rect 19057 48184 19062 48240
rect 19118 48184 22374 48240
rect 22430 48184 22435 48240
rect 19057 48182 22435 48184
rect 19057 48179 19123 48182
rect 22369 48179 22435 48182
rect 24485 48242 24551 48245
rect 28165 48242 28231 48245
rect 28809 48242 28875 48245
rect 29637 48244 29703 48245
rect 29637 48242 29684 48244
rect 24485 48240 28875 48242
rect 24485 48184 24490 48240
rect 24546 48184 28170 48240
rect 28226 48184 28814 48240
rect 28870 48184 28875 48240
rect 24485 48182 28875 48184
rect 29592 48240 29684 48242
rect 29592 48184 29642 48240
rect 29592 48182 29684 48184
rect 24485 48179 24551 48182
rect 28165 48179 28231 48182
rect 28809 48179 28875 48182
rect 29637 48180 29684 48182
rect 29748 48180 29754 48244
rect 29913 48242 29979 48245
rect 30046 48242 30052 48244
rect 29913 48240 30052 48242
rect 29913 48184 29918 48240
rect 29974 48184 30052 48240
rect 29913 48182 30052 48184
rect 29637 48179 29703 48180
rect 29913 48179 29979 48182
rect 30046 48180 30052 48182
rect 30116 48180 30122 48244
rect 27337 48106 27403 48109
rect 29729 48106 29795 48109
rect 30741 48106 30807 48109
rect 27337 48104 30807 48106
rect 27337 48048 27342 48104
rect 27398 48048 29734 48104
rect 29790 48048 30746 48104
rect 30802 48048 30807 48104
rect 27337 48046 30807 48048
rect 27337 48043 27403 48046
rect 29729 48043 29795 48046
rect 30741 48043 30807 48046
rect 26417 47970 26483 47973
rect 29453 47970 29519 47973
rect 26417 47968 29519 47970
rect 26417 47912 26422 47968
rect 26478 47912 29458 47968
rect 29514 47912 29519 47968
rect 26417 47910 29519 47912
rect 26417 47907 26483 47910
rect 29453 47907 29519 47910
rect 4208 47904 4528 47905
rect 4208 47840 4216 47904
rect 4280 47840 4296 47904
rect 4360 47840 4376 47904
rect 4440 47840 4456 47904
rect 4520 47840 4528 47904
rect 4208 47839 4528 47840
rect 34928 47904 35248 47905
rect 34928 47840 34936 47904
rect 35000 47840 35016 47904
rect 35080 47840 35096 47904
rect 35160 47840 35176 47904
rect 35240 47840 35248 47904
rect 34928 47839 35248 47840
rect 21357 47834 21423 47837
rect 24853 47834 24919 47837
rect 21357 47832 24919 47834
rect 21357 47776 21362 47832
rect 21418 47776 24858 47832
rect 24914 47776 24919 47832
rect 21357 47774 24919 47776
rect 21357 47771 21423 47774
rect 24853 47771 24919 47774
rect 26601 47834 26667 47837
rect 29085 47834 29151 47837
rect 26601 47832 29151 47834
rect 26601 47776 26606 47832
rect 26662 47776 29090 47832
rect 29146 47776 29151 47832
rect 26601 47774 29151 47776
rect 26601 47771 26667 47774
rect 29085 47771 29151 47774
rect 28349 47698 28415 47701
rect 32397 47698 32463 47701
rect 28349 47696 32463 47698
rect 28349 47640 28354 47696
rect 28410 47640 32402 47696
rect 32458 47640 32463 47696
rect 28349 47638 32463 47640
rect 28349 47635 28415 47638
rect 32397 47635 32463 47638
rect 25313 47426 25379 47429
rect 30649 47426 30715 47429
rect 25313 47424 30715 47426
rect 25313 47368 25318 47424
rect 25374 47368 30654 47424
rect 30710 47368 30715 47424
rect 25313 47366 30715 47368
rect 25313 47363 25379 47366
rect 30649 47363 30715 47366
rect 19568 47360 19888 47361
rect 19568 47296 19576 47360
rect 19640 47296 19656 47360
rect 19720 47296 19736 47360
rect 19800 47296 19816 47360
rect 19880 47296 19888 47360
rect 19568 47295 19888 47296
rect 20989 47290 21055 47293
rect 24209 47290 24275 47293
rect 20989 47288 24275 47290
rect 20989 47232 20994 47288
rect 21050 47232 24214 47288
rect 24270 47232 24275 47288
rect 20989 47230 24275 47232
rect 20989 47227 21055 47230
rect 24209 47227 24275 47230
rect 25221 47290 25287 47293
rect 30925 47290 30991 47293
rect 25221 47288 30991 47290
rect 25221 47232 25226 47288
rect 25282 47232 30930 47288
rect 30986 47232 30991 47288
rect 25221 47230 30991 47232
rect 25221 47227 25287 47230
rect 30925 47227 30991 47230
rect 21173 47154 21239 47157
rect 23565 47154 23631 47157
rect 21173 47152 23631 47154
rect 21173 47096 21178 47152
rect 21234 47096 23570 47152
rect 23626 47096 23631 47152
rect 21173 47094 23631 47096
rect 21173 47091 21239 47094
rect 23565 47091 23631 47094
rect 27153 47154 27219 47157
rect 31109 47154 31175 47157
rect 27153 47152 31175 47154
rect 27153 47096 27158 47152
rect 27214 47096 31114 47152
rect 31170 47096 31175 47152
rect 27153 47094 31175 47096
rect 27153 47091 27219 47094
rect 31109 47091 31175 47094
rect 32029 47154 32095 47157
rect 33133 47154 33199 47157
rect 32029 47152 33199 47154
rect 32029 47096 32034 47152
rect 32090 47096 33138 47152
rect 33194 47096 33199 47152
rect 32029 47094 33199 47096
rect 32029 47091 32095 47094
rect 33133 47091 33199 47094
rect 0 47018 800 47048
rect 3509 47018 3575 47021
rect 0 47016 3575 47018
rect 0 46960 3514 47016
rect 3570 46960 3575 47016
rect 0 46958 3575 46960
rect 0 46928 800 46958
rect 3509 46955 3575 46958
rect 3693 47018 3759 47021
rect 6269 47018 6335 47021
rect 3693 47016 6335 47018
rect 3693 46960 3698 47016
rect 3754 46960 6274 47016
rect 6330 46960 6335 47016
rect 3693 46958 6335 46960
rect 3693 46955 3759 46958
rect 6269 46955 6335 46958
rect 19977 47018 20043 47021
rect 20294 47018 20300 47020
rect 19977 47016 20300 47018
rect 19977 46960 19982 47016
rect 20038 46960 20300 47016
rect 19977 46958 20300 46960
rect 19977 46955 20043 46958
rect 20294 46956 20300 46958
rect 20364 46956 20370 47020
rect 21909 47018 21975 47021
rect 23749 47018 23815 47021
rect 24485 47018 24551 47021
rect 21909 47016 24551 47018
rect 21909 46960 21914 47016
rect 21970 46960 23754 47016
rect 23810 46960 24490 47016
rect 24546 46960 24551 47016
rect 21909 46958 24551 46960
rect 21909 46955 21975 46958
rect 23749 46955 23815 46958
rect 24485 46955 24551 46958
rect 25589 47018 25655 47021
rect 27521 47018 27587 47021
rect 25589 47016 27587 47018
rect 25589 46960 25594 47016
rect 25650 46960 27526 47016
rect 27582 46960 27587 47016
rect 25589 46958 27587 46960
rect 25589 46955 25655 46958
rect 27521 46955 27587 46958
rect 28206 46956 28212 47020
rect 28276 47018 28282 47020
rect 28349 47018 28415 47021
rect 28993 47018 29059 47021
rect 28276 47016 28415 47018
rect 28276 46960 28354 47016
rect 28410 46960 28415 47016
rect 28276 46958 28415 46960
rect 28276 46956 28282 46958
rect 28349 46955 28415 46958
rect 28950 47016 29059 47018
rect 28950 46960 28998 47016
rect 29054 46960 29059 47016
rect 28950 46955 29059 46960
rect 32673 47018 32739 47021
rect 34605 47018 34671 47021
rect 32673 47016 34671 47018
rect 32673 46960 32678 47016
rect 32734 46960 34610 47016
rect 34666 46960 34671 47016
rect 32673 46958 34671 46960
rect 32673 46955 32739 46958
rect 34605 46955 34671 46958
rect 35617 47018 35683 47021
rect 39200 47018 40000 47048
rect 35617 47016 40000 47018
rect 35617 46960 35622 47016
rect 35678 46960 40000 47016
rect 35617 46958 40000 46960
rect 35617 46955 35683 46958
rect 12801 46882 12867 46885
rect 15653 46882 15719 46885
rect 16849 46882 16915 46885
rect 12801 46880 16915 46882
rect 12801 46824 12806 46880
rect 12862 46824 15658 46880
rect 15714 46824 16854 46880
rect 16910 46824 16915 46880
rect 12801 46822 16915 46824
rect 12801 46819 12867 46822
rect 15653 46819 15719 46822
rect 16849 46819 16915 46822
rect 20069 46882 20135 46885
rect 22461 46882 22527 46885
rect 20069 46880 22527 46882
rect 20069 46824 20074 46880
rect 20130 46824 22466 46880
rect 22522 46824 22527 46880
rect 20069 46822 22527 46824
rect 20069 46819 20135 46822
rect 22461 46819 22527 46822
rect 27245 46882 27311 46885
rect 28950 46882 29010 46955
rect 39200 46928 40000 46958
rect 27245 46880 29010 46882
rect 27245 46824 27250 46880
rect 27306 46824 29010 46880
rect 27245 46822 29010 46824
rect 27245 46819 27311 46822
rect 4208 46816 4528 46817
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 46751 4528 46752
rect 34928 46816 35248 46817
rect 34928 46752 34936 46816
rect 35000 46752 35016 46816
rect 35080 46752 35096 46816
rect 35160 46752 35176 46816
rect 35240 46752 35248 46816
rect 34928 46751 35248 46752
rect 29177 46610 29243 46613
rect 30557 46610 30623 46613
rect 29177 46608 30623 46610
rect 29177 46552 29182 46608
rect 29238 46552 30562 46608
rect 30618 46552 30623 46608
rect 29177 46550 30623 46552
rect 29177 46547 29243 46550
rect 30557 46547 30623 46550
rect 17033 46474 17099 46477
rect 20846 46474 20852 46476
rect 17033 46472 20852 46474
rect 17033 46416 17038 46472
rect 17094 46416 20852 46472
rect 17033 46414 20852 46416
rect 17033 46411 17099 46414
rect 20846 46412 20852 46414
rect 20916 46412 20922 46476
rect 0 46338 800 46368
rect 1761 46338 1827 46341
rect 0 46336 1827 46338
rect 0 46280 1766 46336
rect 1822 46280 1827 46336
rect 0 46278 1827 46280
rect 0 46248 800 46278
rect 1761 46275 1827 46278
rect 11421 46338 11487 46341
rect 13629 46338 13695 46341
rect 11421 46336 13695 46338
rect 11421 46280 11426 46336
rect 11482 46280 13634 46336
rect 13690 46280 13695 46336
rect 11421 46278 13695 46280
rect 11421 46275 11487 46278
rect 13629 46275 13695 46278
rect 25773 46338 25839 46341
rect 26877 46338 26943 46341
rect 25773 46336 26943 46338
rect 25773 46280 25778 46336
rect 25834 46280 26882 46336
rect 26938 46280 26943 46336
rect 25773 46278 26943 46280
rect 25773 46275 25839 46278
rect 26877 46275 26943 46278
rect 28901 46338 28967 46341
rect 29269 46338 29335 46341
rect 32121 46338 32187 46341
rect 28901 46336 32187 46338
rect 28901 46280 28906 46336
rect 28962 46280 29274 46336
rect 29330 46280 32126 46336
rect 32182 46280 32187 46336
rect 28901 46278 32187 46280
rect 28901 46275 28967 46278
rect 29269 46275 29335 46278
rect 32121 46275 32187 46278
rect 19568 46272 19888 46273
rect 19568 46208 19576 46272
rect 19640 46208 19656 46272
rect 19720 46208 19736 46272
rect 19800 46208 19816 46272
rect 19880 46208 19888 46272
rect 19568 46207 19888 46208
rect 3049 46202 3115 46205
rect 8845 46202 8911 46205
rect 3049 46200 8911 46202
rect 3049 46144 3054 46200
rect 3110 46144 8850 46200
rect 8906 46144 8911 46200
rect 3049 46142 8911 46144
rect 3049 46139 3115 46142
rect 8845 46139 8911 46142
rect 15694 46140 15700 46204
rect 15764 46202 15770 46204
rect 19333 46202 19399 46205
rect 15764 46200 19399 46202
rect 15764 46144 19338 46200
rect 19394 46144 19399 46200
rect 15764 46142 19399 46144
rect 15764 46140 15770 46142
rect 19333 46139 19399 46142
rect 28942 46140 28948 46204
rect 29012 46202 29018 46204
rect 32213 46202 32279 46205
rect 29012 46200 32279 46202
rect 29012 46144 32218 46200
rect 32274 46144 32279 46200
rect 29012 46142 32279 46144
rect 29012 46140 29018 46142
rect 32213 46139 32279 46142
rect 33041 46202 33107 46205
rect 34789 46202 34855 46205
rect 33041 46200 34855 46202
rect 33041 46144 33046 46200
rect 33102 46144 34794 46200
rect 34850 46144 34855 46200
rect 33041 46142 34855 46144
rect 33041 46139 33107 46142
rect 34789 46139 34855 46142
rect 1301 46066 1367 46069
rect 18045 46066 18111 46069
rect 1301 46064 18111 46066
rect 1301 46008 1306 46064
rect 1362 46008 18050 46064
rect 18106 46008 18111 46064
rect 1301 46006 18111 46008
rect 1301 46003 1367 46006
rect 18045 46003 18111 46006
rect 27429 46066 27495 46069
rect 28349 46066 28415 46069
rect 31109 46066 31175 46069
rect 27429 46064 31175 46066
rect 27429 46008 27434 46064
rect 27490 46008 28354 46064
rect 28410 46008 31114 46064
rect 31170 46008 31175 46064
rect 27429 46006 31175 46008
rect 27429 46003 27495 46006
rect 28349 46003 28415 46006
rect 31109 46003 31175 46006
rect 26233 45930 26299 45933
rect 26190 45928 26299 45930
rect 26190 45872 26238 45928
rect 26294 45872 26299 45928
rect 26190 45867 26299 45872
rect 27521 45930 27587 45933
rect 28073 45930 28139 45933
rect 32397 45930 32463 45933
rect 27521 45928 32463 45930
rect 27521 45872 27526 45928
rect 27582 45872 28078 45928
rect 28134 45872 32402 45928
rect 32458 45872 32463 45928
rect 27521 45870 32463 45872
rect 27521 45867 27587 45870
rect 28073 45867 28139 45870
rect 32397 45867 32463 45870
rect 25405 45794 25471 45797
rect 26190 45794 26250 45867
rect 28942 45794 28948 45796
rect 25405 45792 28948 45794
rect 25405 45736 25410 45792
rect 25466 45736 28948 45792
rect 25405 45734 28948 45736
rect 25405 45731 25471 45734
rect 28942 45732 28948 45734
rect 29012 45732 29018 45796
rect 4208 45728 4528 45729
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 45663 4528 45664
rect 34928 45728 35248 45729
rect 34928 45664 34936 45728
rect 35000 45664 35016 45728
rect 35080 45664 35096 45728
rect 35160 45664 35176 45728
rect 35240 45664 35248 45728
rect 34928 45663 35248 45664
rect 23933 45658 23999 45661
rect 29085 45658 29151 45661
rect 39200 45658 40000 45688
rect 23933 45656 29151 45658
rect 23933 45600 23938 45656
rect 23994 45600 29090 45656
rect 29146 45600 29151 45656
rect 23933 45598 29151 45600
rect 23933 45595 23999 45598
rect 29085 45595 29151 45598
rect 37782 45598 40000 45658
rect 14457 45522 14523 45525
rect 15561 45522 15627 45525
rect 14457 45520 15627 45522
rect 14457 45464 14462 45520
rect 14518 45464 15566 45520
rect 15622 45464 15627 45520
rect 14457 45462 15627 45464
rect 14457 45459 14523 45462
rect 15561 45459 15627 45462
rect 37641 45522 37707 45525
rect 37782 45522 37842 45598
rect 39200 45568 40000 45598
rect 37641 45520 37842 45522
rect 37641 45464 37646 45520
rect 37702 45464 37842 45520
rect 37641 45462 37842 45464
rect 37641 45459 37707 45462
rect 9857 45386 9923 45389
rect 27797 45386 27863 45389
rect 9857 45384 27863 45386
rect 9857 45328 9862 45384
rect 9918 45328 27802 45384
rect 27858 45328 27863 45384
rect 9857 45326 27863 45328
rect 9857 45323 9923 45326
rect 27797 45323 27863 45326
rect 19568 45184 19888 45185
rect 19568 45120 19576 45184
rect 19640 45120 19656 45184
rect 19720 45120 19736 45184
rect 19800 45120 19816 45184
rect 19880 45120 19888 45184
rect 19568 45119 19888 45120
rect 0 44978 800 45008
rect 8109 44978 8175 44981
rect 0 44976 8175 44978
rect 0 44920 8114 44976
rect 8170 44920 8175 44976
rect 0 44918 8175 44920
rect 0 44888 800 44918
rect 8109 44915 8175 44918
rect 28533 44978 28599 44981
rect 31201 44978 31267 44981
rect 28533 44976 31267 44978
rect 28533 44920 28538 44976
rect 28594 44920 31206 44976
rect 31262 44920 31267 44976
rect 28533 44918 31267 44920
rect 28533 44915 28599 44918
rect 31201 44915 31267 44918
rect 32949 44978 33015 44981
rect 39200 44978 40000 45008
rect 32949 44976 40000 44978
rect 32949 44920 32954 44976
rect 33010 44920 40000 44976
rect 32949 44918 40000 44920
rect 32949 44915 33015 44918
rect 39200 44888 40000 44918
rect 28625 44842 28691 44845
rect 31109 44842 31175 44845
rect 28625 44840 31175 44842
rect 28625 44784 28630 44840
rect 28686 44784 31114 44840
rect 31170 44784 31175 44840
rect 28625 44782 31175 44784
rect 28625 44779 28691 44782
rect 31109 44779 31175 44782
rect 25957 44706 26023 44709
rect 29085 44706 29151 44709
rect 25957 44704 29151 44706
rect 25957 44648 25962 44704
rect 26018 44648 29090 44704
rect 29146 44648 29151 44704
rect 25957 44646 29151 44648
rect 25957 44643 26023 44646
rect 29085 44643 29151 44646
rect 29729 44706 29795 44709
rect 31845 44706 31911 44709
rect 29729 44704 31911 44706
rect 29729 44648 29734 44704
rect 29790 44648 31850 44704
rect 31906 44648 31911 44704
rect 29729 44646 31911 44648
rect 29729 44643 29795 44646
rect 31845 44643 31911 44646
rect 4208 44640 4528 44641
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 44575 4528 44576
rect 34928 44640 35248 44641
rect 34928 44576 34936 44640
rect 35000 44576 35016 44640
rect 35080 44576 35096 44640
rect 35160 44576 35176 44640
rect 35240 44576 35248 44640
rect 34928 44575 35248 44576
rect 27889 44570 27955 44573
rect 31569 44570 31635 44573
rect 27889 44568 31635 44570
rect 27889 44512 27894 44568
rect 27950 44512 31574 44568
rect 31630 44512 31635 44568
rect 27889 44510 31635 44512
rect 27889 44507 27955 44510
rect 31569 44507 31635 44510
rect 17769 44434 17835 44437
rect 23565 44434 23631 44437
rect 17769 44432 23631 44434
rect 17769 44376 17774 44432
rect 17830 44376 23570 44432
rect 23626 44376 23631 44432
rect 17769 44374 23631 44376
rect 17769 44371 17835 44374
rect 23565 44371 23631 44374
rect 2037 44298 2103 44301
rect 8293 44298 8359 44301
rect 2037 44296 8359 44298
rect 2037 44240 2042 44296
rect 2098 44240 8298 44296
rect 8354 44240 8359 44296
rect 2037 44238 8359 44240
rect 2037 44235 2103 44238
rect 8293 44235 8359 44238
rect 24025 44298 24091 44301
rect 25957 44298 26023 44301
rect 26417 44298 26483 44301
rect 30741 44298 30807 44301
rect 24025 44296 30807 44298
rect 24025 44240 24030 44296
rect 24086 44240 25962 44296
rect 26018 44240 26422 44296
rect 26478 44240 30746 44296
rect 30802 44240 30807 44296
rect 24025 44238 30807 44240
rect 24025 44235 24091 44238
rect 25957 44235 26023 44238
rect 26417 44235 26483 44238
rect 30741 44235 30807 44238
rect 25497 44162 25563 44165
rect 29637 44162 29703 44165
rect 25497 44160 29703 44162
rect 25497 44104 25502 44160
rect 25558 44104 29642 44160
rect 29698 44104 29703 44160
rect 25497 44102 29703 44104
rect 25497 44099 25563 44102
rect 29637 44099 29703 44102
rect 19568 44096 19888 44097
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 44031 19888 44032
rect 24669 44026 24735 44029
rect 26325 44026 26391 44029
rect 28717 44026 28783 44029
rect 24669 44024 28783 44026
rect 24669 43968 24674 44024
rect 24730 43968 26330 44024
rect 26386 43968 28722 44024
rect 28778 43968 28783 44024
rect 24669 43966 28783 43968
rect 24669 43963 24735 43966
rect 26325 43963 26391 43966
rect 28717 43963 28783 43966
rect 28574 43890 28580 43892
rect 4064 43830 28580 43890
rect 0 43618 800 43648
rect 4064 43618 4124 43830
rect 28574 43828 28580 43830
rect 28644 43828 28650 43892
rect 9121 43754 9187 43757
rect 26601 43754 26667 43757
rect 9121 43752 26667 43754
rect 9121 43696 9126 43752
rect 9182 43696 26606 43752
rect 26662 43696 26667 43752
rect 9121 43694 26667 43696
rect 9121 43691 9187 43694
rect 26601 43691 26667 43694
rect 0 43558 4124 43618
rect 35341 43618 35407 43621
rect 39200 43618 40000 43648
rect 35341 43616 40000 43618
rect 35341 43560 35346 43616
rect 35402 43560 40000 43616
rect 35341 43558 40000 43560
rect 0 43528 800 43558
rect 35341 43555 35407 43558
rect 4208 43552 4528 43553
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 43487 4528 43488
rect 34928 43552 35248 43553
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 39200 43528 40000 43558
rect 34928 43487 35248 43488
rect 3049 43346 3115 43349
rect 27153 43346 27219 43349
rect 3049 43344 27219 43346
rect 3049 43288 3054 43344
rect 3110 43288 27158 43344
rect 27214 43288 27219 43344
rect 3049 43286 27219 43288
rect 3049 43283 3115 43286
rect 27153 43283 27219 43286
rect 19241 43210 19307 43213
rect 24669 43210 24735 43213
rect 19241 43208 24735 43210
rect 19241 43152 19246 43208
rect 19302 43152 24674 43208
rect 24730 43152 24735 43208
rect 19241 43150 24735 43152
rect 19241 43147 19307 43150
rect 24669 43147 24735 43150
rect 19568 43008 19888 43009
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 42943 19888 42944
rect 29453 42938 29519 42941
rect 34513 42938 34579 42941
rect 29453 42936 34579 42938
rect 29453 42880 29458 42936
rect 29514 42880 34518 42936
rect 34574 42880 34579 42936
rect 29453 42878 34579 42880
rect 29453 42875 29519 42878
rect 34513 42875 34579 42878
rect 29453 42802 29519 42805
rect 31385 42802 31451 42805
rect 35157 42802 35223 42805
rect 29453 42800 35223 42802
rect 29453 42744 29458 42800
rect 29514 42744 31390 42800
rect 31446 42744 35162 42800
rect 35218 42744 35223 42800
rect 29453 42742 35223 42744
rect 29453 42739 29519 42742
rect 31385 42739 31451 42742
rect 35157 42739 35223 42742
rect 12709 42666 12775 42669
rect 27838 42666 27844 42668
rect 12709 42664 27844 42666
rect 12709 42608 12714 42664
rect 12770 42608 27844 42664
rect 12709 42606 27844 42608
rect 12709 42603 12775 42606
rect 27838 42604 27844 42606
rect 27908 42604 27914 42668
rect 28717 42666 28783 42669
rect 34789 42666 34855 42669
rect 28717 42664 34855 42666
rect 28717 42608 28722 42664
rect 28778 42608 34794 42664
rect 34850 42608 34855 42664
rect 28717 42606 34855 42608
rect 28717 42603 28783 42606
rect 34789 42603 34855 42606
rect 4208 42464 4528 42465
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 42399 4528 42400
rect 34928 42464 35248 42465
rect 34928 42400 34936 42464
rect 35000 42400 35016 42464
rect 35080 42400 35096 42464
rect 35160 42400 35176 42464
rect 35240 42400 35248 42464
rect 34928 42399 35248 42400
rect 8845 42394 8911 42397
rect 18873 42394 18939 42397
rect 8845 42392 18939 42394
rect 8845 42336 8850 42392
rect 8906 42336 18878 42392
rect 18934 42336 18939 42392
rect 8845 42334 18939 42336
rect 8845 42331 8911 42334
rect 18873 42331 18939 42334
rect 28073 42394 28139 42397
rect 30833 42394 30899 42397
rect 28073 42392 30899 42394
rect 28073 42336 28078 42392
rect 28134 42336 30838 42392
rect 30894 42336 30899 42392
rect 28073 42334 30899 42336
rect 28073 42331 28139 42334
rect 30833 42331 30899 42334
rect 0 42258 800 42288
rect 39200 42258 40000 42288
rect 0 42198 1410 42258
rect 0 42168 800 42198
rect 1350 41714 1410 42198
rect 39070 42198 40000 42258
rect 19568 41920 19888 41921
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 41855 19888 41856
rect 5717 41850 5783 41853
rect 8937 41850 9003 41853
rect 5717 41848 9003 41850
rect 5717 41792 5722 41848
rect 5778 41792 8942 41848
rect 8998 41792 9003 41848
rect 5717 41790 9003 41792
rect 5717 41787 5783 41790
rect 8937 41787 9003 41790
rect 14365 41852 14431 41853
rect 28257 41852 28323 41853
rect 14365 41848 14412 41852
rect 14476 41850 14482 41852
rect 28206 41850 28212 41852
rect 14365 41792 14370 41848
rect 14365 41788 14412 41792
rect 14476 41790 14522 41850
rect 28166 41790 28212 41850
rect 28276 41848 28323 41852
rect 28318 41792 28323 41848
rect 14476 41788 14482 41790
rect 28206 41788 28212 41790
rect 28276 41788 28323 41792
rect 14365 41787 14431 41788
rect 28257 41787 28323 41788
rect 27521 41714 27587 41717
rect 1350 41712 27587 41714
rect 1350 41656 27526 41712
rect 27582 41656 27587 41712
rect 1350 41654 27587 41656
rect 27521 41651 27587 41654
rect 23749 41578 23815 41581
rect 39070 41578 39130 42198
rect 39200 42168 40000 42198
rect 23749 41576 39130 41578
rect 23749 41520 23754 41576
rect 23810 41520 39130 41576
rect 23749 41518 39130 41520
rect 23749 41515 23815 41518
rect 23381 41442 23447 41445
rect 23841 41442 23907 41445
rect 24853 41442 24919 41445
rect 23381 41440 24919 41442
rect 23381 41384 23386 41440
rect 23442 41384 23846 41440
rect 23902 41384 24858 41440
rect 24914 41384 24919 41440
rect 23381 41382 24919 41384
rect 23381 41379 23447 41382
rect 23841 41379 23907 41382
rect 24853 41379 24919 41382
rect 27245 41442 27311 41445
rect 27705 41442 27771 41445
rect 29545 41442 29611 41445
rect 27245 41440 29611 41442
rect 27245 41384 27250 41440
rect 27306 41384 27710 41440
rect 27766 41384 29550 41440
rect 29606 41384 29611 41440
rect 27245 41382 29611 41384
rect 27245 41379 27311 41382
rect 27705 41379 27771 41382
rect 29545 41379 29611 41382
rect 4208 41376 4528 41377
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 41311 4528 41312
rect 34928 41376 35248 41377
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 34928 41311 35248 41312
rect 29678 41244 29684 41308
rect 29748 41306 29754 41308
rect 29821 41306 29887 41309
rect 29748 41304 29887 41306
rect 29748 41248 29826 41304
rect 29882 41248 29887 41304
rect 29748 41246 29887 41248
rect 29748 41244 29754 41246
rect 29821 41243 29887 41246
rect 28349 41170 28415 41173
rect 35617 41170 35683 41173
rect 28349 41168 35683 41170
rect 28349 41112 28354 41168
rect 28410 41112 35622 41168
rect 35678 41112 35683 41168
rect 28349 41110 35683 41112
rect 28349 41107 28415 41110
rect 35617 41107 35683 41110
rect 21357 41034 21423 41037
rect 23473 41034 23539 41037
rect 21357 41032 23539 41034
rect 21357 40976 21362 41032
rect 21418 40976 23478 41032
rect 23534 40976 23539 41032
rect 21357 40974 23539 40976
rect 21357 40971 21423 40974
rect 23473 40971 23539 40974
rect 0 40898 800 40928
rect 3877 40898 3943 40901
rect 0 40896 3943 40898
rect 0 40840 3882 40896
rect 3938 40840 3943 40896
rect 0 40838 3943 40840
rect 0 40808 800 40838
rect 3877 40835 3943 40838
rect 12249 40898 12315 40901
rect 17309 40898 17375 40901
rect 12249 40896 17375 40898
rect 12249 40840 12254 40896
rect 12310 40840 17314 40896
rect 17370 40840 17375 40896
rect 12249 40838 17375 40840
rect 12249 40835 12315 40838
rect 17309 40835 17375 40838
rect 24761 40898 24827 40901
rect 29729 40898 29795 40901
rect 24761 40896 29795 40898
rect 24761 40840 24766 40896
rect 24822 40840 29734 40896
rect 29790 40840 29795 40896
rect 24761 40838 29795 40840
rect 24761 40835 24827 40838
rect 29729 40835 29795 40838
rect 34513 40898 34579 40901
rect 39200 40898 40000 40928
rect 34513 40896 40000 40898
rect 34513 40840 34518 40896
rect 34574 40840 40000 40896
rect 34513 40838 40000 40840
rect 34513 40835 34579 40838
rect 19568 40832 19888 40833
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 39200 40808 40000 40838
rect 19568 40767 19888 40768
rect 3785 40762 3851 40765
rect 19241 40762 19307 40765
rect 3785 40760 19307 40762
rect 3785 40704 3790 40760
rect 3846 40704 19246 40760
rect 19302 40704 19307 40760
rect 3785 40702 19307 40704
rect 3785 40699 3851 40702
rect 19241 40699 19307 40702
rect 24761 40762 24827 40765
rect 35525 40762 35591 40765
rect 24761 40760 35591 40762
rect 24761 40704 24766 40760
rect 24822 40704 35530 40760
rect 35586 40704 35591 40760
rect 24761 40702 35591 40704
rect 24761 40699 24827 40702
rect 35525 40699 35591 40702
rect 1945 40626 2011 40629
rect 3969 40626 4035 40629
rect 1945 40624 4035 40626
rect 1945 40568 1950 40624
rect 2006 40568 3974 40624
rect 4030 40568 4035 40624
rect 1945 40566 4035 40568
rect 1945 40563 2011 40566
rect 3969 40563 4035 40566
rect 17861 40626 17927 40629
rect 20713 40626 20779 40629
rect 35341 40626 35407 40629
rect 17861 40624 20779 40626
rect 17861 40568 17866 40624
rect 17922 40568 20718 40624
rect 20774 40568 20779 40624
rect 17861 40566 20779 40568
rect 17861 40563 17927 40566
rect 20713 40563 20779 40566
rect 22740 40624 35407 40626
rect 22740 40568 35346 40624
rect 35402 40568 35407 40624
rect 22740 40566 35407 40568
rect 13670 40428 13676 40492
rect 13740 40490 13746 40492
rect 22740 40490 22800 40566
rect 35341 40563 35407 40566
rect 13740 40456 22018 40490
rect 22142 40456 22800 40490
rect 13740 40430 22800 40456
rect 13740 40428 13746 40430
rect 21958 40396 22202 40430
rect 12617 40354 12683 40357
rect 13169 40354 13235 40357
rect 13997 40354 14063 40357
rect 12617 40352 14063 40354
rect 12617 40296 12622 40352
rect 12678 40296 13174 40352
rect 13230 40296 14002 40352
rect 14058 40296 14063 40352
rect 12617 40294 14063 40296
rect 12617 40291 12683 40294
rect 13169 40291 13235 40294
rect 13997 40291 14063 40294
rect 4208 40288 4528 40289
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 40223 4528 40224
rect 34928 40288 35248 40289
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 34928 40223 35248 40224
rect 17309 40218 17375 40221
rect 28717 40218 28783 40221
rect 17309 40216 28783 40218
rect 17309 40160 17314 40216
rect 17370 40160 28722 40216
rect 28778 40160 28783 40216
rect 17309 40158 28783 40160
rect 17309 40155 17375 40158
rect 28717 40155 28783 40158
rect 16481 40082 16547 40085
rect 18229 40082 18295 40085
rect 16481 40080 18295 40082
rect 16481 40024 16486 40080
rect 16542 40024 18234 40080
rect 18290 40024 18295 40080
rect 16481 40022 18295 40024
rect 16481 40019 16547 40022
rect 18229 40019 18295 40022
rect 25405 40082 25471 40085
rect 28257 40082 28323 40085
rect 25405 40080 28323 40082
rect 25405 40024 25410 40080
rect 25466 40024 28262 40080
rect 28318 40024 28323 40080
rect 25405 40022 28323 40024
rect 25405 40019 25471 40022
rect 28257 40019 28323 40022
rect 10225 39946 10291 39949
rect 13077 39946 13143 39949
rect 10225 39944 13143 39946
rect 10225 39888 10230 39944
rect 10286 39888 13082 39944
rect 13138 39888 13143 39944
rect 10225 39886 13143 39888
rect 10225 39883 10291 39886
rect 13077 39883 13143 39886
rect 17861 39946 17927 39949
rect 19701 39946 19767 39949
rect 17861 39944 19767 39946
rect 17861 39888 17866 39944
rect 17922 39888 19706 39944
rect 19762 39888 19767 39944
rect 17861 39886 19767 39888
rect 17861 39883 17927 39886
rect 19701 39883 19767 39886
rect 14825 39810 14891 39813
rect 18597 39810 18663 39813
rect 14825 39808 18663 39810
rect 14825 39752 14830 39808
rect 14886 39752 18602 39808
rect 18658 39752 18663 39808
rect 14825 39750 18663 39752
rect 14825 39747 14891 39750
rect 18597 39747 18663 39750
rect 19568 39744 19888 39745
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 19568 39679 19888 39680
rect 4061 39674 4127 39677
rect 19057 39674 19123 39677
rect 4061 39672 19123 39674
rect 4061 39616 4066 39672
rect 4122 39616 19062 39672
rect 19118 39616 19123 39672
rect 4061 39614 19123 39616
rect 4061 39611 4127 39614
rect 19057 39611 19123 39614
rect 0 39538 800 39568
rect 1577 39538 1643 39541
rect 0 39536 1643 39538
rect 0 39480 1582 39536
rect 1638 39480 1643 39536
rect 0 39478 1643 39480
rect 0 39448 800 39478
rect 1577 39475 1643 39478
rect 34789 39538 34855 39541
rect 39200 39538 40000 39568
rect 34789 39536 40000 39538
rect 34789 39480 34794 39536
rect 34850 39480 40000 39536
rect 34789 39478 40000 39480
rect 34789 39475 34855 39478
rect 39200 39448 40000 39478
rect 3877 39402 3943 39405
rect 9397 39402 9463 39405
rect 3877 39400 9463 39402
rect 3877 39344 3882 39400
rect 3938 39344 9402 39400
rect 9458 39344 9463 39400
rect 3877 39342 9463 39344
rect 3877 39339 3943 39342
rect 9397 39339 9463 39342
rect 4208 39200 4528 39201
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 39135 4528 39136
rect 34928 39200 35248 39201
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 39135 35248 39136
rect 16665 38858 16731 38861
rect 21633 38858 21699 38861
rect 16665 38856 21699 38858
rect 16665 38800 16670 38856
rect 16726 38800 21638 38856
rect 21694 38800 21699 38856
rect 16665 38798 21699 38800
rect 16665 38795 16731 38798
rect 21633 38795 21699 38798
rect 25773 38858 25839 38861
rect 26969 38858 27035 38861
rect 25773 38856 27035 38858
rect 25773 38800 25778 38856
rect 25834 38800 26974 38856
rect 27030 38800 27035 38856
rect 25773 38798 27035 38800
rect 25773 38795 25839 38798
rect 26969 38795 27035 38798
rect 15878 38660 15884 38724
rect 15948 38722 15954 38724
rect 18689 38722 18755 38725
rect 15948 38720 18755 38722
rect 15948 38664 18694 38720
rect 18750 38664 18755 38720
rect 15948 38662 18755 38664
rect 15948 38660 15954 38662
rect 18689 38659 18755 38662
rect 23105 38722 23171 38725
rect 26141 38722 26207 38725
rect 23105 38720 26207 38722
rect 23105 38664 23110 38720
rect 23166 38664 26146 38720
rect 26202 38664 26207 38720
rect 23105 38662 26207 38664
rect 23105 38659 23171 38662
rect 26141 38659 26207 38662
rect 19568 38656 19888 38657
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 19568 38591 19888 38592
rect 15101 38586 15167 38589
rect 16849 38586 16915 38589
rect 15101 38584 16915 38586
rect 15101 38528 15106 38584
rect 15162 38528 16854 38584
rect 16910 38528 16915 38584
rect 15101 38526 16915 38528
rect 15101 38523 15167 38526
rect 16849 38523 16915 38526
rect 14365 38450 14431 38453
rect 16757 38450 16823 38453
rect 28073 38452 28139 38453
rect 14365 38448 16823 38450
rect 14365 38392 14370 38448
rect 14426 38392 16762 38448
rect 16818 38392 16823 38448
rect 14365 38390 16823 38392
rect 14365 38387 14431 38390
rect 16757 38387 16823 38390
rect 28022 38388 28028 38452
rect 28092 38450 28139 38452
rect 28092 38448 28184 38450
rect 28134 38392 28184 38448
rect 28092 38390 28184 38392
rect 28092 38388 28139 38390
rect 28073 38387 28139 38388
rect 13537 38314 13603 38317
rect 16481 38314 16547 38317
rect 18781 38314 18847 38317
rect 13537 38312 18847 38314
rect 13537 38256 13542 38312
rect 13598 38256 16486 38312
rect 16542 38256 18786 38312
rect 18842 38256 18847 38312
rect 13537 38254 18847 38256
rect 13537 38251 13603 38254
rect 16481 38251 16547 38254
rect 18781 38251 18847 38254
rect 21081 38314 21147 38317
rect 34697 38314 34763 38317
rect 21081 38312 34763 38314
rect 21081 38256 21086 38312
rect 21142 38256 34702 38312
rect 34758 38256 34763 38312
rect 21081 38254 34763 38256
rect 21081 38251 21147 38254
rect 34697 38251 34763 38254
rect 0 38178 800 38208
rect 2773 38178 2839 38181
rect 0 38176 2839 38178
rect 0 38120 2778 38176
rect 2834 38120 2839 38176
rect 0 38118 2839 38120
rect 0 38088 800 38118
rect 2773 38115 2839 38118
rect 35617 38178 35683 38181
rect 39200 38178 40000 38208
rect 35617 38176 40000 38178
rect 35617 38120 35622 38176
rect 35678 38120 40000 38176
rect 35617 38118 40000 38120
rect 35617 38115 35683 38118
rect 4208 38112 4528 38113
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 38047 4528 38048
rect 34928 38112 35248 38113
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 39200 38088 40000 38118
rect 34928 38047 35248 38048
rect 17401 38042 17467 38045
rect 19793 38042 19859 38045
rect 17401 38040 19859 38042
rect 17401 37984 17406 38040
rect 17462 37984 19798 38040
rect 19854 37984 19859 38040
rect 17401 37982 19859 37984
rect 17401 37979 17467 37982
rect 19793 37979 19859 37982
rect 21633 38042 21699 38045
rect 27838 38042 27844 38044
rect 21633 38040 27844 38042
rect 21633 37984 21638 38040
rect 21694 37984 27844 38040
rect 21633 37982 27844 37984
rect 21633 37979 21699 37982
rect 27838 37980 27844 37982
rect 27908 38042 27914 38044
rect 30465 38042 30531 38045
rect 27908 38040 30531 38042
rect 27908 37984 30470 38040
rect 30526 37984 30531 38040
rect 27908 37982 30531 37984
rect 27908 37980 27914 37982
rect 30465 37979 30531 37982
rect 3509 37906 3575 37909
rect 14825 37906 14891 37909
rect 3509 37904 14891 37906
rect 3509 37848 3514 37904
rect 3570 37848 14830 37904
rect 14886 37848 14891 37904
rect 3509 37846 14891 37848
rect 3509 37843 3575 37846
rect 14825 37843 14891 37846
rect 15009 37906 15075 37909
rect 16573 37906 16639 37909
rect 18321 37906 18387 37909
rect 15009 37904 18387 37906
rect 15009 37848 15014 37904
rect 15070 37848 16578 37904
rect 16634 37848 18326 37904
rect 18382 37848 18387 37904
rect 15009 37846 18387 37848
rect 15009 37843 15075 37846
rect 16573 37843 16639 37846
rect 18321 37843 18387 37846
rect 18597 37906 18663 37909
rect 20989 37906 21055 37909
rect 21541 37906 21607 37909
rect 18597 37904 21607 37906
rect 18597 37848 18602 37904
rect 18658 37848 20994 37904
rect 21050 37848 21546 37904
rect 21602 37848 21607 37904
rect 18597 37846 21607 37848
rect 18597 37843 18663 37846
rect 20989 37843 21055 37846
rect 21541 37843 21607 37846
rect 15469 37770 15535 37773
rect 16941 37770 17007 37773
rect 17166 37770 17172 37772
rect 15469 37768 17172 37770
rect 15469 37712 15474 37768
rect 15530 37712 16946 37768
rect 17002 37712 17172 37768
rect 15469 37710 17172 37712
rect 15469 37707 15535 37710
rect 16941 37707 17007 37710
rect 17166 37708 17172 37710
rect 17236 37708 17242 37772
rect 18965 37770 19031 37773
rect 22737 37770 22803 37773
rect 18965 37768 22803 37770
rect 18965 37712 18970 37768
rect 19026 37712 22742 37768
rect 22798 37712 22803 37768
rect 18965 37710 22803 37712
rect 18965 37707 19031 37710
rect 22737 37707 22803 37710
rect 20069 37634 20135 37637
rect 23749 37634 23815 37637
rect 20069 37632 23815 37634
rect 20069 37576 20074 37632
rect 20130 37576 23754 37632
rect 23810 37576 23815 37632
rect 20069 37574 23815 37576
rect 20069 37571 20135 37574
rect 23749 37571 23815 37574
rect 19568 37568 19888 37569
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 37503 19888 37504
rect 15101 37498 15167 37501
rect 16941 37498 17007 37501
rect 15101 37496 17007 37498
rect 15101 37440 15106 37496
rect 15162 37440 16946 37496
rect 17002 37440 17007 37496
rect 15101 37438 17007 37440
rect 15101 37435 15167 37438
rect 16941 37435 17007 37438
rect 17309 37498 17375 37501
rect 20805 37498 20871 37501
rect 26785 37498 26851 37501
rect 17309 37496 19442 37498
rect 17309 37440 17314 37496
rect 17370 37440 19442 37496
rect 17309 37438 19442 37440
rect 17309 37435 17375 37438
rect 3693 37362 3759 37365
rect 11329 37362 11395 37365
rect 3693 37360 11395 37362
rect 3693 37304 3698 37360
rect 3754 37304 11334 37360
rect 11390 37304 11395 37360
rect 3693 37302 11395 37304
rect 3693 37299 3759 37302
rect 11329 37299 11395 37302
rect 13721 37362 13787 37365
rect 18413 37362 18479 37365
rect 13721 37360 18479 37362
rect 13721 37304 13726 37360
rect 13782 37304 18418 37360
rect 18474 37304 18479 37360
rect 13721 37302 18479 37304
rect 19382 37362 19442 37438
rect 20805 37496 26851 37498
rect 20805 37440 20810 37496
rect 20866 37440 26790 37496
rect 26846 37440 26851 37496
rect 20805 37438 26851 37440
rect 20805 37435 20871 37438
rect 26785 37435 26851 37438
rect 21633 37362 21699 37365
rect 19382 37360 21699 37362
rect 19382 37304 21638 37360
rect 21694 37304 21699 37360
rect 19382 37302 21699 37304
rect 13721 37299 13787 37302
rect 18413 37299 18479 37302
rect 21633 37299 21699 37302
rect 24342 37300 24348 37364
rect 24412 37362 24418 37364
rect 24485 37362 24551 37365
rect 24412 37360 24551 37362
rect 24412 37304 24490 37360
rect 24546 37304 24551 37360
rect 24412 37302 24551 37304
rect 24412 37300 24418 37302
rect 24485 37299 24551 37302
rect 29453 37362 29519 37365
rect 31293 37362 31359 37365
rect 29453 37360 31359 37362
rect 29453 37304 29458 37360
rect 29514 37304 31298 37360
rect 31354 37304 31359 37360
rect 29453 37302 31359 37304
rect 29453 37299 29519 37302
rect 31293 37299 31359 37302
rect 16849 37226 16915 37229
rect 20253 37226 20319 37229
rect 16849 37224 20319 37226
rect 16849 37168 16854 37224
rect 16910 37168 20258 37224
rect 20314 37168 20319 37224
rect 16849 37166 20319 37168
rect 16849 37163 16915 37166
rect 20253 37163 20319 37166
rect 20897 37226 20963 37229
rect 22277 37226 22343 37229
rect 20897 37224 22343 37226
rect 20897 37168 20902 37224
rect 20958 37168 22282 37224
rect 22338 37168 22343 37224
rect 20897 37166 22343 37168
rect 20897 37163 20963 37166
rect 22277 37163 22343 37166
rect 28809 37226 28875 37229
rect 35525 37226 35591 37229
rect 28809 37224 35591 37226
rect 28809 37168 28814 37224
rect 28870 37168 35530 37224
rect 35586 37168 35591 37224
rect 28809 37166 35591 37168
rect 28809 37163 28875 37166
rect 35525 37163 35591 37166
rect 14089 37090 14155 37093
rect 14733 37090 14799 37093
rect 18781 37090 18847 37093
rect 14089 37088 18847 37090
rect 14089 37032 14094 37088
rect 14150 37032 14738 37088
rect 14794 37032 18786 37088
rect 18842 37032 18847 37088
rect 14089 37030 18847 37032
rect 14089 37027 14155 37030
rect 14733 37027 14799 37030
rect 18781 37027 18847 37030
rect 4208 37024 4528 37025
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36959 4528 36960
rect 34928 37024 35248 37025
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36959 35248 36960
rect 9029 36954 9095 36957
rect 13997 36954 14063 36957
rect 9029 36952 14063 36954
rect 9029 36896 9034 36952
rect 9090 36896 14002 36952
rect 14058 36896 14063 36952
rect 9029 36894 14063 36896
rect 9029 36891 9095 36894
rect 13997 36891 14063 36894
rect 0 36818 800 36848
rect 3049 36818 3115 36821
rect 0 36816 3115 36818
rect 0 36760 3054 36816
rect 3110 36760 3115 36816
rect 0 36758 3115 36760
rect 0 36728 800 36758
rect 3049 36755 3115 36758
rect 12985 36818 13051 36821
rect 16205 36818 16271 36821
rect 12985 36816 16271 36818
rect 12985 36760 12990 36816
rect 13046 36760 16210 36816
rect 16266 36760 16271 36816
rect 12985 36758 16271 36760
rect 12985 36755 13051 36758
rect 16205 36755 16271 36758
rect 22829 36818 22895 36821
rect 28073 36818 28139 36821
rect 22829 36816 28139 36818
rect 22829 36760 22834 36816
rect 22890 36760 28078 36816
rect 28134 36760 28139 36816
rect 22829 36758 28139 36760
rect 22829 36755 22895 36758
rect 28073 36755 28139 36758
rect 32581 36818 32647 36821
rect 39200 36818 40000 36848
rect 32581 36816 40000 36818
rect 32581 36760 32586 36816
rect 32642 36760 40000 36816
rect 32581 36758 40000 36760
rect 32581 36755 32647 36758
rect 39200 36728 40000 36758
rect 10961 36682 11027 36685
rect 14917 36682 14983 36685
rect 15929 36682 15995 36685
rect 10961 36680 15995 36682
rect 10961 36624 10966 36680
rect 11022 36624 14922 36680
rect 14978 36624 15934 36680
rect 15990 36624 15995 36680
rect 10961 36622 15995 36624
rect 10961 36619 11027 36622
rect 14917 36619 14983 36622
rect 15929 36619 15995 36622
rect 25681 36682 25747 36685
rect 33041 36682 33107 36685
rect 25681 36680 33107 36682
rect 25681 36624 25686 36680
rect 25742 36624 33046 36680
rect 33102 36624 33107 36680
rect 25681 36622 33107 36624
rect 25681 36619 25747 36622
rect 33041 36619 33107 36622
rect 2957 36546 3023 36549
rect 8661 36546 8727 36549
rect 2957 36544 8727 36546
rect 2957 36488 2962 36544
rect 3018 36488 8666 36544
rect 8722 36488 8727 36544
rect 2957 36486 8727 36488
rect 2957 36483 3023 36486
rect 8661 36483 8727 36486
rect 13537 36546 13603 36549
rect 14181 36546 14247 36549
rect 15193 36546 15259 36549
rect 13537 36544 15259 36546
rect 13537 36488 13542 36544
rect 13598 36488 14186 36544
rect 14242 36488 15198 36544
rect 15254 36488 15259 36544
rect 13537 36486 15259 36488
rect 13537 36483 13603 36486
rect 14181 36483 14247 36486
rect 15193 36483 15259 36486
rect 19568 36480 19888 36481
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 36415 19888 36416
rect 9305 36410 9371 36413
rect 15193 36410 15259 36413
rect 9305 36408 15259 36410
rect 9305 36352 9310 36408
rect 9366 36352 15198 36408
rect 15254 36352 15259 36408
rect 9305 36350 15259 36352
rect 9305 36347 9371 36350
rect 15193 36347 15259 36350
rect 17125 36410 17191 36413
rect 19333 36410 19399 36413
rect 17125 36408 19399 36410
rect 17125 36352 17130 36408
rect 17186 36352 19338 36408
rect 19394 36352 19399 36408
rect 17125 36350 19399 36352
rect 17125 36347 17191 36350
rect 19333 36347 19399 36350
rect 27429 36410 27495 36413
rect 29545 36410 29611 36413
rect 27429 36408 29611 36410
rect 27429 36352 27434 36408
rect 27490 36352 29550 36408
rect 29606 36352 29611 36408
rect 27429 36350 29611 36352
rect 27429 36347 27495 36350
rect 29545 36347 29611 36350
rect 11329 36274 11395 36277
rect 15285 36274 15351 36277
rect 16665 36274 16731 36277
rect 11329 36272 16731 36274
rect 11329 36216 11334 36272
rect 11390 36216 15290 36272
rect 15346 36216 16670 36272
rect 16726 36216 16731 36272
rect 11329 36214 16731 36216
rect 11329 36211 11395 36214
rect 15285 36211 15351 36214
rect 16665 36211 16731 36214
rect 17861 36274 17927 36277
rect 18597 36274 18663 36277
rect 20897 36274 20963 36277
rect 17861 36272 20963 36274
rect 17861 36216 17866 36272
rect 17922 36216 18602 36272
rect 18658 36216 20902 36272
rect 20958 36216 20963 36272
rect 17861 36214 20963 36216
rect 17861 36211 17927 36214
rect 18597 36211 18663 36214
rect 20897 36211 20963 36214
rect 23238 36212 23244 36276
rect 23308 36274 23314 36276
rect 23381 36274 23447 36277
rect 23308 36272 23447 36274
rect 23308 36216 23386 36272
rect 23442 36216 23447 36272
rect 23308 36214 23447 36216
rect 23308 36212 23314 36214
rect 23381 36211 23447 36214
rect 3877 36138 3943 36141
rect 9622 36138 9628 36140
rect 3877 36136 9628 36138
rect 3877 36080 3882 36136
rect 3938 36080 9628 36136
rect 3877 36078 9628 36080
rect 3877 36075 3943 36078
rect 9622 36076 9628 36078
rect 9692 36076 9698 36140
rect 18045 36138 18111 36141
rect 22369 36138 22435 36141
rect 18045 36136 22435 36138
rect 18045 36080 18050 36136
rect 18106 36080 22374 36136
rect 22430 36080 22435 36136
rect 18045 36078 22435 36080
rect 18045 36075 18111 36078
rect 22369 36075 22435 36078
rect 12249 36002 12315 36005
rect 16481 36002 16547 36005
rect 19333 36002 19399 36005
rect 12249 36000 19399 36002
rect 12249 35944 12254 36000
rect 12310 35944 16486 36000
rect 16542 35944 19338 36000
rect 19394 35944 19399 36000
rect 12249 35942 19399 35944
rect 12249 35939 12315 35942
rect 16481 35939 16547 35942
rect 19333 35939 19399 35942
rect 4208 35936 4528 35937
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 35871 4528 35872
rect 34928 35936 35248 35937
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 35871 35248 35872
rect 10777 35866 10843 35869
rect 15929 35866 15995 35869
rect 16665 35866 16731 35869
rect 10777 35864 16731 35866
rect 10777 35808 10782 35864
rect 10838 35808 15934 35864
rect 15990 35808 16670 35864
rect 16726 35808 16731 35864
rect 10777 35806 16731 35808
rect 10777 35803 10843 35806
rect 15929 35803 15995 35806
rect 16665 35803 16731 35806
rect 19149 35866 19215 35869
rect 22645 35866 22711 35869
rect 19149 35864 22711 35866
rect 19149 35808 19154 35864
rect 19210 35808 22650 35864
rect 22706 35808 22711 35864
rect 19149 35806 22711 35808
rect 19149 35803 19215 35806
rect 22645 35803 22711 35806
rect 27061 35866 27127 35869
rect 28533 35866 28599 35869
rect 27061 35864 28599 35866
rect 27061 35808 27066 35864
rect 27122 35808 28538 35864
rect 28594 35808 28599 35864
rect 27061 35806 28599 35808
rect 27061 35803 27127 35806
rect 28533 35803 28599 35806
rect 10961 35730 11027 35733
rect 16297 35730 16363 35733
rect 10961 35728 16363 35730
rect 10961 35672 10966 35728
rect 11022 35672 16302 35728
rect 16358 35672 16363 35728
rect 10961 35670 16363 35672
rect 10961 35667 11027 35670
rect 16297 35667 16363 35670
rect 16757 35730 16823 35733
rect 21081 35730 21147 35733
rect 16757 35728 21147 35730
rect 16757 35672 16762 35728
rect 16818 35672 21086 35728
rect 21142 35672 21147 35728
rect 16757 35670 21147 35672
rect 16757 35667 16823 35670
rect 21081 35667 21147 35670
rect 11697 35594 11763 35597
rect 14365 35594 14431 35597
rect 11697 35592 14431 35594
rect 11697 35536 11702 35592
rect 11758 35536 14370 35592
rect 14426 35536 14431 35592
rect 11697 35534 14431 35536
rect 11697 35531 11763 35534
rect 14365 35531 14431 35534
rect 16573 35594 16639 35597
rect 20989 35594 21055 35597
rect 16573 35592 21055 35594
rect 16573 35536 16578 35592
rect 16634 35536 20994 35592
rect 21050 35536 21055 35592
rect 16573 35534 21055 35536
rect 16573 35531 16639 35534
rect 20989 35531 21055 35534
rect 0 35458 800 35488
rect 3785 35458 3851 35461
rect 0 35456 3851 35458
rect 0 35400 3790 35456
rect 3846 35400 3851 35456
rect 0 35398 3851 35400
rect 0 35368 800 35398
rect 3785 35395 3851 35398
rect 14641 35458 14707 35461
rect 17125 35458 17191 35461
rect 14641 35456 17191 35458
rect 14641 35400 14646 35456
rect 14702 35400 17130 35456
rect 17186 35400 17191 35456
rect 14641 35398 17191 35400
rect 14641 35395 14707 35398
rect 17125 35395 17191 35398
rect 35433 35458 35499 35461
rect 39200 35458 40000 35488
rect 35433 35456 40000 35458
rect 35433 35400 35438 35456
rect 35494 35400 40000 35456
rect 35433 35398 40000 35400
rect 35433 35395 35499 35398
rect 19568 35392 19888 35393
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 39200 35368 40000 35398
rect 19568 35327 19888 35328
rect 8937 35186 9003 35189
rect 11145 35186 11211 35189
rect 14641 35186 14707 35189
rect 8937 35184 14707 35186
rect 8937 35128 8942 35184
rect 8998 35128 11150 35184
rect 11206 35128 14646 35184
rect 14702 35128 14707 35184
rect 8937 35126 14707 35128
rect 8937 35123 9003 35126
rect 11145 35123 11211 35126
rect 14641 35123 14707 35126
rect 15193 35186 15259 35189
rect 16573 35186 16639 35189
rect 19333 35186 19399 35189
rect 15193 35184 19399 35186
rect 15193 35128 15198 35184
rect 15254 35128 16578 35184
rect 16634 35128 19338 35184
rect 19394 35128 19399 35184
rect 15193 35126 19399 35128
rect 15193 35123 15259 35126
rect 16573 35123 16639 35126
rect 19333 35123 19399 35126
rect 11881 35050 11947 35053
rect 14958 35050 14964 35052
rect 11881 35048 14964 35050
rect 11881 34992 11886 35048
rect 11942 34992 14964 35048
rect 11881 34990 14964 34992
rect 11881 34987 11947 34990
rect 14958 34988 14964 34990
rect 15028 34988 15034 35052
rect 16205 35050 16271 35053
rect 20069 35050 20135 35053
rect 16205 35048 20135 35050
rect 16205 34992 16210 35048
rect 16266 34992 20074 35048
rect 20130 34992 20135 35048
rect 16205 34990 20135 34992
rect 16205 34987 16271 34990
rect 20069 34987 20135 34990
rect 10133 34914 10199 34917
rect 16389 34914 16455 34917
rect 20069 34914 20135 34917
rect 10133 34912 20135 34914
rect 10133 34856 10138 34912
rect 10194 34856 16394 34912
rect 16450 34856 20074 34912
rect 20130 34856 20135 34912
rect 10133 34854 20135 34856
rect 10133 34851 10199 34854
rect 16389 34851 16455 34854
rect 20069 34851 20135 34854
rect 20897 34914 20963 34917
rect 23841 34914 23907 34917
rect 20897 34912 23907 34914
rect 20897 34856 20902 34912
rect 20958 34856 23846 34912
rect 23902 34856 23907 34912
rect 20897 34854 23907 34856
rect 20897 34851 20963 34854
rect 23841 34851 23907 34854
rect 4208 34848 4528 34849
rect 0 34778 800 34808
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 34783 4528 34784
rect 34928 34848 35248 34849
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 34783 35248 34784
rect 3877 34778 3943 34781
rect 0 34776 3943 34778
rect 0 34720 3882 34776
rect 3938 34720 3943 34776
rect 0 34718 3943 34720
rect 0 34688 800 34718
rect 3877 34715 3943 34718
rect 10041 34778 10107 34781
rect 14222 34778 14228 34780
rect 10041 34776 14228 34778
rect 10041 34720 10046 34776
rect 10102 34720 14228 34776
rect 10041 34718 14228 34720
rect 10041 34715 10107 34718
rect 14222 34716 14228 34718
rect 14292 34778 14298 34780
rect 14917 34778 14983 34781
rect 14292 34776 14983 34778
rect 14292 34720 14922 34776
rect 14978 34720 14983 34776
rect 14292 34718 14983 34720
rect 14292 34716 14298 34718
rect 14917 34715 14983 34718
rect 16297 34778 16363 34781
rect 19609 34778 19675 34781
rect 16297 34776 19675 34778
rect 16297 34720 16302 34776
rect 16358 34720 19614 34776
rect 19670 34720 19675 34776
rect 16297 34718 19675 34720
rect 16297 34715 16363 34718
rect 19609 34715 19675 34718
rect 24669 34778 24735 34781
rect 25865 34778 25931 34781
rect 24669 34776 25931 34778
rect 24669 34720 24674 34776
rect 24730 34720 25870 34776
rect 25926 34720 25931 34776
rect 24669 34718 25931 34720
rect 24669 34715 24735 34718
rect 25865 34715 25931 34718
rect 12801 34642 12867 34645
rect 13905 34644 13971 34645
rect 13118 34642 13124 34644
rect 12801 34640 13124 34642
rect 12801 34584 12806 34640
rect 12862 34584 13124 34640
rect 12801 34582 13124 34584
rect 12801 34579 12867 34582
rect 13118 34580 13124 34582
rect 13188 34580 13194 34644
rect 13854 34642 13860 34644
rect 13814 34582 13860 34642
rect 13924 34640 13971 34644
rect 13966 34584 13971 34640
rect 13854 34580 13860 34582
rect 13924 34580 13971 34584
rect 13905 34579 13971 34580
rect 14825 34642 14891 34645
rect 16389 34642 16455 34645
rect 18321 34642 18387 34645
rect 20805 34642 20871 34645
rect 14825 34640 16314 34642
rect 14825 34584 14830 34640
rect 14886 34584 16314 34640
rect 14825 34582 16314 34584
rect 14825 34579 14891 34582
rect 8334 34444 8340 34508
rect 8404 34506 8410 34508
rect 8477 34506 8543 34509
rect 8404 34504 8543 34506
rect 8404 34448 8482 34504
rect 8538 34448 8543 34504
rect 8404 34446 8543 34448
rect 16254 34506 16314 34582
rect 16389 34640 20871 34642
rect 16389 34584 16394 34640
rect 16450 34584 18326 34640
rect 18382 34584 20810 34640
rect 20866 34584 20871 34640
rect 16389 34582 20871 34584
rect 16389 34579 16455 34582
rect 18321 34579 18387 34582
rect 20805 34579 20871 34582
rect 21357 34642 21423 34645
rect 25037 34642 25103 34645
rect 21357 34640 25103 34642
rect 21357 34584 21362 34640
rect 21418 34584 25042 34640
rect 25098 34584 25103 34640
rect 21357 34582 25103 34584
rect 21357 34579 21423 34582
rect 25037 34579 25103 34582
rect 16757 34506 16823 34509
rect 16254 34504 16823 34506
rect 16254 34448 16762 34504
rect 16818 34448 16823 34504
rect 16254 34446 16823 34448
rect 8404 34444 8410 34446
rect 8477 34443 8543 34446
rect 16757 34443 16823 34446
rect 17769 34506 17835 34509
rect 20529 34506 20595 34509
rect 20897 34506 20963 34509
rect 17769 34504 20963 34506
rect 17769 34448 17774 34504
rect 17830 34448 20534 34504
rect 20590 34448 20902 34504
rect 20958 34448 20963 34504
rect 17769 34446 20963 34448
rect 17769 34443 17835 34446
rect 20529 34443 20595 34446
rect 20897 34443 20963 34446
rect 14958 34308 14964 34372
rect 15028 34370 15034 34372
rect 16798 34370 16804 34372
rect 15028 34310 16804 34370
rect 15028 34308 15034 34310
rect 16798 34308 16804 34310
rect 16868 34370 16874 34372
rect 17953 34370 18019 34373
rect 16868 34368 18019 34370
rect 16868 34312 17958 34368
rect 18014 34312 18019 34368
rect 16868 34310 18019 34312
rect 16868 34308 16874 34310
rect 17953 34307 18019 34310
rect 19977 34370 20043 34373
rect 20662 34370 20668 34372
rect 19977 34368 20668 34370
rect 19977 34312 19982 34368
rect 20038 34312 20668 34368
rect 19977 34310 20668 34312
rect 19977 34307 20043 34310
rect 20662 34308 20668 34310
rect 20732 34370 20738 34372
rect 22093 34370 22159 34373
rect 20732 34368 22159 34370
rect 20732 34312 22098 34368
rect 22154 34312 22159 34368
rect 20732 34310 22159 34312
rect 20732 34308 20738 34310
rect 22093 34307 22159 34310
rect 19568 34304 19888 34305
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 34239 19888 34240
rect 12566 34172 12572 34236
rect 12636 34234 12642 34236
rect 19333 34234 19399 34237
rect 12636 34232 19399 34234
rect 12636 34176 19338 34232
rect 19394 34176 19399 34232
rect 12636 34174 19399 34176
rect 12636 34172 12642 34174
rect 19333 34171 19399 34174
rect 20110 34172 20116 34236
rect 20180 34234 20186 34236
rect 20345 34234 20411 34237
rect 20180 34232 20411 34234
rect 20180 34176 20350 34232
rect 20406 34176 20411 34232
rect 20180 34174 20411 34176
rect 20180 34172 20186 34174
rect 20345 34171 20411 34174
rect 27613 34234 27679 34237
rect 35433 34234 35499 34237
rect 27613 34232 35499 34234
rect 27613 34176 27618 34232
rect 27674 34176 35438 34232
rect 35494 34176 35499 34232
rect 27613 34174 35499 34176
rect 27613 34171 27679 34174
rect 35433 34171 35499 34174
rect 10593 34098 10659 34101
rect 13537 34098 13603 34101
rect 10593 34096 13603 34098
rect 10593 34040 10598 34096
rect 10654 34040 13542 34096
rect 13598 34040 13603 34096
rect 10593 34038 13603 34040
rect 10593 34035 10659 34038
rect 13537 34035 13603 34038
rect 15929 34098 15995 34101
rect 17953 34098 18019 34101
rect 15929 34096 18019 34098
rect 15929 34040 15934 34096
rect 15990 34040 17958 34096
rect 18014 34040 18019 34096
rect 15929 34038 18019 34040
rect 15929 34035 15995 34038
rect 17953 34035 18019 34038
rect 32397 34098 32463 34101
rect 39200 34098 40000 34128
rect 32397 34096 40000 34098
rect 32397 34040 32402 34096
rect 32458 34040 40000 34096
rect 32397 34038 40000 34040
rect 32397 34035 32463 34038
rect 39200 34008 40000 34038
rect 8569 33962 8635 33965
rect 10961 33962 11027 33965
rect 8569 33960 11027 33962
rect 8569 33904 8574 33960
rect 8630 33904 10966 33960
rect 11022 33904 11027 33960
rect 8569 33902 11027 33904
rect 8569 33899 8635 33902
rect 10961 33899 11027 33902
rect 11881 33962 11947 33965
rect 14825 33962 14891 33965
rect 11881 33960 14891 33962
rect 11881 33904 11886 33960
rect 11942 33904 14830 33960
rect 14886 33904 14891 33960
rect 11881 33902 14891 33904
rect 11881 33899 11947 33902
rect 14825 33899 14891 33902
rect 15837 33962 15903 33965
rect 19425 33962 19491 33965
rect 15837 33960 19491 33962
rect 15837 33904 15842 33960
rect 15898 33904 19430 33960
rect 19486 33904 19491 33960
rect 15837 33902 19491 33904
rect 15837 33899 15903 33902
rect 19425 33899 19491 33902
rect 19609 33962 19675 33965
rect 25313 33962 25379 33965
rect 19609 33960 25379 33962
rect 19609 33904 19614 33960
rect 19670 33904 25318 33960
rect 25374 33904 25379 33960
rect 19609 33902 25379 33904
rect 19609 33899 19675 33902
rect 25313 33899 25379 33902
rect 6729 33826 6795 33829
rect 8477 33826 8543 33829
rect 6729 33824 8543 33826
rect 6729 33768 6734 33824
rect 6790 33768 8482 33824
rect 8538 33768 8543 33824
rect 6729 33766 8543 33768
rect 6729 33763 6795 33766
rect 8477 33763 8543 33766
rect 9397 33826 9463 33829
rect 11513 33826 11579 33829
rect 16849 33826 16915 33829
rect 9397 33824 16915 33826
rect 9397 33768 9402 33824
rect 9458 33768 11518 33824
rect 11574 33768 16854 33824
rect 16910 33768 16915 33824
rect 9397 33766 16915 33768
rect 9397 33763 9463 33766
rect 11513 33763 11579 33766
rect 16849 33763 16915 33766
rect 21725 33826 21791 33829
rect 27429 33826 27495 33829
rect 21725 33824 27495 33826
rect 21725 33768 21730 33824
rect 21786 33768 27434 33824
rect 27490 33768 27495 33824
rect 21725 33766 27495 33768
rect 21725 33763 21791 33766
rect 27429 33763 27495 33766
rect 4208 33760 4528 33761
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 33695 4528 33696
rect 34928 33760 35248 33761
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 33695 35248 33696
rect 10501 33690 10567 33693
rect 12801 33690 12867 33693
rect 10501 33688 12867 33690
rect 10501 33632 10506 33688
rect 10562 33632 12806 33688
rect 12862 33632 12867 33688
rect 10501 33630 12867 33632
rect 10501 33627 10567 33630
rect 12801 33627 12867 33630
rect 13537 33690 13603 33693
rect 14365 33690 14431 33693
rect 13537 33688 14431 33690
rect 13537 33632 13542 33688
rect 13598 33632 14370 33688
rect 14426 33632 14431 33688
rect 13537 33630 14431 33632
rect 13537 33627 13603 33630
rect 14365 33627 14431 33630
rect 14825 33690 14891 33693
rect 16062 33690 16068 33692
rect 14825 33688 16068 33690
rect 14825 33632 14830 33688
rect 14886 33632 16068 33688
rect 14825 33630 16068 33632
rect 14825 33627 14891 33630
rect 16062 33628 16068 33630
rect 16132 33690 16138 33692
rect 18689 33690 18755 33693
rect 20713 33690 20779 33693
rect 16132 33688 20779 33690
rect 16132 33632 18694 33688
rect 18750 33632 20718 33688
rect 20774 33632 20779 33688
rect 16132 33630 20779 33632
rect 16132 33628 16138 33630
rect 18689 33627 18755 33630
rect 20713 33627 20779 33630
rect 21633 33690 21699 33693
rect 25589 33690 25655 33693
rect 26049 33690 26115 33693
rect 30649 33690 30715 33693
rect 21633 33688 30715 33690
rect 21633 33632 21638 33688
rect 21694 33632 25594 33688
rect 25650 33632 26054 33688
rect 26110 33632 30654 33688
rect 30710 33632 30715 33688
rect 21633 33630 30715 33632
rect 21633 33627 21699 33630
rect 25589 33627 25655 33630
rect 26049 33627 26115 33630
rect 30649 33627 30715 33630
rect 9581 33554 9647 33557
rect 12525 33554 12591 33557
rect 9581 33552 12591 33554
rect 9581 33496 9586 33552
rect 9642 33496 12530 33552
rect 12586 33496 12591 33552
rect 9581 33494 12591 33496
rect 9581 33491 9647 33494
rect 12525 33491 12591 33494
rect 18321 33554 18387 33557
rect 22461 33554 22527 33557
rect 18321 33552 22527 33554
rect 18321 33496 18326 33552
rect 18382 33496 22466 33552
rect 22522 33496 22527 33552
rect 18321 33494 22527 33496
rect 18321 33491 18387 33494
rect 22461 33491 22527 33494
rect 0 33418 800 33448
rect 11881 33418 11947 33421
rect 14273 33418 14339 33421
rect 0 33328 858 33418
rect 11881 33416 14339 33418
rect 11881 33360 11886 33416
rect 11942 33360 14278 33416
rect 14334 33360 14339 33416
rect 11881 33358 14339 33360
rect 11881 33355 11947 33358
rect 14273 33355 14339 33358
rect 14641 33418 14707 33421
rect 16297 33418 16363 33421
rect 20989 33418 21055 33421
rect 14641 33416 15348 33418
rect 14641 33360 14646 33416
rect 14702 33360 15348 33416
rect 14641 33358 15348 33360
rect 14641 33355 14707 33358
rect 798 33010 858 33328
rect 15288 33282 15348 33358
rect 16297 33416 21055 33418
rect 16297 33360 16302 33416
rect 16358 33360 20994 33416
rect 21050 33360 21055 33416
rect 16297 33358 21055 33360
rect 16297 33355 16363 33358
rect 20989 33355 21055 33358
rect 22001 33418 22067 33421
rect 25037 33418 25103 33421
rect 22001 33416 25103 33418
rect 22001 33360 22006 33416
rect 22062 33360 25042 33416
rect 25098 33360 25103 33416
rect 22001 33358 25103 33360
rect 22001 33355 22067 33358
rect 25037 33355 25103 33358
rect 35525 33418 35591 33421
rect 39200 33418 40000 33448
rect 35525 33416 40000 33418
rect 35525 33360 35530 33416
rect 35586 33360 40000 33416
rect 35525 33358 40000 33360
rect 35525 33355 35591 33358
rect 39200 33328 40000 33358
rect 19149 33282 19215 33285
rect 15288 33280 19215 33282
rect 15288 33224 19154 33280
rect 19210 33224 19215 33280
rect 15288 33222 19215 33224
rect 19149 33219 19215 33222
rect 20529 33282 20595 33285
rect 23105 33282 23171 33285
rect 20529 33280 23171 33282
rect 20529 33224 20534 33280
rect 20590 33224 23110 33280
rect 23166 33224 23171 33280
rect 20529 33222 23171 33224
rect 20529 33219 20595 33222
rect 23105 33219 23171 33222
rect 19568 33216 19888 33217
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 33151 19888 33152
rect 8753 33146 8819 33149
rect 13486 33146 13492 33148
rect 8753 33144 13492 33146
rect 8753 33088 8758 33144
rect 8814 33088 13492 33144
rect 8753 33086 13492 33088
rect 8753 33083 8819 33086
rect 13486 33084 13492 33086
rect 13556 33146 13562 33148
rect 13905 33146 13971 33149
rect 13556 33144 13971 33146
rect 13556 33088 13910 33144
rect 13966 33088 13971 33144
rect 13556 33086 13971 33088
rect 13556 33084 13562 33086
rect 13905 33083 13971 33086
rect 20713 33146 20779 33149
rect 21449 33146 21515 33149
rect 20713 33144 21515 33146
rect 20713 33088 20718 33144
rect 20774 33088 21454 33144
rect 21510 33088 21515 33144
rect 20713 33086 21515 33088
rect 20713 33083 20779 33086
rect 21449 33083 21515 33086
rect 9857 33010 9923 33013
rect 798 33008 9923 33010
rect 798 32952 9862 33008
rect 9918 32952 9923 33008
rect 798 32950 9923 32952
rect 9857 32947 9923 32950
rect 11145 33010 11211 33013
rect 11421 33010 11487 33013
rect 11145 33008 11487 33010
rect 11145 32952 11150 33008
rect 11206 32952 11426 33008
rect 11482 32952 11487 33008
rect 11145 32950 11487 32952
rect 11145 32947 11211 32950
rect 11421 32947 11487 32950
rect 12157 33010 12223 33013
rect 17677 33010 17743 33013
rect 12157 33008 17743 33010
rect 12157 32952 12162 33008
rect 12218 32952 17682 33008
rect 17738 32952 17743 33008
rect 12157 32950 17743 32952
rect 12157 32947 12223 32950
rect 17677 32947 17743 32950
rect 17953 33010 18019 33013
rect 18689 33010 18755 33013
rect 25589 33010 25655 33013
rect 17953 33008 25655 33010
rect 17953 32952 17958 33008
rect 18014 32952 18694 33008
rect 18750 32952 25594 33008
rect 25650 32952 25655 33008
rect 17953 32950 25655 32952
rect 17953 32947 18019 32950
rect 18689 32947 18755 32950
rect 25589 32947 25655 32950
rect 28901 33010 28967 33013
rect 32673 33010 32739 33013
rect 28901 33008 32739 33010
rect 28901 32952 28906 33008
rect 28962 32952 32678 33008
rect 32734 32952 32739 33008
rect 28901 32950 32739 32952
rect 28901 32947 28967 32950
rect 32673 32947 32739 32950
rect 8109 32874 8175 32877
rect 11053 32874 11119 32877
rect 11697 32874 11763 32877
rect 12709 32874 12775 32877
rect 8109 32872 11119 32874
rect 8109 32816 8114 32872
rect 8170 32816 11058 32872
rect 11114 32816 11119 32872
rect 8109 32814 11119 32816
rect 8109 32811 8175 32814
rect 11053 32811 11119 32814
rect 11286 32872 12775 32874
rect 11286 32816 11702 32872
rect 11758 32816 12714 32872
rect 12770 32816 12775 32872
rect 11286 32814 12775 32816
rect 7741 32738 7807 32741
rect 8569 32738 8635 32741
rect 8753 32738 8819 32741
rect 11286 32738 11346 32814
rect 11697 32811 11763 32814
rect 12709 32811 12775 32814
rect 13077 32874 13143 32877
rect 18045 32874 18111 32877
rect 13077 32872 18111 32874
rect 13077 32816 13082 32872
rect 13138 32816 18050 32872
rect 18106 32816 18111 32872
rect 13077 32814 18111 32816
rect 13077 32811 13143 32814
rect 18045 32811 18111 32814
rect 18781 32874 18847 32877
rect 23657 32874 23723 32877
rect 18781 32872 23723 32874
rect 18781 32816 18786 32872
rect 18842 32816 23662 32872
rect 23718 32816 23723 32872
rect 18781 32814 23723 32816
rect 18781 32811 18847 32814
rect 23657 32811 23723 32814
rect 7741 32736 11346 32738
rect 7741 32680 7746 32736
rect 7802 32680 8574 32736
rect 8630 32680 8758 32736
rect 8814 32680 11346 32736
rect 7741 32678 11346 32680
rect 12065 32738 12131 32741
rect 15285 32738 15351 32741
rect 12065 32736 15351 32738
rect 12065 32680 12070 32736
rect 12126 32680 15290 32736
rect 15346 32680 15351 32736
rect 12065 32678 15351 32680
rect 7741 32675 7807 32678
rect 8569 32675 8635 32678
rect 8753 32675 8819 32678
rect 12065 32675 12131 32678
rect 15285 32675 15351 32678
rect 20805 32738 20871 32741
rect 21173 32738 21239 32741
rect 20805 32736 21239 32738
rect 20805 32680 20810 32736
rect 20866 32680 21178 32736
rect 21234 32680 21239 32736
rect 20805 32678 21239 32680
rect 20805 32675 20871 32678
rect 21173 32675 21239 32678
rect 4208 32672 4528 32673
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 32607 4528 32608
rect 34928 32672 35248 32673
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 32607 35248 32608
rect 9213 32602 9279 32605
rect 9581 32602 9647 32605
rect 10869 32602 10935 32605
rect 9213 32600 10935 32602
rect 9213 32544 9218 32600
rect 9274 32544 9586 32600
rect 9642 32544 10874 32600
rect 10930 32544 10935 32600
rect 9213 32542 10935 32544
rect 9213 32539 9279 32542
rect 9581 32539 9647 32542
rect 10869 32539 10935 32542
rect 11697 32602 11763 32605
rect 16021 32602 16087 32605
rect 11697 32600 16087 32602
rect 11697 32544 11702 32600
rect 11758 32544 16026 32600
rect 16082 32544 16087 32600
rect 11697 32542 16087 32544
rect 11697 32539 11763 32542
rect 16021 32539 16087 32542
rect 18781 32602 18847 32605
rect 21725 32602 21791 32605
rect 18781 32600 21791 32602
rect 18781 32544 18786 32600
rect 18842 32544 21730 32600
rect 21786 32544 21791 32600
rect 18781 32542 21791 32544
rect 18781 32539 18847 32542
rect 21725 32539 21791 32542
rect 10961 32466 11027 32469
rect 15326 32466 15332 32468
rect 10961 32464 15332 32466
rect 10961 32408 10966 32464
rect 11022 32408 15332 32464
rect 10961 32406 15332 32408
rect 10961 32403 11027 32406
rect 15326 32404 15332 32406
rect 15396 32404 15402 32468
rect 18321 32466 18387 32469
rect 24853 32466 24919 32469
rect 18321 32464 24919 32466
rect 18321 32408 18326 32464
rect 18382 32408 24858 32464
rect 24914 32408 24919 32464
rect 18321 32406 24919 32408
rect 18321 32403 18387 32406
rect 24853 32403 24919 32406
rect 10869 32330 10935 32333
rect 15837 32330 15903 32333
rect 21541 32330 21607 32333
rect 10869 32328 15903 32330
rect 10869 32272 10874 32328
rect 10930 32272 15842 32328
rect 15898 32272 15903 32328
rect 10869 32270 15903 32272
rect 10869 32267 10935 32270
rect 15837 32267 15903 32270
rect 20854 32328 21607 32330
rect 20854 32272 21546 32328
rect 21602 32272 21607 32328
rect 20854 32270 21607 32272
rect 9673 32194 9739 32197
rect 11605 32194 11671 32197
rect 9673 32192 11671 32194
rect 9673 32136 9678 32192
rect 9734 32136 11610 32192
rect 11666 32136 11671 32192
rect 9673 32134 11671 32136
rect 9673 32131 9739 32134
rect 11605 32131 11671 32134
rect 11881 32194 11947 32197
rect 16573 32194 16639 32197
rect 11881 32192 16639 32194
rect 11881 32136 11886 32192
rect 11942 32136 16578 32192
rect 16634 32136 16639 32192
rect 11881 32134 16639 32136
rect 11881 32131 11947 32134
rect 16573 32131 16639 32134
rect 20621 32194 20687 32197
rect 20854 32194 20914 32270
rect 21541 32267 21607 32270
rect 23238 32268 23244 32332
rect 23308 32330 23314 32332
rect 23933 32330 23999 32333
rect 23308 32328 23999 32330
rect 23308 32272 23938 32328
rect 23994 32272 23999 32328
rect 23308 32270 23999 32272
rect 23308 32268 23314 32270
rect 23933 32267 23999 32270
rect 24209 32330 24275 32333
rect 26785 32330 26851 32333
rect 26969 32330 27035 32333
rect 24209 32328 27035 32330
rect 24209 32272 24214 32328
rect 24270 32272 26790 32328
rect 26846 32272 26974 32328
rect 27030 32272 27035 32328
rect 24209 32270 27035 32272
rect 24209 32267 24275 32270
rect 26785 32267 26851 32270
rect 26969 32267 27035 32270
rect 20621 32192 20914 32194
rect 20621 32136 20626 32192
rect 20682 32136 20914 32192
rect 20621 32134 20914 32136
rect 20989 32194 21055 32197
rect 22921 32194 22987 32197
rect 20989 32192 22987 32194
rect 20989 32136 20994 32192
rect 21050 32136 22926 32192
rect 22982 32136 22987 32192
rect 20989 32134 22987 32136
rect 20621 32131 20687 32134
rect 20989 32131 21055 32134
rect 22921 32131 22987 32134
rect 23657 32194 23723 32197
rect 23790 32194 23796 32196
rect 23657 32192 23796 32194
rect 23657 32136 23662 32192
rect 23718 32136 23796 32192
rect 23657 32134 23796 32136
rect 23657 32131 23723 32134
rect 23790 32132 23796 32134
rect 23860 32132 23866 32196
rect 19568 32128 19888 32129
rect 0 32058 800 32088
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 32063 19888 32064
rect 3325 32058 3391 32061
rect 0 32056 3391 32058
rect 0 32000 3330 32056
rect 3386 32000 3391 32056
rect 0 31998 3391 32000
rect 0 31968 800 31998
rect 3325 31995 3391 31998
rect 12249 32058 12315 32061
rect 13813 32058 13879 32061
rect 14825 32058 14891 32061
rect 18781 32058 18847 32061
rect 12249 32056 13879 32058
rect 12249 32000 12254 32056
rect 12310 32000 13818 32056
rect 13874 32000 13879 32056
rect 12249 31998 13879 32000
rect 12249 31995 12315 31998
rect 13813 31995 13879 31998
rect 14230 32056 18847 32058
rect 14230 32000 14830 32056
rect 14886 32000 18786 32056
rect 18842 32000 18847 32056
rect 14230 31998 18847 32000
rect 7557 31922 7623 31925
rect 9857 31922 9923 31925
rect 7557 31920 9923 31922
rect 7557 31864 7562 31920
rect 7618 31864 9862 31920
rect 9918 31864 9923 31920
rect 7557 31862 9923 31864
rect 7557 31859 7623 31862
rect 9857 31859 9923 31862
rect 7649 31786 7715 31789
rect 11329 31786 11395 31789
rect 14230 31786 14290 31998
rect 14825 31995 14891 31998
rect 18781 31995 18847 31998
rect 22921 32058 22987 32061
rect 23289 32058 23355 32061
rect 26325 32058 26391 32061
rect 22921 32056 23122 32058
rect 22921 32000 22926 32056
rect 22982 32000 23122 32056
rect 22921 31998 23122 32000
rect 22921 31995 22987 31998
rect 14365 31922 14431 31925
rect 18321 31922 18387 31925
rect 22829 31922 22895 31925
rect 14365 31920 22895 31922
rect 14365 31864 14370 31920
rect 14426 31864 18326 31920
rect 18382 31864 22834 31920
rect 22890 31864 22895 31920
rect 14365 31862 22895 31864
rect 23062 31922 23122 31998
rect 23289 32056 26391 32058
rect 23289 32000 23294 32056
rect 23350 32000 26330 32056
rect 26386 32000 26391 32056
rect 23289 31998 26391 32000
rect 23289 31995 23355 31998
rect 26325 31995 26391 31998
rect 28073 32058 28139 32061
rect 39200 32058 40000 32088
rect 28073 32056 40000 32058
rect 28073 32000 28078 32056
rect 28134 32000 40000 32056
rect 28073 31998 40000 32000
rect 28073 31995 28139 31998
rect 39200 31968 40000 31998
rect 25589 31922 25655 31925
rect 23062 31920 25655 31922
rect 23062 31864 25594 31920
rect 25650 31864 25655 31920
rect 23062 31862 25655 31864
rect 14365 31859 14431 31862
rect 18321 31859 18387 31862
rect 22829 31859 22895 31862
rect 25589 31859 25655 31862
rect 7649 31784 11395 31786
rect 7649 31728 7654 31784
rect 7710 31728 11334 31784
rect 11390 31728 11395 31784
rect 7649 31726 11395 31728
rect 7649 31723 7715 31726
rect 11329 31723 11395 31726
rect 13678 31726 14290 31786
rect 14917 31786 14983 31789
rect 15101 31786 15167 31789
rect 14917 31784 15167 31786
rect 14917 31728 14922 31784
rect 14978 31728 15106 31784
rect 15162 31728 15167 31784
rect 14917 31726 15167 31728
rect 10593 31650 10659 31653
rect 12893 31650 12959 31653
rect 10593 31648 12959 31650
rect 10593 31592 10598 31648
rect 10654 31592 12898 31648
rect 12954 31592 12959 31648
rect 10593 31590 12959 31592
rect 10593 31587 10659 31590
rect 12893 31587 12959 31590
rect 13261 31650 13327 31653
rect 13678 31650 13738 31726
rect 14917 31723 14983 31726
rect 15101 31723 15167 31726
rect 15837 31786 15903 31789
rect 16021 31786 16087 31789
rect 18229 31786 18295 31789
rect 15837 31784 18295 31786
rect 15837 31728 15842 31784
rect 15898 31728 16026 31784
rect 16082 31728 18234 31784
rect 18290 31728 18295 31784
rect 15837 31726 18295 31728
rect 15837 31723 15903 31726
rect 16021 31723 16087 31726
rect 18229 31723 18295 31726
rect 18413 31786 18479 31789
rect 20989 31786 21055 31789
rect 18413 31784 21055 31786
rect 18413 31728 18418 31784
rect 18474 31728 20994 31784
rect 21050 31728 21055 31784
rect 18413 31726 21055 31728
rect 18413 31723 18479 31726
rect 20989 31723 21055 31726
rect 26417 31786 26483 31789
rect 28901 31786 28967 31789
rect 30557 31786 30623 31789
rect 26417 31784 30623 31786
rect 26417 31728 26422 31784
rect 26478 31728 28906 31784
rect 28962 31728 30562 31784
rect 30618 31728 30623 31784
rect 26417 31726 30623 31728
rect 26417 31723 26483 31726
rect 28901 31723 28967 31726
rect 30557 31723 30623 31726
rect 14273 31652 14339 31653
rect 16021 31652 16087 31653
rect 14222 31650 14228 31652
rect 13261 31648 13738 31650
rect 13261 31592 13266 31648
rect 13322 31592 13738 31648
rect 13261 31590 13738 31592
rect 14182 31590 14228 31650
rect 14292 31648 14339 31652
rect 14334 31592 14339 31648
rect 13261 31587 13327 31590
rect 14222 31588 14228 31590
rect 14292 31588 14339 31592
rect 14958 31588 14964 31652
rect 15028 31650 15034 31652
rect 15326 31650 15332 31652
rect 15028 31590 15332 31650
rect 15028 31588 15034 31590
rect 15326 31588 15332 31590
rect 15396 31588 15402 31652
rect 16021 31650 16068 31652
rect 15976 31648 16068 31650
rect 15976 31592 16026 31648
rect 15976 31590 16068 31592
rect 16021 31588 16068 31590
rect 16132 31588 16138 31652
rect 16757 31650 16823 31653
rect 22921 31650 22987 31653
rect 16254 31648 22987 31650
rect 16254 31592 16762 31648
rect 16818 31592 22926 31648
rect 22982 31592 22987 31648
rect 16254 31590 22987 31592
rect 14273 31587 14339 31588
rect 16021 31587 16087 31588
rect 4208 31584 4528 31585
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 31519 4528 31520
rect 9489 31514 9555 31517
rect 12249 31514 12315 31517
rect 9489 31512 12315 31514
rect 9489 31456 9494 31512
rect 9550 31456 12254 31512
rect 12310 31456 12315 31512
rect 9489 31454 12315 31456
rect 9489 31451 9555 31454
rect 12249 31451 12315 31454
rect 15101 31514 15167 31517
rect 16254 31514 16314 31590
rect 16757 31587 16823 31590
rect 22921 31587 22987 31590
rect 23238 31588 23244 31652
rect 23308 31650 23314 31652
rect 23565 31650 23631 31653
rect 23308 31648 23631 31650
rect 23308 31592 23570 31648
rect 23626 31592 23631 31648
rect 23308 31590 23631 31592
rect 23308 31588 23314 31590
rect 23565 31587 23631 31590
rect 27153 31650 27219 31653
rect 27521 31650 27587 31653
rect 27153 31648 27587 31650
rect 27153 31592 27158 31648
rect 27214 31592 27526 31648
rect 27582 31592 27587 31648
rect 27153 31590 27587 31592
rect 27153 31587 27219 31590
rect 27521 31587 27587 31590
rect 34928 31584 35248 31585
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 31519 35248 31520
rect 15101 31512 16314 31514
rect 15101 31456 15106 31512
rect 15162 31456 16314 31512
rect 15101 31454 16314 31456
rect 16849 31514 16915 31517
rect 18505 31514 18571 31517
rect 19885 31514 19951 31517
rect 16849 31512 19951 31514
rect 16849 31456 16854 31512
rect 16910 31456 18510 31512
rect 18566 31456 19890 31512
rect 19946 31456 19951 31512
rect 16849 31454 19951 31456
rect 15101 31451 15167 31454
rect 16849 31451 16915 31454
rect 18505 31451 18571 31454
rect 19885 31451 19951 31454
rect 23749 31514 23815 31517
rect 28717 31514 28783 31517
rect 23749 31512 28783 31514
rect 23749 31456 23754 31512
rect 23810 31456 28722 31512
rect 28778 31456 28783 31512
rect 23749 31454 28783 31456
rect 23749 31451 23815 31454
rect 28717 31451 28783 31454
rect 15469 31378 15535 31381
rect 18873 31378 18939 31381
rect 15469 31376 18939 31378
rect 15469 31320 15474 31376
rect 15530 31320 18878 31376
rect 18934 31320 18939 31376
rect 15469 31318 18939 31320
rect 15469 31315 15535 31318
rect 18873 31315 18939 31318
rect 21449 31378 21515 31381
rect 21582 31378 21588 31380
rect 21449 31376 21588 31378
rect 21449 31320 21454 31376
rect 21510 31320 21588 31376
rect 21449 31318 21588 31320
rect 21449 31315 21515 31318
rect 21582 31316 21588 31318
rect 21652 31316 21658 31380
rect 25037 31378 25103 31381
rect 26509 31378 26575 31381
rect 27245 31378 27311 31381
rect 25037 31376 27311 31378
rect 25037 31320 25042 31376
rect 25098 31320 26514 31376
rect 26570 31320 27250 31376
rect 27306 31320 27311 31376
rect 25037 31318 27311 31320
rect 25037 31315 25103 31318
rect 26509 31315 26575 31318
rect 27245 31315 27311 31318
rect 7005 31242 7071 31245
rect 10777 31242 10843 31245
rect 11973 31242 12039 31245
rect 7005 31240 12039 31242
rect 7005 31184 7010 31240
rect 7066 31184 10782 31240
rect 10838 31184 11978 31240
rect 12034 31184 12039 31240
rect 7005 31182 12039 31184
rect 7005 31179 7071 31182
rect 10777 31179 10843 31182
rect 11973 31179 12039 31182
rect 12157 31242 12223 31245
rect 19609 31242 19675 31245
rect 19885 31242 19951 31245
rect 12157 31240 19951 31242
rect 12157 31184 12162 31240
rect 12218 31184 19614 31240
rect 19670 31184 19890 31240
rect 19946 31184 19951 31240
rect 12157 31182 19951 31184
rect 12157 31179 12223 31182
rect 19609 31179 19675 31182
rect 19885 31179 19951 31182
rect 23105 31242 23171 31245
rect 23105 31240 25376 31242
rect 23105 31184 23110 31240
rect 23166 31184 25376 31240
rect 23105 31182 25376 31184
rect 23105 31179 23171 31182
rect 25316 31109 25376 31182
rect 7465 31106 7531 31109
rect 8017 31106 8083 31109
rect 10961 31106 11027 31109
rect 7465 31104 11027 31106
rect 7465 31048 7470 31104
rect 7526 31048 8022 31104
rect 8078 31048 10966 31104
rect 11022 31048 11027 31104
rect 7465 31046 11027 31048
rect 7465 31043 7531 31046
rect 8017 31043 8083 31046
rect 10961 31043 11027 31046
rect 12249 31106 12315 31109
rect 16389 31106 16455 31109
rect 12249 31104 16455 31106
rect 12249 31048 12254 31104
rect 12310 31048 16394 31104
rect 16450 31048 16455 31104
rect 12249 31046 16455 31048
rect 12249 31043 12315 31046
rect 16389 31043 16455 31046
rect 20345 31106 20411 31109
rect 24853 31106 24919 31109
rect 20345 31104 24919 31106
rect 20345 31048 20350 31104
rect 20406 31048 24858 31104
rect 24914 31048 24919 31104
rect 20345 31046 24919 31048
rect 20345 31043 20411 31046
rect 24853 31043 24919 31046
rect 25313 31104 25379 31109
rect 25313 31048 25318 31104
rect 25374 31048 25379 31104
rect 25313 31043 25379 31048
rect 19568 31040 19888 31041
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 30975 19888 30976
rect 12525 30972 12591 30973
rect 12525 30968 12572 30972
rect 12636 30970 12642 30972
rect 12525 30912 12530 30968
rect 12525 30908 12572 30912
rect 12636 30910 12682 30970
rect 12636 30908 12642 30910
rect 12525 30907 12591 30908
rect 7741 30834 7807 30837
rect 11237 30834 11303 30837
rect 7741 30832 11303 30834
rect 7741 30776 7746 30832
rect 7802 30776 11242 30832
rect 11298 30776 11303 30832
rect 7741 30774 11303 30776
rect 7741 30771 7807 30774
rect 11237 30771 11303 30774
rect 11881 30834 11947 30837
rect 14825 30834 14891 30837
rect 15745 30834 15811 30837
rect 11881 30832 15811 30834
rect 11881 30776 11886 30832
rect 11942 30776 14830 30832
rect 14886 30776 15750 30832
rect 15806 30776 15811 30832
rect 11881 30774 15811 30776
rect 11881 30771 11947 30774
rect 14825 30771 14891 30774
rect 15745 30771 15811 30774
rect 19977 30834 20043 30837
rect 26601 30834 26667 30837
rect 19977 30832 26667 30834
rect 19977 30776 19982 30832
rect 20038 30776 26606 30832
rect 26662 30776 26667 30832
rect 19977 30774 26667 30776
rect 19977 30771 20043 30774
rect 26601 30771 26667 30774
rect 28533 30834 28599 30837
rect 28533 30832 39130 30834
rect 28533 30776 28538 30832
rect 28594 30776 39130 30832
rect 28533 30774 39130 30776
rect 28533 30771 28599 30774
rect 0 30698 800 30728
rect 4061 30698 4127 30701
rect 0 30696 4127 30698
rect 0 30640 4066 30696
rect 4122 30640 4127 30696
rect 0 30638 4127 30640
rect 0 30608 800 30638
rect 4061 30635 4127 30638
rect 9489 30698 9555 30701
rect 11789 30698 11855 30701
rect 12709 30698 12775 30701
rect 9489 30696 11855 30698
rect 9489 30640 9494 30696
rect 9550 30640 11794 30696
rect 11850 30640 11855 30696
rect 9489 30638 11855 30640
rect 9489 30635 9555 30638
rect 11789 30635 11855 30638
rect 12022 30696 12775 30698
rect 12022 30640 12714 30696
rect 12770 30640 12775 30696
rect 12022 30638 12775 30640
rect 9581 30562 9647 30565
rect 12022 30562 12082 30638
rect 12709 30635 12775 30638
rect 12893 30698 12959 30701
rect 13118 30698 13124 30700
rect 12893 30696 13124 30698
rect 12893 30640 12898 30696
rect 12954 30640 13124 30696
rect 12893 30638 13124 30640
rect 12893 30635 12959 30638
rect 13118 30636 13124 30638
rect 13188 30636 13194 30700
rect 13486 30636 13492 30700
rect 13556 30698 13562 30700
rect 14917 30698 14983 30701
rect 18597 30698 18663 30701
rect 13556 30696 14983 30698
rect 13556 30640 14922 30696
rect 14978 30640 14983 30696
rect 13556 30638 14983 30640
rect 13556 30636 13562 30638
rect 14917 30635 14983 30638
rect 17542 30696 18663 30698
rect 17542 30640 18602 30696
rect 18658 30640 18663 30696
rect 17542 30638 18663 30640
rect 13077 30562 13143 30565
rect 9581 30560 12082 30562
rect 9581 30504 9586 30560
rect 9642 30504 12082 30560
rect 9581 30502 12082 30504
rect 12206 30560 13143 30562
rect 12206 30504 13082 30560
rect 13138 30504 13143 30560
rect 12206 30502 13143 30504
rect 9581 30499 9647 30502
rect 4208 30496 4528 30497
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 30431 4528 30432
rect 10961 30426 11027 30429
rect 12206 30426 12266 30502
rect 13077 30499 13143 30502
rect 13537 30562 13603 30565
rect 17542 30562 17602 30638
rect 18597 30635 18663 30638
rect 19057 30698 19123 30701
rect 21357 30698 21423 30701
rect 19057 30696 21423 30698
rect 19057 30640 19062 30696
rect 19118 30640 21362 30696
rect 21418 30640 21423 30696
rect 19057 30638 21423 30640
rect 19057 30635 19123 30638
rect 21357 30635 21423 30638
rect 22001 30698 22067 30701
rect 25405 30698 25471 30701
rect 22001 30696 25471 30698
rect 22001 30640 22006 30696
rect 22062 30640 25410 30696
rect 25466 30640 25471 30696
rect 22001 30638 25471 30640
rect 39070 30698 39130 30774
rect 39200 30698 40000 30728
rect 39070 30638 40000 30698
rect 22001 30635 22067 30638
rect 25405 30635 25471 30638
rect 39200 30608 40000 30638
rect 13537 30560 17602 30562
rect 13537 30504 13542 30560
rect 13598 30504 17602 30560
rect 13537 30502 17602 30504
rect 17677 30562 17743 30565
rect 18413 30562 18479 30565
rect 17677 30560 18479 30562
rect 17677 30504 17682 30560
rect 17738 30504 18418 30560
rect 18474 30504 18479 30560
rect 17677 30502 18479 30504
rect 13537 30499 13603 30502
rect 17677 30499 17743 30502
rect 18413 30499 18479 30502
rect 21449 30562 21515 30565
rect 21449 30560 23306 30562
rect 21449 30504 21454 30560
rect 21510 30504 23306 30560
rect 21449 30502 23306 30504
rect 21449 30499 21515 30502
rect 10961 30424 12266 30426
rect 10961 30368 10966 30424
rect 11022 30368 12266 30424
rect 10961 30366 12266 30368
rect 17217 30426 17283 30429
rect 17585 30426 17651 30429
rect 17217 30424 17651 30426
rect 17217 30368 17222 30424
rect 17278 30368 17590 30424
rect 17646 30368 17651 30424
rect 17217 30366 17651 30368
rect 10961 30363 11027 30366
rect 17217 30363 17283 30366
rect 17585 30363 17651 30366
rect 18045 30426 18111 30429
rect 20713 30426 20779 30429
rect 18045 30424 20779 30426
rect 18045 30368 18050 30424
rect 18106 30368 20718 30424
rect 20774 30368 20779 30424
rect 18045 30366 20779 30368
rect 18045 30363 18111 30366
rect 20713 30363 20779 30366
rect 21265 30426 21331 30429
rect 21950 30426 21956 30428
rect 21265 30424 21956 30426
rect 21265 30368 21270 30424
rect 21326 30368 21956 30424
rect 21265 30366 21956 30368
rect 21265 30363 21331 30366
rect 21950 30364 21956 30366
rect 22020 30364 22026 30428
rect 22134 30364 22140 30428
rect 22204 30426 22210 30428
rect 22553 30426 22619 30429
rect 22204 30424 22619 30426
rect 22204 30368 22558 30424
rect 22614 30368 22619 30424
rect 22204 30366 22619 30368
rect 23246 30426 23306 30502
rect 34928 30496 35248 30497
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 30431 35248 30432
rect 23246 30366 23536 30426
rect 22204 30364 22210 30366
rect 22553 30363 22619 30366
rect 23476 30293 23536 30366
rect 3325 30290 3391 30293
rect 7649 30290 7715 30293
rect 3325 30288 7715 30290
rect 3325 30232 3330 30288
rect 3386 30232 7654 30288
rect 7710 30232 7715 30288
rect 3325 30230 7715 30232
rect 3325 30227 3391 30230
rect 7649 30227 7715 30230
rect 12617 30290 12683 30293
rect 12750 30290 12756 30292
rect 12617 30288 12756 30290
rect 12617 30232 12622 30288
rect 12678 30232 12756 30288
rect 12617 30230 12756 30232
rect 12617 30227 12683 30230
rect 12750 30228 12756 30230
rect 12820 30228 12826 30292
rect 18229 30290 18295 30293
rect 19241 30290 19307 30293
rect 13678 30288 19307 30290
rect 13678 30232 18234 30288
rect 18290 30232 19246 30288
rect 19302 30232 19307 30288
rect 13678 30230 19307 30232
rect 10869 30154 10935 30157
rect 13678 30154 13738 30230
rect 18229 30227 18295 30230
rect 19241 30227 19307 30230
rect 23473 30288 23539 30293
rect 23473 30232 23478 30288
rect 23534 30232 23539 30288
rect 23473 30227 23539 30232
rect 24025 30290 24091 30293
rect 24945 30290 25011 30293
rect 24025 30288 25011 30290
rect 24025 30232 24030 30288
rect 24086 30232 24950 30288
rect 25006 30232 25011 30288
rect 24025 30230 25011 30232
rect 24025 30227 24091 30230
rect 24945 30227 25011 30230
rect 26233 30290 26299 30293
rect 28993 30290 29059 30293
rect 26233 30288 29059 30290
rect 26233 30232 26238 30288
rect 26294 30232 28998 30288
rect 29054 30232 29059 30288
rect 26233 30230 29059 30232
rect 26233 30227 26299 30230
rect 28993 30227 29059 30230
rect 10869 30152 13738 30154
rect 10869 30096 10874 30152
rect 10930 30096 13738 30152
rect 10869 30094 13738 30096
rect 18781 30154 18847 30157
rect 25681 30154 25747 30157
rect 18781 30152 25747 30154
rect 18781 30096 18786 30152
rect 18842 30096 25686 30152
rect 25742 30096 25747 30152
rect 18781 30094 25747 30096
rect 10869 30091 10935 30094
rect 18781 30091 18847 30094
rect 25681 30091 25747 30094
rect 25865 30154 25931 30157
rect 27838 30154 27844 30156
rect 25865 30152 27844 30154
rect 25865 30096 25870 30152
rect 25926 30096 27844 30152
rect 25865 30094 27844 30096
rect 25865 30091 25931 30094
rect 27838 30092 27844 30094
rect 27908 30154 27914 30156
rect 28073 30154 28139 30157
rect 27908 30152 28139 30154
rect 27908 30096 28078 30152
rect 28134 30096 28139 30152
rect 27908 30094 28139 30096
rect 27908 30092 27914 30094
rect 28073 30091 28139 30094
rect 7557 30018 7623 30021
rect 11881 30018 11947 30021
rect 15837 30018 15903 30021
rect 16757 30018 16823 30021
rect 7557 30016 16823 30018
rect 7557 29960 7562 30016
rect 7618 29960 11886 30016
rect 11942 29960 15842 30016
rect 15898 29960 16762 30016
rect 16818 29960 16823 30016
rect 7557 29958 16823 29960
rect 7557 29955 7623 29958
rect 11881 29955 11947 29958
rect 15837 29955 15903 29958
rect 16757 29955 16823 29958
rect 20069 30018 20135 30021
rect 22093 30018 22159 30021
rect 20069 30016 22159 30018
rect 20069 29960 20074 30016
rect 20130 29960 22098 30016
rect 22154 29960 22159 30016
rect 20069 29958 22159 29960
rect 20069 29955 20135 29958
rect 22093 29955 22159 29958
rect 22553 30018 22619 30021
rect 22870 30018 22876 30020
rect 22553 30016 22876 30018
rect 22553 29960 22558 30016
rect 22614 29960 22876 30016
rect 22553 29958 22876 29960
rect 22553 29955 22619 29958
rect 22870 29956 22876 29958
rect 22940 29956 22946 30020
rect 24669 30018 24735 30021
rect 27245 30018 27311 30021
rect 24669 30016 27311 30018
rect 24669 29960 24674 30016
rect 24730 29960 27250 30016
rect 27306 29960 27311 30016
rect 24669 29958 27311 29960
rect 24669 29955 24735 29958
rect 27245 29955 27311 29958
rect 19568 29952 19888 29953
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 29887 19888 29888
rect 10961 29882 11027 29885
rect 15469 29882 15535 29885
rect 10961 29880 15535 29882
rect 10961 29824 10966 29880
rect 11022 29824 15474 29880
rect 15530 29824 15535 29880
rect 10961 29822 15535 29824
rect 10961 29819 11027 29822
rect 15469 29819 15535 29822
rect 20805 29882 20871 29885
rect 23933 29882 23999 29885
rect 20805 29880 23999 29882
rect 20805 29824 20810 29880
rect 20866 29824 23938 29880
rect 23994 29824 23999 29880
rect 20805 29822 23999 29824
rect 20805 29819 20871 29822
rect 23933 29819 23999 29822
rect 24761 29882 24827 29885
rect 26233 29882 26299 29885
rect 24761 29880 26299 29882
rect 24761 29824 24766 29880
rect 24822 29824 26238 29880
rect 26294 29824 26299 29880
rect 24761 29822 26299 29824
rect 24761 29819 24827 29822
rect 26233 29819 26299 29822
rect 9121 29746 9187 29749
rect 12065 29746 12131 29749
rect 21173 29746 21239 29749
rect 23841 29746 23907 29749
rect 26417 29746 26483 29749
rect 9121 29744 12818 29746
rect 9121 29688 9126 29744
rect 9182 29688 12070 29744
rect 12126 29688 12818 29744
rect 9121 29686 12818 29688
rect 9121 29683 9187 29686
rect 12065 29683 12131 29686
rect 10961 29610 11027 29613
rect 12433 29610 12499 29613
rect 10961 29608 12499 29610
rect 10961 29552 10966 29608
rect 11022 29552 12438 29608
rect 12494 29552 12499 29608
rect 10961 29550 12499 29552
rect 12758 29610 12818 29686
rect 21173 29744 26483 29746
rect 21173 29688 21178 29744
rect 21234 29688 23846 29744
rect 23902 29688 26422 29744
rect 26478 29688 26483 29744
rect 21173 29686 26483 29688
rect 21173 29683 21239 29686
rect 23841 29683 23907 29686
rect 26417 29683 26483 29686
rect 14181 29610 14247 29613
rect 12758 29608 14247 29610
rect 12758 29552 14186 29608
rect 14242 29552 14247 29608
rect 12758 29550 14247 29552
rect 10961 29547 11027 29550
rect 12433 29547 12499 29550
rect 14181 29547 14247 29550
rect 14825 29610 14891 29613
rect 15101 29610 15167 29613
rect 21541 29610 21607 29613
rect 23657 29610 23723 29613
rect 28165 29610 28231 29613
rect 14825 29608 16866 29610
rect 14825 29552 14830 29608
rect 14886 29552 15106 29608
rect 15162 29552 16866 29608
rect 14825 29550 16866 29552
rect 14825 29547 14891 29550
rect 15101 29547 15167 29550
rect 9949 29474 10015 29477
rect 12617 29474 12683 29477
rect 16573 29474 16639 29477
rect 9949 29472 16639 29474
rect 9949 29416 9954 29472
rect 10010 29416 12622 29472
rect 12678 29416 16578 29472
rect 16634 29416 16639 29472
rect 9949 29414 16639 29416
rect 16806 29474 16866 29550
rect 21541 29608 28231 29610
rect 21541 29552 21546 29608
rect 21602 29552 23662 29608
rect 23718 29552 28170 29608
rect 28226 29552 28231 29608
rect 21541 29550 28231 29552
rect 21541 29547 21607 29550
rect 23657 29547 23723 29550
rect 28165 29547 28231 29550
rect 18965 29474 19031 29477
rect 26969 29474 27035 29477
rect 16806 29472 27035 29474
rect 16806 29416 18970 29472
rect 19026 29416 26974 29472
rect 27030 29416 27035 29472
rect 16806 29414 27035 29416
rect 9949 29411 10015 29414
rect 12617 29411 12683 29414
rect 16573 29411 16639 29414
rect 18965 29411 19031 29414
rect 26969 29411 27035 29414
rect 4208 29408 4528 29409
rect 0 29338 800 29368
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 29343 4528 29344
rect 34928 29408 35248 29409
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 29343 35248 29344
rect 1853 29338 1919 29341
rect 0 29336 1919 29338
rect 0 29280 1858 29336
rect 1914 29280 1919 29336
rect 0 29278 1919 29280
rect 0 29248 800 29278
rect 1853 29275 1919 29278
rect 8201 29336 8267 29341
rect 8201 29280 8206 29336
rect 8262 29280 8267 29336
rect 8201 29275 8267 29280
rect 9581 29338 9647 29341
rect 11329 29338 11395 29341
rect 9581 29336 11395 29338
rect 9581 29280 9586 29336
rect 9642 29280 11334 29336
rect 11390 29280 11395 29336
rect 9581 29278 11395 29280
rect 9581 29275 9647 29278
rect 11329 29275 11395 29278
rect 11881 29338 11947 29341
rect 15101 29338 15167 29341
rect 11881 29336 15167 29338
rect 11881 29280 11886 29336
rect 11942 29280 15106 29336
rect 15162 29280 15167 29336
rect 11881 29278 15167 29280
rect 11881 29275 11947 29278
rect 15101 29275 15167 29278
rect 19977 29338 20043 29341
rect 23105 29338 23171 29341
rect 19977 29336 23171 29338
rect 19977 29280 19982 29336
rect 20038 29280 23110 29336
rect 23166 29280 23171 29336
rect 19977 29278 23171 29280
rect 19977 29275 20043 29278
rect 23105 29275 23171 29278
rect 35566 29276 35572 29340
rect 35636 29338 35642 29340
rect 39200 29338 40000 29368
rect 35636 29278 40000 29338
rect 35636 29276 35642 29278
rect 8204 29205 8264 29275
rect 39200 29248 40000 29278
rect 8201 29200 8267 29205
rect 8385 29204 8451 29205
rect 8201 29144 8206 29200
rect 8262 29144 8267 29200
rect 8201 29139 8267 29144
rect 8334 29140 8340 29204
rect 8404 29202 8451 29204
rect 10869 29202 10935 29205
rect 13261 29202 13327 29205
rect 13813 29202 13879 29205
rect 8404 29200 8496 29202
rect 8446 29144 8496 29200
rect 8404 29142 8496 29144
rect 10869 29200 13879 29202
rect 10869 29144 10874 29200
rect 10930 29144 13266 29200
rect 13322 29144 13818 29200
rect 13874 29144 13879 29200
rect 10869 29142 13879 29144
rect 8404 29140 8451 29142
rect 8385 29139 8451 29140
rect 10869 29139 10935 29142
rect 13261 29139 13327 29142
rect 13813 29139 13879 29142
rect 14089 29202 14155 29205
rect 14222 29202 14228 29204
rect 14089 29200 14228 29202
rect 14089 29144 14094 29200
rect 14150 29144 14228 29200
rect 14089 29142 14228 29144
rect 14089 29139 14155 29142
rect 14222 29140 14228 29142
rect 14292 29140 14298 29204
rect 14590 29140 14596 29204
rect 14660 29202 14666 29204
rect 16798 29202 16804 29204
rect 14660 29142 16804 29202
rect 14660 29140 14666 29142
rect 16798 29140 16804 29142
rect 16868 29202 16874 29204
rect 19149 29202 19215 29205
rect 16868 29200 19215 29202
rect 16868 29144 19154 29200
rect 19210 29144 19215 29200
rect 16868 29142 19215 29144
rect 16868 29140 16874 29142
rect 19149 29139 19215 29142
rect 19517 29202 19583 29205
rect 22318 29202 22324 29204
rect 19517 29200 22324 29202
rect 19517 29144 19522 29200
rect 19578 29144 22324 29200
rect 19517 29142 22324 29144
rect 19517 29139 19583 29142
rect 22318 29140 22324 29142
rect 22388 29140 22394 29204
rect 10869 29066 10935 29069
rect 15561 29066 15627 29069
rect 10869 29064 15627 29066
rect 10869 29008 10874 29064
rect 10930 29008 15566 29064
rect 15622 29008 15627 29064
rect 10869 29006 15627 29008
rect 10869 29003 10935 29006
rect 15561 29003 15627 29006
rect 17125 29066 17191 29069
rect 22277 29066 22343 29069
rect 17125 29064 22343 29066
rect 17125 29008 17130 29064
rect 17186 29008 22282 29064
rect 22338 29008 22343 29064
rect 17125 29006 22343 29008
rect 17125 29003 17191 29006
rect 22277 29003 22343 29006
rect 22461 29066 22527 29069
rect 26509 29066 26575 29069
rect 22461 29064 26575 29066
rect 22461 29008 22466 29064
rect 22522 29008 26514 29064
rect 26570 29008 26575 29064
rect 22461 29006 26575 29008
rect 22461 29003 22527 29006
rect 26509 29003 26575 29006
rect 4061 28930 4127 28933
rect 7557 28930 7623 28933
rect 8109 28930 8175 28933
rect 4061 28928 7623 28930
rect 4061 28872 4066 28928
rect 4122 28872 7562 28928
rect 7618 28872 7623 28928
rect 4061 28870 7623 28872
rect 4061 28867 4127 28870
rect 7557 28867 7623 28870
rect 7974 28928 8175 28930
rect 7974 28872 8114 28928
rect 8170 28872 8175 28928
rect 7974 28870 8175 28872
rect 7974 28658 8034 28870
rect 8109 28867 8175 28870
rect 8293 28928 8359 28933
rect 8293 28872 8298 28928
rect 8354 28872 8359 28928
rect 8293 28867 8359 28872
rect 8477 28928 8543 28933
rect 8477 28872 8482 28928
rect 8538 28872 8543 28928
rect 8477 28867 8543 28872
rect 10593 28930 10659 28933
rect 13353 28930 13419 28933
rect 10593 28928 13419 28930
rect 10593 28872 10598 28928
rect 10654 28872 13358 28928
rect 13414 28872 13419 28928
rect 10593 28870 13419 28872
rect 10593 28867 10659 28870
rect 13353 28867 13419 28870
rect 13905 28930 13971 28933
rect 16665 28930 16731 28933
rect 13905 28928 16731 28930
rect 13905 28872 13910 28928
rect 13966 28872 16670 28928
rect 16726 28872 16731 28928
rect 13905 28870 16731 28872
rect 13905 28867 13971 28870
rect 16665 28867 16731 28870
rect 17033 28930 17099 28933
rect 19241 28930 19307 28933
rect 17033 28928 19307 28930
rect 17033 28872 17038 28928
rect 17094 28872 19246 28928
rect 19302 28872 19307 28928
rect 17033 28870 19307 28872
rect 17033 28867 17099 28870
rect 19241 28867 19307 28870
rect 8109 28794 8175 28797
rect 8296 28794 8356 28867
rect 8109 28792 8356 28794
rect 8109 28736 8114 28792
rect 8170 28736 8356 28792
rect 8109 28734 8356 28736
rect 8109 28731 8175 28734
rect 8201 28658 8267 28661
rect 7974 28656 8267 28658
rect 7974 28600 8206 28656
rect 8262 28600 8267 28656
rect 7974 28598 8267 28600
rect 8480 28658 8540 28867
rect 19568 28864 19888 28865
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 28799 19888 28800
rect 9673 28794 9739 28797
rect 18413 28794 18479 28797
rect 9673 28792 18479 28794
rect 9673 28736 9678 28792
rect 9734 28736 18418 28792
rect 18474 28736 18479 28792
rect 9673 28734 18479 28736
rect 9673 28731 9739 28734
rect 18413 28731 18479 28734
rect 22134 28732 22140 28796
rect 22204 28794 22210 28796
rect 23105 28794 23171 28797
rect 23749 28796 23815 28797
rect 23749 28794 23796 28796
rect 22204 28792 23171 28794
rect 22204 28736 23110 28792
rect 23166 28736 23171 28792
rect 22204 28734 23171 28736
rect 23704 28792 23796 28794
rect 23860 28794 23866 28796
rect 28993 28794 29059 28797
rect 23860 28792 29059 28794
rect 23704 28736 23754 28792
rect 23860 28736 28998 28792
rect 29054 28736 29059 28792
rect 23704 28734 23796 28736
rect 22204 28732 22210 28734
rect 23105 28731 23171 28734
rect 23749 28732 23796 28734
rect 23860 28734 29059 28736
rect 23860 28732 23866 28734
rect 23749 28731 23815 28732
rect 28993 28731 29059 28734
rect 8937 28658 9003 28661
rect 8480 28656 9003 28658
rect 8480 28600 8942 28656
rect 8998 28600 9003 28656
rect 8480 28598 9003 28600
rect 8201 28595 8267 28598
rect 8937 28595 9003 28598
rect 10501 28658 10567 28661
rect 10961 28658 11027 28661
rect 15101 28658 15167 28661
rect 10501 28656 15167 28658
rect 10501 28600 10506 28656
rect 10562 28600 10966 28656
rect 11022 28600 15106 28656
rect 15162 28600 15167 28656
rect 10501 28598 15167 28600
rect 10501 28595 10567 28598
rect 10961 28595 11027 28598
rect 15101 28595 15167 28598
rect 18873 28658 18939 28661
rect 20110 28658 20116 28660
rect 18873 28656 20116 28658
rect 18873 28600 18878 28656
rect 18934 28600 20116 28656
rect 18873 28598 20116 28600
rect 18873 28595 18939 28598
rect 20110 28596 20116 28598
rect 20180 28596 20186 28660
rect 21265 28658 21331 28661
rect 28073 28658 28139 28661
rect 29269 28658 29335 28661
rect 21265 28656 29335 28658
rect 21265 28600 21270 28656
rect 21326 28600 28078 28656
rect 28134 28600 29274 28656
rect 29330 28600 29335 28656
rect 21265 28598 29335 28600
rect 21265 28595 21331 28598
rect 28073 28595 28139 28598
rect 29269 28595 29335 28598
rect 10317 28522 10383 28525
rect 12801 28522 12867 28525
rect 10317 28520 12867 28522
rect 10317 28464 10322 28520
rect 10378 28464 12806 28520
rect 12862 28464 12867 28520
rect 10317 28462 12867 28464
rect 10317 28459 10383 28462
rect 12801 28459 12867 28462
rect 16614 28460 16620 28524
rect 16684 28522 16690 28524
rect 17585 28522 17651 28525
rect 16684 28520 17651 28522
rect 16684 28464 17590 28520
rect 17646 28464 17651 28520
rect 16684 28462 17651 28464
rect 16684 28460 16690 28462
rect 17585 28459 17651 28462
rect 17769 28522 17835 28525
rect 20713 28522 20779 28525
rect 17769 28520 20779 28522
rect 17769 28464 17774 28520
rect 17830 28464 20718 28520
rect 20774 28464 20779 28520
rect 17769 28462 20779 28464
rect 17769 28459 17835 28462
rect 20713 28459 20779 28462
rect 20989 28522 21055 28525
rect 21766 28522 21772 28524
rect 20989 28520 21772 28522
rect 20989 28464 20994 28520
rect 21050 28464 21772 28520
rect 20989 28462 21772 28464
rect 20989 28459 21055 28462
rect 21766 28460 21772 28462
rect 21836 28460 21842 28524
rect 22093 28522 22159 28525
rect 26417 28522 26483 28525
rect 22093 28520 26483 28522
rect 22093 28464 22098 28520
rect 22154 28464 26422 28520
rect 26478 28464 26483 28520
rect 22093 28462 26483 28464
rect 22093 28459 22159 28462
rect 26417 28459 26483 28462
rect 9489 28386 9555 28389
rect 15653 28386 15719 28389
rect 9489 28384 15719 28386
rect 9489 28328 9494 28384
rect 9550 28328 15658 28384
rect 15714 28328 15719 28384
rect 9489 28326 15719 28328
rect 9489 28323 9555 28326
rect 15653 28323 15719 28326
rect 18873 28386 18939 28389
rect 19885 28386 19951 28389
rect 22829 28386 22895 28389
rect 24117 28386 24183 28389
rect 26785 28386 26851 28389
rect 18873 28384 22895 28386
rect 18873 28328 18878 28384
rect 18934 28328 19890 28384
rect 19946 28328 22834 28384
rect 22890 28328 22895 28384
rect 18873 28326 22895 28328
rect 18873 28323 18939 28326
rect 19885 28323 19951 28326
rect 22829 28323 22895 28326
rect 23062 28384 26851 28386
rect 23062 28328 24122 28384
rect 24178 28328 26790 28384
rect 26846 28328 26851 28384
rect 23062 28326 26851 28328
rect 4208 28320 4528 28321
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 28255 4528 28256
rect 9121 28250 9187 28253
rect 13445 28250 13511 28253
rect 14038 28250 14044 28252
rect 9121 28248 14044 28250
rect 9121 28192 9126 28248
rect 9182 28192 13450 28248
rect 13506 28192 14044 28248
rect 9121 28190 14044 28192
rect 9121 28187 9187 28190
rect 13445 28187 13511 28190
rect 14038 28188 14044 28190
rect 14108 28250 14114 28252
rect 14181 28250 14247 28253
rect 14108 28248 14247 28250
rect 14108 28192 14186 28248
rect 14242 28192 14247 28248
rect 14108 28190 14247 28192
rect 14108 28188 14114 28190
rect 14181 28187 14247 28190
rect 20478 28188 20484 28252
rect 20548 28250 20554 28252
rect 21950 28250 21956 28252
rect 20548 28190 21956 28250
rect 20548 28188 20554 28190
rect 21950 28188 21956 28190
rect 22020 28188 22026 28252
rect 23062 28250 23122 28326
rect 24117 28323 24183 28326
rect 26785 28323 26851 28326
rect 34928 28320 35248 28321
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34928 28255 35248 28256
rect 22924 28190 23122 28250
rect 23933 28252 23999 28253
rect 23933 28248 23980 28252
rect 24044 28250 24050 28252
rect 23933 28192 23938 28248
rect 18781 28114 18847 28117
rect 21725 28114 21791 28117
rect 22924 28114 22984 28190
rect 23933 28188 23980 28192
rect 24044 28190 24090 28250
rect 24044 28188 24050 28190
rect 23933 28187 23999 28188
rect 18781 28112 22984 28114
rect 18781 28056 18786 28112
rect 18842 28056 21730 28112
rect 21786 28056 22984 28112
rect 18781 28054 22984 28056
rect 23105 28114 23171 28117
rect 28165 28114 28231 28117
rect 23105 28112 28231 28114
rect 23105 28056 23110 28112
rect 23166 28056 28170 28112
rect 28226 28056 28231 28112
rect 23105 28054 28231 28056
rect 18781 28051 18847 28054
rect 21725 28051 21791 28054
rect 23105 28051 23171 28054
rect 28165 28051 28231 28054
rect 28901 28114 28967 28117
rect 29453 28114 29519 28117
rect 32765 28114 32831 28117
rect 28901 28112 32831 28114
rect 28901 28056 28906 28112
rect 28962 28056 29458 28112
rect 29514 28056 32770 28112
rect 32826 28056 32831 28112
rect 28901 28054 32831 28056
rect 28901 28051 28967 28054
rect 29453 28051 29519 28054
rect 32765 28051 32831 28054
rect 0 27978 800 28008
rect 3693 27978 3759 27981
rect 0 27976 3759 27978
rect 0 27920 3698 27976
rect 3754 27920 3759 27976
rect 0 27918 3759 27920
rect 0 27888 800 27918
rect 3693 27915 3759 27918
rect 8937 27978 9003 27981
rect 10777 27978 10843 27981
rect 8937 27976 10843 27978
rect 8937 27920 8942 27976
rect 8998 27920 10782 27976
rect 10838 27920 10843 27976
rect 8937 27918 10843 27920
rect 8937 27915 9003 27918
rect 10777 27915 10843 27918
rect 15929 27978 15995 27981
rect 20253 27978 20319 27981
rect 20662 27978 20668 27980
rect 15929 27976 20178 27978
rect 15929 27920 15934 27976
rect 15990 27920 20178 27976
rect 15929 27918 20178 27920
rect 15929 27915 15995 27918
rect 8017 27842 8083 27845
rect 10225 27842 10291 27845
rect 8017 27840 10291 27842
rect 8017 27784 8022 27840
rect 8078 27784 10230 27840
rect 10286 27784 10291 27840
rect 8017 27782 10291 27784
rect 8017 27779 8083 27782
rect 10225 27779 10291 27782
rect 13445 27842 13511 27845
rect 14365 27842 14431 27845
rect 13445 27840 14431 27842
rect 13445 27784 13450 27840
rect 13506 27784 14370 27840
rect 14426 27784 14431 27840
rect 13445 27782 14431 27784
rect 20118 27842 20178 27918
rect 20253 27976 20668 27978
rect 20253 27920 20258 27976
rect 20314 27920 20668 27976
rect 20253 27918 20668 27920
rect 20253 27915 20319 27918
rect 20662 27916 20668 27918
rect 20732 27916 20738 27980
rect 20805 27978 20871 27981
rect 23381 27978 23447 27981
rect 20805 27976 23447 27978
rect 20805 27920 20810 27976
rect 20866 27920 23386 27976
rect 23442 27920 23447 27976
rect 20805 27918 23447 27920
rect 20805 27915 20871 27918
rect 23381 27915 23447 27918
rect 29729 27978 29795 27981
rect 39200 27978 40000 28008
rect 29729 27976 40000 27978
rect 29729 27920 29734 27976
rect 29790 27920 40000 27976
rect 29729 27918 40000 27920
rect 29729 27915 29795 27918
rect 39200 27888 40000 27918
rect 21449 27844 21515 27845
rect 21398 27842 21404 27844
rect 20118 27782 21404 27842
rect 21468 27842 21515 27844
rect 21468 27840 21560 27842
rect 21510 27784 21560 27840
rect 13445 27779 13511 27782
rect 14365 27779 14431 27782
rect 21398 27780 21404 27782
rect 21468 27782 21560 27784
rect 21468 27780 21515 27782
rect 21449 27779 21515 27780
rect 19568 27776 19888 27777
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 19568 27711 19888 27712
rect 9857 27706 9923 27709
rect 17585 27706 17651 27709
rect 19425 27706 19491 27709
rect 9857 27704 19491 27706
rect 9857 27648 9862 27704
rect 9918 27648 17590 27704
rect 17646 27648 19430 27704
rect 19486 27648 19491 27704
rect 9857 27646 19491 27648
rect 9857 27643 9923 27646
rect 17585 27643 17651 27646
rect 19425 27643 19491 27646
rect 20253 27706 20319 27709
rect 21173 27706 21239 27709
rect 29453 27706 29519 27709
rect 20253 27704 29519 27706
rect 20253 27648 20258 27704
rect 20314 27648 21178 27704
rect 21234 27648 29458 27704
rect 29514 27648 29519 27704
rect 20253 27646 29519 27648
rect 20253 27643 20319 27646
rect 21173 27643 21239 27646
rect 29453 27643 29519 27646
rect 10501 27570 10567 27573
rect 12985 27570 13051 27573
rect 10501 27568 13051 27570
rect 10501 27512 10506 27568
rect 10562 27512 12990 27568
rect 13046 27512 13051 27568
rect 10501 27510 13051 27512
rect 10501 27507 10567 27510
rect 12985 27507 13051 27510
rect 21265 27570 21331 27573
rect 22185 27570 22251 27573
rect 21265 27568 22251 27570
rect 21265 27512 21270 27568
rect 21326 27512 22190 27568
rect 22246 27512 22251 27568
rect 21265 27510 22251 27512
rect 21265 27507 21331 27510
rect 22185 27507 22251 27510
rect 22318 27508 22324 27572
rect 22388 27570 22394 27572
rect 23289 27570 23355 27573
rect 22388 27568 23355 27570
rect 22388 27512 23294 27568
rect 23350 27512 23355 27568
rect 22388 27510 23355 27512
rect 22388 27508 22394 27510
rect 23289 27507 23355 27510
rect 34053 27570 34119 27573
rect 34697 27570 34763 27573
rect 34053 27568 34763 27570
rect 34053 27512 34058 27568
rect 34114 27512 34702 27568
rect 34758 27512 34763 27568
rect 34053 27510 34763 27512
rect 34053 27507 34119 27510
rect 34697 27507 34763 27510
rect 10133 27434 10199 27437
rect 13997 27434 14063 27437
rect 10133 27432 14063 27434
rect 10133 27376 10138 27432
rect 10194 27376 14002 27432
rect 14058 27376 14063 27432
rect 10133 27374 14063 27376
rect 10133 27371 10199 27374
rect 13997 27371 14063 27374
rect 14457 27434 14523 27437
rect 18045 27434 18111 27437
rect 14457 27432 18111 27434
rect 14457 27376 14462 27432
rect 14518 27376 18050 27432
rect 18106 27376 18111 27432
rect 14457 27374 18111 27376
rect 14457 27371 14523 27374
rect 18045 27371 18111 27374
rect 18965 27434 19031 27437
rect 26049 27434 26115 27437
rect 18965 27432 26115 27434
rect 18965 27376 18970 27432
rect 19026 27376 26054 27432
rect 26110 27376 26115 27432
rect 18965 27374 26115 27376
rect 18965 27371 19031 27374
rect 26049 27371 26115 27374
rect 27797 27434 27863 27437
rect 28993 27434 29059 27437
rect 27797 27432 29059 27434
rect 27797 27376 27802 27432
rect 27858 27376 28998 27432
rect 29054 27376 29059 27432
rect 27797 27374 29059 27376
rect 27797 27371 27863 27374
rect 28993 27371 29059 27374
rect 29637 27434 29703 27437
rect 35341 27434 35407 27437
rect 29637 27432 35407 27434
rect 29637 27376 29642 27432
rect 29698 27376 35346 27432
rect 35402 27376 35407 27432
rect 29637 27374 35407 27376
rect 29637 27371 29703 27374
rect 35341 27371 35407 27374
rect 14089 27300 14155 27301
rect 14038 27298 14044 27300
rect 13998 27238 14044 27298
rect 14108 27296 14155 27300
rect 14150 27240 14155 27296
rect 14038 27236 14044 27238
rect 14108 27236 14155 27240
rect 14089 27235 14155 27236
rect 17585 27298 17651 27301
rect 18689 27298 18755 27301
rect 21725 27298 21791 27301
rect 17585 27296 21791 27298
rect 17585 27240 17590 27296
rect 17646 27240 18694 27296
rect 18750 27240 21730 27296
rect 21786 27240 21791 27296
rect 17585 27238 21791 27240
rect 17585 27235 17651 27238
rect 18689 27235 18755 27238
rect 21725 27235 21791 27238
rect 22134 27236 22140 27300
rect 22204 27298 22210 27300
rect 27797 27298 27863 27301
rect 22204 27296 27863 27298
rect 22204 27240 27802 27296
rect 27858 27240 27863 27296
rect 22204 27238 27863 27240
rect 22204 27236 22210 27238
rect 27797 27235 27863 27238
rect 4208 27232 4528 27233
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 27167 4528 27168
rect 34928 27232 35248 27233
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34928 27167 35248 27168
rect 17166 27100 17172 27164
rect 17236 27162 17242 27164
rect 19425 27162 19491 27165
rect 17236 27160 19491 27162
rect 17236 27104 19430 27160
rect 19486 27104 19491 27160
rect 17236 27102 19491 27104
rect 17236 27100 17242 27102
rect 19425 27099 19491 27102
rect 22277 27162 22343 27165
rect 23289 27164 23355 27165
rect 22277 27160 22938 27162
rect 22277 27104 22282 27160
rect 22338 27104 22938 27160
rect 22277 27102 22938 27104
rect 22277 27099 22343 27102
rect 9121 27026 9187 27029
rect 13537 27026 13603 27029
rect 16573 27026 16639 27029
rect 9121 27024 13603 27026
rect 9121 26968 9126 27024
rect 9182 26968 13542 27024
rect 13598 26968 13603 27024
rect 9121 26966 13603 26968
rect 9121 26963 9187 26966
rect 13537 26963 13603 26966
rect 14046 27024 16639 27026
rect 14046 26968 16578 27024
rect 16634 26968 16639 27024
rect 14046 26966 16639 26968
rect 10869 26890 10935 26893
rect 14046 26890 14106 26966
rect 16573 26963 16639 26966
rect 16941 27026 17007 27029
rect 22737 27026 22803 27029
rect 16941 27024 22803 27026
rect 16941 26968 16946 27024
rect 17002 26968 22742 27024
rect 22798 26968 22803 27024
rect 16941 26966 22803 26968
rect 22878 27026 22938 27102
rect 23238 27100 23244 27164
rect 23308 27162 23355 27164
rect 28349 27162 28415 27165
rect 23308 27160 28415 27162
rect 23350 27104 28354 27160
rect 28410 27104 28415 27160
rect 23308 27102 28415 27104
rect 23308 27100 23355 27102
rect 23289 27099 23355 27100
rect 28349 27099 28415 27102
rect 25037 27026 25103 27029
rect 25405 27026 25471 27029
rect 22878 27024 25471 27026
rect 22878 26968 25042 27024
rect 25098 26968 25410 27024
rect 25466 26968 25471 27024
rect 22878 26966 25471 26968
rect 16941 26963 17007 26966
rect 22737 26963 22803 26966
rect 25037 26963 25103 26966
rect 25405 26963 25471 26966
rect 10869 26888 14106 26890
rect 10869 26832 10874 26888
rect 10930 26832 14106 26888
rect 10869 26830 14106 26832
rect 10869 26827 10935 26830
rect 14222 26828 14228 26892
rect 14292 26890 14298 26892
rect 14958 26890 14964 26892
rect 14292 26830 14964 26890
rect 14292 26828 14298 26830
rect 14958 26828 14964 26830
rect 15028 26828 15034 26892
rect 19425 26890 19491 26893
rect 20621 26890 20687 26893
rect 25773 26890 25839 26893
rect 28073 26890 28139 26893
rect 19425 26888 20178 26890
rect 19425 26832 19430 26888
rect 19486 26832 20178 26888
rect 19425 26830 20178 26832
rect 19425 26827 19491 26830
rect 7097 26754 7163 26757
rect 7230 26754 7236 26756
rect 7097 26752 7236 26754
rect 7097 26696 7102 26752
rect 7158 26696 7236 26752
rect 7097 26694 7236 26696
rect 7097 26691 7163 26694
rect 7230 26692 7236 26694
rect 7300 26692 7306 26756
rect 19568 26688 19888 26689
rect 0 26618 800 26648
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 26623 19888 26624
rect 1577 26618 1643 26621
rect 0 26616 1643 26618
rect 0 26560 1582 26616
rect 1638 26560 1643 26616
rect 0 26558 1643 26560
rect 0 26528 800 26558
rect 1577 26555 1643 26558
rect 11329 26618 11395 26621
rect 14641 26618 14707 26621
rect 11329 26616 14707 26618
rect 11329 26560 11334 26616
rect 11390 26560 14646 26616
rect 14702 26560 14707 26616
rect 11329 26558 14707 26560
rect 20118 26618 20178 26830
rect 20621 26888 28139 26890
rect 20621 26832 20626 26888
rect 20682 26832 25778 26888
rect 25834 26832 28078 26888
rect 28134 26832 28139 26888
rect 20621 26830 28139 26832
rect 20621 26827 20687 26830
rect 25773 26827 25839 26830
rect 28073 26827 28139 26830
rect 28809 26890 28875 26893
rect 30465 26890 30531 26893
rect 28809 26888 30531 26890
rect 28809 26832 28814 26888
rect 28870 26832 30470 26888
rect 30526 26832 30531 26888
rect 28809 26830 30531 26832
rect 28809 26827 28875 26830
rect 30465 26827 30531 26830
rect 21449 26754 21515 26757
rect 24761 26754 24827 26757
rect 21449 26752 24827 26754
rect 21449 26696 21454 26752
rect 21510 26696 24766 26752
rect 24822 26696 24827 26752
rect 21449 26694 24827 26696
rect 21449 26691 21515 26694
rect 24761 26691 24827 26694
rect 24485 26618 24551 26621
rect 20118 26616 24551 26618
rect 20118 26560 24490 26616
rect 24546 26560 24551 26616
rect 20118 26558 24551 26560
rect 11329 26555 11395 26558
rect 14641 26555 14707 26558
rect 24485 26555 24551 26558
rect 24669 26618 24735 26621
rect 25773 26618 25839 26621
rect 28441 26618 28507 26621
rect 24669 26616 28507 26618
rect 24669 26560 24674 26616
rect 24730 26560 25778 26616
rect 25834 26560 28446 26616
rect 28502 26560 28507 26616
rect 24669 26558 28507 26560
rect 24669 26555 24735 26558
rect 25773 26555 25839 26558
rect 28441 26555 28507 26558
rect 34462 26556 34468 26620
rect 34532 26618 34538 26620
rect 39200 26618 40000 26648
rect 34532 26558 40000 26618
rect 34532 26556 34538 26558
rect 39200 26528 40000 26558
rect 8477 26482 8543 26485
rect 11237 26482 11303 26485
rect 11513 26482 11579 26485
rect 8477 26480 11579 26482
rect 8477 26424 8482 26480
rect 8538 26424 11242 26480
rect 11298 26424 11518 26480
rect 11574 26424 11579 26480
rect 8477 26422 11579 26424
rect 8477 26419 8543 26422
rect 11237 26419 11303 26422
rect 11513 26419 11579 26422
rect 13077 26482 13143 26485
rect 13302 26482 13308 26484
rect 13077 26480 13308 26482
rect 13077 26424 13082 26480
rect 13138 26424 13308 26480
rect 13077 26422 13308 26424
rect 13077 26419 13143 26422
rect 13302 26420 13308 26422
rect 13372 26420 13378 26484
rect 18965 26482 19031 26485
rect 20897 26482 20963 26485
rect 18965 26480 20963 26482
rect 18965 26424 18970 26480
rect 19026 26424 20902 26480
rect 20958 26424 20963 26480
rect 18965 26422 20963 26424
rect 18965 26419 19031 26422
rect 20897 26419 20963 26422
rect 21449 26482 21515 26485
rect 25497 26482 25563 26485
rect 28533 26482 28599 26485
rect 21449 26480 25563 26482
rect 21449 26424 21454 26480
rect 21510 26424 25502 26480
rect 25558 26424 25563 26480
rect 21449 26422 25563 26424
rect 21449 26419 21515 26422
rect 25497 26419 25563 26422
rect 27294 26480 28599 26482
rect 27294 26424 28538 26480
rect 28594 26424 28599 26480
rect 27294 26422 28599 26424
rect 4061 26346 4127 26349
rect 6678 26346 6684 26348
rect 4061 26344 6684 26346
rect 4061 26288 4066 26344
rect 4122 26288 6684 26344
rect 4061 26286 6684 26288
rect 4061 26283 4127 26286
rect 6678 26284 6684 26286
rect 6748 26284 6754 26348
rect 9857 26346 9923 26349
rect 12893 26346 12959 26349
rect 13169 26348 13235 26349
rect 9857 26344 12959 26346
rect 9857 26288 9862 26344
rect 9918 26288 12898 26344
rect 12954 26288 12959 26344
rect 9857 26286 12959 26288
rect 9857 26283 9923 26286
rect 12893 26283 12959 26286
rect 13118 26284 13124 26348
rect 13188 26346 13235 26348
rect 22553 26346 22619 26349
rect 22829 26346 22895 26349
rect 13188 26344 13280 26346
rect 13230 26288 13280 26344
rect 13188 26286 13280 26288
rect 22553 26344 22895 26346
rect 22553 26288 22558 26344
rect 22614 26288 22834 26344
rect 22890 26288 22895 26344
rect 22553 26286 22895 26288
rect 13188 26284 13235 26286
rect 13169 26283 13235 26284
rect 22553 26283 22619 26286
rect 22829 26283 22895 26286
rect 23381 26346 23447 26349
rect 23933 26346 23999 26349
rect 23381 26344 23999 26346
rect 23381 26288 23386 26344
rect 23442 26288 23938 26344
rect 23994 26288 23999 26344
rect 23381 26286 23999 26288
rect 23381 26283 23447 26286
rect 23933 26283 23999 26286
rect 24209 26346 24275 26349
rect 26785 26346 26851 26349
rect 27294 26346 27354 26422
rect 28533 26419 28599 26422
rect 24209 26344 27354 26346
rect 24209 26288 24214 26344
rect 24270 26288 26790 26344
rect 26846 26288 27354 26344
rect 24209 26286 27354 26288
rect 27613 26346 27679 26349
rect 33501 26346 33567 26349
rect 27613 26344 33567 26346
rect 27613 26288 27618 26344
rect 27674 26288 33506 26344
rect 33562 26288 33567 26344
rect 27613 26286 33567 26288
rect 24209 26283 24275 26286
rect 26785 26283 26851 26286
rect 27613 26283 27679 26286
rect 33501 26283 33567 26286
rect 35801 26346 35867 26349
rect 36353 26346 36419 26349
rect 35801 26344 36419 26346
rect 35801 26288 35806 26344
rect 35862 26288 36358 26344
rect 36414 26288 36419 26344
rect 35801 26286 36419 26288
rect 35801 26283 35867 26286
rect 36353 26283 36419 26286
rect 13997 26210 14063 26213
rect 16757 26210 16823 26213
rect 13997 26208 16823 26210
rect 13997 26152 14002 26208
rect 14058 26152 16762 26208
rect 16818 26152 16823 26208
rect 13997 26150 16823 26152
rect 13997 26147 14063 26150
rect 16757 26147 16823 26150
rect 19609 26210 19675 26213
rect 25037 26210 25103 26213
rect 19609 26208 25103 26210
rect 19609 26152 19614 26208
rect 19670 26152 25042 26208
rect 25098 26152 25103 26208
rect 19609 26150 25103 26152
rect 19609 26147 19675 26150
rect 25037 26147 25103 26150
rect 4208 26144 4528 26145
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 26079 4528 26080
rect 34928 26144 35248 26145
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34928 26079 35248 26080
rect 16297 26074 16363 26077
rect 20897 26074 20963 26077
rect 16297 26072 20963 26074
rect 16297 26016 16302 26072
rect 16358 26016 20902 26072
rect 20958 26016 20963 26072
rect 16297 26014 20963 26016
rect 16297 26011 16363 26014
rect 20897 26011 20963 26014
rect 21081 26074 21147 26077
rect 25313 26074 25379 26077
rect 21081 26072 25379 26074
rect 21081 26016 21086 26072
rect 21142 26016 25318 26072
rect 25374 26016 25379 26072
rect 21081 26014 25379 26016
rect 21081 26011 21147 26014
rect 25313 26011 25379 26014
rect 11513 25938 11579 25941
rect 17309 25938 17375 25941
rect 11513 25936 17375 25938
rect 11513 25880 11518 25936
rect 11574 25880 17314 25936
rect 17370 25880 17375 25936
rect 11513 25878 17375 25880
rect 11513 25875 11579 25878
rect 17309 25875 17375 25878
rect 19149 25938 19215 25941
rect 24853 25938 24919 25941
rect 19149 25936 24919 25938
rect 19149 25880 19154 25936
rect 19210 25880 24858 25936
rect 24914 25880 24919 25936
rect 19149 25878 24919 25880
rect 19149 25875 19215 25878
rect 24853 25875 24919 25878
rect 12157 25802 12223 25805
rect 16205 25802 16271 25805
rect 12157 25800 16271 25802
rect 12157 25744 12162 25800
rect 12218 25744 16210 25800
rect 16266 25744 16271 25800
rect 12157 25742 16271 25744
rect 12157 25739 12223 25742
rect 16205 25739 16271 25742
rect 18689 25802 18755 25805
rect 20989 25802 21055 25805
rect 18689 25800 21055 25802
rect 18689 25744 18694 25800
rect 18750 25744 20994 25800
rect 21050 25744 21055 25800
rect 18689 25742 21055 25744
rect 18689 25739 18755 25742
rect 20989 25739 21055 25742
rect 22829 25802 22895 25805
rect 25865 25802 25931 25805
rect 22829 25800 25931 25802
rect 22829 25744 22834 25800
rect 22890 25744 25870 25800
rect 25926 25744 25931 25800
rect 22829 25742 25931 25744
rect 22829 25739 22895 25742
rect 25865 25739 25931 25742
rect 12617 25666 12683 25669
rect 18781 25666 18847 25669
rect 12617 25664 18847 25666
rect 12617 25608 12622 25664
rect 12678 25608 18786 25664
rect 18842 25608 18847 25664
rect 12617 25606 18847 25608
rect 12617 25603 12683 25606
rect 18781 25603 18847 25606
rect 20805 25666 20871 25669
rect 23289 25666 23355 25669
rect 20805 25664 23355 25666
rect 20805 25608 20810 25664
rect 20866 25608 23294 25664
rect 23350 25608 23355 25664
rect 20805 25606 23355 25608
rect 20805 25603 20871 25606
rect 23289 25603 23355 25606
rect 19568 25600 19888 25601
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 25535 19888 25536
rect 9305 25530 9371 25533
rect 11329 25530 11395 25533
rect 15653 25530 15719 25533
rect 9305 25528 15719 25530
rect 9305 25472 9310 25528
rect 9366 25472 11334 25528
rect 11390 25472 15658 25528
rect 15714 25472 15719 25528
rect 9305 25470 15719 25472
rect 9305 25467 9371 25470
rect 11329 25467 11395 25470
rect 15653 25467 15719 25470
rect 21265 25530 21331 25533
rect 25313 25530 25379 25533
rect 21265 25528 25379 25530
rect 21265 25472 21270 25528
rect 21326 25472 25318 25528
rect 25374 25472 25379 25528
rect 21265 25470 25379 25472
rect 21265 25467 21331 25470
rect 25313 25467 25379 25470
rect 11973 25394 12039 25397
rect 22185 25394 22251 25397
rect 22921 25396 22987 25397
rect 11973 25392 22251 25394
rect 11973 25336 11978 25392
rect 12034 25336 22190 25392
rect 22246 25336 22251 25392
rect 11973 25334 22251 25336
rect 11973 25331 12039 25334
rect 22185 25331 22251 25334
rect 22870 25332 22876 25396
rect 22940 25394 22987 25396
rect 22940 25392 23032 25394
rect 22982 25336 23032 25392
rect 22940 25334 23032 25336
rect 22940 25332 22987 25334
rect 22921 25331 22987 25332
rect 0 25258 800 25288
rect 3509 25258 3575 25261
rect 0 25256 3575 25258
rect 0 25200 3514 25256
rect 3570 25200 3575 25256
rect 0 25198 3575 25200
rect 0 25168 800 25198
rect 3509 25195 3575 25198
rect 4061 25258 4127 25261
rect 9673 25258 9739 25261
rect 4061 25256 9739 25258
rect 4061 25200 4066 25256
rect 4122 25200 9678 25256
rect 9734 25200 9739 25256
rect 4061 25198 9739 25200
rect 4061 25195 4127 25198
rect 9673 25195 9739 25198
rect 14457 25258 14523 25261
rect 17217 25258 17283 25261
rect 14457 25256 17283 25258
rect 14457 25200 14462 25256
rect 14518 25200 17222 25256
rect 17278 25200 17283 25256
rect 14457 25198 17283 25200
rect 14457 25195 14523 25198
rect 17217 25195 17283 25198
rect 17585 25258 17651 25261
rect 19793 25258 19859 25261
rect 23841 25258 23907 25261
rect 17585 25256 23907 25258
rect 17585 25200 17590 25256
rect 17646 25200 19798 25256
rect 19854 25200 23846 25256
rect 23902 25200 23907 25256
rect 17585 25198 23907 25200
rect 17585 25195 17651 25198
rect 19793 25195 19859 25198
rect 23841 25195 23907 25198
rect 34462 25196 34468 25260
rect 34532 25258 34538 25260
rect 39200 25258 40000 25288
rect 34532 25198 40000 25258
rect 34532 25196 34538 25198
rect 39200 25168 40000 25198
rect 14641 25124 14707 25125
rect 14590 25122 14596 25124
rect 14550 25062 14596 25122
rect 14660 25120 14707 25124
rect 14702 25064 14707 25120
rect 14590 25060 14596 25062
rect 14660 25060 14707 25064
rect 14641 25059 14707 25060
rect 16481 25122 16547 25125
rect 22185 25122 22251 25125
rect 23238 25122 23244 25124
rect 16481 25120 21834 25122
rect 16481 25064 16486 25120
rect 16542 25064 21834 25120
rect 16481 25062 21834 25064
rect 16481 25059 16547 25062
rect 4208 25056 4528 25057
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 24991 4528 24992
rect 14549 24986 14615 24989
rect 18689 24986 18755 24989
rect 20437 24986 20503 24989
rect 14549 24984 20503 24986
rect 14549 24928 14554 24984
rect 14610 24928 18694 24984
rect 18750 24928 20442 24984
rect 20498 24928 20503 24984
rect 14549 24926 20503 24928
rect 14549 24923 14615 24926
rect 18689 24923 18755 24926
rect 20437 24923 20503 24926
rect 12801 24850 12867 24853
rect 13670 24850 13676 24852
rect 12801 24848 13676 24850
rect 12801 24792 12806 24848
rect 12862 24792 13676 24848
rect 12801 24790 13676 24792
rect 12801 24787 12867 24790
rect 13670 24788 13676 24790
rect 13740 24788 13746 24852
rect 15101 24850 15167 24853
rect 16757 24850 16823 24853
rect 17033 24850 17099 24853
rect 20805 24850 20871 24853
rect 15101 24848 16823 24850
rect 15101 24792 15106 24848
rect 15162 24792 16762 24848
rect 16818 24792 16823 24848
rect 15101 24790 16823 24792
rect 15101 24787 15167 24790
rect 16757 24787 16823 24790
rect 16990 24848 20871 24850
rect 16990 24792 17038 24848
rect 17094 24792 20810 24848
rect 20866 24792 20871 24848
rect 16990 24790 20871 24792
rect 16990 24787 17099 24790
rect 20805 24787 20871 24790
rect 14733 24714 14799 24717
rect 16990 24714 17050 24787
rect 14733 24712 17050 24714
rect 14733 24656 14738 24712
rect 14794 24656 17050 24712
rect 14733 24654 17050 24656
rect 17677 24714 17743 24717
rect 20437 24714 20503 24717
rect 21081 24714 21147 24717
rect 17677 24712 21147 24714
rect 17677 24656 17682 24712
rect 17738 24656 20442 24712
rect 20498 24656 21086 24712
rect 21142 24656 21147 24712
rect 17677 24654 21147 24656
rect 21774 24714 21834 25062
rect 22185 25120 23244 25122
rect 22185 25064 22190 25120
rect 22246 25064 23244 25120
rect 22185 25062 23244 25064
rect 22185 25059 22251 25062
rect 23238 25060 23244 25062
rect 23308 25060 23314 25124
rect 34928 25056 35248 25057
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 24991 35248 24992
rect 24669 24850 24735 24853
rect 26233 24850 26299 24853
rect 24669 24848 26299 24850
rect 24669 24792 24674 24848
rect 24730 24792 26238 24848
rect 26294 24792 26299 24848
rect 24669 24790 26299 24792
rect 24669 24787 24735 24790
rect 26233 24787 26299 24790
rect 25221 24714 25287 24717
rect 21774 24712 25287 24714
rect 21774 24656 25226 24712
rect 25282 24656 25287 24712
rect 21774 24654 25287 24656
rect 14733 24651 14799 24654
rect 17677 24651 17743 24654
rect 20437 24651 20503 24654
rect 21081 24651 21147 24654
rect 25221 24651 25287 24654
rect 13629 24578 13695 24581
rect 16665 24578 16731 24581
rect 13629 24576 16731 24578
rect 13629 24520 13634 24576
rect 13690 24520 16670 24576
rect 16726 24520 16731 24576
rect 13629 24518 16731 24520
rect 13629 24515 13695 24518
rect 16665 24515 16731 24518
rect 21582 24516 21588 24580
rect 21652 24578 21658 24580
rect 23749 24578 23815 24581
rect 21652 24576 23815 24578
rect 21652 24520 23754 24576
rect 23810 24520 23815 24576
rect 21652 24518 23815 24520
rect 21652 24516 21658 24518
rect 23749 24515 23815 24518
rect 19568 24512 19888 24513
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 19568 24447 19888 24448
rect 13905 24442 13971 24445
rect 14089 24442 14155 24445
rect 15837 24442 15903 24445
rect 13905 24440 15903 24442
rect 13905 24384 13910 24440
rect 13966 24384 14094 24440
rect 14150 24384 15842 24440
rect 15898 24384 15903 24440
rect 13905 24382 15903 24384
rect 13905 24379 13971 24382
rect 14089 24379 14155 24382
rect 15837 24379 15903 24382
rect 22001 24442 22067 24445
rect 23841 24442 23907 24445
rect 22001 24440 23907 24442
rect 22001 24384 22006 24440
rect 22062 24384 23846 24440
rect 23902 24384 23907 24440
rect 22001 24382 23907 24384
rect 22001 24379 22067 24382
rect 23841 24379 23907 24382
rect 17585 24306 17651 24309
rect 19425 24306 19491 24309
rect 23749 24306 23815 24309
rect 17585 24304 19491 24306
rect 17585 24248 17590 24304
rect 17646 24248 19430 24304
rect 19486 24248 19491 24304
rect 17585 24246 19491 24248
rect 17585 24243 17651 24246
rect 19425 24243 19491 24246
rect 19566 24304 23815 24306
rect 19566 24248 23754 24304
rect 23810 24248 23815 24304
rect 19566 24246 23815 24248
rect 13077 24170 13143 24173
rect 17769 24170 17835 24173
rect 13077 24168 17835 24170
rect 13077 24112 13082 24168
rect 13138 24112 17774 24168
rect 17830 24112 17835 24168
rect 13077 24110 17835 24112
rect 13077 24107 13143 24110
rect 17769 24107 17835 24110
rect 18229 24170 18295 24173
rect 19566 24170 19626 24246
rect 23749 24243 23815 24246
rect 21449 24172 21515 24173
rect 21398 24170 21404 24172
rect 18229 24168 19626 24170
rect 18229 24112 18234 24168
rect 18290 24112 19626 24168
rect 18229 24110 19626 24112
rect 21358 24110 21404 24170
rect 21468 24168 21515 24172
rect 21510 24112 21515 24168
rect 18229 24107 18295 24110
rect 21398 24108 21404 24110
rect 21468 24108 21515 24112
rect 21449 24107 21515 24108
rect 26141 24170 26207 24173
rect 26141 24168 35404 24170
rect 26141 24112 26146 24168
rect 26202 24112 35404 24168
rect 26141 24110 35404 24112
rect 26141 24107 26207 24110
rect 8109 24034 8175 24037
rect 15101 24034 15167 24037
rect 17309 24034 17375 24037
rect 8109 24032 15026 24034
rect 8109 23976 8114 24032
rect 8170 23976 15026 24032
rect 8109 23974 15026 23976
rect 8109 23971 8175 23974
rect 4208 23968 4528 23969
rect 0 23898 800 23928
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 23903 4528 23904
rect 4061 23898 4127 23901
rect 0 23896 4127 23898
rect 0 23840 4066 23896
rect 4122 23840 4127 23896
rect 0 23838 4127 23840
rect 0 23808 800 23838
rect 4061 23835 4127 23838
rect 7833 23762 7899 23765
rect 8937 23762 9003 23765
rect 12341 23762 12407 23765
rect 14549 23762 14615 23765
rect 7833 23760 14615 23762
rect 7833 23704 7838 23760
rect 7894 23704 8942 23760
rect 8998 23704 12346 23760
rect 12402 23704 14554 23760
rect 14610 23704 14615 23760
rect 7833 23702 14615 23704
rect 14966 23762 15026 23974
rect 15101 24032 17375 24034
rect 15101 23976 15106 24032
rect 15162 23976 17314 24032
rect 17370 23976 17375 24032
rect 15101 23974 17375 23976
rect 15101 23971 15167 23974
rect 17309 23971 17375 23974
rect 17769 24034 17835 24037
rect 20069 24034 20135 24037
rect 17769 24032 20135 24034
rect 17769 23976 17774 24032
rect 17830 23976 20074 24032
rect 20130 23976 20135 24032
rect 17769 23974 20135 23976
rect 17769 23971 17835 23974
rect 20069 23971 20135 23974
rect 21541 24034 21607 24037
rect 25405 24034 25471 24037
rect 21541 24032 25471 24034
rect 21541 23976 21546 24032
rect 21602 23976 25410 24032
rect 25466 23976 25471 24032
rect 21541 23974 25471 23976
rect 21541 23971 21607 23974
rect 25405 23971 25471 23974
rect 34928 23968 35248 23969
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 23903 35248 23904
rect 15101 23898 15167 23901
rect 18321 23898 18387 23901
rect 15101 23896 18387 23898
rect 15101 23840 15106 23896
rect 15162 23840 18326 23896
rect 18382 23840 18387 23896
rect 15101 23838 18387 23840
rect 15101 23835 15167 23838
rect 18321 23835 18387 23838
rect 19241 23898 19307 23901
rect 23657 23898 23723 23901
rect 19241 23896 23723 23898
rect 19241 23840 19246 23896
rect 19302 23840 23662 23896
rect 23718 23840 23723 23896
rect 19241 23838 23723 23840
rect 35344 23898 35404 24110
rect 39200 23898 40000 23928
rect 35344 23838 40000 23898
rect 19241 23835 19307 23838
rect 23657 23835 23723 23838
rect 39200 23808 40000 23838
rect 16614 23762 16620 23764
rect 14966 23702 16620 23762
rect 7833 23699 7899 23702
rect 8937 23699 9003 23702
rect 12341 23699 12407 23702
rect 14549 23699 14615 23702
rect 16614 23700 16620 23702
rect 16684 23700 16690 23764
rect 23657 23762 23723 23765
rect 26417 23762 26483 23765
rect 23657 23760 26483 23762
rect 23657 23704 23662 23760
rect 23718 23704 26422 23760
rect 26478 23704 26483 23760
rect 23657 23702 26483 23704
rect 23657 23699 23723 23702
rect 26417 23699 26483 23702
rect 14038 23564 14044 23628
rect 14108 23626 14114 23628
rect 21541 23626 21607 23629
rect 21950 23626 21956 23628
rect 14108 23624 21956 23626
rect 14108 23568 21546 23624
rect 21602 23568 21956 23624
rect 14108 23566 21956 23568
rect 14108 23564 14114 23566
rect 21541 23563 21607 23566
rect 21950 23564 21956 23566
rect 22020 23564 22026 23628
rect 22829 23626 22895 23629
rect 33777 23626 33843 23629
rect 22829 23624 33843 23626
rect 22829 23568 22834 23624
rect 22890 23568 33782 23624
rect 33838 23568 33843 23624
rect 22829 23566 33843 23568
rect 22829 23563 22895 23566
rect 33777 23563 33843 23566
rect 19568 23424 19888 23425
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 23359 19888 23360
rect 2681 23354 2747 23357
rect 798 23352 2747 23354
rect 798 23296 2686 23352
rect 2742 23296 2747 23352
rect 798 23294 2747 23296
rect 798 23248 858 23294
rect 2681 23291 2747 23294
rect 3141 23354 3207 23357
rect 9673 23354 9739 23357
rect 11789 23354 11855 23357
rect 3141 23352 11855 23354
rect 3141 23296 3146 23352
rect 3202 23296 9678 23352
rect 9734 23296 11794 23352
rect 11850 23296 11855 23352
rect 3141 23294 11855 23296
rect 3141 23291 3207 23294
rect 9673 23291 9739 23294
rect 11789 23291 11855 23294
rect 13997 23354 14063 23357
rect 15285 23354 15351 23357
rect 13997 23352 15351 23354
rect 13997 23296 14002 23352
rect 14058 23296 15290 23352
rect 15346 23296 15351 23352
rect 13997 23294 15351 23296
rect 13997 23291 14063 23294
rect 15285 23291 15351 23294
rect 26417 23354 26483 23357
rect 29085 23354 29151 23357
rect 26417 23352 29151 23354
rect 26417 23296 26422 23352
rect 26478 23296 29090 23352
rect 29146 23296 29151 23352
rect 26417 23294 29151 23296
rect 26417 23291 26483 23294
rect 29085 23291 29151 23294
rect 0 23158 858 23248
rect 17033 23218 17099 23221
rect 21173 23218 21239 23221
rect 17033 23216 21239 23218
rect 17033 23160 17038 23216
rect 17094 23160 21178 23216
rect 21234 23160 21239 23216
rect 17033 23158 21239 23160
rect 0 23128 800 23158
rect 17033 23155 17099 23158
rect 21173 23155 21239 23158
rect 23238 23156 23244 23220
rect 23308 23218 23314 23220
rect 24669 23218 24735 23221
rect 23308 23216 24735 23218
rect 23308 23160 24674 23216
rect 24730 23160 24735 23216
rect 23308 23158 24735 23160
rect 23308 23156 23314 23158
rect 24669 23155 24735 23158
rect 19149 23082 19215 23085
rect 20069 23082 20135 23085
rect 19149 23080 20135 23082
rect 19149 23024 19154 23080
rect 19210 23024 20074 23080
rect 20130 23024 20135 23080
rect 19149 23022 20135 23024
rect 19149 23019 19215 23022
rect 20069 23019 20135 23022
rect 21633 23082 21699 23085
rect 22001 23082 22067 23085
rect 22829 23082 22895 23085
rect 21633 23080 22895 23082
rect 21633 23024 21638 23080
rect 21694 23024 22006 23080
rect 22062 23024 22834 23080
rect 22890 23024 22895 23080
rect 21633 23022 22895 23024
rect 21633 23019 21699 23022
rect 22001 23019 22067 23022
rect 22829 23019 22895 23022
rect 23289 23082 23355 23085
rect 24485 23082 24551 23085
rect 27429 23082 27495 23085
rect 23289 23080 27495 23082
rect 23289 23024 23294 23080
rect 23350 23024 24490 23080
rect 24546 23024 27434 23080
rect 27490 23024 27495 23080
rect 23289 23022 27495 23024
rect 23289 23019 23355 23022
rect 24485 23019 24551 23022
rect 27429 23019 27495 23022
rect 12525 22946 12591 22949
rect 21541 22946 21607 22949
rect 12525 22944 21607 22946
rect 12525 22888 12530 22944
rect 12586 22888 21546 22944
rect 21602 22888 21607 22944
rect 12525 22886 21607 22888
rect 12525 22883 12591 22886
rect 21541 22883 21607 22886
rect 4208 22880 4528 22881
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 22815 4528 22816
rect 34928 22880 35248 22881
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 22815 35248 22816
rect 12157 22810 12223 22813
rect 14641 22810 14707 22813
rect 12157 22808 14707 22810
rect 12157 22752 12162 22808
rect 12218 22752 14646 22808
rect 14702 22752 14707 22808
rect 12157 22750 14707 22752
rect 12157 22747 12223 22750
rect 14641 22747 14707 22750
rect 14825 22810 14891 22813
rect 24025 22810 24091 22813
rect 14825 22808 24091 22810
rect 14825 22752 14830 22808
rect 14886 22752 24030 22808
rect 24086 22752 24091 22808
rect 14825 22750 24091 22752
rect 14825 22747 14891 22750
rect 24025 22747 24091 22750
rect 13169 22674 13235 22677
rect 15929 22674 15995 22677
rect 17493 22674 17559 22677
rect 13169 22672 17559 22674
rect 13169 22616 13174 22672
rect 13230 22616 15934 22672
rect 15990 22616 17498 22672
rect 17554 22616 17559 22672
rect 13169 22614 17559 22616
rect 13169 22611 13235 22614
rect 15929 22611 15995 22614
rect 17493 22611 17559 22614
rect 21449 22674 21515 22677
rect 22001 22674 22067 22677
rect 21449 22672 22067 22674
rect 21449 22616 21454 22672
rect 21510 22616 22006 22672
rect 22062 22616 22067 22672
rect 21449 22614 22067 22616
rect 21449 22611 21515 22614
rect 22001 22611 22067 22614
rect 23841 22674 23907 22677
rect 26601 22674 26667 22677
rect 29177 22674 29243 22677
rect 23841 22672 26667 22674
rect 23841 22616 23846 22672
rect 23902 22616 26606 22672
rect 26662 22616 26667 22672
rect 23841 22614 26667 22616
rect 23841 22611 23907 22614
rect 26601 22611 26667 22614
rect 26742 22672 29243 22674
rect 26742 22616 29182 22672
rect 29238 22616 29243 22672
rect 26742 22614 29243 22616
rect 18321 22538 18387 22541
rect 21173 22538 21239 22541
rect 18321 22536 21239 22538
rect 18321 22480 18326 22536
rect 18382 22480 21178 22536
rect 21234 22480 21239 22536
rect 18321 22478 21239 22480
rect 18321 22475 18387 22478
rect 21173 22475 21239 22478
rect 23105 22538 23171 22541
rect 26742 22538 26802 22614
rect 29177 22611 29243 22614
rect 23105 22536 26802 22538
rect 23105 22480 23110 22536
rect 23166 22480 26802 22536
rect 23105 22478 26802 22480
rect 28993 22538 29059 22541
rect 39200 22538 40000 22568
rect 28993 22536 40000 22538
rect 28993 22480 28998 22536
rect 29054 22480 40000 22536
rect 28993 22478 40000 22480
rect 23105 22475 23171 22478
rect 28993 22475 29059 22478
rect 39200 22448 40000 22478
rect 12433 22402 12499 22405
rect 14733 22402 14799 22405
rect 18505 22402 18571 22405
rect 12433 22400 18571 22402
rect 12433 22344 12438 22400
rect 12494 22344 14738 22400
rect 14794 22344 18510 22400
rect 18566 22344 18571 22400
rect 12433 22342 18571 22344
rect 12433 22339 12499 22342
rect 14733 22339 14799 22342
rect 18505 22339 18571 22342
rect 21173 22402 21239 22405
rect 24301 22402 24367 22405
rect 21173 22400 24367 22402
rect 21173 22344 21178 22400
rect 21234 22344 24306 22400
rect 24362 22344 24367 22400
rect 21173 22342 24367 22344
rect 21173 22339 21239 22342
rect 24301 22339 24367 22342
rect 19568 22336 19888 22337
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 22271 19888 22272
rect 10041 22266 10107 22269
rect 18781 22266 18847 22269
rect 10041 22264 18847 22266
rect 10041 22208 10046 22264
rect 10102 22208 18786 22264
rect 18842 22208 18847 22264
rect 10041 22206 18847 22208
rect 10041 22203 10107 22206
rect 18781 22203 18847 22206
rect 20437 22266 20503 22269
rect 22921 22266 22987 22269
rect 20437 22264 22987 22266
rect 20437 22208 20442 22264
rect 20498 22208 22926 22264
rect 22982 22208 22987 22264
rect 20437 22206 22987 22208
rect 20437 22203 20503 22206
rect 22921 22203 22987 22206
rect 15193 22130 15259 22133
rect 18597 22130 18663 22133
rect 20345 22130 20411 22133
rect 15193 22128 20411 22130
rect 15193 22072 15198 22128
rect 15254 22072 18602 22128
rect 18658 22072 20350 22128
rect 20406 22072 20411 22128
rect 15193 22070 20411 22072
rect 15193 22067 15259 22070
rect 18597 22067 18663 22070
rect 20345 22067 20411 22070
rect 8845 21994 8911 21997
rect 4064 21992 8911 21994
rect 4064 21936 8850 21992
rect 8906 21936 8911 21992
rect 4064 21934 8911 21936
rect 0 21858 800 21888
rect 4064 21858 4124 21934
rect 8845 21931 8911 21934
rect 18413 21994 18479 21997
rect 19885 21994 19951 21997
rect 18413 21992 19951 21994
rect 18413 21936 18418 21992
rect 18474 21936 19890 21992
rect 19946 21936 19951 21992
rect 18413 21934 19951 21936
rect 18413 21931 18479 21934
rect 19885 21931 19951 21934
rect 23381 21994 23447 21997
rect 23381 21992 35404 21994
rect 23381 21936 23386 21992
rect 23442 21936 35404 21992
rect 23381 21934 35404 21936
rect 23381 21931 23447 21934
rect 0 21798 4124 21858
rect 6269 21858 6335 21861
rect 11605 21858 11671 21861
rect 6269 21856 11671 21858
rect 6269 21800 6274 21856
rect 6330 21800 11610 21856
rect 11666 21800 11671 21856
rect 6269 21798 11671 21800
rect 0 21768 800 21798
rect 6269 21795 6335 21798
rect 11605 21795 11671 21798
rect 15561 21858 15627 21861
rect 21909 21858 21975 21861
rect 24485 21858 24551 21861
rect 15561 21856 24551 21858
rect 15561 21800 15566 21856
rect 15622 21800 21914 21856
rect 21970 21800 24490 21856
rect 24546 21800 24551 21856
rect 15561 21798 24551 21800
rect 35344 21858 35404 21934
rect 39200 21858 40000 21888
rect 35344 21798 40000 21858
rect 15561 21795 15627 21798
rect 21909 21795 21975 21798
rect 24485 21795 24551 21798
rect 4208 21792 4528 21793
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 21727 4528 21728
rect 34928 21792 35248 21793
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 39200 21768 40000 21798
rect 34928 21727 35248 21728
rect 18781 21722 18847 21725
rect 21357 21722 21423 21725
rect 18781 21720 21423 21722
rect 18781 21664 18786 21720
rect 18842 21664 21362 21720
rect 21418 21664 21423 21720
rect 18781 21662 21423 21664
rect 18781 21659 18847 21662
rect 21357 21659 21423 21662
rect 19149 21586 19215 21589
rect 19609 21586 19675 21589
rect 19149 21584 19675 21586
rect 19149 21528 19154 21584
rect 19210 21528 19614 21584
rect 19670 21528 19675 21584
rect 19149 21526 19675 21528
rect 19149 21523 19215 21526
rect 19609 21523 19675 21526
rect 10961 21450 11027 21453
rect 13077 21450 13143 21453
rect 10961 21448 13143 21450
rect 10961 21392 10966 21448
rect 11022 21392 13082 21448
rect 13138 21392 13143 21448
rect 10961 21390 13143 21392
rect 10961 21387 11027 21390
rect 13077 21387 13143 21390
rect 20437 21450 20503 21453
rect 27153 21450 27219 21453
rect 20437 21448 27219 21450
rect 20437 21392 20442 21448
rect 20498 21392 27158 21448
rect 27214 21392 27219 21448
rect 20437 21390 27219 21392
rect 20437 21387 20503 21390
rect 27153 21387 27219 21390
rect 19568 21248 19888 21249
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 21183 19888 21184
rect 18781 21042 18847 21045
rect 21081 21042 21147 21045
rect 18781 21040 21147 21042
rect 18781 20984 18786 21040
rect 18842 20984 21086 21040
rect 21142 20984 21147 21040
rect 18781 20982 21147 20984
rect 18781 20979 18847 20982
rect 21081 20979 21147 20982
rect 16665 20906 16731 20909
rect 18965 20906 19031 20909
rect 16665 20904 19031 20906
rect 16665 20848 16670 20904
rect 16726 20848 18970 20904
rect 19026 20848 19031 20904
rect 16665 20846 19031 20848
rect 16665 20843 16731 20846
rect 18965 20843 19031 20846
rect 15878 20770 15884 20772
rect 11332 20710 15884 20770
rect 4208 20704 4528 20705
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 20639 4528 20640
rect 0 20498 800 20528
rect 0 20438 4906 20498
rect 0 20408 800 20438
rect 4846 20362 4906 20438
rect 11332 20362 11392 20710
rect 15878 20708 15884 20710
rect 15948 20708 15954 20772
rect 34928 20704 35248 20705
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 20639 35248 20640
rect 14273 20634 14339 20637
rect 15561 20634 15627 20637
rect 14273 20632 15627 20634
rect 14273 20576 14278 20632
rect 14334 20576 15566 20632
rect 15622 20576 15627 20632
rect 14273 20574 15627 20576
rect 14273 20571 14339 20574
rect 15561 20571 15627 20574
rect 22185 20634 22251 20637
rect 31477 20634 31543 20637
rect 22185 20632 31543 20634
rect 22185 20576 22190 20632
rect 22246 20576 31482 20632
rect 31538 20576 31543 20632
rect 22185 20574 31543 20576
rect 22185 20571 22251 20574
rect 31477 20571 31543 20574
rect 13905 20498 13971 20501
rect 19517 20498 19583 20501
rect 13905 20496 19583 20498
rect 13905 20440 13910 20496
rect 13966 20440 19522 20496
rect 19578 20440 19583 20496
rect 13905 20438 19583 20440
rect 13905 20435 13971 20438
rect 19517 20435 19583 20438
rect 35617 20498 35683 20501
rect 39200 20498 40000 20528
rect 35617 20496 40000 20498
rect 35617 20440 35622 20496
rect 35678 20440 40000 20496
rect 35617 20438 40000 20440
rect 35617 20435 35683 20438
rect 39200 20408 40000 20438
rect 4846 20302 11392 20362
rect 11881 20362 11947 20365
rect 15653 20362 15719 20365
rect 11881 20360 15719 20362
rect 11881 20304 11886 20360
rect 11942 20304 15658 20360
rect 15714 20304 15719 20360
rect 11881 20302 15719 20304
rect 11881 20299 11947 20302
rect 15653 20299 15719 20302
rect 31109 20362 31175 20365
rect 37733 20362 37799 20365
rect 31109 20360 37799 20362
rect 31109 20304 31114 20360
rect 31170 20304 37738 20360
rect 37794 20304 37799 20360
rect 31109 20302 37799 20304
rect 31109 20299 31175 20302
rect 37733 20299 37799 20302
rect 19568 20160 19888 20161
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 20095 19888 20096
rect 9029 19954 9095 19957
rect 22461 19954 22527 19957
rect 9029 19952 22527 19954
rect 9029 19896 9034 19952
rect 9090 19896 22466 19952
rect 22522 19896 22527 19952
rect 9029 19894 22527 19896
rect 9029 19891 9095 19894
rect 22461 19891 22527 19894
rect 24710 19892 24716 19956
rect 24780 19954 24786 19956
rect 35433 19954 35499 19957
rect 24780 19952 35499 19954
rect 24780 19896 35438 19952
rect 35494 19896 35499 19952
rect 24780 19894 35499 19896
rect 24780 19892 24786 19894
rect 35433 19891 35499 19894
rect 18137 19818 18203 19821
rect 21081 19818 21147 19821
rect 18137 19816 21147 19818
rect 18137 19760 18142 19816
rect 18198 19760 21086 19816
rect 21142 19760 21147 19816
rect 18137 19758 21147 19760
rect 18137 19755 18203 19758
rect 21081 19755 21147 19758
rect 4208 19616 4528 19617
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 19551 4528 19552
rect 34928 19616 35248 19617
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 19551 35248 19552
rect 13629 19546 13695 19549
rect 14457 19546 14523 19549
rect 21633 19546 21699 19549
rect 13629 19544 21699 19546
rect 13629 19488 13634 19544
rect 13690 19488 14462 19544
rect 14518 19488 21638 19544
rect 21694 19488 21699 19544
rect 13629 19486 21699 19488
rect 13629 19483 13695 19486
rect 14457 19483 14523 19486
rect 21633 19483 21699 19486
rect 4613 19410 4679 19413
rect 6085 19410 6151 19413
rect 4613 19408 6151 19410
rect 4613 19352 4618 19408
rect 4674 19352 6090 19408
rect 6146 19352 6151 19408
rect 4613 19350 6151 19352
rect 4613 19347 4679 19350
rect 6085 19347 6151 19350
rect 12985 19410 13051 19413
rect 17309 19410 17375 19413
rect 12985 19408 17375 19410
rect 12985 19352 12990 19408
rect 13046 19352 17314 19408
rect 17370 19352 17375 19408
rect 12985 19350 17375 19352
rect 12985 19347 13051 19350
rect 17309 19347 17375 19350
rect 19149 19274 19215 19277
rect 23841 19274 23907 19277
rect 19149 19272 23907 19274
rect 19149 19216 19154 19272
rect 19210 19216 23846 19272
rect 23902 19216 23907 19272
rect 19149 19214 23907 19216
rect 19149 19211 19215 19214
rect 23841 19211 23907 19214
rect 0 19138 800 19168
rect 1761 19138 1827 19141
rect 0 19136 1827 19138
rect 0 19080 1766 19136
rect 1822 19080 1827 19136
rect 0 19078 1827 19080
rect 0 19048 800 19078
rect 1761 19075 1827 19078
rect 2865 19138 2931 19141
rect 4429 19138 4495 19141
rect 2865 19136 4495 19138
rect 2865 19080 2870 19136
rect 2926 19080 4434 19136
rect 4490 19080 4495 19136
rect 2865 19078 4495 19080
rect 2865 19075 2931 19078
rect 4429 19075 4495 19078
rect 22737 19138 22803 19141
rect 39200 19138 40000 19168
rect 22737 19136 40000 19138
rect 22737 19080 22742 19136
rect 22798 19080 40000 19136
rect 22737 19078 40000 19080
rect 22737 19075 22803 19078
rect 19568 19072 19888 19073
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 39200 19048 40000 19078
rect 19568 19007 19888 19008
rect 13721 18866 13787 18869
rect 16297 18866 16363 18869
rect 13721 18864 16363 18866
rect 13721 18808 13726 18864
rect 13782 18808 16302 18864
rect 16358 18808 16363 18864
rect 13721 18806 16363 18808
rect 13721 18803 13787 18806
rect 16297 18803 16363 18806
rect 24945 18594 25011 18597
rect 30097 18594 30163 18597
rect 24945 18592 30163 18594
rect 24945 18536 24950 18592
rect 25006 18536 30102 18592
rect 30158 18536 30163 18592
rect 24945 18534 30163 18536
rect 24945 18531 25011 18534
rect 30097 18531 30163 18534
rect 4208 18528 4528 18529
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 18463 4528 18464
rect 34928 18528 35248 18529
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 18463 35248 18464
rect 14457 18458 14523 18461
rect 17953 18458 18019 18461
rect 14457 18456 18019 18458
rect 14457 18400 14462 18456
rect 14518 18400 17958 18456
rect 18014 18400 18019 18456
rect 14457 18398 18019 18400
rect 14457 18395 14523 18398
rect 17953 18395 18019 18398
rect 11421 18186 11487 18189
rect 11421 18184 12082 18186
rect 11421 18128 11426 18184
rect 11482 18128 12082 18184
rect 11421 18126 12082 18128
rect 11421 18123 11487 18126
rect 3877 18050 3943 18053
rect 11881 18050 11947 18053
rect 3877 18048 11947 18050
rect 3877 17992 3882 18048
rect 3938 17992 11886 18048
rect 11942 17992 11947 18048
rect 3877 17990 11947 17992
rect 12022 18050 12082 18126
rect 14825 18050 14891 18053
rect 15561 18050 15627 18053
rect 12022 18048 15627 18050
rect 12022 17992 14830 18048
rect 14886 17992 15566 18048
rect 15622 17992 15627 18048
rect 12022 17990 15627 17992
rect 3877 17987 3943 17990
rect 11881 17987 11947 17990
rect 14825 17987 14891 17990
rect 15561 17987 15627 17990
rect 19568 17984 19888 17985
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 17919 19888 17920
rect 9673 17914 9739 17917
rect 1350 17912 9739 17914
rect 1350 17856 9678 17912
rect 9734 17856 9739 17912
rect 1350 17854 9739 17856
rect 0 17778 800 17808
rect 1350 17778 1410 17854
rect 9673 17851 9739 17854
rect 20069 17914 20135 17917
rect 20478 17914 20484 17916
rect 20069 17912 20484 17914
rect 20069 17856 20074 17912
rect 20130 17856 20484 17912
rect 20069 17854 20484 17856
rect 20069 17851 20135 17854
rect 20478 17852 20484 17854
rect 20548 17852 20554 17916
rect 21030 17852 21036 17916
rect 21100 17914 21106 17916
rect 22185 17914 22251 17917
rect 21100 17912 22251 17914
rect 21100 17856 22190 17912
rect 22246 17856 22251 17912
rect 21100 17854 22251 17856
rect 21100 17852 21106 17854
rect 22185 17851 22251 17854
rect 27061 17914 27127 17917
rect 34513 17914 34579 17917
rect 27061 17912 34579 17914
rect 27061 17856 27066 17912
rect 27122 17856 34518 17912
rect 34574 17856 34579 17912
rect 27061 17854 34579 17856
rect 27061 17851 27127 17854
rect 34513 17851 34579 17854
rect 0 17718 1410 17778
rect 4889 17778 4955 17781
rect 8385 17778 8451 17781
rect 4889 17776 8451 17778
rect 4889 17720 4894 17776
rect 4950 17720 8390 17776
rect 8446 17720 8451 17776
rect 4889 17718 8451 17720
rect 0 17688 800 17718
rect 4889 17715 4955 17718
rect 8385 17715 8451 17718
rect 35249 17778 35315 17781
rect 39200 17778 40000 17808
rect 35249 17776 40000 17778
rect 35249 17720 35254 17776
rect 35310 17720 40000 17776
rect 35249 17718 40000 17720
rect 35249 17715 35315 17718
rect 39200 17688 40000 17718
rect 4208 17440 4528 17441
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 17375 4528 17376
rect 34928 17440 35248 17441
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 17375 35248 17376
rect 24117 17234 24183 17237
rect 28993 17234 29059 17237
rect 24117 17232 29059 17234
rect 24117 17176 24122 17232
rect 24178 17176 28998 17232
rect 29054 17176 29059 17232
rect 24117 17174 29059 17176
rect 24117 17171 24183 17174
rect 28993 17171 29059 17174
rect 1393 16962 1459 16965
rect 4889 16962 4955 16965
rect 1393 16960 4955 16962
rect 1393 16904 1398 16960
rect 1454 16904 4894 16960
rect 4950 16904 4955 16960
rect 1393 16902 4955 16904
rect 1393 16899 1459 16902
rect 4889 16899 4955 16902
rect 19568 16896 19888 16897
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 16831 19888 16832
rect 2221 16554 2287 16557
rect 19149 16554 19215 16557
rect 21214 16554 21220 16556
rect 2221 16552 7666 16554
rect 2221 16496 2226 16552
rect 2282 16496 7666 16552
rect 2221 16494 7666 16496
rect 2221 16491 2287 16494
rect 0 16418 800 16448
rect 7606 16418 7666 16494
rect 19149 16552 21220 16554
rect 19149 16496 19154 16552
rect 19210 16496 21220 16552
rect 19149 16494 21220 16496
rect 19149 16491 19215 16494
rect 21214 16492 21220 16494
rect 21284 16492 21290 16556
rect 22645 16418 22711 16421
rect 0 16358 4124 16418
rect 7606 16416 22711 16418
rect 7606 16360 22650 16416
rect 22706 16360 22711 16416
rect 7606 16358 22711 16360
rect 0 16328 800 16358
rect 4064 16146 4124 16358
rect 22645 16355 22711 16358
rect 35341 16418 35407 16421
rect 39200 16418 40000 16448
rect 35341 16416 40000 16418
rect 35341 16360 35346 16416
rect 35402 16360 40000 16416
rect 35341 16358 40000 16360
rect 35341 16355 35407 16358
rect 4208 16352 4528 16353
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 16287 4528 16288
rect 34928 16352 35248 16353
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 39200 16328 40000 16358
rect 34928 16287 35248 16288
rect 7925 16282 7991 16285
rect 10225 16282 10291 16285
rect 7925 16280 10291 16282
rect 7925 16224 7930 16280
rect 7986 16224 10230 16280
rect 10286 16224 10291 16280
rect 7925 16222 10291 16224
rect 7925 16219 7991 16222
rect 10225 16219 10291 16222
rect 11973 16146 12039 16149
rect 4064 16144 12039 16146
rect 4064 16088 11978 16144
rect 12034 16088 12039 16144
rect 4064 16086 12039 16088
rect 11973 16083 12039 16086
rect 28625 15874 28691 15877
rect 37365 15874 37431 15877
rect 28625 15872 37431 15874
rect 28625 15816 28630 15872
rect 28686 15816 37370 15872
rect 37426 15816 37431 15872
rect 28625 15814 37431 15816
rect 28625 15811 28691 15814
rect 37365 15811 37431 15814
rect 19568 15808 19888 15809
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 15743 19888 15744
rect 15377 15738 15443 15741
rect 18045 15738 18111 15741
rect 15377 15736 18111 15738
rect 15377 15680 15382 15736
rect 15438 15680 18050 15736
rect 18106 15680 18111 15736
rect 15377 15678 18111 15680
rect 15377 15675 15443 15678
rect 18045 15675 18111 15678
rect 20846 15540 20852 15604
rect 20916 15602 20922 15604
rect 21173 15602 21239 15605
rect 20916 15600 21239 15602
rect 20916 15544 21178 15600
rect 21234 15544 21239 15600
rect 20916 15542 21239 15544
rect 20916 15540 20922 15542
rect 21173 15539 21239 15542
rect 20161 15466 20227 15469
rect 24853 15466 24919 15469
rect 20161 15464 24919 15466
rect 20161 15408 20166 15464
rect 20222 15408 24858 15464
rect 24914 15408 24919 15464
rect 20161 15406 24919 15408
rect 20161 15403 20227 15406
rect 24853 15403 24919 15406
rect 1577 15330 1643 15333
rect 1534 15328 1643 15330
rect 1534 15272 1582 15328
rect 1638 15272 1643 15328
rect 1534 15267 1643 15272
rect 0 15058 800 15088
rect 1534 15058 1594 15267
rect 4208 15264 4528 15265
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 15199 4528 15200
rect 34928 15264 35248 15265
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 15199 35248 15200
rect 18321 15194 18387 15197
rect 22502 15194 22508 15196
rect 18321 15192 22508 15194
rect 18321 15136 18326 15192
rect 18382 15136 22508 15192
rect 18321 15134 22508 15136
rect 18321 15131 18387 15134
rect 22502 15132 22508 15134
rect 22572 15132 22578 15196
rect 24526 15132 24532 15196
rect 24596 15194 24602 15196
rect 29637 15194 29703 15197
rect 24596 15192 29703 15194
rect 24596 15136 29642 15192
rect 29698 15136 29703 15192
rect 24596 15134 29703 15136
rect 24596 15132 24602 15134
rect 29637 15131 29703 15134
rect 0 14998 1594 15058
rect 3417 15058 3483 15061
rect 10593 15058 10659 15061
rect 13813 15060 13879 15061
rect 13813 15058 13860 15060
rect 3417 15056 10659 15058
rect 3417 15000 3422 15056
rect 3478 15000 10598 15056
rect 10654 15000 10659 15056
rect 3417 14998 10659 15000
rect 13768 15056 13860 15058
rect 13768 15000 13818 15056
rect 13768 14998 13860 15000
rect 0 14968 800 14998
rect 3417 14995 3483 14998
rect 10593 14995 10659 14998
rect 13813 14996 13860 14998
rect 13924 14996 13930 15060
rect 30281 15058 30347 15061
rect 37457 15058 37523 15061
rect 39200 15058 40000 15088
rect 30281 15056 37523 15058
rect 30281 15000 30286 15056
rect 30342 15000 37462 15056
rect 37518 15000 37523 15056
rect 30281 14998 37523 15000
rect 13813 14995 13879 14996
rect 30281 14995 30347 14998
rect 37457 14995 37523 14998
rect 37598 14998 40000 15058
rect 19568 14720 19888 14721
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 14655 19888 14656
rect 11697 14514 11763 14517
rect 15285 14514 15351 14517
rect 11697 14512 15351 14514
rect 11697 14456 11702 14512
rect 11758 14456 15290 14512
rect 15346 14456 15351 14512
rect 11697 14454 15351 14456
rect 11697 14451 11763 14454
rect 15285 14451 15351 14454
rect 18965 14514 19031 14517
rect 26325 14514 26391 14517
rect 18965 14512 26391 14514
rect 18965 14456 18970 14512
rect 19026 14456 26330 14512
rect 26386 14456 26391 14512
rect 18965 14454 26391 14456
rect 18965 14451 19031 14454
rect 26325 14451 26391 14454
rect 18321 14378 18387 14381
rect 21265 14378 21331 14381
rect 18321 14376 21331 14378
rect 18321 14320 18326 14376
rect 18382 14320 21270 14376
rect 21326 14320 21331 14376
rect 18321 14318 21331 14320
rect 18321 14315 18387 14318
rect 21265 14315 21331 14318
rect 23197 14242 23263 14245
rect 22694 14240 23263 14242
rect 22694 14184 23202 14240
rect 23258 14184 23263 14240
rect 22694 14182 23263 14184
rect 4208 14176 4528 14177
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 14111 4528 14112
rect 22001 13970 22067 13973
rect 22694 13970 22754 14182
rect 23197 14179 23263 14182
rect 34928 14176 35248 14177
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 14111 35248 14112
rect 22001 13968 22754 13970
rect 22001 13912 22006 13968
rect 22062 13912 22754 13968
rect 22001 13910 22754 13912
rect 23105 13970 23171 13973
rect 25129 13970 25195 13973
rect 23105 13968 25195 13970
rect 23105 13912 23110 13968
rect 23166 13912 25134 13968
rect 25190 13912 25195 13968
rect 23105 13910 25195 13912
rect 22001 13907 22067 13910
rect 23105 13907 23171 13910
rect 25129 13907 25195 13910
rect 1945 13834 2011 13837
rect 4705 13834 4771 13837
rect 1945 13832 4771 13834
rect 1945 13776 1950 13832
rect 2006 13776 4710 13832
rect 4766 13776 4771 13832
rect 1945 13774 4771 13776
rect 1945 13771 2011 13774
rect 4705 13771 4771 13774
rect 22461 13834 22527 13837
rect 37598 13834 37658 14998
rect 39200 14968 40000 14998
rect 22461 13832 37658 13834
rect 22461 13776 22466 13832
rect 22522 13776 37658 13832
rect 22461 13774 37658 13776
rect 22461 13771 22527 13774
rect 0 13698 800 13728
rect 2773 13698 2839 13701
rect 0 13696 2839 13698
rect 0 13640 2778 13696
rect 2834 13640 2839 13696
rect 0 13638 2839 13640
rect 0 13608 800 13638
rect 2773 13635 2839 13638
rect 34513 13698 34579 13701
rect 39200 13698 40000 13728
rect 34513 13696 40000 13698
rect 34513 13640 34518 13696
rect 34574 13640 40000 13696
rect 34513 13638 40000 13640
rect 34513 13635 34579 13638
rect 19568 13632 19888 13633
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 39200 13608 40000 13638
rect 19568 13567 19888 13568
rect 22093 13562 22159 13565
rect 35617 13562 35683 13565
rect 22093 13560 35683 13562
rect 22093 13504 22098 13560
rect 22154 13504 35622 13560
rect 35678 13504 35683 13560
rect 22093 13502 35683 13504
rect 22093 13499 22159 13502
rect 35617 13499 35683 13502
rect 3325 13426 3391 13429
rect 14774 13426 14780 13428
rect 3325 13424 14780 13426
rect 3325 13368 3330 13424
rect 3386 13368 14780 13424
rect 3325 13366 14780 13368
rect 3325 13363 3391 13366
rect 14774 13364 14780 13366
rect 14844 13364 14850 13428
rect 16481 13426 16547 13429
rect 23473 13426 23539 13429
rect 16481 13424 23539 13426
rect 16481 13368 16486 13424
rect 16542 13368 23478 13424
rect 23534 13368 23539 13424
rect 16481 13366 23539 13368
rect 16481 13363 16547 13366
rect 23473 13363 23539 13366
rect 14406 13228 14412 13292
rect 14476 13290 14482 13292
rect 37549 13290 37615 13293
rect 14476 13288 37615 13290
rect 14476 13232 37554 13288
rect 37610 13232 37615 13288
rect 14476 13230 37615 13232
rect 14476 13228 14482 13230
rect 37549 13227 37615 13230
rect 4208 13088 4528 13089
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 13023 4528 13024
rect 34928 13088 35248 13089
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 34928 13023 35248 13024
rect 19568 12544 19888 12545
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 19568 12479 19888 12480
rect 9622 12412 9628 12476
rect 9692 12474 9698 12476
rect 15694 12474 15700 12476
rect 9692 12414 15700 12474
rect 9692 12412 9698 12414
rect 15694 12412 15700 12414
rect 15764 12412 15770 12476
rect 32121 12474 32187 12477
rect 33133 12474 33199 12477
rect 32121 12472 33199 12474
rect 32121 12416 32126 12472
rect 32182 12416 33138 12472
rect 33194 12416 33199 12472
rect 32121 12414 33199 12416
rect 32121 12411 32187 12414
rect 33133 12411 33199 12414
rect 0 12338 800 12368
rect 2773 12338 2839 12341
rect 0 12336 2839 12338
rect 0 12280 2778 12336
rect 2834 12280 2839 12336
rect 0 12278 2839 12280
rect 0 12248 800 12278
rect 2773 12275 2839 12278
rect 3693 12338 3759 12341
rect 13169 12338 13235 12341
rect 39200 12338 40000 12368
rect 3693 12336 13235 12338
rect 3693 12280 3698 12336
rect 3754 12280 13174 12336
rect 13230 12280 13235 12336
rect 3693 12278 13235 12280
rect 3693 12275 3759 12278
rect 13169 12275 13235 12278
rect 39070 12278 40000 12338
rect 28942 12140 28948 12204
rect 29012 12202 29018 12204
rect 39070 12202 39130 12278
rect 39200 12248 40000 12278
rect 29012 12142 39130 12202
rect 29012 12140 29018 12142
rect 4208 12000 4528 12001
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 11935 4528 11936
rect 34928 12000 35248 12001
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 34928 11935 35248 11936
rect 2773 11794 2839 11797
rect 9622 11794 9628 11796
rect 2773 11792 9628 11794
rect 2773 11736 2778 11792
rect 2834 11736 9628 11792
rect 2773 11734 9628 11736
rect 2773 11731 2839 11734
rect 9622 11732 9628 11734
rect 9692 11732 9698 11796
rect 0 11658 800 11688
rect 3325 11658 3391 11661
rect 0 11656 3391 11658
rect 0 11600 3330 11656
rect 3386 11600 3391 11656
rect 0 11598 3391 11600
rect 0 11568 800 11598
rect 3325 11595 3391 11598
rect 19568 11456 19888 11457
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 11391 19888 11392
rect 22645 11250 22711 11253
rect 28942 11250 28948 11252
rect 22645 11248 28948 11250
rect 22645 11192 22650 11248
rect 22706 11192 28948 11248
rect 22645 11190 28948 11192
rect 22645 11187 22711 11190
rect 28942 11188 28948 11190
rect 29012 11188 29018 11252
rect 23933 11114 23999 11117
rect 30005 11114 30071 11117
rect 23933 11112 30071 11114
rect 23933 11056 23938 11112
rect 23994 11056 30010 11112
rect 30066 11056 30071 11112
rect 23933 11054 30071 11056
rect 23933 11051 23999 11054
rect 30005 11051 30071 11054
rect 35433 10978 35499 10981
rect 39200 10978 40000 11008
rect 35433 10976 40000 10978
rect 35433 10920 35438 10976
rect 35494 10920 40000 10976
rect 35433 10918 40000 10920
rect 35433 10915 35499 10918
rect 4208 10912 4528 10913
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 10847 4528 10848
rect 34928 10912 35248 10913
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 39200 10888 40000 10918
rect 34928 10847 35248 10848
rect 2681 10570 2747 10573
rect 26877 10570 26943 10573
rect 2681 10568 26943 10570
rect 2681 10512 2686 10568
rect 2742 10512 26882 10568
rect 26938 10512 26943 10568
rect 2681 10510 26943 10512
rect 2681 10507 2747 10510
rect 26877 10507 26943 10510
rect 19568 10368 19888 10369
rect 0 10298 800 10328
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 10303 19888 10304
rect 3877 10298 3943 10301
rect 0 10296 3943 10298
rect 0 10240 3882 10296
rect 3938 10240 3943 10296
rect 0 10238 3943 10240
rect 0 10208 800 10238
rect 3877 10235 3943 10238
rect 19977 10298 20043 10301
rect 39200 10298 40000 10328
rect 19977 10296 40000 10298
rect 19977 10240 19982 10296
rect 20038 10240 40000 10296
rect 19977 10238 40000 10240
rect 19977 10235 20043 10238
rect 39200 10208 40000 10238
rect 2037 10162 2103 10165
rect 7097 10162 7163 10165
rect 2037 10160 7163 10162
rect 2037 10104 2042 10160
rect 2098 10104 7102 10160
rect 7158 10104 7163 10160
rect 2037 10102 7163 10104
rect 2037 10099 2103 10102
rect 7097 10099 7163 10102
rect 3141 10026 3207 10029
rect 22093 10026 22159 10029
rect 3141 10024 22159 10026
rect 3141 9968 3146 10024
rect 3202 9968 22098 10024
rect 22154 9968 22159 10024
rect 3141 9966 22159 9968
rect 3141 9963 3207 9966
rect 22093 9963 22159 9966
rect 4208 9824 4528 9825
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 9759 4528 9760
rect 34928 9824 35248 9825
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 34928 9759 35248 9760
rect 16113 9754 16179 9757
rect 17033 9754 17099 9757
rect 24342 9754 24348 9756
rect 16113 9752 17099 9754
rect 16113 9696 16118 9752
rect 16174 9696 17038 9752
rect 17094 9696 17099 9752
rect 16113 9694 17099 9696
rect 16113 9691 16179 9694
rect 17033 9691 17099 9694
rect 19888 9694 24348 9754
rect 19425 9482 19491 9485
rect 19888 9482 19948 9694
rect 24342 9692 24348 9694
rect 24412 9692 24418 9756
rect 30281 9754 30347 9757
rect 30281 9752 30482 9754
rect 30281 9696 30286 9752
rect 30342 9696 30482 9752
rect 30281 9694 30482 9696
rect 30281 9691 30347 9694
rect 30422 9620 30482 9694
rect 30414 9556 30420 9620
rect 30484 9556 30490 9620
rect 19425 9480 19948 9482
rect 19425 9424 19430 9480
rect 19486 9424 19948 9480
rect 19425 9422 19948 9424
rect 19425 9419 19491 9422
rect 19568 9280 19888 9281
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 9215 19888 9216
rect 8293 9074 8359 9077
rect 18505 9074 18571 9077
rect 8293 9072 18571 9074
rect 8293 9016 8298 9072
rect 8354 9016 18510 9072
rect 18566 9016 18571 9072
rect 8293 9014 18571 9016
rect 8293 9011 8359 9014
rect 18505 9011 18571 9014
rect 18873 9074 18939 9077
rect 36353 9074 36419 9077
rect 18873 9072 36419 9074
rect 18873 9016 18878 9072
rect 18934 9016 36358 9072
rect 36414 9016 36419 9072
rect 18873 9014 36419 9016
rect 18873 9011 18939 9014
rect 36353 9011 36419 9014
rect 0 8938 800 8968
rect 1577 8938 1643 8941
rect 39200 8938 40000 8968
rect 0 8936 1643 8938
rect 0 8880 1582 8936
rect 1638 8880 1643 8936
rect 0 8878 1643 8880
rect 0 8848 800 8878
rect 1577 8875 1643 8878
rect 39070 8878 40000 8938
rect 4208 8736 4528 8737
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 8671 4528 8672
rect 34928 8736 35248 8737
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 8671 35248 8672
rect 13261 8530 13327 8533
rect 15561 8530 15627 8533
rect 13261 8528 15627 8530
rect 13261 8472 13266 8528
rect 13322 8472 15566 8528
rect 15622 8472 15627 8528
rect 13261 8470 15627 8472
rect 13261 8467 13327 8470
rect 15561 8467 15627 8470
rect 7189 8394 7255 8397
rect 39070 8394 39130 8878
rect 39200 8848 40000 8878
rect 7189 8392 39130 8394
rect 7189 8336 7194 8392
rect 7250 8336 39130 8392
rect 7189 8334 39130 8336
rect 7189 8331 7255 8334
rect 19568 8192 19888 8193
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 8127 19888 8128
rect 1393 7850 1459 7853
rect 24669 7850 24735 7853
rect 1393 7848 24735 7850
rect 1393 7792 1398 7848
rect 1454 7792 24674 7848
rect 24730 7792 24735 7848
rect 1393 7790 24735 7792
rect 1393 7787 1459 7790
rect 24669 7787 24735 7790
rect 26509 7850 26575 7853
rect 26509 7848 35450 7850
rect 26509 7792 26514 7848
rect 26570 7792 35450 7848
rect 26509 7790 35450 7792
rect 26509 7787 26575 7790
rect 24393 7714 24459 7717
rect 25773 7714 25839 7717
rect 24393 7712 25839 7714
rect 24393 7656 24398 7712
rect 24454 7656 25778 7712
rect 25834 7656 25839 7712
rect 24393 7654 25839 7656
rect 24393 7651 24459 7654
rect 25773 7651 25839 7654
rect 4208 7648 4528 7649
rect 0 7578 800 7608
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 7583 4528 7584
rect 34928 7648 35248 7649
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 7583 35248 7584
rect 5993 7578 6059 7581
rect 20294 7578 20300 7580
rect 0 7518 3986 7578
rect 0 7488 800 7518
rect 3926 7306 3986 7518
rect 5993 7576 20300 7578
rect 5993 7520 5998 7576
rect 6054 7520 20300 7576
rect 5993 7518 20300 7520
rect 5993 7515 6059 7518
rect 20294 7516 20300 7518
rect 20364 7516 20370 7580
rect 25037 7578 25103 7581
rect 26693 7578 26759 7581
rect 34513 7578 34579 7581
rect 25037 7576 26759 7578
rect 25037 7520 25042 7576
rect 25098 7520 26698 7576
rect 26754 7520 26759 7576
rect 25037 7518 26759 7520
rect 25037 7515 25103 7518
rect 26693 7515 26759 7518
rect 26926 7576 34579 7578
rect 26926 7520 34518 7576
rect 34574 7520 34579 7576
rect 26926 7518 34579 7520
rect 35390 7578 35450 7790
rect 39200 7578 40000 7608
rect 35390 7518 40000 7578
rect 23473 7442 23539 7445
rect 26926 7442 26986 7518
rect 34513 7515 34579 7518
rect 39200 7488 40000 7518
rect 23473 7440 26986 7442
rect 23473 7384 23478 7440
rect 23534 7384 26986 7440
rect 23473 7382 26986 7384
rect 23473 7379 23539 7382
rect 12341 7306 12407 7309
rect 3926 7304 12407 7306
rect 3926 7248 12346 7304
rect 12402 7248 12407 7304
rect 3926 7246 12407 7248
rect 12341 7243 12407 7246
rect 13445 7306 13511 7309
rect 23841 7306 23907 7309
rect 13445 7304 23907 7306
rect 13445 7248 13450 7304
rect 13506 7248 23846 7304
rect 23902 7248 23907 7304
rect 13445 7246 23907 7248
rect 13445 7243 13511 7246
rect 23841 7243 23907 7246
rect 19568 7104 19888 7105
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 7039 19888 7040
rect 4061 6898 4127 6901
rect 19425 6898 19491 6901
rect 4061 6896 19491 6898
rect 4061 6840 4066 6896
rect 4122 6840 19430 6896
rect 19486 6840 19491 6896
rect 4061 6838 19491 6840
rect 4061 6835 4127 6838
rect 19425 6835 19491 6838
rect 24945 6898 25011 6901
rect 26141 6898 26207 6901
rect 24945 6896 26207 6898
rect 24945 6840 24950 6896
rect 25006 6840 26146 6896
rect 26202 6840 26207 6896
rect 24945 6838 26207 6840
rect 24945 6835 25011 6838
rect 26141 6835 26207 6838
rect 4208 6560 4528 6561
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 6495 4528 6496
rect 34928 6560 35248 6561
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 6495 35248 6496
rect 7833 6354 7899 6357
rect 25957 6354 26023 6357
rect 7833 6352 26023 6354
rect 7833 6296 7838 6352
rect 7894 6296 25962 6352
rect 26018 6296 26023 6352
rect 7833 6294 26023 6296
rect 7833 6291 7899 6294
rect 25957 6291 26023 6294
rect 36261 6354 36327 6357
rect 36261 6352 37658 6354
rect 36261 6296 36266 6352
rect 36322 6296 37658 6352
rect 36261 6294 37658 6296
rect 36261 6291 36327 6294
rect 0 6218 800 6248
rect 4061 6218 4127 6221
rect 0 6216 4127 6218
rect 0 6160 4066 6216
rect 4122 6160 4127 6216
rect 0 6158 4127 6160
rect 0 6128 800 6158
rect 4061 6155 4127 6158
rect 4797 6218 4863 6221
rect 27981 6218 28047 6221
rect 37365 6218 37431 6221
rect 4797 6216 37431 6218
rect 4797 6160 4802 6216
rect 4858 6160 27986 6216
rect 28042 6160 37370 6216
rect 37426 6160 37431 6216
rect 4797 6158 37431 6160
rect 37598 6218 37658 6294
rect 39200 6218 40000 6248
rect 37598 6158 40000 6218
rect 4797 6155 4863 6158
rect 27981 6155 28047 6158
rect 37365 6155 37431 6158
rect 39200 6128 40000 6158
rect 19568 6016 19888 6017
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 5951 19888 5952
rect 26141 5674 26207 5677
rect 35985 5674 36051 5677
rect 26141 5672 36051 5674
rect 26141 5616 26146 5672
rect 26202 5616 35990 5672
rect 36046 5616 36051 5672
rect 26141 5614 36051 5616
rect 26141 5611 26207 5614
rect 35985 5611 36051 5614
rect 13629 5538 13695 5541
rect 14733 5538 14799 5541
rect 13629 5536 14799 5538
rect 13629 5480 13634 5536
rect 13690 5480 14738 5536
rect 14794 5480 14799 5536
rect 13629 5478 14799 5480
rect 13629 5475 13695 5478
rect 14733 5475 14799 5478
rect 4208 5472 4528 5473
rect 4208 5408 4216 5472
rect 4280 5408 4296 5472
rect 4360 5408 4376 5472
rect 4440 5408 4456 5472
rect 4520 5408 4528 5472
rect 4208 5407 4528 5408
rect 34928 5472 35248 5473
rect 34928 5408 34936 5472
rect 35000 5408 35016 5472
rect 35080 5408 35096 5472
rect 35160 5408 35176 5472
rect 35240 5408 35248 5472
rect 34928 5407 35248 5408
rect 16021 5266 16087 5269
rect 32673 5266 32739 5269
rect 16021 5264 32739 5266
rect 16021 5208 16026 5264
rect 16082 5208 32678 5264
rect 32734 5208 32739 5264
rect 16021 5206 32739 5208
rect 16021 5203 16087 5206
rect 32673 5203 32739 5206
rect 3509 5130 3575 5133
rect 23013 5130 23079 5133
rect 3509 5128 23079 5130
rect 3509 5072 3514 5128
rect 3570 5072 23018 5128
rect 23074 5072 23079 5128
rect 3509 5070 23079 5072
rect 3509 5067 3575 5070
rect 23013 5067 23079 5070
rect 19568 4928 19888 4929
rect 0 4858 800 4888
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 19568 4863 19888 4864
rect 3417 4858 3483 4861
rect 13997 4860 14063 4861
rect 13997 4858 14044 4860
rect 0 4856 3483 4858
rect 0 4800 3422 4856
rect 3478 4800 3483 4856
rect 0 4798 3483 4800
rect 13952 4856 14044 4858
rect 13952 4800 14002 4856
rect 13952 4798 14044 4800
rect 0 4768 800 4798
rect 3417 4795 3483 4798
rect 13997 4796 14044 4798
rect 14108 4796 14114 4860
rect 28942 4796 28948 4860
rect 29012 4858 29018 4860
rect 39200 4858 40000 4888
rect 29012 4798 40000 4858
rect 29012 4796 29018 4798
rect 13997 4795 14063 4796
rect 39200 4768 40000 4798
rect 9622 4524 9628 4588
rect 9692 4586 9698 4588
rect 17902 4586 17908 4588
rect 9692 4526 17908 4586
rect 9692 4524 9698 4526
rect 17902 4524 17908 4526
rect 17972 4524 17978 4588
rect 4208 4384 4528 4385
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 4319 4528 4320
rect 34928 4384 35248 4385
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 4319 35248 4320
rect 9581 4316 9647 4317
rect 9581 4312 9628 4316
rect 9692 4314 9698 4316
rect 9581 4256 9586 4312
rect 9581 4252 9628 4256
rect 9692 4254 9774 4314
rect 9692 4252 9698 4254
rect 17902 4252 17908 4316
rect 17972 4314 17978 4316
rect 19241 4314 19307 4317
rect 17972 4312 19307 4314
rect 17972 4256 19246 4312
rect 19302 4256 19307 4312
rect 17972 4254 19307 4256
rect 17972 4252 17978 4254
rect 9581 4251 9647 4252
rect 19241 4251 19307 4254
rect 19425 4314 19491 4317
rect 28942 4314 28948 4316
rect 19425 4312 28948 4314
rect 19425 4256 19430 4312
rect 19486 4256 28948 4312
rect 19425 4254 28948 4256
rect 19425 4251 19491 4254
rect 28942 4252 28948 4254
rect 29012 4252 29018 4316
rect 14273 4044 14339 4045
rect 14222 4042 14228 4044
rect 14182 3982 14228 4042
rect 14292 4040 14339 4044
rect 14334 3984 14339 4040
rect 14222 3980 14228 3982
rect 14292 3980 14339 3984
rect 14273 3979 14339 3980
rect 15837 4042 15903 4045
rect 17033 4042 17099 4045
rect 15837 4040 17099 4042
rect 15837 3984 15842 4040
rect 15898 3984 17038 4040
rect 17094 3984 17099 4040
rect 15837 3982 17099 3984
rect 15837 3979 15903 3982
rect 17033 3979 17099 3982
rect 19568 3840 19888 3841
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 3775 19888 3776
rect 0 3498 800 3528
rect 3693 3498 3759 3501
rect 0 3496 3759 3498
rect 0 3440 3698 3496
rect 3754 3440 3759 3496
rect 0 3438 3759 3440
rect 0 3408 800 3438
rect 3693 3435 3759 3438
rect 35801 3498 35867 3501
rect 39200 3498 40000 3528
rect 35801 3496 40000 3498
rect 35801 3440 35806 3496
rect 35862 3440 40000 3496
rect 35801 3438 40000 3440
rect 35801 3435 35867 3438
rect 39200 3408 40000 3438
rect 18229 3362 18295 3365
rect 19425 3362 19491 3365
rect 18229 3360 19491 3362
rect 18229 3304 18234 3360
rect 18290 3304 19430 3360
rect 19486 3304 19491 3360
rect 18229 3302 19491 3304
rect 18229 3299 18295 3302
rect 19425 3299 19491 3302
rect 4208 3296 4528 3297
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 3231 4528 3232
rect 34928 3296 35248 3297
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 3231 35248 3232
rect 19568 2752 19888 2753
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2687 19888 2688
rect 28441 2684 28507 2685
rect 28390 2682 28396 2684
rect 28350 2622 28396 2682
rect 28460 2680 28507 2684
rect 28502 2624 28507 2680
rect 28390 2620 28396 2622
rect 28460 2620 28507 2624
rect 28441 2619 28507 2620
rect 23749 2410 23815 2413
rect 3374 2408 23815 2410
rect 3374 2352 23754 2408
rect 23810 2352 23815 2408
rect 3374 2350 23815 2352
rect 0 2138 800 2168
rect 3374 2138 3434 2350
rect 23749 2347 23815 2350
rect 18965 2274 19031 2277
rect 31293 2274 31359 2277
rect 18965 2272 31359 2274
rect 18965 2216 18970 2272
rect 19026 2216 31298 2272
rect 31354 2216 31359 2272
rect 18965 2214 31359 2216
rect 18965 2211 19031 2214
rect 31293 2211 31359 2214
rect 4208 2208 4528 2209
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2143 4528 2144
rect 34928 2208 35248 2209
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2143 35248 2144
rect 39200 2138 40000 2168
rect 0 2078 3434 2138
rect 35390 2078 40000 2138
rect 0 2048 800 2078
rect 29637 2002 29703 2005
rect 35390 2002 35450 2078
rect 39200 2048 40000 2078
rect 29637 2000 35450 2002
rect 29637 1944 29642 2000
rect 29698 1944 35450 2000
rect 29637 1942 35450 1944
rect 29637 1939 29703 1942
rect 30373 916 30439 917
rect 30373 914 30420 916
rect 30328 912 30420 914
rect 30328 856 30378 912
rect 30328 854 30420 856
rect 30373 852 30420 854
rect 30484 852 30490 916
rect 30373 851 30439 852
rect 0 778 800 808
rect 3417 778 3483 781
rect 39200 778 40000 808
rect 0 776 3483 778
rect 0 720 3422 776
rect 3478 720 3483 776
rect 0 718 3483 720
rect 0 688 800 718
rect 3417 715 3483 718
rect 39070 718 40000 778
rect 22737 234 22803 237
rect 39070 234 39130 718
rect 39200 688 40000 718
rect 22737 232 39130 234
rect 22737 176 22742 232
rect 22798 176 39130 232
rect 22737 174 39130 176
rect 22737 171 22803 174
<< via3 >>
rect 19576 77820 19640 77824
rect 19576 77764 19580 77820
rect 19580 77764 19636 77820
rect 19636 77764 19640 77820
rect 19576 77760 19640 77764
rect 19656 77820 19720 77824
rect 19656 77764 19660 77820
rect 19660 77764 19716 77820
rect 19716 77764 19720 77820
rect 19656 77760 19720 77764
rect 19736 77820 19800 77824
rect 19736 77764 19740 77820
rect 19740 77764 19796 77820
rect 19796 77764 19800 77820
rect 19736 77760 19800 77764
rect 19816 77820 19880 77824
rect 19816 77764 19820 77820
rect 19820 77764 19876 77820
rect 19876 77764 19880 77820
rect 19816 77760 19880 77764
rect 4216 77276 4280 77280
rect 4216 77220 4220 77276
rect 4220 77220 4276 77276
rect 4276 77220 4280 77276
rect 4216 77216 4280 77220
rect 4296 77276 4360 77280
rect 4296 77220 4300 77276
rect 4300 77220 4356 77276
rect 4356 77220 4360 77276
rect 4296 77216 4360 77220
rect 4376 77276 4440 77280
rect 4376 77220 4380 77276
rect 4380 77220 4436 77276
rect 4436 77220 4440 77276
rect 4376 77216 4440 77220
rect 4456 77276 4520 77280
rect 4456 77220 4460 77276
rect 4460 77220 4516 77276
rect 4516 77220 4520 77276
rect 4456 77216 4520 77220
rect 34936 77276 35000 77280
rect 34936 77220 34940 77276
rect 34940 77220 34996 77276
rect 34996 77220 35000 77276
rect 34936 77216 35000 77220
rect 35016 77276 35080 77280
rect 35016 77220 35020 77276
rect 35020 77220 35076 77276
rect 35076 77220 35080 77276
rect 35016 77216 35080 77220
rect 35096 77276 35160 77280
rect 35096 77220 35100 77276
rect 35100 77220 35156 77276
rect 35156 77220 35160 77276
rect 35096 77216 35160 77220
rect 35176 77276 35240 77280
rect 35176 77220 35180 77276
rect 35180 77220 35236 77276
rect 35236 77220 35240 77276
rect 35176 77216 35240 77220
rect 19576 76732 19640 76736
rect 19576 76676 19580 76732
rect 19580 76676 19636 76732
rect 19636 76676 19640 76732
rect 19576 76672 19640 76676
rect 19656 76732 19720 76736
rect 19656 76676 19660 76732
rect 19660 76676 19716 76732
rect 19716 76676 19720 76732
rect 19656 76672 19720 76676
rect 19736 76732 19800 76736
rect 19736 76676 19740 76732
rect 19740 76676 19796 76732
rect 19796 76676 19800 76732
rect 19736 76672 19800 76676
rect 19816 76732 19880 76736
rect 19816 76676 19820 76732
rect 19820 76676 19876 76732
rect 19876 76676 19880 76732
rect 19816 76672 19880 76676
rect 4216 76188 4280 76192
rect 4216 76132 4220 76188
rect 4220 76132 4276 76188
rect 4276 76132 4280 76188
rect 4216 76128 4280 76132
rect 4296 76188 4360 76192
rect 4296 76132 4300 76188
rect 4300 76132 4356 76188
rect 4356 76132 4360 76188
rect 4296 76128 4360 76132
rect 4376 76188 4440 76192
rect 4376 76132 4380 76188
rect 4380 76132 4436 76188
rect 4436 76132 4440 76188
rect 4376 76128 4440 76132
rect 4456 76188 4520 76192
rect 4456 76132 4460 76188
rect 4460 76132 4516 76188
rect 4516 76132 4520 76188
rect 4456 76128 4520 76132
rect 34936 76188 35000 76192
rect 34936 76132 34940 76188
rect 34940 76132 34996 76188
rect 34996 76132 35000 76188
rect 34936 76128 35000 76132
rect 35016 76188 35080 76192
rect 35016 76132 35020 76188
rect 35020 76132 35076 76188
rect 35076 76132 35080 76188
rect 35016 76128 35080 76132
rect 35096 76188 35160 76192
rect 35096 76132 35100 76188
rect 35100 76132 35156 76188
rect 35156 76132 35160 76188
rect 35096 76128 35160 76132
rect 35176 76188 35240 76192
rect 35176 76132 35180 76188
rect 35180 76132 35236 76188
rect 35236 76132 35240 76188
rect 35176 76128 35240 76132
rect 19576 75644 19640 75648
rect 19576 75588 19580 75644
rect 19580 75588 19636 75644
rect 19636 75588 19640 75644
rect 19576 75584 19640 75588
rect 19656 75644 19720 75648
rect 19656 75588 19660 75644
rect 19660 75588 19716 75644
rect 19716 75588 19720 75644
rect 19656 75584 19720 75588
rect 19736 75644 19800 75648
rect 19736 75588 19740 75644
rect 19740 75588 19796 75644
rect 19796 75588 19800 75644
rect 19736 75584 19800 75588
rect 19816 75644 19880 75648
rect 19816 75588 19820 75644
rect 19820 75588 19876 75644
rect 19876 75588 19880 75644
rect 19816 75584 19880 75588
rect 4216 75100 4280 75104
rect 4216 75044 4220 75100
rect 4220 75044 4276 75100
rect 4276 75044 4280 75100
rect 4216 75040 4280 75044
rect 4296 75100 4360 75104
rect 4296 75044 4300 75100
rect 4300 75044 4356 75100
rect 4356 75044 4360 75100
rect 4296 75040 4360 75044
rect 4376 75100 4440 75104
rect 4376 75044 4380 75100
rect 4380 75044 4436 75100
rect 4436 75044 4440 75100
rect 4376 75040 4440 75044
rect 4456 75100 4520 75104
rect 4456 75044 4460 75100
rect 4460 75044 4516 75100
rect 4516 75044 4520 75100
rect 4456 75040 4520 75044
rect 34936 75100 35000 75104
rect 34936 75044 34940 75100
rect 34940 75044 34996 75100
rect 34996 75044 35000 75100
rect 34936 75040 35000 75044
rect 35016 75100 35080 75104
rect 35016 75044 35020 75100
rect 35020 75044 35076 75100
rect 35076 75044 35080 75100
rect 35016 75040 35080 75044
rect 35096 75100 35160 75104
rect 35096 75044 35100 75100
rect 35100 75044 35156 75100
rect 35156 75044 35160 75100
rect 35096 75040 35160 75044
rect 35176 75100 35240 75104
rect 35176 75044 35180 75100
rect 35180 75044 35236 75100
rect 35236 75044 35240 75100
rect 35176 75040 35240 75044
rect 19576 74556 19640 74560
rect 19576 74500 19580 74556
rect 19580 74500 19636 74556
rect 19636 74500 19640 74556
rect 19576 74496 19640 74500
rect 19656 74556 19720 74560
rect 19656 74500 19660 74556
rect 19660 74500 19716 74556
rect 19716 74500 19720 74556
rect 19656 74496 19720 74500
rect 19736 74556 19800 74560
rect 19736 74500 19740 74556
rect 19740 74500 19796 74556
rect 19796 74500 19800 74556
rect 19736 74496 19800 74500
rect 19816 74556 19880 74560
rect 19816 74500 19820 74556
rect 19820 74500 19876 74556
rect 19876 74500 19880 74556
rect 19816 74496 19880 74500
rect 4216 74012 4280 74016
rect 4216 73956 4220 74012
rect 4220 73956 4276 74012
rect 4276 73956 4280 74012
rect 4216 73952 4280 73956
rect 4296 74012 4360 74016
rect 4296 73956 4300 74012
rect 4300 73956 4356 74012
rect 4356 73956 4360 74012
rect 4296 73952 4360 73956
rect 4376 74012 4440 74016
rect 4376 73956 4380 74012
rect 4380 73956 4436 74012
rect 4436 73956 4440 74012
rect 4376 73952 4440 73956
rect 4456 74012 4520 74016
rect 4456 73956 4460 74012
rect 4460 73956 4516 74012
rect 4516 73956 4520 74012
rect 4456 73952 4520 73956
rect 34936 74012 35000 74016
rect 34936 73956 34940 74012
rect 34940 73956 34996 74012
rect 34996 73956 35000 74012
rect 34936 73952 35000 73956
rect 35016 74012 35080 74016
rect 35016 73956 35020 74012
rect 35020 73956 35076 74012
rect 35076 73956 35080 74012
rect 35016 73952 35080 73956
rect 35096 74012 35160 74016
rect 35096 73956 35100 74012
rect 35100 73956 35156 74012
rect 35156 73956 35160 74012
rect 35096 73952 35160 73956
rect 35176 74012 35240 74016
rect 35176 73956 35180 74012
rect 35180 73956 35236 74012
rect 35236 73956 35240 74012
rect 35176 73952 35240 73956
rect 19576 73468 19640 73472
rect 19576 73412 19580 73468
rect 19580 73412 19636 73468
rect 19636 73412 19640 73468
rect 19576 73408 19640 73412
rect 19656 73468 19720 73472
rect 19656 73412 19660 73468
rect 19660 73412 19716 73468
rect 19716 73412 19720 73468
rect 19656 73408 19720 73412
rect 19736 73468 19800 73472
rect 19736 73412 19740 73468
rect 19740 73412 19796 73468
rect 19796 73412 19800 73468
rect 19736 73408 19800 73412
rect 19816 73468 19880 73472
rect 19816 73412 19820 73468
rect 19820 73412 19876 73468
rect 19876 73412 19880 73468
rect 19816 73408 19880 73412
rect 28948 73204 29012 73268
rect 4216 72924 4280 72928
rect 4216 72868 4220 72924
rect 4220 72868 4276 72924
rect 4276 72868 4280 72924
rect 4216 72864 4280 72868
rect 4296 72924 4360 72928
rect 4296 72868 4300 72924
rect 4300 72868 4356 72924
rect 4356 72868 4360 72924
rect 4296 72864 4360 72868
rect 4376 72924 4440 72928
rect 4376 72868 4380 72924
rect 4380 72868 4436 72924
rect 4436 72868 4440 72924
rect 4376 72864 4440 72868
rect 4456 72924 4520 72928
rect 4456 72868 4460 72924
rect 4460 72868 4516 72924
rect 4516 72868 4520 72924
rect 4456 72864 4520 72868
rect 28948 72932 29012 72996
rect 34936 72924 35000 72928
rect 34936 72868 34940 72924
rect 34940 72868 34996 72924
rect 34996 72868 35000 72924
rect 34936 72864 35000 72868
rect 35016 72924 35080 72928
rect 35016 72868 35020 72924
rect 35020 72868 35076 72924
rect 35076 72868 35080 72924
rect 35016 72864 35080 72868
rect 35096 72924 35160 72928
rect 35096 72868 35100 72924
rect 35100 72868 35156 72924
rect 35156 72868 35160 72924
rect 35096 72864 35160 72868
rect 35176 72924 35240 72928
rect 35176 72868 35180 72924
rect 35180 72868 35236 72924
rect 35236 72868 35240 72924
rect 35176 72864 35240 72868
rect 19576 72380 19640 72384
rect 19576 72324 19580 72380
rect 19580 72324 19636 72380
rect 19636 72324 19640 72380
rect 19576 72320 19640 72324
rect 19656 72380 19720 72384
rect 19656 72324 19660 72380
rect 19660 72324 19716 72380
rect 19716 72324 19720 72380
rect 19656 72320 19720 72324
rect 19736 72380 19800 72384
rect 19736 72324 19740 72380
rect 19740 72324 19796 72380
rect 19796 72324 19800 72380
rect 19736 72320 19800 72324
rect 19816 72380 19880 72384
rect 19816 72324 19820 72380
rect 19820 72324 19876 72380
rect 19876 72324 19880 72380
rect 19816 72320 19880 72324
rect 21036 71904 21100 71908
rect 21036 71848 21086 71904
rect 21086 71848 21100 71904
rect 21036 71844 21100 71848
rect 4216 71836 4280 71840
rect 4216 71780 4220 71836
rect 4220 71780 4276 71836
rect 4276 71780 4280 71836
rect 4216 71776 4280 71780
rect 4296 71836 4360 71840
rect 4296 71780 4300 71836
rect 4300 71780 4356 71836
rect 4356 71780 4360 71836
rect 4296 71776 4360 71780
rect 4376 71836 4440 71840
rect 4376 71780 4380 71836
rect 4380 71780 4436 71836
rect 4436 71780 4440 71836
rect 4376 71776 4440 71780
rect 4456 71836 4520 71840
rect 4456 71780 4460 71836
rect 4460 71780 4516 71836
rect 4516 71780 4520 71836
rect 4456 71776 4520 71780
rect 34936 71836 35000 71840
rect 34936 71780 34940 71836
rect 34940 71780 34996 71836
rect 34996 71780 35000 71836
rect 34936 71776 35000 71780
rect 35016 71836 35080 71840
rect 35016 71780 35020 71836
rect 35020 71780 35076 71836
rect 35076 71780 35080 71836
rect 35016 71776 35080 71780
rect 35096 71836 35160 71840
rect 35096 71780 35100 71836
rect 35100 71780 35156 71836
rect 35156 71780 35160 71836
rect 35096 71776 35160 71780
rect 35176 71836 35240 71840
rect 35176 71780 35180 71836
rect 35180 71780 35236 71836
rect 35236 71780 35240 71836
rect 35176 71776 35240 71780
rect 19576 71292 19640 71296
rect 19576 71236 19580 71292
rect 19580 71236 19636 71292
rect 19636 71236 19640 71292
rect 19576 71232 19640 71236
rect 19656 71292 19720 71296
rect 19656 71236 19660 71292
rect 19660 71236 19716 71292
rect 19716 71236 19720 71292
rect 19656 71232 19720 71236
rect 19736 71292 19800 71296
rect 19736 71236 19740 71292
rect 19740 71236 19796 71292
rect 19796 71236 19800 71292
rect 19736 71232 19800 71236
rect 19816 71292 19880 71296
rect 19816 71236 19820 71292
rect 19820 71236 19876 71292
rect 19876 71236 19880 71292
rect 19816 71232 19880 71236
rect 4216 70748 4280 70752
rect 4216 70692 4220 70748
rect 4220 70692 4276 70748
rect 4276 70692 4280 70748
rect 4216 70688 4280 70692
rect 4296 70748 4360 70752
rect 4296 70692 4300 70748
rect 4300 70692 4356 70748
rect 4356 70692 4360 70748
rect 4296 70688 4360 70692
rect 4376 70748 4440 70752
rect 4376 70692 4380 70748
rect 4380 70692 4436 70748
rect 4436 70692 4440 70748
rect 4376 70688 4440 70692
rect 4456 70748 4520 70752
rect 4456 70692 4460 70748
rect 4460 70692 4516 70748
rect 4516 70692 4520 70748
rect 4456 70688 4520 70692
rect 34936 70748 35000 70752
rect 34936 70692 34940 70748
rect 34940 70692 34996 70748
rect 34996 70692 35000 70748
rect 34936 70688 35000 70692
rect 35016 70748 35080 70752
rect 35016 70692 35020 70748
rect 35020 70692 35076 70748
rect 35076 70692 35080 70748
rect 35016 70688 35080 70692
rect 35096 70748 35160 70752
rect 35096 70692 35100 70748
rect 35100 70692 35156 70748
rect 35156 70692 35160 70748
rect 35096 70688 35160 70692
rect 35176 70748 35240 70752
rect 35176 70692 35180 70748
rect 35180 70692 35236 70748
rect 35236 70692 35240 70748
rect 35176 70688 35240 70692
rect 19576 70204 19640 70208
rect 19576 70148 19580 70204
rect 19580 70148 19636 70204
rect 19636 70148 19640 70204
rect 19576 70144 19640 70148
rect 19656 70204 19720 70208
rect 19656 70148 19660 70204
rect 19660 70148 19716 70204
rect 19716 70148 19720 70204
rect 19656 70144 19720 70148
rect 19736 70204 19800 70208
rect 19736 70148 19740 70204
rect 19740 70148 19796 70204
rect 19796 70148 19800 70204
rect 19736 70144 19800 70148
rect 19816 70204 19880 70208
rect 19816 70148 19820 70204
rect 19820 70148 19876 70204
rect 19876 70148 19880 70204
rect 19816 70144 19880 70148
rect 4216 69660 4280 69664
rect 4216 69604 4220 69660
rect 4220 69604 4276 69660
rect 4276 69604 4280 69660
rect 4216 69600 4280 69604
rect 4296 69660 4360 69664
rect 4296 69604 4300 69660
rect 4300 69604 4356 69660
rect 4356 69604 4360 69660
rect 4296 69600 4360 69604
rect 4376 69660 4440 69664
rect 4376 69604 4380 69660
rect 4380 69604 4436 69660
rect 4436 69604 4440 69660
rect 4376 69600 4440 69604
rect 4456 69660 4520 69664
rect 4456 69604 4460 69660
rect 4460 69604 4516 69660
rect 4516 69604 4520 69660
rect 4456 69600 4520 69604
rect 34936 69660 35000 69664
rect 34936 69604 34940 69660
rect 34940 69604 34996 69660
rect 34996 69604 35000 69660
rect 34936 69600 35000 69604
rect 35016 69660 35080 69664
rect 35016 69604 35020 69660
rect 35020 69604 35076 69660
rect 35076 69604 35080 69660
rect 35016 69600 35080 69604
rect 35096 69660 35160 69664
rect 35096 69604 35100 69660
rect 35100 69604 35156 69660
rect 35156 69604 35160 69660
rect 35096 69600 35160 69604
rect 35176 69660 35240 69664
rect 35176 69604 35180 69660
rect 35180 69604 35236 69660
rect 35236 69604 35240 69660
rect 35176 69600 35240 69604
rect 19576 69116 19640 69120
rect 19576 69060 19580 69116
rect 19580 69060 19636 69116
rect 19636 69060 19640 69116
rect 19576 69056 19640 69060
rect 19656 69116 19720 69120
rect 19656 69060 19660 69116
rect 19660 69060 19716 69116
rect 19716 69060 19720 69116
rect 19656 69056 19720 69060
rect 19736 69116 19800 69120
rect 19736 69060 19740 69116
rect 19740 69060 19796 69116
rect 19796 69060 19800 69116
rect 19736 69056 19800 69060
rect 19816 69116 19880 69120
rect 19816 69060 19820 69116
rect 19820 69060 19876 69116
rect 19876 69060 19880 69116
rect 19816 69056 19880 69060
rect 30052 68988 30116 69052
rect 4216 68572 4280 68576
rect 4216 68516 4220 68572
rect 4220 68516 4276 68572
rect 4276 68516 4280 68572
rect 4216 68512 4280 68516
rect 4296 68572 4360 68576
rect 4296 68516 4300 68572
rect 4300 68516 4356 68572
rect 4356 68516 4360 68572
rect 4296 68512 4360 68516
rect 4376 68572 4440 68576
rect 4376 68516 4380 68572
rect 4380 68516 4436 68572
rect 4436 68516 4440 68572
rect 4376 68512 4440 68516
rect 4456 68572 4520 68576
rect 4456 68516 4460 68572
rect 4460 68516 4516 68572
rect 4516 68516 4520 68572
rect 4456 68512 4520 68516
rect 34936 68572 35000 68576
rect 34936 68516 34940 68572
rect 34940 68516 34996 68572
rect 34996 68516 35000 68572
rect 34936 68512 35000 68516
rect 35016 68572 35080 68576
rect 35016 68516 35020 68572
rect 35020 68516 35076 68572
rect 35076 68516 35080 68572
rect 35016 68512 35080 68516
rect 35096 68572 35160 68576
rect 35096 68516 35100 68572
rect 35100 68516 35156 68572
rect 35156 68516 35160 68572
rect 35096 68512 35160 68516
rect 35176 68572 35240 68576
rect 35176 68516 35180 68572
rect 35180 68516 35236 68572
rect 35236 68516 35240 68572
rect 35176 68512 35240 68516
rect 28948 68308 29012 68372
rect 19576 68028 19640 68032
rect 19576 67972 19580 68028
rect 19580 67972 19636 68028
rect 19636 67972 19640 68028
rect 19576 67968 19640 67972
rect 19656 68028 19720 68032
rect 19656 67972 19660 68028
rect 19660 67972 19716 68028
rect 19716 67972 19720 68028
rect 19656 67968 19720 67972
rect 19736 68028 19800 68032
rect 19736 67972 19740 68028
rect 19740 67972 19796 68028
rect 19796 67972 19800 68028
rect 19736 67968 19800 67972
rect 19816 68028 19880 68032
rect 19816 67972 19820 68028
rect 19820 67972 19876 68028
rect 19876 67972 19880 68028
rect 19816 67968 19880 67972
rect 28948 67900 29012 67964
rect 4216 67484 4280 67488
rect 4216 67428 4220 67484
rect 4220 67428 4276 67484
rect 4276 67428 4280 67484
rect 4216 67424 4280 67428
rect 4296 67484 4360 67488
rect 4296 67428 4300 67484
rect 4300 67428 4356 67484
rect 4356 67428 4360 67484
rect 4296 67424 4360 67428
rect 4376 67484 4440 67488
rect 4376 67428 4380 67484
rect 4380 67428 4436 67484
rect 4436 67428 4440 67484
rect 4376 67424 4440 67428
rect 4456 67484 4520 67488
rect 4456 67428 4460 67484
rect 4460 67428 4516 67484
rect 4516 67428 4520 67484
rect 4456 67424 4520 67428
rect 34936 67484 35000 67488
rect 34936 67428 34940 67484
rect 34940 67428 34996 67484
rect 34996 67428 35000 67484
rect 34936 67424 35000 67428
rect 35016 67484 35080 67488
rect 35016 67428 35020 67484
rect 35020 67428 35076 67484
rect 35076 67428 35080 67484
rect 35016 67424 35080 67428
rect 35096 67484 35160 67488
rect 35096 67428 35100 67484
rect 35100 67428 35156 67484
rect 35156 67428 35160 67484
rect 35096 67424 35160 67428
rect 35176 67484 35240 67488
rect 35176 67428 35180 67484
rect 35180 67428 35236 67484
rect 35236 67428 35240 67484
rect 35176 67424 35240 67428
rect 28396 67084 28460 67148
rect 19576 66940 19640 66944
rect 19576 66884 19580 66940
rect 19580 66884 19636 66940
rect 19636 66884 19640 66940
rect 19576 66880 19640 66884
rect 19656 66940 19720 66944
rect 19656 66884 19660 66940
rect 19660 66884 19716 66940
rect 19716 66884 19720 66940
rect 19656 66880 19720 66884
rect 19736 66940 19800 66944
rect 19736 66884 19740 66940
rect 19740 66884 19796 66940
rect 19796 66884 19800 66940
rect 19736 66880 19800 66884
rect 19816 66940 19880 66944
rect 19816 66884 19820 66940
rect 19820 66884 19876 66940
rect 19876 66884 19880 66940
rect 19816 66880 19880 66884
rect 4216 66396 4280 66400
rect 4216 66340 4220 66396
rect 4220 66340 4276 66396
rect 4276 66340 4280 66396
rect 4216 66336 4280 66340
rect 4296 66396 4360 66400
rect 4296 66340 4300 66396
rect 4300 66340 4356 66396
rect 4356 66340 4360 66396
rect 4296 66336 4360 66340
rect 4376 66396 4440 66400
rect 4376 66340 4380 66396
rect 4380 66340 4436 66396
rect 4436 66340 4440 66396
rect 4376 66336 4440 66340
rect 4456 66396 4520 66400
rect 4456 66340 4460 66396
rect 4460 66340 4516 66396
rect 4516 66340 4520 66396
rect 4456 66336 4520 66340
rect 34936 66396 35000 66400
rect 34936 66340 34940 66396
rect 34940 66340 34996 66396
rect 34996 66340 35000 66396
rect 34936 66336 35000 66340
rect 35016 66396 35080 66400
rect 35016 66340 35020 66396
rect 35020 66340 35076 66396
rect 35076 66340 35080 66396
rect 35016 66336 35080 66340
rect 35096 66396 35160 66400
rect 35096 66340 35100 66396
rect 35100 66340 35156 66396
rect 35156 66340 35160 66396
rect 35096 66336 35160 66340
rect 35176 66396 35240 66400
rect 35176 66340 35180 66396
rect 35180 66340 35236 66396
rect 35236 66340 35240 66396
rect 35176 66336 35240 66340
rect 19576 65852 19640 65856
rect 19576 65796 19580 65852
rect 19580 65796 19636 65852
rect 19636 65796 19640 65852
rect 19576 65792 19640 65796
rect 19656 65852 19720 65856
rect 19656 65796 19660 65852
rect 19660 65796 19716 65852
rect 19716 65796 19720 65852
rect 19656 65792 19720 65796
rect 19736 65852 19800 65856
rect 19736 65796 19740 65852
rect 19740 65796 19796 65852
rect 19796 65796 19800 65852
rect 19736 65792 19800 65796
rect 19816 65852 19880 65856
rect 19816 65796 19820 65852
rect 19820 65796 19876 65852
rect 19876 65796 19880 65852
rect 19816 65792 19880 65796
rect 4216 65308 4280 65312
rect 4216 65252 4220 65308
rect 4220 65252 4276 65308
rect 4276 65252 4280 65308
rect 4216 65248 4280 65252
rect 4296 65308 4360 65312
rect 4296 65252 4300 65308
rect 4300 65252 4356 65308
rect 4356 65252 4360 65308
rect 4296 65248 4360 65252
rect 4376 65308 4440 65312
rect 4376 65252 4380 65308
rect 4380 65252 4436 65308
rect 4436 65252 4440 65308
rect 4376 65248 4440 65252
rect 4456 65308 4520 65312
rect 4456 65252 4460 65308
rect 4460 65252 4516 65308
rect 4516 65252 4520 65308
rect 4456 65248 4520 65252
rect 34936 65308 35000 65312
rect 34936 65252 34940 65308
rect 34940 65252 34996 65308
rect 34996 65252 35000 65308
rect 34936 65248 35000 65252
rect 35016 65308 35080 65312
rect 35016 65252 35020 65308
rect 35020 65252 35076 65308
rect 35076 65252 35080 65308
rect 35016 65248 35080 65252
rect 35096 65308 35160 65312
rect 35096 65252 35100 65308
rect 35100 65252 35156 65308
rect 35156 65252 35160 65308
rect 35096 65248 35160 65252
rect 35176 65308 35240 65312
rect 35176 65252 35180 65308
rect 35180 65252 35236 65308
rect 35236 65252 35240 65308
rect 35176 65248 35240 65252
rect 19576 64764 19640 64768
rect 19576 64708 19580 64764
rect 19580 64708 19636 64764
rect 19636 64708 19640 64764
rect 19576 64704 19640 64708
rect 19656 64764 19720 64768
rect 19656 64708 19660 64764
rect 19660 64708 19716 64764
rect 19716 64708 19720 64764
rect 19656 64704 19720 64708
rect 19736 64764 19800 64768
rect 19736 64708 19740 64764
rect 19740 64708 19796 64764
rect 19796 64708 19800 64764
rect 19736 64704 19800 64708
rect 19816 64764 19880 64768
rect 19816 64708 19820 64764
rect 19820 64708 19876 64764
rect 19876 64708 19880 64764
rect 19816 64704 19880 64708
rect 4216 64220 4280 64224
rect 4216 64164 4220 64220
rect 4220 64164 4276 64220
rect 4276 64164 4280 64220
rect 4216 64160 4280 64164
rect 4296 64220 4360 64224
rect 4296 64164 4300 64220
rect 4300 64164 4356 64220
rect 4356 64164 4360 64220
rect 4296 64160 4360 64164
rect 4376 64220 4440 64224
rect 4376 64164 4380 64220
rect 4380 64164 4436 64220
rect 4436 64164 4440 64220
rect 4376 64160 4440 64164
rect 4456 64220 4520 64224
rect 4456 64164 4460 64220
rect 4460 64164 4516 64220
rect 4516 64164 4520 64220
rect 4456 64160 4520 64164
rect 34936 64220 35000 64224
rect 34936 64164 34940 64220
rect 34940 64164 34996 64220
rect 34996 64164 35000 64220
rect 34936 64160 35000 64164
rect 35016 64220 35080 64224
rect 35016 64164 35020 64220
rect 35020 64164 35076 64220
rect 35076 64164 35080 64220
rect 35016 64160 35080 64164
rect 35096 64220 35160 64224
rect 35096 64164 35100 64220
rect 35100 64164 35156 64220
rect 35156 64164 35160 64220
rect 35096 64160 35160 64164
rect 35176 64220 35240 64224
rect 35176 64164 35180 64220
rect 35180 64164 35236 64220
rect 35236 64164 35240 64220
rect 35176 64160 35240 64164
rect 19576 63676 19640 63680
rect 19576 63620 19580 63676
rect 19580 63620 19636 63676
rect 19636 63620 19640 63676
rect 19576 63616 19640 63620
rect 19656 63676 19720 63680
rect 19656 63620 19660 63676
rect 19660 63620 19716 63676
rect 19716 63620 19720 63676
rect 19656 63616 19720 63620
rect 19736 63676 19800 63680
rect 19736 63620 19740 63676
rect 19740 63620 19796 63676
rect 19796 63620 19800 63676
rect 19736 63616 19800 63620
rect 19816 63676 19880 63680
rect 19816 63620 19820 63676
rect 19820 63620 19876 63676
rect 19876 63620 19880 63676
rect 19816 63616 19880 63620
rect 4216 63132 4280 63136
rect 4216 63076 4220 63132
rect 4220 63076 4276 63132
rect 4276 63076 4280 63132
rect 4216 63072 4280 63076
rect 4296 63132 4360 63136
rect 4296 63076 4300 63132
rect 4300 63076 4356 63132
rect 4356 63076 4360 63132
rect 4296 63072 4360 63076
rect 4376 63132 4440 63136
rect 4376 63076 4380 63132
rect 4380 63076 4436 63132
rect 4436 63076 4440 63132
rect 4376 63072 4440 63076
rect 4456 63132 4520 63136
rect 4456 63076 4460 63132
rect 4460 63076 4516 63132
rect 4516 63076 4520 63132
rect 4456 63072 4520 63076
rect 34936 63132 35000 63136
rect 34936 63076 34940 63132
rect 34940 63076 34996 63132
rect 34996 63076 35000 63132
rect 34936 63072 35000 63076
rect 35016 63132 35080 63136
rect 35016 63076 35020 63132
rect 35020 63076 35076 63132
rect 35076 63076 35080 63132
rect 35016 63072 35080 63076
rect 35096 63132 35160 63136
rect 35096 63076 35100 63132
rect 35100 63076 35156 63132
rect 35156 63076 35160 63132
rect 35096 63072 35160 63076
rect 35176 63132 35240 63136
rect 35176 63076 35180 63132
rect 35180 63076 35236 63132
rect 35236 63076 35240 63132
rect 35176 63072 35240 63076
rect 22508 62732 22572 62796
rect 19576 62588 19640 62592
rect 19576 62532 19580 62588
rect 19580 62532 19636 62588
rect 19636 62532 19640 62588
rect 19576 62528 19640 62532
rect 19656 62588 19720 62592
rect 19656 62532 19660 62588
rect 19660 62532 19716 62588
rect 19716 62532 19720 62588
rect 19656 62528 19720 62532
rect 19736 62588 19800 62592
rect 19736 62532 19740 62588
rect 19740 62532 19796 62588
rect 19796 62532 19800 62588
rect 19736 62528 19800 62532
rect 19816 62588 19880 62592
rect 19816 62532 19820 62588
rect 19820 62532 19876 62588
rect 19876 62532 19880 62588
rect 19816 62528 19880 62532
rect 28028 62188 28092 62252
rect 4216 62044 4280 62048
rect 4216 61988 4220 62044
rect 4220 61988 4276 62044
rect 4276 61988 4280 62044
rect 4216 61984 4280 61988
rect 4296 62044 4360 62048
rect 4296 61988 4300 62044
rect 4300 61988 4356 62044
rect 4356 61988 4360 62044
rect 4296 61984 4360 61988
rect 4376 62044 4440 62048
rect 4376 61988 4380 62044
rect 4380 61988 4436 62044
rect 4436 61988 4440 62044
rect 4376 61984 4440 61988
rect 4456 62044 4520 62048
rect 4456 61988 4460 62044
rect 4460 61988 4516 62044
rect 4516 61988 4520 62044
rect 4456 61984 4520 61988
rect 34936 62044 35000 62048
rect 34936 61988 34940 62044
rect 34940 61988 34996 62044
rect 34996 61988 35000 62044
rect 34936 61984 35000 61988
rect 35016 62044 35080 62048
rect 35016 61988 35020 62044
rect 35020 61988 35076 62044
rect 35076 61988 35080 62044
rect 35016 61984 35080 61988
rect 35096 62044 35160 62048
rect 35096 61988 35100 62044
rect 35100 61988 35156 62044
rect 35156 61988 35160 62044
rect 35096 61984 35160 61988
rect 35176 62044 35240 62048
rect 35176 61988 35180 62044
rect 35180 61988 35236 62044
rect 35236 61988 35240 62044
rect 35176 61984 35240 61988
rect 19576 61500 19640 61504
rect 19576 61444 19580 61500
rect 19580 61444 19636 61500
rect 19636 61444 19640 61500
rect 19576 61440 19640 61444
rect 19656 61500 19720 61504
rect 19656 61444 19660 61500
rect 19660 61444 19716 61500
rect 19716 61444 19720 61500
rect 19656 61440 19720 61444
rect 19736 61500 19800 61504
rect 19736 61444 19740 61500
rect 19740 61444 19796 61500
rect 19796 61444 19800 61500
rect 19736 61440 19800 61444
rect 19816 61500 19880 61504
rect 19816 61444 19820 61500
rect 19820 61444 19876 61500
rect 19876 61444 19880 61500
rect 19816 61440 19880 61444
rect 4216 60956 4280 60960
rect 4216 60900 4220 60956
rect 4220 60900 4276 60956
rect 4276 60900 4280 60956
rect 4216 60896 4280 60900
rect 4296 60956 4360 60960
rect 4296 60900 4300 60956
rect 4300 60900 4356 60956
rect 4356 60900 4360 60956
rect 4296 60896 4360 60900
rect 4376 60956 4440 60960
rect 4376 60900 4380 60956
rect 4380 60900 4436 60956
rect 4436 60900 4440 60956
rect 4376 60896 4440 60900
rect 4456 60956 4520 60960
rect 4456 60900 4460 60956
rect 4460 60900 4516 60956
rect 4516 60900 4520 60956
rect 4456 60896 4520 60900
rect 34936 60956 35000 60960
rect 34936 60900 34940 60956
rect 34940 60900 34996 60956
rect 34996 60900 35000 60956
rect 34936 60896 35000 60900
rect 35016 60956 35080 60960
rect 35016 60900 35020 60956
rect 35020 60900 35076 60956
rect 35076 60900 35080 60956
rect 35016 60896 35080 60900
rect 35096 60956 35160 60960
rect 35096 60900 35100 60956
rect 35100 60900 35156 60956
rect 35156 60900 35160 60956
rect 35096 60896 35160 60900
rect 35176 60956 35240 60960
rect 35176 60900 35180 60956
rect 35180 60900 35236 60956
rect 35236 60900 35240 60956
rect 35176 60896 35240 60900
rect 19576 60412 19640 60416
rect 19576 60356 19580 60412
rect 19580 60356 19636 60412
rect 19636 60356 19640 60412
rect 19576 60352 19640 60356
rect 19656 60412 19720 60416
rect 19656 60356 19660 60412
rect 19660 60356 19716 60412
rect 19716 60356 19720 60412
rect 19656 60352 19720 60356
rect 19736 60412 19800 60416
rect 19736 60356 19740 60412
rect 19740 60356 19796 60412
rect 19796 60356 19800 60412
rect 19736 60352 19800 60356
rect 19816 60412 19880 60416
rect 19816 60356 19820 60412
rect 19820 60356 19876 60412
rect 19876 60356 19880 60412
rect 19816 60352 19880 60356
rect 4216 59868 4280 59872
rect 4216 59812 4220 59868
rect 4220 59812 4276 59868
rect 4276 59812 4280 59868
rect 4216 59808 4280 59812
rect 4296 59868 4360 59872
rect 4296 59812 4300 59868
rect 4300 59812 4356 59868
rect 4356 59812 4360 59868
rect 4296 59808 4360 59812
rect 4376 59868 4440 59872
rect 4376 59812 4380 59868
rect 4380 59812 4436 59868
rect 4436 59812 4440 59868
rect 4376 59808 4440 59812
rect 4456 59868 4520 59872
rect 4456 59812 4460 59868
rect 4460 59812 4516 59868
rect 4516 59812 4520 59868
rect 4456 59808 4520 59812
rect 34936 59868 35000 59872
rect 34936 59812 34940 59868
rect 34940 59812 34996 59868
rect 34996 59812 35000 59868
rect 34936 59808 35000 59812
rect 35016 59868 35080 59872
rect 35016 59812 35020 59868
rect 35020 59812 35076 59868
rect 35076 59812 35080 59868
rect 35016 59808 35080 59812
rect 35096 59868 35160 59872
rect 35096 59812 35100 59868
rect 35100 59812 35156 59868
rect 35156 59812 35160 59868
rect 35096 59808 35160 59812
rect 35176 59868 35240 59872
rect 35176 59812 35180 59868
rect 35180 59812 35236 59868
rect 35236 59812 35240 59868
rect 35176 59808 35240 59812
rect 19576 59324 19640 59328
rect 19576 59268 19580 59324
rect 19580 59268 19636 59324
rect 19636 59268 19640 59324
rect 19576 59264 19640 59268
rect 19656 59324 19720 59328
rect 19656 59268 19660 59324
rect 19660 59268 19716 59324
rect 19716 59268 19720 59324
rect 19656 59264 19720 59268
rect 19736 59324 19800 59328
rect 19736 59268 19740 59324
rect 19740 59268 19796 59324
rect 19796 59268 19800 59324
rect 19736 59264 19800 59268
rect 19816 59324 19880 59328
rect 19816 59268 19820 59324
rect 19820 59268 19876 59324
rect 19876 59268 19880 59324
rect 19816 59264 19880 59268
rect 4216 58780 4280 58784
rect 4216 58724 4220 58780
rect 4220 58724 4276 58780
rect 4276 58724 4280 58780
rect 4216 58720 4280 58724
rect 4296 58780 4360 58784
rect 4296 58724 4300 58780
rect 4300 58724 4356 58780
rect 4356 58724 4360 58780
rect 4296 58720 4360 58724
rect 4376 58780 4440 58784
rect 4376 58724 4380 58780
rect 4380 58724 4436 58780
rect 4436 58724 4440 58780
rect 4376 58720 4440 58724
rect 4456 58780 4520 58784
rect 4456 58724 4460 58780
rect 4460 58724 4516 58780
rect 4516 58724 4520 58780
rect 4456 58720 4520 58724
rect 34936 58780 35000 58784
rect 34936 58724 34940 58780
rect 34940 58724 34996 58780
rect 34996 58724 35000 58780
rect 34936 58720 35000 58724
rect 35016 58780 35080 58784
rect 35016 58724 35020 58780
rect 35020 58724 35076 58780
rect 35076 58724 35080 58780
rect 35016 58720 35080 58724
rect 35096 58780 35160 58784
rect 35096 58724 35100 58780
rect 35100 58724 35156 58780
rect 35156 58724 35160 58780
rect 35096 58720 35160 58724
rect 35176 58780 35240 58784
rect 35176 58724 35180 58780
rect 35180 58724 35236 58780
rect 35236 58724 35240 58780
rect 35176 58720 35240 58724
rect 19576 58236 19640 58240
rect 19576 58180 19580 58236
rect 19580 58180 19636 58236
rect 19636 58180 19640 58236
rect 19576 58176 19640 58180
rect 19656 58236 19720 58240
rect 19656 58180 19660 58236
rect 19660 58180 19716 58236
rect 19716 58180 19720 58236
rect 19656 58176 19720 58180
rect 19736 58236 19800 58240
rect 19736 58180 19740 58236
rect 19740 58180 19796 58236
rect 19796 58180 19800 58236
rect 19736 58176 19800 58180
rect 19816 58236 19880 58240
rect 19816 58180 19820 58236
rect 19820 58180 19876 58236
rect 19876 58180 19880 58236
rect 19816 58176 19880 58180
rect 4216 57692 4280 57696
rect 4216 57636 4220 57692
rect 4220 57636 4276 57692
rect 4276 57636 4280 57692
rect 4216 57632 4280 57636
rect 4296 57692 4360 57696
rect 4296 57636 4300 57692
rect 4300 57636 4356 57692
rect 4356 57636 4360 57692
rect 4296 57632 4360 57636
rect 4376 57692 4440 57696
rect 4376 57636 4380 57692
rect 4380 57636 4436 57692
rect 4436 57636 4440 57692
rect 4376 57632 4440 57636
rect 4456 57692 4520 57696
rect 4456 57636 4460 57692
rect 4460 57636 4516 57692
rect 4516 57636 4520 57692
rect 4456 57632 4520 57636
rect 34936 57692 35000 57696
rect 34936 57636 34940 57692
rect 34940 57636 34996 57692
rect 34996 57636 35000 57692
rect 34936 57632 35000 57636
rect 35016 57692 35080 57696
rect 35016 57636 35020 57692
rect 35020 57636 35076 57692
rect 35076 57636 35080 57692
rect 35016 57632 35080 57636
rect 35096 57692 35160 57696
rect 35096 57636 35100 57692
rect 35100 57636 35156 57692
rect 35156 57636 35160 57692
rect 35096 57632 35160 57636
rect 35176 57692 35240 57696
rect 35176 57636 35180 57692
rect 35180 57636 35236 57692
rect 35236 57636 35240 57692
rect 35176 57632 35240 57636
rect 19576 57148 19640 57152
rect 19576 57092 19580 57148
rect 19580 57092 19636 57148
rect 19636 57092 19640 57148
rect 19576 57088 19640 57092
rect 19656 57148 19720 57152
rect 19656 57092 19660 57148
rect 19660 57092 19716 57148
rect 19716 57092 19720 57148
rect 19656 57088 19720 57092
rect 19736 57148 19800 57152
rect 19736 57092 19740 57148
rect 19740 57092 19796 57148
rect 19796 57092 19800 57148
rect 19736 57088 19800 57092
rect 19816 57148 19880 57152
rect 19816 57092 19820 57148
rect 19820 57092 19876 57148
rect 19876 57092 19880 57148
rect 19816 57088 19880 57092
rect 4216 56604 4280 56608
rect 4216 56548 4220 56604
rect 4220 56548 4276 56604
rect 4276 56548 4280 56604
rect 4216 56544 4280 56548
rect 4296 56604 4360 56608
rect 4296 56548 4300 56604
rect 4300 56548 4356 56604
rect 4356 56548 4360 56604
rect 4296 56544 4360 56548
rect 4376 56604 4440 56608
rect 4376 56548 4380 56604
rect 4380 56548 4436 56604
rect 4436 56548 4440 56604
rect 4376 56544 4440 56548
rect 4456 56604 4520 56608
rect 4456 56548 4460 56604
rect 4460 56548 4516 56604
rect 4516 56548 4520 56604
rect 4456 56544 4520 56548
rect 34936 56604 35000 56608
rect 34936 56548 34940 56604
rect 34940 56548 34996 56604
rect 34996 56548 35000 56604
rect 34936 56544 35000 56548
rect 35016 56604 35080 56608
rect 35016 56548 35020 56604
rect 35020 56548 35076 56604
rect 35076 56548 35080 56604
rect 35016 56544 35080 56548
rect 35096 56604 35160 56608
rect 35096 56548 35100 56604
rect 35100 56548 35156 56604
rect 35156 56548 35160 56604
rect 35096 56544 35160 56548
rect 35176 56604 35240 56608
rect 35176 56548 35180 56604
rect 35180 56548 35236 56604
rect 35236 56548 35240 56604
rect 35176 56544 35240 56548
rect 19576 56060 19640 56064
rect 19576 56004 19580 56060
rect 19580 56004 19636 56060
rect 19636 56004 19640 56060
rect 19576 56000 19640 56004
rect 19656 56060 19720 56064
rect 19656 56004 19660 56060
rect 19660 56004 19716 56060
rect 19716 56004 19720 56060
rect 19656 56000 19720 56004
rect 19736 56060 19800 56064
rect 19736 56004 19740 56060
rect 19740 56004 19796 56060
rect 19796 56004 19800 56060
rect 19736 56000 19800 56004
rect 19816 56060 19880 56064
rect 19816 56004 19820 56060
rect 19820 56004 19876 56060
rect 19876 56004 19880 56060
rect 19816 56000 19880 56004
rect 4216 55516 4280 55520
rect 4216 55460 4220 55516
rect 4220 55460 4276 55516
rect 4276 55460 4280 55516
rect 4216 55456 4280 55460
rect 4296 55516 4360 55520
rect 4296 55460 4300 55516
rect 4300 55460 4356 55516
rect 4356 55460 4360 55516
rect 4296 55456 4360 55460
rect 4376 55516 4440 55520
rect 4376 55460 4380 55516
rect 4380 55460 4436 55516
rect 4436 55460 4440 55516
rect 4376 55456 4440 55460
rect 4456 55516 4520 55520
rect 4456 55460 4460 55516
rect 4460 55460 4516 55516
rect 4516 55460 4520 55516
rect 4456 55456 4520 55460
rect 34936 55516 35000 55520
rect 34936 55460 34940 55516
rect 34940 55460 34996 55516
rect 34996 55460 35000 55516
rect 34936 55456 35000 55460
rect 35016 55516 35080 55520
rect 35016 55460 35020 55516
rect 35020 55460 35076 55516
rect 35076 55460 35080 55516
rect 35016 55456 35080 55460
rect 35096 55516 35160 55520
rect 35096 55460 35100 55516
rect 35100 55460 35156 55516
rect 35156 55460 35160 55516
rect 35096 55456 35160 55460
rect 35176 55516 35240 55520
rect 35176 55460 35180 55516
rect 35180 55460 35236 55516
rect 35236 55460 35240 55516
rect 35176 55456 35240 55460
rect 19576 54972 19640 54976
rect 19576 54916 19580 54972
rect 19580 54916 19636 54972
rect 19636 54916 19640 54972
rect 19576 54912 19640 54916
rect 19656 54972 19720 54976
rect 19656 54916 19660 54972
rect 19660 54916 19716 54972
rect 19716 54916 19720 54972
rect 19656 54912 19720 54916
rect 19736 54972 19800 54976
rect 19736 54916 19740 54972
rect 19740 54916 19796 54972
rect 19796 54916 19800 54972
rect 19736 54912 19800 54916
rect 19816 54972 19880 54976
rect 19816 54916 19820 54972
rect 19820 54916 19876 54972
rect 19876 54916 19880 54972
rect 19816 54912 19880 54916
rect 4216 54428 4280 54432
rect 4216 54372 4220 54428
rect 4220 54372 4276 54428
rect 4276 54372 4280 54428
rect 4216 54368 4280 54372
rect 4296 54428 4360 54432
rect 4296 54372 4300 54428
rect 4300 54372 4356 54428
rect 4356 54372 4360 54428
rect 4296 54368 4360 54372
rect 4376 54428 4440 54432
rect 4376 54372 4380 54428
rect 4380 54372 4436 54428
rect 4436 54372 4440 54428
rect 4376 54368 4440 54372
rect 4456 54428 4520 54432
rect 4456 54372 4460 54428
rect 4460 54372 4516 54428
rect 4516 54372 4520 54428
rect 4456 54368 4520 54372
rect 34936 54428 35000 54432
rect 34936 54372 34940 54428
rect 34940 54372 34996 54428
rect 34996 54372 35000 54428
rect 34936 54368 35000 54372
rect 35016 54428 35080 54432
rect 35016 54372 35020 54428
rect 35020 54372 35076 54428
rect 35076 54372 35080 54428
rect 35016 54368 35080 54372
rect 35096 54428 35160 54432
rect 35096 54372 35100 54428
rect 35100 54372 35156 54428
rect 35156 54372 35160 54428
rect 35096 54368 35160 54372
rect 35176 54428 35240 54432
rect 35176 54372 35180 54428
rect 35180 54372 35236 54428
rect 35236 54372 35240 54428
rect 35176 54368 35240 54372
rect 24716 54164 24780 54228
rect 21772 54028 21836 54092
rect 14780 53952 14844 53956
rect 14780 53896 14794 53952
rect 14794 53896 14844 53952
rect 14780 53892 14844 53896
rect 24532 53952 24596 53956
rect 24532 53896 24546 53952
rect 24546 53896 24596 53952
rect 24532 53892 24596 53896
rect 19576 53884 19640 53888
rect 19576 53828 19580 53884
rect 19580 53828 19636 53884
rect 19636 53828 19640 53884
rect 19576 53824 19640 53828
rect 19656 53884 19720 53888
rect 19656 53828 19660 53884
rect 19660 53828 19716 53884
rect 19716 53828 19720 53884
rect 19656 53824 19720 53828
rect 19736 53884 19800 53888
rect 19736 53828 19740 53884
rect 19740 53828 19796 53884
rect 19796 53828 19800 53884
rect 19736 53824 19800 53828
rect 19816 53884 19880 53888
rect 19816 53828 19820 53884
rect 19820 53828 19876 53884
rect 19876 53828 19880 53884
rect 19816 53824 19880 53828
rect 4216 53340 4280 53344
rect 4216 53284 4220 53340
rect 4220 53284 4276 53340
rect 4276 53284 4280 53340
rect 4216 53280 4280 53284
rect 4296 53340 4360 53344
rect 4296 53284 4300 53340
rect 4300 53284 4356 53340
rect 4356 53284 4360 53340
rect 4296 53280 4360 53284
rect 4376 53340 4440 53344
rect 4376 53284 4380 53340
rect 4380 53284 4436 53340
rect 4436 53284 4440 53340
rect 4376 53280 4440 53284
rect 4456 53340 4520 53344
rect 4456 53284 4460 53340
rect 4460 53284 4516 53340
rect 4516 53284 4520 53340
rect 4456 53280 4520 53284
rect 34936 53340 35000 53344
rect 34936 53284 34940 53340
rect 34940 53284 34996 53340
rect 34996 53284 35000 53340
rect 34936 53280 35000 53284
rect 35016 53340 35080 53344
rect 35016 53284 35020 53340
rect 35020 53284 35076 53340
rect 35076 53284 35080 53340
rect 35016 53280 35080 53284
rect 35096 53340 35160 53344
rect 35096 53284 35100 53340
rect 35100 53284 35156 53340
rect 35156 53284 35160 53340
rect 35096 53280 35160 53284
rect 35176 53340 35240 53344
rect 35176 53284 35180 53340
rect 35180 53284 35236 53340
rect 35236 53284 35240 53340
rect 35176 53280 35240 53284
rect 19576 52796 19640 52800
rect 19576 52740 19580 52796
rect 19580 52740 19636 52796
rect 19636 52740 19640 52796
rect 19576 52736 19640 52740
rect 19656 52796 19720 52800
rect 19656 52740 19660 52796
rect 19660 52740 19716 52796
rect 19716 52740 19720 52796
rect 19656 52736 19720 52740
rect 19736 52796 19800 52800
rect 19736 52740 19740 52796
rect 19740 52740 19796 52796
rect 19796 52740 19800 52796
rect 19736 52736 19800 52740
rect 19816 52796 19880 52800
rect 19816 52740 19820 52796
rect 19820 52740 19876 52796
rect 19876 52740 19880 52796
rect 19816 52736 19880 52740
rect 4216 52252 4280 52256
rect 4216 52196 4220 52252
rect 4220 52196 4276 52252
rect 4276 52196 4280 52252
rect 4216 52192 4280 52196
rect 4296 52252 4360 52256
rect 4296 52196 4300 52252
rect 4300 52196 4356 52252
rect 4356 52196 4360 52252
rect 4296 52192 4360 52196
rect 4376 52252 4440 52256
rect 4376 52196 4380 52252
rect 4380 52196 4436 52252
rect 4436 52196 4440 52252
rect 4376 52192 4440 52196
rect 4456 52252 4520 52256
rect 4456 52196 4460 52252
rect 4460 52196 4516 52252
rect 4516 52196 4520 52252
rect 4456 52192 4520 52196
rect 34936 52252 35000 52256
rect 34936 52196 34940 52252
rect 34940 52196 34996 52252
rect 34996 52196 35000 52252
rect 34936 52192 35000 52196
rect 35016 52252 35080 52256
rect 35016 52196 35020 52252
rect 35020 52196 35076 52252
rect 35076 52196 35080 52252
rect 35016 52192 35080 52196
rect 35096 52252 35160 52256
rect 35096 52196 35100 52252
rect 35100 52196 35156 52252
rect 35156 52196 35160 52252
rect 35096 52192 35160 52196
rect 35176 52252 35240 52256
rect 35176 52196 35180 52252
rect 35180 52196 35236 52252
rect 35236 52196 35240 52252
rect 35176 52192 35240 52196
rect 19576 51708 19640 51712
rect 19576 51652 19580 51708
rect 19580 51652 19636 51708
rect 19636 51652 19640 51708
rect 19576 51648 19640 51652
rect 19656 51708 19720 51712
rect 19656 51652 19660 51708
rect 19660 51652 19716 51708
rect 19716 51652 19720 51708
rect 19656 51648 19720 51652
rect 19736 51708 19800 51712
rect 19736 51652 19740 51708
rect 19740 51652 19796 51708
rect 19796 51652 19800 51708
rect 19736 51648 19800 51652
rect 19816 51708 19880 51712
rect 19816 51652 19820 51708
rect 19820 51652 19876 51708
rect 19876 51652 19880 51708
rect 19816 51648 19880 51652
rect 27844 51308 27908 51372
rect 28580 51172 28644 51236
rect 29132 51172 29196 51236
rect 4216 51164 4280 51168
rect 4216 51108 4220 51164
rect 4220 51108 4276 51164
rect 4276 51108 4280 51164
rect 4216 51104 4280 51108
rect 4296 51164 4360 51168
rect 4296 51108 4300 51164
rect 4300 51108 4356 51164
rect 4356 51108 4360 51164
rect 4296 51104 4360 51108
rect 4376 51164 4440 51168
rect 4376 51108 4380 51164
rect 4380 51108 4436 51164
rect 4436 51108 4440 51164
rect 4376 51104 4440 51108
rect 4456 51164 4520 51168
rect 4456 51108 4460 51164
rect 4460 51108 4516 51164
rect 4516 51108 4520 51164
rect 4456 51104 4520 51108
rect 34936 51164 35000 51168
rect 34936 51108 34940 51164
rect 34940 51108 34996 51164
rect 34996 51108 35000 51164
rect 34936 51104 35000 51108
rect 35016 51164 35080 51168
rect 35016 51108 35020 51164
rect 35020 51108 35076 51164
rect 35076 51108 35080 51164
rect 35016 51104 35080 51108
rect 35096 51164 35160 51168
rect 35096 51108 35100 51164
rect 35100 51108 35156 51164
rect 35156 51108 35160 51164
rect 35096 51104 35160 51108
rect 35176 51164 35240 51168
rect 35176 51108 35180 51164
rect 35180 51108 35236 51164
rect 35236 51108 35240 51164
rect 35176 51104 35240 51108
rect 21772 50824 21836 50828
rect 21772 50768 21822 50824
rect 21822 50768 21836 50824
rect 21772 50764 21836 50768
rect 19576 50620 19640 50624
rect 19576 50564 19580 50620
rect 19580 50564 19636 50620
rect 19636 50564 19640 50620
rect 19576 50560 19640 50564
rect 19656 50620 19720 50624
rect 19656 50564 19660 50620
rect 19660 50564 19716 50620
rect 19716 50564 19720 50620
rect 19656 50560 19720 50564
rect 19736 50620 19800 50624
rect 19736 50564 19740 50620
rect 19740 50564 19796 50620
rect 19796 50564 19800 50620
rect 19736 50560 19800 50564
rect 19816 50620 19880 50624
rect 19816 50564 19820 50620
rect 19820 50564 19876 50620
rect 19876 50564 19880 50620
rect 19816 50560 19880 50564
rect 4216 50076 4280 50080
rect 4216 50020 4220 50076
rect 4220 50020 4276 50076
rect 4276 50020 4280 50076
rect 4216 50016 4280 50020
rect 4296 50076 4360 50080
rect 4296 50020 4300 50076
rect 4300 50020 4356 50076
rect 4356 50020 4360 50076
rect 4296 50016 4360 50020
rect 4376 50076 4440 50080
rect 4376 50020 4380 50076
rect 4380 50020 4436 50076
rect 4436 50020 4440 50076
rect 4376 50016 4440 50020
rect 4456 50076 4520 50080
rect 4456 50020 4460 50076
rect 4460 50020 4516 50076
rect 4516 50020 4520 50076
rect 4456 50016 4520 50020
rect 34936 50076 35000 50080
rect 34936 50020 34940 50076
rect 34940 50020 34996 50076
rect 34996 50020 35000 50076
rect 34936 50016 35000 50020
rect 35016 50076 35080 50080
rect 35016 50020 35020 50076
rect 35020 50020 35076 50076
rect 35076 50020 35080 50076
rect 35016 50016 35080 50020
rect 35096 50076 35160 50080
rect 35096 50020 35100 50076
rect 35100 50020 35156 50076
rect 35156 50020 35160 50076
rect 35096 50016 35160 50020
rect 35176 50076 35240 50080
rect 35176 50020 35180 50076
rect 35180 50020 35236 50076
rect 35236 50020 35240 50076
rect 35176 50016 35240 50020
rect 21220 49676 21284 49740
rect 19576 49532 19640 49536
rect 19576 49476 19580 49532
rect 19580 49476 19636 49532
rect 19636 49476 19640 49532
rect 19576 49472 19640 49476
rect 19656 49532 19720 49536
rect 19656 49476 19660 49532
rect 19660 49476 19716 49532
rect 19716 49476 19720 49532
rect 19656 49472 19720 49476
rect 19736 49532 19800 49536
rect 19736 49476 19740 49532
rect 19740 49476 19796 49532
rect 19796 49476 19800 49532
rect 19736 49472 19800 49476
rect 19816 49532 19880 49536
rect 19816 49476 19820 49532
rect 19820 49476 19876 49532
rect 19876 49476 19880 49532
rect 19816 49472 19880 49476
rect 29132 49464 29196 49468
rect 29132 49408 29146 49464
rect 29146 49408 29196 49464
rect 29132 49404 29196 49408
rect 4216 48988 4280 48992
rect 4216 48932 4220 48988
rect 4220 48932 4276 48988
rect 4276 48932 4280 48988
rect 4216 48928 4280 48932
rect 4296 48988 4360 48992
rect 4296 48932 4300 48988
rect 4300 48932 4356 48988
rect 4356 48932 4360 48988
rect 4296 48928 4360 48932
rect 4376 48988 4440 48992
rect 4376 48932 4380 48988
rect 4380 48932 4436 48988
rect 4436 48932 4440 48988
rect 4376 48928 4440 48932
rect 4456 48988 4520 48992
rect 4456 48932 4460 48988
rect 4460 48932 4516 48988
rect 4516 48932 4520 48988
rect 4456 48928 4520 48932
rect 34936 48988 35000 48992
rect 34936 48932 34940 48988
rect 34940 48932 34996 48988
rect 34996 48932 35000 48988
rect 34936 48928 35000 48932
rect 35016 48988 35080 48992
rect 35016 48932 35020 48988
rect 35020 48932 35076 48988
rect 35076 48932 35080 48988
rect 35016 48928 35080 48932
rect 35096 48988 35160 48992
rect 35096 48932 35100 48988
rect 35100 48932 35156 48988
rect 35156 48932 35160 48988
rect 35096 48928 35160 48932
rect 35176 48988 35240 48992
rect 35176 48932 35180 48988
rect 35180 48932 35236 48988
rect 35236 48932 35240 48988
rect 35176 48928 35240 48932
rect 19576 48444 19640 48448
rect 19576 48388 19580 48444
rect 19580 48388 19636 48444
rect 19636 48388 19640 48444
rect 19576 48384 19640 48388
rect 19656 48444 19720 48448
rect 19656 48388 19660 48444
rect 19660 48388 19716 48444
rect 19716 48388 19720 48444
rect 19656 48384 19720 48388
rect 19736 48444 19800 48448
rect 19736 48388 19740 48444
rect 19740 48388 19796 48444
rect 19796 48388 19800 48444
rect 19736 48384 19800 48388
rect 19816 48444 19880 48448
rect 19816 48388 19820 48444
rect 19820 48388 19876 48444
rect 19876 48388 19880 48444
rect 19816 48384 19880 48388
rect 29684 48240 29748 48244
rect 29684 48184 29698 48240
rect 29698 48184 29748 48240
rect 29684 48180 29748 48184
rect 30052 48180 30116 48244
rect 4216 47900 4280 47904
rect 4216 47844 4220 47900
rect 4220 47844 4276 47900
rect 4276 47844 4280 47900
rect 4216 47840 4280 47844
rect 4296 47900 4360 47904
rect 4296 47844 4300 47900
rect 4300 47844 4356 47900
rect 4356 47844 4360 47900
rect 4296 47840 4360 47844
rect 4376 47900 4440 47904
rect 4376 47844 4380 47900
rect 4380 47844 4436 47900
rect 4436 47844 4440 47900
rect 4376 47840 4440 47844
rect 4456 47900 4520 47904
rect 4456 47844 4460 47900
rect 4460 47844 4516 47900
rect 4516 47844 4520 47900
rect 4456 47840 4520 47844
rect 34936 47900 35000 47904
rect 34936 47844 34940 47900
rect 34940 47844 34996 47900
rect 34996 47844 35000 47900
rect 34936 47840 35000 47844
rect 35016 47900 35080 47904
rect 35016 47844 35020 47900
rect 35020 47844 35076 47900
rect 35076 47844 35080 47900
rect 35016 47840 35080 47844
rect 35096 47900 35160 47904
rect 35096 47844 35100 47900
rect 35100 47844 35156 47900
rect 35156 47844 35160 47900
rect 35096 47840 35160 47844
rect 35176 47900 35240 47904
rect 35176 47844 35180 47900
rect 35180 47844 35236 47900
rect 35236 47844 35240 47900
rect 35176 47840 35240 47844
rect 19576 47356 19640 47360
rect 19576 47300 19580 47356
rect 19580 47300 19636 47356
rect 19636 47300 19640 47356
rect 19576 47296 19640 47300
rect 19656 47356 19720 47360
rect 19656 47300 19660 47356
rect 19660 47300 19716 47356
rect 19716 47300 19720 47356
rect 19656 47296 19720 47300
rect 19736 47356 19800 47360
rect 19736 47300 19740 47356
rect 19740 47300 19796 47356
rect 19796 47300 19800 47356
rect 19736 47296 19800 47300
rect 19816 47356 19880 47360
rect 19816 47300 19820 47356
rect 19820 47300 19876 47356
rect 19876 47300 19880 47356
rect 19816 47296 19880 47300
rect 20300 46956 20364 47020
rect 28212 46956 28276 47020
rect 4216 46812 4280 46816
rect 4216 46756 4220 46812
rect 4220 46756 4276 46812
rect 4276 46756 4280 46812
rect 4216 46752 4280 46756
rect 4296 46812 4360 46816
rect 4296 46756 4300 46812
rect 4300 46756 4356 46812
rect 4356 46756 4360 46812
rect 4296 46752 4360 46756
rect 4376 46812 4440 46816
rect 4376 46756 4380 46812
rect 4380 46756 4436 46812
rect 4436 46756 4440 46812
rect 4376 46752 4440 46756
rect 4456 46812 4520 46816
rect 4456 46756 4460 46812
rect 4460 46756 4516 46812
rect 4516 46756 4520 46812
rect 4456 46752 4520 46756
rect 34936 46812 35000 46816
rect 34936 46756 34940 46812
rect 34940 46756 34996 46812
rect 34996 46756 35000 46812
rect 34936 46752 35000 46756
rect 35016 46812 35080 46816
rect 35016 46756 35020 46812
rect 35020 46756 35076 46812
rect 35076 46756 35080 46812
rect 35016 46752 35080 46756
rect 35096 46812 35160 46816
rect 35096 46756 35100 46812
rect 35100 46756 35156 46812
rect 35156 46756 35160 46812
rect 35096 46752 35160 46756
rect 35176 46812 35240 46816
rect 35176 46756 35180 46812
rect 35180 46756 35236 46812
rect 35236 46756 35240 46812
rect 35176 46752 35240 46756
rect 20852 46412 20916 46476
rect 19576 46268 19640 46272
rect 19576 46212 19580 46268
rect 19580 46212 19636 46268
rect 19636 46212 19640 46268
rect 19576 46208 19640 46212
rect 19656 46268 19720 46272
rect 19656 46212 19660 46268
rect 19660 46212 19716 46268
rect 19716 46212 19720 46268
rect 19656 46208 19720 46212
rect 19736 46268 19800 46272
rect 19736 46212 19740 46268
rect 19740 46212 19796 46268
rect 19796 46212 19800 46268
rect 19736 46208 19800 46212
rect 19816 46268 19880 46272
rect 19816 46212 19820 46268
rect 19820 46212 19876 46268
rect 19876 46212 19880 46268
rect 19816 46208 19880 46212
rect 15700 46140 15764 46204
rect 28948 46140 29012 46204
rect 28948 45732 29012 45796
rect 4216 45724 4280 45728
rect 4216 45668 4220 45724
rect 4220 45668 4276 45724
rect 4276 45668 4280 45724
rect 4216 45664 4280 45668
rect 4296 45724 4360 45728
rect 4296 45668 4300 45724
rect 4300 45668 4356 45724
rect 4356 45668 4360 45724
rect 4296 45664 4360 45668
rect 4376 45724 4440 45728
rect 4376 45668 4380 45724
rect 4380 45668 4436 45724
rect 4436 45668 4440 45724
rect 4376 45664 4440 45668
rect 4456 45724 4520 45728
rect 4456 45668 4460 45724
rect 4460 45668 4516 45724
rect 4516 45668 4520 45724
rect 4456 45664 4520 45668
rect 34936 45724 35000 45728
rect 34936 45668 34940 45724
rect 34940 45668 34996 45724
rect 34996 45668 35000 45724
rect 34936 45664 35000 45668
rect 35016 45724 35080 45728
rect 35016 45668 35020 45724
rect 35020 45668 35076 45724
rect 35076 45668 35080 45724
rect 35016 45664 35080 45668
rect 35096 45724 35160 45728
rect 35096 45668 35100 45724
rect 35100 45668 35156 45724
rect 35156 45668 35160 45724
rect 35096 45664 35160 45668
rect 35176 45724 35240 45728
rect 35176 45668 35180 45724
rect 35180 45668 35236 45724
rect 35236 45668 35240 45724
rect 35176 45664 35240 45668
rect 19576 45180 19640 45184
rect 19576 45124 19580 45180
rect 19580 45124 19636 45180
rect 19636 45124 19640 45180
rect 19576 45120 19640 45124
rect 19656 45180 19720 45184
rect 19656 45124 19660 45180
rect 19660 45124 19716 45180
rect 19716 45124 19720 45180
rect 19656 45120 19720 45124
rect 19736 45180 19800 45184
rect 19736 45124 19740 45180
rect 19740 45124 19796 45180
rect 19796 45124 19800 45180
rect 19736 45120 19800 45124
rect 19816 45180 19880 45184
rect 19816 45124 19820 45180
rect 19820 45124 19876 45180
rect 19876 45124 19880 45180
rect 19816 45120 19880 45124
rect 4216 44636 4280 44640
rect 4216 44580 4220 44636
rect 4220 44580 4276 44636
rect 4276 44580 4280 44636
rect 4216 44576 4280 44580
rect 4296 44636 4360 44640
rect 4296 44580 4300 44636
rect 4300 44580 4356 44636
rect 4356 44580 4360 44636
rect 4296 44576 4360 44580
rect 4376 44636 4440 44640
rect 4376 44580 4380 44636
rect 4380 44580 4436 44636
rect 4436 44580 4440 44636
rect 4376 44576 4440 44580
rect 4456 44636 4520 44640
rect 4456 44580 4460 44636
rect 4460 44580 4516 44636
rect 4516 44580 4520 44636
rect 4456 44576 4520 44580
rect 34936 44636 35000 44640
rect 34936 44580 34940 44636
rect 34940 44580 34996 44636
rect 34996 44580 35000 44636
rect 34936 44576 35000 44580
rect 35016 44636 35080 44640
rect 35016 44580 35020 44636
rect 35020 44580 35076 44636
rect 35076 44580 35080 44636
rect 35016 44576 35080 44580
rect 35096 44636 35160 44640
rect 35096 44580 35100 44636
rect 35100 44580 35156 44636
rect 35156 44580 35160 44636
rect 35096 44576 35160 44580
rect 35176 44636 35240 44640
rect 35176 44580 35180 44636
rect 35180 44580 35236 44636
rect 35236 44580 35240 44636
rect 35176 44576 35240 44580
rect 19576 44092 19640 44096
rect 19576 44036 19580 44092
rect 19580 44036 19636 44092
rect 19636 44036 19640 44092
rect 19576 44032 19640 44036
rect 19656 44092 19720 44096
rect 19656 44036 19660 44092
rect 19660 44036 19716 44092
rect 19716 44036 19720 44092
rect 19656 44032 19720 44036
rect 19736 44092 19800 44096
rect 19736 44036 19740 44092
rect 19740 44036 19796 44092
rect 19796 44036 19800 44092
rect 19736 44032 19800 44036
rect 19816 44092 19880 44096
rect 19816 44036 19820 44092
rect 19820 44036 19876 44092
rect 19876 44036 19880 44092
rect 19816 44032 19880 44036
rect 28580 43828 28644 43892
rect 4216 43548 4280 43552
rect 4216 43492 4220 43548
rect 4220 43492 4276 43548
rect 4276 43492 4280 43548
rect 4216 43488 4280 43492
rect 4296 43548 4360 43552
rect 4296 43492 4300 43548
rect 4300 43492 4356 43548
rect 4356 43492 4360 43548
rect 4296 43488 4360 43492
rect 4376 43548 4440 43552
rect 4376 43492 4380 43548
rect 4380 43492 4436 43548
rect 4436 43492 4440 43548
rect 4376 43488 4440 43492
rect 4456 43548 4520 43552
rect 4456 43492 4460 43548
rect 4460 43492 4516 43548
rect 4516 43492 4520 43548
rect 4456 43488 4520 43492
rect 34936 43548 35000 43552
rect 34936 43492 34940 43548
rect 34940 43492 34996 43548
rect 34996 43492 35000 43548
rect 34936 43488 35000 43492
rect 35016 43548 35080 43552
rect 35016 43492 35020 43548
rect 35020 43492 35076 43548
rect 35076 43492 35080 43548
rect 35016 43488 35080 43492
rect 35096 43548 35160 43552
rect 35096 43492 35100 43548
rect 35100 43492 35156 43548
rect 35156 43492 35160 43548
rect 35096 43488 35160 43492
rect 35176 43548 35240 43552
rect 35176 43492 35180 43548
rect 35180 43492 35236 43548
rect 35236 43492 35240 43548
rect 35176 43488 35240 43492
rect 19576 43004 19640 43008
rect 19576 42948 19580 43004
rect 19580 42948 19636 43004
rect 19636 42948 19640 43004
rect 19576 42944 19640 42948
rect 19656 43004 19720 43008
rect 19656 42948 19660 43004
rect 19660 42948 19716 43004
rect 19716 42948 19720 43004
rect 19656 42944 19720 42948
rect 19736 43004 19800 43008
rect 19736 42948 19740 43004
rect 19740 42948 19796 43004
rect 19796 42948 19800 43004
rect 19736 42944 19800 42948
rect 19816 43004 19880 43008
rect 19816 42948 19820 43004
rect 19820 42948 19876 43004
rect 19876 42948 19880 43004
rect 19816 42944 19880 42948
rect 27844 42604 27908 42668
rect 4216 42460 4280 42464
rect 4216 42404 4220 42460
rect 4220 42404 4276 42460
rect 4276 42404 4280 42460
rect 4216 42400 4280 42404
rect 4296 42460 4360 42464
rect 4296 42404 4300 42460
rect 4300 42404 4356 42460
rect 4356 42404 4360 42460
rect 4296 42400 4360 42404
rect 4376 42460 4440 42464
rect 4376 42404 4380 42460
rect 4380 42404 4436 42460
rect 4436 42404 4440 42460
rect 4376 42400 4440 42404
rect 4456 42460 4520 42464
rect 4456 42404 4460 42460
rect 4460 42404 4516 42460
rect 4516 42404 4520 42460
rect 4456 42400 4520 42404
rect 34936 42460 35000 42464
rect 34936 42404 34940 42460
rect 34940 42404 34996 42460
rect 34996 42404 35000 42460
rect 34936 42400 35000 42404
rect 35016 42460 35080 42464
rect 35016 42404 35020 42460
rect 35020 42404 35076 42460
rect 35076 42404 35080 42460
rect 35016 42400 35080 42404
rect 35096 42460 35160 42464
rect 35096 42404 35100 42460
rect 35100 42404 35156 42460
rect 35156 42404 35160 42460
rect 35096 42400 35160 42404
rect 35176 42460 35240 42464
rect 35176 42404 35180 42460
rect 35180 42404 35236 42460
rect 35236 42404 35240 42460
rect 35176 42400 35240 42404
rect 19576 41916 19640 41920
rect 19576 41860 19580 41916
rect 19580 41860 19636 41916
rect 19636 41860 19640 41916
rect 19576 41856 19640 41860
rect 19656 41916 19720 41920
rect 19656 41860 19660 41916
rect 19660 41860 19716 41916
rect 19716 41860 19720 41916
rect 19656 41856 19720 41860
rect 19736 41916 19800 41920
rect 19736 41860 19740 41916
rect 19740 41860 19796 41916
rect 19796 41860 19800 41916
rect 19736 41856 19800 41860
rect 19816 41916 19880 41920
rect 19816 41860 19820 41916
rect 19820 41860 19876 41916
rect 19876 41860 19880 41916
rect 19816 41856 19880 41860
rect 14412 41848 14476 41852
rect 14412 41792 14426 41848
rect 14426 41792 14476 41848
rect 14412 41788 14476 41792
rect 28212 41848 28276 41852
rect 28212 41792 28262 41848
rect 28262 41792 28276 41848
rect 28212 41788 28276 41792
rect 4216 41372 4280 41376
rect 4216 41316 4220 41372
rect 4220 41316 4276 41372
rect 4276 41316 4280 41372
rect 4216 41312 4280 41316
rect 4296 41372 4360 41376
rect 4296 41316 4300 41372
rect 4300 41316 4356 41372
rect 4356 41316 4360 41372
rect 4296 41312 4360 41316
rect 4376 41372 4440 41376
rect 4376 41316 4380 41372
rect 4380 41316 4436 41372
rect 4436 41316 4440 41372
rect 4376 41312 4440 41316
rect 4456 41372 4520 41376
rect 4456 41316 4460 41372
rect 4460 41316 4516 41372
rect 4516 41316 4520 41372
rect 4456 41312 4520 41316
rect 34936 41372 35000 41376
rect 34936 41316 34940 41372
rect 34940 41316 34996 41372
rect 34996 41316 35000 41372
rect 34936 41312 35000 41316
rect 35016 41372 35080 41376
rect 35016 41316 35020 41372
rect 35020 41316 35076 41372
rect 35076 41316 35080 41372
rect 35016 41312 35080 41316
rect 35096 41372 35160 41376
rect 35096 41316 35100 41372
rect 35100 41316 35156 41372
rect 35156 41316 35160 41372
rect 35096 41312 35160 41316
rect 35176 41372 35240 41376
rect 35176 41316 35180 41372
rect 35180 41316 35236 41372
rect 35236 41316 35240 41372
rect 35176 41312 35240 41316
rect 29684 41244 29748 41308
rect 19576 40828 19640 40832
rect 19576 40772 19580 40828
rect 19580 40772 19636 40828
rect 19636 40772 19640 40828
rect 19576 40768 19640 40772
rect 19656 40828 19720 40832
rect 19656 40772 19660 40828
rect 19660 40772 19716 40828
rect 19716 40772 19720 40828
rect 19656 40768 19720 40772
rect 19736 40828 19800 40832
rect 19736 40772 19740 40828
rect 19740 40772 19796 40828
rect 19796 40772 19800 40828
rect 19736 40768 19800 40772
rect 19816 40828 19880 40832
rect 19816 40772 19820 40828
rect 19820 40772 19876 40828
rect 19876 40772 19880 40828
rect 19816 40768 19880 40772
rect 13676 40428 13740 40492
rect 4216 40284 4280 40288
rect 4216 40228 4220 40284
rect 4220 40228 4276 40284
rect 4276 40228 4280 40284
rect 4216 40224 4280 40228
rect 4296 40284 4360 40288
rect 4296 40228 4300 40284
rect 4300 40228 4356 40284
rect 4356 40228 4360 40284
rect 4296 40224 4360 40228
rect 4376 40284 4440 40288
rect 4376 40228 4380 40284
rect 4380 40228 4436 40284
rect 4436 40228 4440 40284
rect 4376 40224 4440 40228
rect 4456 40284 4520 40288
rect 4456 40228 4460 40284
rect 4460 40228 4516 40284
rect 4516 40228 4520 40284
rect 4456 40224 4520 40228
rect 34936 40284 35000 40288
rect 34936 40228 34940 40284
rect 34940 40228 34996 40284
rect 34996 40228 35000 40284
rect 34936 40224 35000 40228
rect 35016 40284 35080 40288
rect 35016 40228 35020 40284
rect 35020 40228 35076 40284
rect 35076 40228 35080 40284
rect 35016 40224 35080 40228
rect 35096 40284 35160 40288
rect 35096 40228 35100 40284
rect 35100 40228 35156 40284
rect 35156 40228 35160 40284
rect 35096 40224 35160 40228
rect 35176 40284 35240 40288
rect 35176 40228 35180 40284
rect 35180 40228 35236 40284
rect 35236 40228 35240 40284
rect 35176 40224 35240 40228
rect 19576 39740 19640 39744
rect 19576 39684 19580 39740
rect 19580 39684 19636 39740
rect 19636 39684 19640 39740
rect 19576 39680 19640 39684
rect 19656 39740 19720 39744
rect 19656 39684 19660 39740
rect 19660 39684 19716 39740
rect 19716 39684 19720 39740
rect 19656 39680 19720 39684
rect 19736 39740 19800 39744
rect 19736 39684 19740 39740
rect 19740 39684 19796 39740
rect 19796 39684 19800 39740
rect 19736 39680 19800 39684
rect 19816 39740 19880 39744
rect 19816 39684 19820 39740
rect 19820 39684 19876 39740
rect 19876 39684 19880 39740
rect 19816 39680 19880 39684
rect 4216 39196 4280 39200
rect 4216 39140 4220 39196
rect 4220 39140 4276 39196
rect 4276 39140 4280 39196
rect 4216 39136 4280 39140
rect 4296 39196 4360 39200
rect 4296 39140 4300 39196
rect 4300 39140 4356 39196
rect 4356 39140 4360 39196
rect 4296 39136 4360 39140
rect 4376 39196 4440 39200
rect 4376 39140 4380 39196
rect 4380 39140 4436 39196
rect 4436 39140 4440 39196
rect 4376 39136 4440 39140
rect 4456 39196 4520 39200
rect 4456 39140 4460 39196
rect 4460 39140 4516 39196
rect 4516 39140 4520 39196
rect 4456 39136 4520 39140
rect 34936 39196 35000 39200
rect 34936 39140 34940 39196
rect 34940 39140 34996 39196
rect 34996 39140 35000 39196
rect 34936 39136 35000 39140
rect 35016 39196 35080 39200
rect 35016 39140 35020 39196
rect 35020 39140 35076 39196
rect 35076 39140 35080 39196
rect 35016 39136 35080 39140
rect 35096 39196 35160 39200
rect 35096 39140 35100 39196
rect 35100 39140 35156 39196
rect 35156 39140 35160 39196
rect 35096 39136 35160 39140
rect 35176 39196 35240 39200
rect 35176 39140 35180 39196
rect 35180 39140 35236 39196
rect 35236 39140 35240 39196
rect 35176 39136 35240 39140
rect 15884 38660 15948 38724
rect 19576 38652 19640 38656
rect 19576 38596 19580 38652
rect 19580 38596 19636 38652
rect 19636 38596 19640 38652
rect 19576 38592 19640 38596
rect 19656 38652 19720 38656
rect 19656 38596 19660 38652
rect 19660 38596 19716 38652
rect 19716 38596 19720 38652
rect 19656 38592 19720 38596
rect 19736 38652 19800 38656
rect 19736 38596 19740 38652
rect 19740 38596 19796 38652
rect 19796 38596 19800 38652
rect 19736 38592 19800 38596
rect 19816 38652 19880 38656
rect 19816 38596 19820 38652
rect 19820 38596 19876 38652
rect 19876 38596 19880 38652
rect 19816 38592 19880 38596
rect 28028 38448 28092 38452
rect 28028 38392 28078 38448
rect 28078 38392 28092 38448
rect 28028 38388 28092 38392
rect 4216 38108 4280 38112
rect 4216 38052 4220 38108
rect 4220 38052 4276 38108
rect 4276 38052 4280 38108
rect 4216 38048 4280 38052
rect 4296 38108 4360 38112
rect 4296 38052 4300 38108
rect 4300 38052 4356 38108
rect 4356 38052 4360 38108
rect 4296 38048 4360 38052
rect 4376 38108 4440 38112
rect 4376 38052 4380 38108
rect 4380 38052 4436 38108
rect 4436 38052 4440 38108
rect 4376 38048 4440 38052
rect 4456 38108 4520 38112
rect 4456 38052 4460 38108
rect 4460 38052 4516 38108
rect 4516 38052 4520 38108
rect 4456 38048 4520 38052
rect 34936 38108 35000 38112
rect 34936 38052 34940 38108
rect 34940 38052 34996 38108
rect 34996 38052 35000 38108
rect 34936 38048 35000 38052
rect 35016 38108 35080 38112
rect 35016 38052 35020 38108
rect 35020 38052 35076 38108
rect 35076 38052 35080 38108
rect 35016 38048 35080 38052
rect 35096 38108 35160 38112
rect 35096 38052 35100 38108
rect 35100 38052 35156 38108
rect 35156 38052 35160 38108
rect 35096 38048 35160 38052
rect 35176 38108 35240 38112
rect 35176 38052 35180 38108
rect 35180 38052 35236 38108
rect 35236 38052 35240 38108
rect 35176 38048 35240 38052
rect 27844 37980 27908 38044
rect 17172 37708 17236 37772
rect 19576 37564 19640 37568
rect 19576 37508 19580 37564
rect 19580 37508 19636 37564
rect 19636 37508 19640 37564
rect 19576 37504 19640 37508
rect 19656 37564 19720 37568
rect 19656 37508 19660 37564
rect 19660 37508 19716 37564
rect 19716 37508 19720 37564
rect 19656 37504 19720 37508
rect 19736 37564 19800 37568
rect 19736 37508 19740 37564
rect 19740 37508 19796 37564
rect 19796 37508 19800 37564
rect 19736 37504 19800 37508
rect 19816 37564 19880 37568
rect 19816 37508 19820 37564
rect 19820 37508 19876 37564
rect 19876 37508 19880 37564
rect 19816 37504 19880 37508
rect 24348 37300 24412 37364
rect 4216 37020 4280 37024
rect 4216 36964 4220 37020
rect 4220 36964 4276 37020
rect 4276 36964 4280 37020
rect 4216 36960 4280 36964
rect 4296 37020 4360 37024
rect 4296 36964 4300 37020
rect 4300 36964 4356 37020
rect 4356 36964 4360 37020
rect 4296 36960 4360 36964
rect 4376 37020 4440 37024
rect 4376 36964 4380 37020
rect 4380 36964 4436 37020
rect 4436 36964 4440 37020
rect 4376 36960 4440 36964
rect 4456 37020 4520 37024
rect 4456 36964 4460 37020
rect 4460 36964 4516 37020
rect 4516 36964 4520 37020
rect 4456 36960 4520 36964
rect 34936 37020 35000 37024
rect 34936 36964 34940 37020
rect 34940 36964 34996 37020
rect 34996 36964 35000 37020
rect 34936 36960 35000 36964
rect 35016 37020 35080 37024
rect 35016 36964 35020 37020
rect 35020 36964 35076 37020
rect 35076 36964 35080 37020
rect 35016 36960 35080 36964
rect 35096 37020 35160 37024
rect 35096 36964 35100 37020
rect 35100 36964 35156 37020
rect 35156 36964 35160 37020
rect 35096 36960 35160 36964
rect 35176 37020 35240 37024
rect 35176 36964 35180 37020
rect 35180 36964 35236 37020
rect 35236 36964 35240 37020
rect 35176 36960 35240 36964
rect 19576 36476 19640 36480
rect 19576 36420 19580 36476
rect 19580 36420 19636 36476
rect 19636 36420 19640 36476
rect 19576 36416 19640 36420
rect 19656 36476 19720 36480
rect 19656 36420 19660 36476
rect 19660 36420 19716 36476
rect 19716 36420 19720 36476
rect 19656 36416 19720 36420
rect 19736 36476 19800 36480
rect 19736 36420 19740 36476
rect 19740 36420 19796 36476
rect 19796 36420 19800 36476
rect 19736 36416 19800 36420
rect 19816 36476 19880 36480
rect 19816 36420 19820 36476
rect 19820 36420 19876 36476
rect 19876 36420 19880 36476
rect 19816 36416 19880 36420
rect 23244 36212 23308 36276
rect 9628 36076 9692 36140
rect 4216 35932 4280 35936
rect 4216 35876 4220 35932
rect 4220 35876 4276 35932
rect 4276 35876 4280 35932
rect 4216 35872 4280 35876
rect 4296 35932 4360 35936
rect 4296 35876 4300 35932
rect 4300 35876 4356 35932
rect 4356 35876 4360 35932
rect 4296 35872 4360 35876
rect 4376 35932 4440 35936
rect 4376 35876 4380 35932
rect 4380 35876 4436 35932
rect 4436 35876 4440 35932
rect 4376 35872 4440 35876
rect 4456 35932 4520 35936
rect 4456 35876 4460 35932
rect 4460 35876 4516 35932
rect 4516 35876 4520 35932
rect 4456 35872 4520 35876
rect 34936 35932 35000 35936
rect 34936 35876 34940 35932
rect 34940 35876 34996 35932
rect 34996 35876 35000 35932
rect 34936 35872 35000 35876
rect 35016 35932 35080 35936
rect 35016 35876 35020 35932
rect 35020 35876 35076 35932
rect 35076 35876 35080 35932
rect 35016 35872 35080 35876
rect 35096 35932 35160 35936
rect 35096 35876 35100 35932
rect 35100 35876 35156 35932
rect 35156 35876 35160 35932
rect 35096 35872 35160 35876
rect 35176 35932 35240 35936
rect 35176 35876 35180 35932
rect 35180 35876 35236 35932
rect 35236 35876 35240 35932
rect 35176 35872 35240 35876
rect 19576 35388 19640 35392
rect 19576 35332 19580 35388
rect 19580 35332 19636 35388
rect 19636 35332 19640 35388
rect 19576 35328 19640 35332
rect 19656 35388 19720 35392
rect 19656 35332 19660 35388
rect 19660 35332 19716 35388
rect 19716 35332 19720 35388
rect 19656 35328 19720 35332
rect 19736 35388 19800 35392
rect 19736 35332 19740 35388
rect 19740 35332 19796 35388
rect 19796 35332 19800 35388
rect 19736 35328 19800 35332
rect 19816 35388 19880 35392
rect 19816 35332 19820 35388
rect 19820 35332 19876 35388
rect 19876 35332 19880 35388
rect 19816 35328 19880 35332
rect 14964 34988 15028 35052
rect 4216 34844 4280 34848
rect 4216 34788 4220 34844
rect 4220 34788 4276 34844
rect 4276 34788 4280 34844
rect 4216 34784 4280 34788
rect 4296 34844 4360 34848
rect 4296 34788 4300 34844
rect 4300 34788 4356 34844
rect 4356 34788 4360 34844
rect 4296 34784 4360 34788
rect 4376 34844 4440 34848
rect 4376 34788 4380 34844
rect 4380 34788 4436 34844
rect 4436 34788 4440 34844
rect 4376 34784 4440 34788
rect 4456 34844 4520 34848
rect 4456 34788 4460 34844
rect 4460 34788 4516 34844
rect 4516 34788 4520 34844
rect 4456 34784 4520 34788
rect 34936 34844 35000 34848
rect 34936 34788 34940 34844
rect 34940 34788 34996 34844
rect 34996 34788 35000 34844
rect 34936 34784 35000 34788
rect 35016 34844 35080 34848
rect 35016 34788 35020 34844
rect 35020 34788 35076 34844
rect 35076 34788 35080 34844
rect 35016 34784 35080 34788
rect 35096 34844 35160 34848
rect 35096 34788 35100 34844
rect 35100 34788 35156 34844
rect 35156 34788 35160 34844
rect 35096 34784 35160 34788
rect 35176 34844 35240 34848
rect 35176 34788 35180 34844
rect 35180 34788 35236 34844
rect 35236 34788 35240 34844
rect 35176 34784 35240 34788
rect 14228 34716 14292 34780
rect 13124 34580 13188 34644
rect 13860 34640 13924 34644
rect 13860 34584 13910 34640
rect 13910 34584 13924 34640
rect 13860 34580 13924 34584
rect 8340 34444 8404 34508
rect 14964 34308 15028 34372
rect 16804 34308 16868 34372
rect 20668 34308 20732 34372
rect 19576 34300 19640 34304
rect 19576 34244 19580 34300
rect 19580 34244 19636 34300
rect 19636 34244 19640 34300
rect 19576 34240 19640 34244
rect 19656 34300 19720 34304
rect 19656 34244 19660 34300
rect 19660 34244 19716 34300
rect 19716 34244 19720 34300
rect 19656 34240 19720 34244
rect 19736 34300 19800 34304
rect 19736 34244 19740 34300
rect 19740 34244 19796 34300
rect 19796 34244 19800 34300
rect 19736 34240 19800 34244
rect 19816 34300 19880 34304
rect 19816 34244 19820 34300
rect 19820 34244 19876 34300
rect 19876 34244 19880 34300
rect 19816 34240 19880 34244
rect 12572 34172 12636 34236
rect 20116 34172 20180 34236
rect 4216 33756 4280 33760
rect 4216 33700 4220 33756
rect 4220 33700 4276 33756
rect 4276 33700 4280 33756
rect 4216 33696 4280 33700
rect 4296 33756 4360 33760
rect 4296 33700 4300 33756
rect 4300 33700 4356 33756
rect 4356 33700 4360 33756
rect 4296 33696 4360 33700
rect 4376 33756 4440 33760
rect 4376 33700 4380 33756
rect 4380 33700 4436 33756
rect 4436 33700 4440 33756
rect 4376 33696 4440 33700
rect 4456 33756 4520 33760
rect 4456 33700 4460 33756
rect 4460 33700 4516 33756
rect 4516 33700 4520 33756
rect 4456 33696 4520 33700
rect 34936 33756 35000 33760
rect 34936 33700 34940 33756
rect 34940 33700 34996 33756
rect 34996 33700 35000 33756
rect 34936 33696 35000 33700
rect 35016 33756 35080 33760
rect 35016 33700 35020 33756
rect 35020 33700 35076 33756
rect 35076 33700 35080 33756
rect 35016 33696 35080 33700
rect 35096 33756 35160 33760
rect 35096 33700 35100 33756
rect 35100 33700 35156 33756
rect 35156 33700 35160 33756
rect 35096 33696 35160 33700
rect 35176 33756 35240 33760
rect 35176 33700 35180 33756
rect 35180 33700 35236 33756
rect 35236 33700 35240 33756
rect 35176 33696 35240 33700
rect 16068 33628 16132 33692
rect 19576 33212 19640 33216
rect 19576 33156 19580 33212
rect 19580 33156 19636 33212
rect 19636 33156 19640 33212
rect 19576 33152 19640 33156
rect 19656 33212 19720 33216
rect 19656 33156 19660 33212
rect 19660 33156 19716 33212
rect 19716 33156 19720 33212
rect 19656 33152 19720 33156
rect 19736 33212 19800 33216
rect 19736 33156 19740 33212
rect 19740 33156 19796 33212
rect 19796 33156 19800 33212
rect 19736 33152 19800 33156
rect 19816 33212 19880 33216
rect 19816 33156 19820 33212
rect 19820 33156 19876 33212
rect 19876 33156 19880 33212
rect 19816 33152 19880 33156
rect 13492 33084 13556 33148
rect 4216 32668 4280 32672
rect 4216 32612 4220 32668
rect 4220 32612 4276 32668
rect 4276 32612 4280 32668
rect 4216 32608 4280 32612
rect 4296 32668 4360 32672
rect 4296 32612 4300 32668
rect 4300 32612 4356 32668
rect 4356 32612 4360 32668
rect 4296 32608 4360 32612
rect 4376 32668 4440 32672
rect 4376 32612 4380 32668
rect 4380 32612 4436 32668
rect 4436 32612 4440 32668
rect 4376 32608 4440 32612
rect 4456 32668 4520 32672
rect 4456 32612 4460 32668
rect 4460 32612 4516 32668
rect 4516 32612 4520 32668
rect 4456 32608 4520 32612
rect 34936 32668 35000 32672
rect 34936 32612 34940 32668
rect 34940 32612 34996 32668
rect 34996 32612 35000 32668
rect 34936 32608 35000 32612
rect 35016 32668 35080 32672
rect 35016 32612 35020 32668
rect 35020 32612 35076 32668
rect 35076 32612 35080 32668
rect 35016 32608 35080 32612
rect 35096 32668 35160 32672
rect 35096 32612 35100 32668
rect 35100 32612 35156 32668
rect 35156 32612 35160 32668
rect 35096 32608 35160 32612
rect 35176 32668 35240 32672
rect 35176 32612 35180 32668
rect 35180 32612 35236 32668
rect 35236 32612 35240 32668
rect 35176 32608 35240 32612
rect 15332 32404 15396 32468
rect 23244 32268 23308 32332
rect 23796 32132 23860 32196
rect 19576 32124 19640 32128
rect 19576 32068 19580 32124
rect 19580 32068 19636 32124
rect 19636 32068 19640 32124
rect 19576 32064 19640 32068
rect 19656 32124 19720 32128
rect 19656 32068 19660 32124
rect 19660 32068 19716 32124
rect 19716 32068 19720 32124
rect 19656 32064 19720 32068
rect 19736 32124 19800 32128
rect 19736 32068 19740 32124
rect 19740 32068 19796 32124
rect 19796 32068 19800 32124
rect 19736 32064 19800 32068
rect 19816 32124 19880 32128
rect 19816 32068 19820 32124
rect 19820 32068 19876 32124
rect 19876 32068 19880 32124
rect 19816 32064 19880 32068
rect 14228 31648 14292 31652
rect 14228 31592 14278 31648
rect 14278 31592 14292 31648
rect 14228 31588 14292 31592
rect 14964 31588 15028 31652
rect 15332 31588 15396 31652
rect 16068 31648 16132 31652
rect 16068 31592 16082 31648
rect 16082 31592 16132 31648
rect 16068 31588 16132 31592
rect 4216 31580 4280 31584
rect 4216 31524 4220 31580
rect 4220 31524 4276 31580
rect 4276 31524 4280 31580
rect 4216 31520 4280 31524
rect 4296 31580 4360 31584
rect 4296 31524 4300 31580
rect 4300 31524 4356 31580
rect 4356 31524 4360 31580
rect 4296 31520 4360 31524
rect 4376 31580 4440 31584
rect 4376 31524 4380 31580
rect 4380 31524 4436 31580
rect 4436 31524 4440 31580
rect 4376 31520 4440 31524
rect 4456 31580 4520 31584
rect 4456 31524 4460 31580
rect 4460 31524 4516 31580
rect 4516 31524 4520 31580
rect 4456 31520 4520 31524
rect 23244 31588 23308 31652
rect 34936 31580 35000 31584
rect 34936 31524 34940 31580
rect 34940 31524 34996 31580
rect 34996 31524 35000 31580
rect 34936 31520 35000 31524
rect 35016 31580 35080 31584
rect 35016 31524 35020 31580
rect 35020 31524 35076 31580
rect 35076 31524 35080 31580
rect 35016 31520 35080 31524
rect 35096 31580 35160 31584
rect 35096 31524 35100 31580
rect 35100 31524 35156 31580
rect 35156 31524 35160 31580
rect 35096 31520 35160 31524
rect 35176 31580 35240 31584
rect 35176 31524 35180 31580
rect 35180 31524 35236 31580
rect 35236 31524 35240 31580
rect 35176 31520 35240 31524
rect 21588 31316 21652 31380
rect 19576 31036 19640 31040
rect 19576 30980 19580 31036
rect 19580 30980 19636 31036
rect 19636 30980 19640 31036
rect 19576 30976 19640 30980
rect 19656 31036 19720 31040
rect 19656 30980 19660 31036
rect 19660 30980 19716 31036
rect 19716 30980 19720 31036
rect 19656 30976 19720 30980
rect 19736 31036 19800 31040
rect 19736 30980 19740 31036
rect 19740 30980 19796 31036
rect 19796 30980 19800 31036
rect 19736 30976 19800 30980
rect 19816 31036 19880 31040
rect 19816 30980 19820 31036
rect 19820 30980 19876 31036
rect 19876 30980 19880 31036
rect 19816 30976 19880 30980
rect 12572 30968 12636 30972
rect 12572 30912 12586 30968
rect 12586 30912 12636 30968
rect 12572 30908 12636 30912
rect 13124 30636 13188 30700
rect 13492 30636 13556 30700
rect 4216 30492 4280 30496
rect 4216 30436 4220 30492
rect 4220 30436 4276 30492
rect 4276 30436 4280 30492
rect 4216 30432 4280 30436
rect 4296 30492 4360 30496
rect 4296 30436 4300 30492
rect 4300 30436 4356 30492
rect 4356 30436 4360 30492
rect 4296 30432 4360 30436
rect 4376 30492 4440 30496
rect 4376 30436 4380 30492
rect 4380 30436 4436 30492
rect 4436 30436 4440 30492
rect 4376 30432 4440 30436
rect 4456 30492 4520 30496
rect 4456 30436 4460 30492
rect 4460 30436 4516 30492
rect 4516 30436 4520 30492
rect 4456 30432 4520 30436
rect 21956 30364 22020 30428
rect 22140 30364 22204 30428
rect 34936 30492 35000 30496
rect 34936 30436 34940 30492
rect 34940 30436 34996 30492
rect 34996 30436 35000 30492
rect 34936 30432 35000 30436
rect 35016 30492 35080 30496
rect 35016 30436 35020 30492
rect 35020 30436 35076 30492
rect 35076 30436 35080 30492
rect 35016 30432 35080 30436
rect 35096 30492 35160 30496
rect 35096 30436 35100 30492
rect 35100 30436 35156 30492
rect 35156 30436 35160 30492
rect 35096 30432 35160 30436
rect 35176 30492 35240 30496
rect 35176 30436 35180 30492
rect 35180 30436 35236 30492
rect 35236 30436 35240 30492
rect 35176 30432 35240 30436
rect 12756 30228 12820 30292
rect 27844 30092 27908 30156
rect 22876 29956 22940 30020
rect 19576 29948 19640 29952
rect 19576 29892 19580 29948
rect 19580 29892 19636 29948
rect 19636 29892 19640 29948
rect 19576 29888 19640 29892
rect 19656 29948 19720 29952
rect 19656 29892 19660 29948
rect 19660 29892 19716 29948
rect 19716 29892 19720 29948
rect 19656 29888 19720 29892
rect 19736 29948 19800 29952
rect 19736 29892 19740 29948
rect 19740 29892 19796 29948
rect 19796 29892 19800 29948
rect 19736 29888 19800 29892
rect 19816 29948 19880 29952
rect 19816 29892 19820 29948
rect 19820 29892 19876 29948
rect 19876 29892 19880 29948
rect 19816 29888 19880 29892
rect 4216 29404 4280 29408
rect 4216 29348 4220 29404
rect 4220 29348 4276 29404
rect 4276 29348 4280 29404
rect 4216 29344 4280 29348
rect 4296 29404 4360 29408
rect 4296 29348 4300 29404
rect 4300 29348 4356 29404
rect 4356 29348 4360 29404
rect 4296 29344 4360 29348
rect 4376 29404 4440 29408
rect 4376 29348 4380 29404
rect 4380 29348 4436 29404
rect 4436 29348 4440 29404
rect 4376 29344 4440 29348
rect 4456 29404 4520 29408
rect 4456 29348 4460 29404
rect 4460 29348 4516 29404
rect 4516 29348 4520 29404
rect 4456 29344 4520 29348
rect 34936 29404 35000 29408
rect 34936 29348 34940 29404
rect 34940 29348 34996 29404
rect 34996 29348 35000 29404
rect 34936 29344 35000 29348
rect 35016 29404 35080 29408
rect 35016 29348 35020 29404
rect 35020 29348 35076 29404
rect 35076 29348 35080 29404
rect 35016 29344 35080 29348
rect 35096 29404 35160 29408
rect 35096 29348 35100 29404
rect 35100 29348 35156 29404
rect 35156 29348 35160 29404
rect 35096 29344 35160 29348
rect 35176 29404 35240 29408
rect 35176 29348 35180 29404
rect 35180 29348 35236 29404
rect 35236 29348 35240 29404
rect 35176 29344 35240 29348
rect 35572 29276 35636 29340
rect 8340 29200 8404 29204
rect 8340 29144 8390 29200
rect 8390 29144 8404 29200
rect 8340 29140 8404 29144
rect 14228 29140 14292 29204
rect 14596 29140 14660 29204
rect 16804 29140 16868 29204
rect 22324 29140 22388 29204
rect 19576 28860 19640 28864
rect 19576 28804 19580 28860
rect 19580 28804 19636 28860
rect 19636 28804 19640 28860
rect 19576 28800 19640 28804
rect 19656 28860 19720 28864
rect 19656 28804 19660 28860
rect 19660 28804 19716 28860
rect 19716 28804 19720 28860
rect 19656 28800 19720 28804
rect 19736 28860 19800 28864
rect 19736 28804 19740 28860
rect 19740 28804 19796 28860
rect 19796 28804 19800 28860
rect 19736 28800 19800 28804
rect 19816 28860 19880 28864
rect 19816 28804 19820 28860
rect 19820 28804 19876 28860
rect 19876 28804 19880 28860
rect 19816 28800 19880 28804
rect 22140 28732 22204 28796
rect 23796 28792 23860 28796
rect 23796 28736 23810 28792
rect 23810 28736 23860 28792
rect 23796 28732 23860 28736
rect 20116 28596 20180 28660
rect 16620 28460 16684 28524
rect 21772 28460 21836 28524
rect 4216 28316 4280 28320
rect 4216 28260 4220 28316
rect 4220 28260 4276 28316
rect 4276 28260 4280 28316
rect 4216 28256 4280 28260
rect 4296 28316 4360 28320
rect 4296 28260 4300 28316
rect 4300 28260 4356 28316
rect 4356 28260 4360 28316
rect 4296 28256 4360 28260
rect 4376 28316 4440 28320
rect 4376 28260 4380 28316
rect 4380 28260 4436 28316
rect 4436 28260 4440 28316
rect 4376 28256 4440 28260
rect 4456 28316 4520 28320
rect 4456 28260 4460 28316
rect 4460 28260 4516 28316
rect 4516 28260 4520 28316
rect 4456 28256 4520 28260
rect 14044 28188 14108 28252
rect 20484 28188 20548 28252
rect 21956 28188 22020 28252
rect 34936 28316 35000 28320
rect 34936 28260 34940 28316
rect 34940 28260 34996 28316
rect 34996 28260 35000 28316
rect 34936 28256 35000 28260
rect 35016 28316 35080 28320
rect 35016 28260 35020 28316
rect 35020 28260 35076 28316
rect 35076 28260 35080 28316
rect 35016 28256 35080 28260
rect 35096 28316 35160 28320
rect 35096 28260 35100 28316
rect 35100 28260 35156 28316
rect 35156 28260 35160 28316
rect 35096 28256 35160 28260
rect 35176 28316 35240 28320
rect 35176 28260 35180 28316
rect 35180 28260 35236 28316
rect 35236 28260 35240 28316
rect 35176 28256 35240 28260
rect 23980 28248 24044 28252
rect 23980 28192 23994 28248
rect 23994 28192 24044 28248
rect 23980 28188 24044 28192
rect 20668 27916 20732 27980
rect 21404 27840 21468 27844
rect 21404 27784 21454 27840
rect 21454 27784 21468 27840
rect 21404 27780 21468 27784
rect 19576 27772 19640 27776
rect 19576 27716 19580 27772
rect 19580 27716 19636 27772
rect 19636 27716 19640 27772
rect 19576 27712 19640 27716
rect 19656 27772 19720 27776
rect 19656 27716 19660 27772
rect 19660 27716 19716 27772
rect 19716 27716 19720 27772
rect 19656 27712 19720 27716
rect 19736 27772 19800 27776
rect 19736 27716 19740 27772
rect 19740 27716 19796 27772
rect 19796 27716 19800 27772
rect 19736 27712 19800 27716
rect 19816 27772 19880 27776
rect 19816 27716 19820 27772
rect 19820 27716 19876 27772
rect 19876 27716 19880 27772
rect 19816 27712 19880 27716
rect 22324 27508 22388 27572
rect 14044 27296 14108 27300
rect 14044 27240 14094 27296
rect 14094 27240 14108 27296
rect 14044 27236 14108 27240
rect 22140 27236 22204 27300
rect 4216 27228 4280 27232
rect 4216 27172 4220 27228
rect 4220 27172 4276 27228
rect 4276 27172 4280 27228
rect 4216 27168 4280 27172
rect 4296 27228 4360 27232
rect 4296 27172 4300 27228
rect 4300 27172 4356 27228
rect 4356 27172 4360 27228
rect 4296 27168 4360 27172
rect 4376 27228 4440 27232
rect 4376 27172 4380 27228
rect 4380 27172 4436 27228
rect 4436 27172 4440 27228
rect 4376 27168 4440 27172
rect 4456 27228 4520 27232
rect 4456 27172 4460 27228
rect 4460 27172 4516 27228
rect 4516 27172 4520 27228
rect 4456 27168 4520 27172
rect 34936 27228 35000 27232
rect 34936 27172 34940 27228
rect 34940 27172 34996 27228
rect 34996 27172 35000 27228
rect 34936 27168 35000 27172
rect 35016 27228 35080 27232
rect 35016 27172 35020 27228
rect 35020 27172 35076 27228
rect 35076 27172 35080 27228
rect 35016 27168 35080 27172
rect 35096 27228 35160 27232
rect 35096 27172 35100 27228
rect 35100 27172 35156 27228
rect 35156 27172 35160 27228
rect 35096 27168 35160 27172
rect 35176 27228 35240 27232
rect 35176 27172 35180 27228
rect 35180 27172 35236 27228
rect 35236 27172 35240 27228
rect 35176 27168 35240 27172
rect 17172 27100 17236 27164
rect 23244 27160 23308 27164
rect 23244 27104 23294 27160
rect 23294 27104 23308 27160
rect 23244 27100 23308 27104
rect 14228 26828 14292 26892
rect 14964 26828 15028 26892
rect 7236 26692 7300 26756
rect 19576 26684 19640 26688
rect 19576 26628 19580 26684
rect 19580 26628 19636 26684
rect 19636 26628 19640 26684
rect 19576 26624 19640 26628
rect 19656 26684 19720 26688
rect 19656 26628 19660 26684
rect 19660 26628 19716 26684
rect 19716 26628 19720 26684
rect 19656 26624 19720 26628
rect 19736 26684 19800 26688
rect 19736 26628 19740 26684
rect 19740 26628 19796 26684
rect 19796 26628 19800 26684
rect 19736 26624 19800 26628
rect 19816 26684 19880 26688
rect 19816 26628 19820 26684
rect 19820 26628 19876 26684
rect 19876 26628 19880 26684
rect 19816 26624 19880 26628
rect 34468 26556 34532 26620
rect 13308 26420 13372 26484
rect 6684 26284 6748 26348
rect 13124 26344 13188 26348
rect 13124 26288 13174 26344
rect 13174 26288 13188 26344
rect 13124 26284 13188 26288
rect 4216 26140 4280 26144
rect 4216 26084 4220 26140
rect 4220 26084 4276 26140
rect 4276 26084 4280 26140
rect 4216 26080 4280 26084
rect 4296 26140 4360 26144
rect 4296 26084 4300 26140
rect 4300 26084 4356 26140
rect 4356 26084 4360 26140
rect 4296 26080 4360 26084
rect 4376 26140 4440 26144
rect 4376 26084 4380 26140
rect 4380 26084 4436 26140
rect 4436 26084 4440 26140
rect 4376 26080 4440 26084
rect 4456 26140 4520 26144
rect 4456 26084 4460 26140
rect 4460 26084 4516 26140
rect 4516 26084 4520 26140
rect 4456 26080 4520 26084
rect 34936 26140 35000 26144
rect 34936 26084 34940 26140
rect 34940 26084 34996 26140
rect 34996 26084 35000 26140
rect 34936 26080 35000 26084
rect 35016 26140 35080 26144
rect 35016 26084 35020 26140
rect 35020 26084 35076 26140
rect 35076 26084 35080 26140
rect 35016 26080 35080 26084
rect 35096 26140 35160 26144
rect 35096 26084 35100 26140
rect 35100 26084 35156 26140
rect 35156 26084 35160 26140
rect 35096 26080 35160 26084
rect 35176 26140 35240 26144
rect 35176 26084 35180 26140
rect 35180 26084 35236 26140
rect 35236 26084 35240 26140
rect 35176 26080 35240 26084
rect 19576 25596 19640 25600
rect 19576 25540 19580 25596
rect 19580 25540 19636 25596
rect 19636 25540 19640 25596
rect 19576 25536 19640 25540
rect 19656 25596 19720 25600
rect 19656 25540 19660 25596
rect 19660 25540 19716 25596
rect 19716 25540 19720 25596
rect 19656 25536 19720 25540
rect 19736 25596 19800 25600
rect 19736 25540 19740 25596
rect 19740 25540 19796 25596
rect 19796 25540 19800 25596
rect 19736 25536 19800 25540
rect 19816 25596 19880 25600
rect 19816 25540 19820 25596
rect 19820 25540 19876 25596
rect 19876 25540 19880 25596
rect 19816 25536 19880 25540
rect 22876 25392 22940 25396
rect 22876 25336 22926 25392
rect 22926 25336 22940 25392
rect 22876 25332 22940 25336
rect 34468 25196 34532 25260
rect 14596 25120 14660 25124
rect 14596 25064 14646 25120
rect 14646 25064 14660 25120
rect 14596 25060 14660 25064
rect 4216 25052 4280 25056
rect 4216 24996 4220 25052
rect 4220 24996 4276 25052
rect 4276 24996 4280 25052
rect 4216 24992 4280 24996
rect 4296 25052 4360 25056
rect 4296 24996 4300 25052
rect 4300 24996 4356 25052
rect 4356 24996 4360 25052
rect 4296 24992 4360 24996
rect 4376 25052 4440 25056
rect 4376 24996 4380 25052
rect 4380 24996 4436 25052
rect 4436 24996 4440 25052
rect 4376 24992 4440 24996
rect 4456 25052 4520 25056
rect 4456 24996 4460 25052
rect 4460 24996 4516 25052
rect 4516 24996 4520 25052
rect 4456 24992 4520 24996
rect 13676 24788 13740 24852
rect 23244 25060 23308 25124
rect 34936 25052 35000 25056
rect 34936 24996 34940 25052
rect 34940 24996 34996 25052
rect 34996 24996 35000 25052
rect 34936 24992 35000 24996
rect 35016 25052 35080 25056
rect 35016 24996 35020 25052
rect 35020 24996 35076 25052
rect 35076 24996 35080 25052
rect 35016 24992 35080 24996
rect 35096 25052 35160 25056
rect 35096 24996 35100 25052
rect 35100 24996 35156 25052
rect 35156 24996 35160 25052
rect 35096 24992 35160 24996
rect 35176 25052 35240 25056
rect 35176 24996 35180 25052
rect 35180 24996 35236 25052
rect 35236 24996 35240 25052
rect 35176 24992 35240 24996
rect 21588 24516 21652 24580
rect 19576 24508 19640 24512
rect 19576 24452 19580 24508
rect 19580 24452 19636 24508
rect 19636 24452 19640 24508
rect 19576 24448 19640 24452
rect 19656 24508 19720 24512
rect 19656 24452 19660 24508
rect 19660 24452 19716 24508
rect 19716 24452 19720 24508
rect 19656 24448 19720 24452
rect 19736 24508 19800 24512
rect 19736 24452 19740 24508
rect 19740 24452 19796 24508
rect 19796 24452 19800 24508
rect 19736 24448 19800 24452
rect 19816 24508 19880 24512
rect 19816 24452 19820 24508
rect 19820 24452 19876 24508
rect 19876 24452 19880 24508
rect 19816 24448 19880 24452
rect 21404 24168 21468 24172
rect 21404 24112 21454 24168
rect 21454 24112 21468 24168
rect 21404 24108 21468 24112
rect 4216 23964 4280 23968
rect 4216 23908 4220 23964
rect 4220 23908 4276 23964
rect 4276 23908 4280 23964
rect 4216 23904 4280 23908
rect 4296 23964 4360 23968
rect 4296 23908 4300 23964
rect 4300 23908 4356 23964
rect 4356 23908 4360 23964
rect 4296 23904 4360 23908
rect 4376 23964 4440 23968
rect 4376 23908 4380 23964
rect 4380 23908 4436 23964
rect 4436 23908 4440 23964
rect 4376 23904 4440 23908
rect 4456 23964 4520 23968
rect 4456 23908 4460 23964
rect 4460 23908 4516 23964
rect 4516 23908 4520 23964
rect 4456 23904 4520 23908
rect 34936 23964 35000 23968
rect 34936 23908 34940 23964
rect 34940 23908 34996 23964
rect 34996 23908 35000 23964
rect 34936 23904 35000 23908
rect 35016 23964 35080 23968
rect 35016 23908 35020 23964
rect 35020 23908 35076 23964
rect 35076 23908 35080 23964
rect 35016 23904 35080 23908
rect 35096 23964 35160 23968
rect 35096 23908 35100 23964
rect 35100 23908 35156 23964
rect 35156 23908 35160 23964
rect 35096 23904 35160 23908
rect 35176 23964 35240 23968
rect 35176 23908 35180 23964
rect 35180 23908 35236 23964
rect 35236 23908 35240 23964
rect 35176 23904 35240 23908
rect 16620 23700 16684 23764
rect 14044 23564 14108 23628
rect 21956 23564 22020 23628
rect 19576 23420 19640 23424
rect 19576 23364 19580 23420
rect 19580 23364 19636 23420
rect 19636 23364 19640 23420
rect 19576 23360 19640 23364
rect 19656 23420 19720 23424
rect 19656 23364 19660 23420
rect 19660 23364 19716 23420
rect 19716 23364 19720 23420
rect 19656 23360 19720 23364
rect 19736 23420 19800 23424
rect 19736 23364 19740 23420
rect 19740 23364 19796 23420
rect 19796 23364 19800 23420
rect 19736 23360 19800 23364
rect 19816 23420 19880 23424
rect 19816 23364 19820 23420
rect 19820 23364 19876 23420
rect 19876 23364 19880 23420
rect 19816 23360 19880 23364
rect 23244 23156 23308 23220
rect 4216 22876 4280 22880
rect 4216 22820 4220 22876
rect 4220 22820 4276 22876
rect 4276 22820 4280 22876
rect 4216 22816 4280 22820
rect 4296 22876 4360 22880
rect 4296 22820 4300 22876
rect 4300 22820 4356 22876
rect 4356 22820 4360 22876
rect 4296 22816 4360 22820
rect 4376 22876 4440 22880
rect 4376 22820 4380 22876
rect 4380 22820 4436 22876
rect 4436 22820 4440 22876
rect 4376 22816 4440 22820
rect 4456 22876 4520 22880
rect 4456 22820 4460 22876
rect 4460 22820 4516 22876
rect 4516 22820 4520 22876
rect 4456 22816 4520 22820
rect 34936 22876 35000 22880
rect 34936 22820 34940 22876
rect 34940 22820 34996 22876
rect 34996 22820 35000 22876
rect 34936 22816 35000 22820
rect 35016 22876 35080 22880
rect 35016 22820 35020 22876
rect 35020 22820 35076 22876
rect 35076 22820 35080 22876
rect 35016 22816 35080 22820
rect 35096 22876 35160 22880
rect 35096 22820 35100 22876
rect 35100 22820 35156 22876
rect 35156 22820 35160 22876
rect 35096 22816 35160 22820
rect 35176 22876 35240 22880
rect 35176 22820 35180 22876
rect 35180 22820 35236 22876
rect 35236 22820 35240 22876
rect 35176 22816 35240 22820
rect 19576 22332 19640 22336
rect 19576 22276 19580 22332
rect 19580 22276 19636 22332
rect 19636 22276 19640 22332
rect 19576 22272 19640 22276
rect 19656 22332 19720 22336
rect 19656 22276 19660 22332
rect 19660 22276 19716 22332
rect 19716 22276 19720 22332
rect 19656 22272 19720 22276
rect 19736 22332 19800 22336
rect 19736 22276 19740 22332
rect 19740 22276 19796 22332
rect 19796 22276 19800 22332
rect 19736 22272 19800 22276
rect 19816 22332 19880 22336
rect 19816 22276 19820 22332
rect 19820 22276 19876 22332
rect 19876 22276 19880 22332
rect 19816 22272 19880 22276
rect 4216 21788 4280 21792
rect 4216 21732 4220 21788
rect 4220 21732 4276 21788
rect 4276 21732 4280 21788
rect 4216 21728 4280 21732
rect 4296 21788 4360 21792
rect 4296 21732 4300 21788
rect 4300 21732 4356 21788
rect 4356 21732 4360 21788
rect 4296 21728 4360 21732
rect 4376 21788 4440 21792
rect 4376 21732 4380 21788
rect 4380 21732 4436 21788
rect 4436 21732 4440 21788
rect 4376 21728 4440 21732
rect 4456 21788 4520 21792
rect 4456 21732 4460 21788
rect 4460 21732 4516 21788
rect 4516 21732 4520 21788
rect 4456 21728 4520 21732
rect 34936 21788 35000 21792
rect 34936 21732 34940 21788
rect 34940 21732 34996 21788
rect 34996 21732 35000 21788
rect 34936 21728 35000 21732
rect 35016 21788 35080 21792
rect 35016 21732 35020 21788
rect 35020 21732 35076 21788
rect 35076 21732 35080 21788
rect 35016 21728 35080 21732
rect 35096 21788 35160 21792
rect 35096 21732 35100 21788
rect 35100 21732 35156 21788
rect 35156 21732 35160 21788
rect 35096 21728 35160 21732
rect 35176 21788 35240 21792
rect 35176 21732 35180 21788
rect 35180 21732 35236 21788
rect 35236 21732 35240 21788
rect 35176 21728 35240 21732
rect 19576 21244 19640 21248
rect 19576 21188 19580 21244
rect 19580 21188 19636 21244
rect 19636 21188 19640 21244
rect 19576 21184 19640 21188
rect 19656 21244 19720 21248
rect 19656 21188 19660 21244
rect 19660 21188 19716 21244
rect 19716 21188 19720 21244
rect 19656 21184 19720 21188
rect 19736 21244 19800 21248
rect 19736 21188 19740 21244
rect 19740 21188 19796 21244
rect 19796 21188 19800 21244
rect 19736 21184 19800 21188
rect 19816 21244 19880 21248
rect 19816 21188 19820 21244
rect 19820 21188 19876 21244
rect 19876 21188 19880 21244
rect 19816 21184 19880 21188
rect 4216 20700 4280 20704
rect 4216 20644 4220 20700
rect 4220 20644 4276 20700
rect 4276 20644 4280 20700
rect 4216 20640 4280 20644
rect 4296 20700 4360 20704
rect 4296 20644 4300 20700
rect 4300 20644 4356 20700
rect 4356 20644 4360 20700
rect 4296 20640 4360 20644
rect 4376 20700 4440 20704
rect 4376 20644 4380 20700
rect 4380 20644 4436 20700
rect 4436 20644 4440 20700
rect 4376 20640 4440 20644
rect 4456 20700 4520 20704
rect 4456 20644 4460 20700
rect 4460 20644 4516 20700
rect 4516 20644 4520 20700
rect 4456 20640 4520 20644
rect 15884 20708 15948 20772
rect 34936 20700 35000 20704
rect 34936 20644 34940 20700
rect 34940 20644 34996 20700
rect 34996 20644 35000 20700
rect 34936 20640 35000 20644
rect 35016 20700 35080 20704
rect 35016 20644 35020 20700
rect 35020 20644 35076 20700
rect 35076 20644 35080 20700
rect 35016 20640 35080 20644
rect 35096 20700 35160 20704
rect 35096 20644 35100 20700
rect 35100 20644 35156 20700
rect 35156 20644 35160 20700
rect 35096 20640 35160 20644
rect 35176 20700 35240 20704
rect 35176 20644 35180 20700
rect 35180 20644 35236 20700
rect 35236 20644 35240 20700
rect 35176 20640 35240 20644
rect 19576 20156 19640 20160
rect 19576 20100 19580 20156
rect 19580 20100 19636 20156
rect 19636 20100 19640 20156
rect 19576 20096 19640 20100
rect 19656 20156 19720 20160
rect 19656 20100 19660 20156
rect 19660 20100 19716 20156
rect 19716 20100 19720 20156
rect 19656 20096 19720 20100
rect 19736 20156 19800 20160
rect 19736 20100 19740 20156
rect 19740 20100 19796 20156
rect 19796 20100 19800 20156
rect 19736 20096 19800 20100
rect 19816 20156 19880 20160
rect 19816 20100 19820 20156
rect 19820 20100 19876 20156
rect 19876 20100 19880 20156
rect 19816 20096 19880 20100
rect 24716 19892 24780 19956
rect 4216 19612 4280 19616
rect 4216 19556 4220 19612
rect 4220 19556 4276 19612
rect 4276 19556 4280 19612
rect 4216 19552 4280 19556
rect 4296 19612 4360 19616
rect 4296 19556 4300 19612
rect 4300 19556 4356 19612
rect 4356 19556 4360 19612
rect 4296 19552 4360 19556
rect 4376 19612 4440 19616
rect 4376 19556 4380 19612
rect 4380 19556 4436 19612
rect 4436 19556 4440 19612
rect 4376 19552 4440 19556
rect 4456 19612 4520 19616
rect 4456 19556 4460 19612
rect 4460 19556 4516 19612
rect 4516 19556 4520 19612
rect 4456 19552 4520 19556
rect 34936 19612 35000 19616
rect 34936 19556 34940 19612
rect 34940 19556 34996 19612
rect 34996 19556 35000 19612
rect 34936 19552 35000 19556
rect 35016 19612 35080 19616
rect 35016 19556 35020 19612
rect 35020 19556 35076 19612
rect 35076 19556 35080 19612
rect 35016 19552 35080 19556
rect 35096 19612 35160 19616
rect 35096 19556 35100 19612
rect 35100 19556 35156 19612
rect 35156 19556 35160 19612
rect 35096 19552 35160 19556
rect 35176 19612 35240 19616
rect 35176 19556 35180 19612
rect 35180 19556 35236 19612
rect 35236 19556 35240 19612
rect 35176 19552 35240 19556
rect 19576 19068 19640 19072
rect 19576 19012 19580 19068
rect 19580 19012 19636 19068
rect 19636 19012 19640 19068
rect 19576 19008 19640 19012
rect 19656 19068 19720 19072
rect 19656 19012 19660 19068
rect 19660 19012 19716 19068
rect 19716 19012 19720 19068
rect 19656 19008 19720 19012
rect 19736 19068 19800 19072
rect 19736 19012 19740 19068
rect 19740 19012 19796 19068
rect 19796 19012 19800 19068
rect 19736 19008 19800 19012
rect 19816 19068 19880 19072
rect 19816 19012 19820 19068
rect 19820 19012 19876 19068
rect 19876 19012 19880 19068
rect 19816 19008 19880 19012
rect 4216 18524 4280 18528
rect 4216 18468 4220 18524
rect 4220 18468 4276 18524
rect 4276 18468 4280 18524
rect 4216 18464 4280 18468
rect 4296 18524 4360 18528
rect 4296 18468 4300 18524
rect 4300 18468 4356 18524
rect 4356 18468 4360 18524
rect 4296 18464 4360 18468
rect 4376 18524 4440 18528
rect 4376 18468 4380 18524
rect 4380 18468 4436 18524
rect 4436 18468 4440 18524
rect 4376 18464 4440 18468
rect 4456 18524 4520 18528
rect 4456 18468 4460 18524
rect 4460 18468 4516 18524
rect 4516 18468 4520 18524
rect 4456 18464 4520 18468
rect 34936 18524 35000 18528
rect 34936 18468 34940 18524
rect 34940 18468 34996 18524
rect 34996 18468 35000 18524
rect 34936 18464 35000 18468
rect 35016 18524 35080 18528
rect 35016 18468 35020 18524
rect 35020 18468 35076 18524
rect 35076 18468 35080 18524
rect 35016 18464 35080 18468
rect 35096 18524 35160 18528
rect 35096 18468 35100 18524
rect 35100 18468 35156 18524
rect 35156 18468 35160 18524
rect 35096 18464 35160 18468
rect 35176 18524 35240 18528
rect 35176 18468 35180 18524
rect 35180 18468 35236 18524
rect 35236 18468 35240 18524
rect 35176 18464 35240 18468
rect 19576 17980 19640 17984
rect 19576 17924 19580 17980
rect 19580 17924 19636 17980
rect 19636 17924 19640 17980
rect 19576 17920 19640 17924
rect 19656 17980 19720 17984
rect 19656 17924 19660 17980
rect 19660 17924 19716 17980
rect 19716 17924 19720 17980
rect 19656 17920 19720 17924
rect 19736 17980 19800 17984
rect 19736 17924 19740 17980
rect 19740 17924 19796 17980
rect 19796 17924 19800 17980
rect 19736 17920 19800 17924
rect 19816 17980 19880 17984
rect 19816 17924 19820 17980
rect 19820 17924 19876 17980
rect 19876 17924 19880 17980
rect 19816 17920 19880 17924
rect 20484 17852 20548 17916
rect 21036 17852 21100 17916
rect 4216 17436 4280 17440
rect 4216 17380 4220 17436
rect 4220 17380 4276 17436
rect 4276 17380 4280 17436
rect 4216 17376 4280 17380
rect 4296 17436 4360 17440
rect 4296 17380 4300 17436
rect 4300 17380 4356 17436
rect 4356 17380 4360 17436
rect 4296 17376 4360 17380
rect 4376 17436 4440 17440
rect 4376 17380 4380 17436
rect 4380 17380 4436 17436
rect 4436 17380 4440 17436
rect 4376 17376 4440 17380
rect 4456 17436 4520 17440
rect 4456 17380 4460 17436
rect 4460 17380 4516 17436
rect 4516 17380 4520 17436
rect 4456 17376 4520 17380
rect 34936 17436 35000 17440
rect 34936 17380 34940 17436
rect 34940 17380 34996 17436
rect 34996 17380 35000 17436
rect 34936 17376 35000 17380
rect 35016 17436 35080 17440
rect 35016 17380 35020 17436
rect 35020 17380 35076 17436
rect 35076 17380 35080 17436
rect 35016 17376 35080 17380
rect 35096 17436 35160 17440
rect 35096 17380 35100 17436
rect 35100 17380 35156 17436
rect 35156 17380 35160 17436
rect 35096 17376 35160 17380
rect 35176 17436 35240 17440
rect 35176 17380 35180 17436
rect 35180 17380 35236 17436
rect 35236 17380 35240 17436
rect 35176 17376 35240 17380
rect 19576 16892 19640 16896
rect 19576 16836 19580 16892
rect 19580 16836 19636 16892
rect 19636 16836 19640 16892
rect 19576 16832 19640 16836
rect 19656 16892 19720 16896
rect 19656 16836 19660 16892
rect 19660 16836 19716 16892
rect 19716 16836 19720 16892
rect 19656 16832 19720 16836
rect 19736 16892 19800 16896
rect 19736 16836 19740 16892
rect 19740 16836 19796 16892
rect 19796 16836 19800 16892
rect 19736 16832 19800 16836
rect 19816 16892 19880 16896
rect 19816 16836 19820 16892
rect 19820 16836 19876 16892
rect 19876 16836 19880 16892
rect 19816 16832 19880 16836
rect 21220 16492 21284 16556
rect 4216 16348 4280 16352
rect 4216 16292 4220 16348
rect 4220 16292 4276 16348
rect 4276 16292 4280 16348
rect 4216 16288 4280 16292
rect 4296 16348 4360 16352
rect 4296 16292 4300 16348
rect 4300 16292 4356 16348
rect 4356 16292 4360 16348
rect 4296 16288 4360 16292
rect 4376 16348 4440 16352
rect 4376 16292 4380 16348
rect 4380 16292 4436 16348
rect 4436 16292 4440 16348
rect 4376 16288 4440 16292
rect 4456 16348 4520 16352
rect 4456 16292 4460 16348
rect 4460 16292 4516 16348
rect 4516 16292 4520 16348
rect 4456 16288 4520 16292
rect 34936 16348 35000 16352
rect 34936 16292 34940 16348
rect 34940 16292 34996 16348
rect 34996 16292 35000 16348
rect 34936 16288 35000 16292
rect 35016 16348 35080 16352
rect 35016 16292 35020 16348
rect 35020 16292 35076 16348
rect 35076 16292 35080 16348
rect 35016 16288 35080 16292
rect 35096 16348 35160 16352
rect 35096 16292 35100 16348
rect 35100 16292 35156 16348
rect 35156 16292 35160 16348
rect 35096 16288 35160 16292
rect 35176 16348 35240 16352
rect 35176 16292 35180 16348
rect 35180 16292 35236 16348
rect 35236 16292 35240 16348
rect 35176 16288 35240 16292
rect 19576 15804 19640 15808
rect 19576 15748 19580 15804
rect 19580 15748 19636 15804
rect 19636 15748 19640 15804
rect 19576 15744 19640 15748
rect 19656 15804 19720 15808
rect 19656 15748 19660 15804
rect 19660 15748 19716 15804
rect 19716 15748 19720 15804
rect 19656 15744 19720 15748
rect 19736 15804 19800 15808
rect 19736 15748 19740 15804
rect 19740 15748 19796 15804
rect 19796 15748 19800 15804
rect 19736 15744 19800 15748
rect 19816 15804 19880 15808
rect 19816 15748 19820 15804
rect 19820 15748 19876 15804
rect 19876 15748 19880 15804
rect 19816 15744 19880 15748
rect 20852 15540 20916 15604
rect 4216 15260 4280 15264
rect 4216 15204 4220 15260
rect 4220 15204 4276 15260
rect 4276 15204 4280 15260
rect 4216 15200 4280 15204
rect 4296 15260 4360 15264
rect 4296 15204 4300 15260
rect 4300 15204 4356 15260
rect 4356 15204 4360 15260
rect 4296 15200 4360 15204
rect 4376 15260 4440 15264
rect 4376 15204 4380 15260
rect 4380 15204 4436 15260
rect 4436 15204 4440 15260
rect 4376 15200 4440 15204
rect 4456 15260 4520 15264
rect 4456 15204 4460 15260
rect 4460 15204 4516 15260
rect 4516 15204 4520 15260
rect 4456 15200 4520 15204
rect 34936 15260 35000 15264
rect 34936 15204 34940 15260
rect 34940 15204 34996 15260
rect 34996 15204 35000 15260
rect 34936 15200 35000 15204
rect 35016 15260 35080 15264
rect 35016 15204 35020 15260
rect 35020 15204 35076 15260
rect 35076 15204 35080 15260
rect 35016 15200 35080 15204
rect 35096 15260 35160 15264
rect 35096 15204 35100 15260
rect 35100 15204 35156 15260
rect 35156 15204 35160 15260
rect 35096 15200 35160 15204
rect 35176 15260 35240 15264
rect 35176 15204 35180 15260
rect 35180 15204 35236 15260
rect 35236 15204 35240 15260
rect 35176 15200 35240 15204
rect 22508 15132 22572 15196
rect 24532 15132 24596 15196
rect 13860 15056 13924 15060
rect 13860 15000 13874 15056
rect 13874 15000 13924 15056
rect 13860 14996 13924 15000
rect 19576 14716 19640 14720
rect 19576 14660 19580 14716
rect 19580 14660 19636 14716
rect 19636 14660 19640 14716
rect 19576 14656 19640 14660
rect 19656 14716 19720 14720
rect 19656 14660 19660 14716
rect 19660 14660 19716 14716
rect 19716 14660 19720 14716
rect 19656 14656 19720 14660
rect 19736 14716 19800 14720
rect 19736 14660 19740 14716
rect 19740 14660 19796 14716
rect 19796 14660 19800 14716
rect 19736 14656 19800 14660
rect 19816 14716 19880 14720
rect 19816 14660 19820 14716
rect 19820 14660 19876 14716
rect 19876 14660 19880 14716
rect 19816 14656 19880 14660
rect 4216 14172 4280 14176
rect 4216 14116 4220 14172
rect 4220 14116 4276 14172
rect 4276 14116 4280 14172
rect 4216 14112 4280 14116
rect 4296 14172 4360 14176
rect 4296 14116 4300 14172
rect 4300 14116 4356 14172
rect 4356 14116 4360 14172
rect 4296 14112 4360 14116
rect 4376 14172 4440 14176
rect 4376 14116 4380 14172
rect 4380 14116 4436 14172
rect 4436 14116 4440 14172
rect 4376 14112 4440 14116
rect 4456 14172 4520 14176
rect 4456 14116 4460 14172
rect 4460 14116 4516 14172
rect 4516 14116 4520 14172
rect 4456 14112 4520 14116
rect 34936 14172 35000 14176
rect 34936 14116 34940 14172
rect 34940 14116 34996 14172
rect 34996 14116 35000 14172
rect 34936 14112 35000 14116
rect 35016 14172 35080 14176
rect 35016 14116 35020 14172
rect 35020 14116 35076 14172
rect 35076 14116 35080 14172
rect 35016 14112 35080 14116
rect 35096 14172 35160 14176
rect 35096 14116 35100 14172
rect 35100 14116 35156 14172
rect 35156 14116 35160 14172
rect 35096 14112 35160 14116
rect 35176 14172 35240 14176
rect 35176 14116 35180 14172
rect 35180 14116 35236 14172
rect 35236 14116 35240 14172
rect 35176 14112 35240 14116
rect 19576 13628 19640 13632
rect 19576 13572 19580 13628
rect 19580 13572 19636 13628
rect 19636 13572 19640 13628
rect 19576 13568 19640 13572
rect 19656 13628 19720 13632
rect 19656 13572 19660 13628
rect 19660 13572 19716 13628
rect 19716 13572 19720 13628
rect 19656 13568 19720 13572
rect 19736 13628 19800 13632
rect 19736 13572 19740 13628
rect 19740 13572 19796 13628
rect 19796 13572 19800 13628
rect 19736 13568 19800 13572
rect 19816 13628 19880 13632
rect 19816 13572 19820 13628
rect 19820 13572 19876 13628
rect 19876 13572 19880 13628
rect 19816 13568 19880 13572
rect 14780 13364 14844 13428
rect 14412 13228 14476 13292
rect 4216 13084 4280 13088
rect 4216 13028 4220 13084
rect 4220 13028 4276 13084
rect 4276 13028 4280 13084
rect 4216 13024 4280 13028
rect 4296 13084 4360 13088
rect 4296 13028 4300 13084
rect 4300 13028 4356 13084
rect 4356 13028 4360 13084
rect 4296 13024 4360 13028
rect 4376 13084 4440 13088
rect 4376 13028 4380 13084
rect 4380 13028 4436 13084
rect 4436 13028 4440 13084
rect 4376 13024 4440 13028
rect 4456 13084 4520 13088
rect 4456 13028 4460 13084
rect 4460 13028 4516 13084
rect 4516 13028 4520 13084
rect 4456 13024 4520 13028
rect 34936 13084 35000 13088
rect 34936 13028 34940 13084
rect 34940 13028 34996 13084
rect 34996 13028 35000 13084
rect 34936 13024 35000 13028
rect 35016 13084 35080 13088
rect 35016 13028 35020 13084
rect 35020 13028 35076 13084
rect 35076 13028 35080 13084
rect 35016 13024 35080 13028
rect 35096 13084 35160 13088
rect 35096 13028 35100 13084
rect 35100 13028 35156 13084
rect 35156 13028 35160 13084
rect 35096 13024 35160 13028
rect 35176 13084 35240 13088
rect 35176 13028 35180 13084
rect 35180 13028 35236 13084
rect 35236 13028 35240 13084
rect 35176 13024 35240 13028
rect 19576 12540 19640 12544
rect 19576 12484 19580 12540
rect 19580 12484 19636 12540
rect 19636 12484 19640 12540
rect 19576 12480 19640 12484
rect 19656 12540 19720 12544
rect 19656 12484 19660 12540
rect 19660 12484 19716 12540
rect 19716 12484 19720 12540
rect 19656 12480 19720 12484
rect 19736 12540 19800 12544
rect 19736 12484 19740 12540
rect 19740 12484 19796 12540
rect 19796 12484 19800 12540
rect 19736 12480 19800 12484
rect 19816 12540 19880 12544
rect 19816 12484 19820 12540
rect 19820 12484 19876 12540
rect 19876 12484 19880 12540
rect 19816 12480 19880 12484
rect 9628 12412 9692 12476
rect 15700 12412 15764 12476
rect 28948 12140 29012 12204
rect 4216 11996 4280 12000
rect 4216 11940 4220 11996
rect 4220 11940 4276 11996
rect 4276 11940 4280 11996
rect 4216 11936 4280 11940
rect 4296 11996 4360 12000
rect 4296 11940 4300 11996
rect 4300 11940 4356 11996
rect 4356 11940 4360 11996
rect 4296 11936 4360 11940
rect 4376 11996 4440 12000
rect 4376 11940 4380 11996
rect 4380 11940 4436 11996
rect 4436 11940 4440 11996
rect 4376 11936 4440 11940
rect 4456 11996 4520 12000
rect 4456 11940 4460 11996
rect 4460 11940 4516 11996
rect 4516 11940 4520 11996
rect 4456 11936 4520 11940
rect 34936 11996 35000 12000
rect 34936 11940 34940 11996
rect 34940 11940 34996 11996
rect 34996 11940 35000 11996
rect 34936 11936 35000 11940
rect 35016 11996 35080 12000
rect 35016 11940 35020 11996
rect 35020 11940 35076 11996
rect 35076 11940 35080 11996
rect 35016 11936 35080 11940
rect 35096 11996 35160 12000
rect 35096 11940 35100 11996
rect 35100 11940 35156 11996
rect 35156 11940 35160 11996
rect 35096 11936 35160 11940
rect 35176 11996 35240 12000
rect 35176 11940 35180 11996
rect 35180 11940 35236 11996
rect 35236 11940 35240 11996
rect 35176 11936 35240 11940
rect 9628 11732 9692 11796
rect 19576 11452 19640 11456
rect 19576 11396 19580 11452
rect 19580 11396 19636 11452
rect 19636 11396 19640 11452
rect 19576 11392 19640 11396
rect 19656 11452 19720 11456
rect 19656 11396 19660 11452
rect 19660 11396 19716 11452
rect 19716 11396 19720 11452
rect 19656 11392 19720 11396
rect 19736 11452 19800 11456
rect 19736 11396 19740 11452
rect 19740 11396 19796 11452
rect 19796 11396 19800 11452
rect 19736 11392 19800 11396
rect 19816 11452 19880 11456
rect 19816 11396 19820 11452
rect 19820 11396 19876 11452
rect 19876 11396 19880 11452
rect 19816 11392 19880 11396
rect 28948 11188 29012 11252
rect 4216 10908 4280 10912
rect 4216 10852 4220 10908
rect 4220 10852 4276 10908
rect 4276 10852 4280 10908
rect 4216 10848 4280 10852
rect 4296 10908 4360 10912
rect 4296 10852 4300 10908
rect 4300 10852 4356 10908
rect 4356 10852 4360 10908
rect 4296 10848 4360 10852
rect 4376 10908 4440 10912
rect 4376 10852 4380 10908
rect 4380 10852 4436 10908
rect 4436 10852 4440 10908
rect 4376 10848 4440 10852
rect 4456 10908 4520 10912
rect 4456 10852 4460 10908
rect 4460 10852 4516 10908
rect 4516 10852 4520 10908
rect 4456 10848 4520 10852
rect 34936 10908 35000 10912
rect 34936 10852 34940 10908
rect 34940 10852 34996 10908
rect 34996 10852 35000 10908
rect 34936 10848 35000 10852
rect 35016 10908 35080 10912
rect 35016 10852 35020 10908
rect 35020 10852 35076 10908
rect 35076 10852 35080 10908
rect 35016 10848 35080 10852
rect 35096 10908 35160 10912
rect 35096 10852 35100 10908
rect 35100 10852 35156 10908
rect 35156 10852 35160 10908
rect 35096 10848 35160 10852
rect 35176 10908 35240 10912
rect 35176 10852 35180 10908
rect 35180 10852 35236 10908
rect 35236 10852 35240 10908
rect 35176 10848 35240 10852
rect 19576 10364 19640 10368
rect 19576 10308 19580 10364
rect 19580 10308 19636 10364
rect 19636 10308 19640 10364
rect 19576 10304 19640 10308
rect 19656 10364 19720 10368
rect 19656 10308 19660 10364
rect 19660 10308 19716 10364
rect 19716 10308 19720 10364
rect 19656 10304 19720 10308
rect 19736 10364 19800 10368
rect 19736 10308 19740 10364
rect 19740 10308 19796 10364
rect 19796 10308 19800 10364
rect 19736 10304 19800 10308
rect 19816 10364 19880 10368
rect 19816 10308 19820 10364
rect 19820 10308 19876 10364
rect 19876 10308 19880 10364
rect 19816 10304 19880 10308
rect 4216 9820 4280 9824
rect 4216 9764 4220 9820
rect 4220 9764 4276 9820
rect 4276 9764 4280 9820
rect 4216 9760 4280 9764
rect 4296 9820 4360 9824
rect 4296 9764 4300 9820
rect 4300 9764 4356 9820
rect 4356 9764 4360 9820
rect 4296 9760 4360 9764
rect 4376 9820 4440 9824
rect 4376 9764 4380 9820
rect 4380 9764 4436 9820
rect 4436 9764 4440 9820
rect 4376 9760 4440 9764
rect 4456 9820 4520 9824
rect 4456 9764 4460 9820
rect 4460 9764 4516 9820
rect 4516 9764 4520 9820
rect 4456 9760 4520 9764
rect 34936 9820 35000 9824
rect 34936 9764 34940 9820
rect 34940 9764 34996 9820
rect 34996 9764 35000 9820
rect 34936 9760 35000 9764
rect 35016 9820 35080 9824
rect 35016 9764 35020 9820
rect 35020 9764 35076 9820
rect 35076 9764 35080 9820
rect 35016 9760 35080 9764
rect 35096 9820 35160 9824
rect 35096 9764 35100 9820
rect 35100 9764 35156 9820
rect 35156 9764 35160 9820
rect 35096 9760 35160 9764
rect 35176 9820 35240 9824
rect 35176 9764 35180 9820
rect 35180 9764 35236 9820
rect 35236 9764 35240 9820
rect 35176 9760 35240 9764
rect 24348 9692 24412 9756
rect 30420 9556 30484 9620
rect 19576 9276 19640 9280
rect 19576 9220 19580 9276
rect 19580 9220 19636 9276
rect 19636 9220 19640 9276
rect 19576 9216 19640 9220
rect 19656 9276 19720 9280
rect 19656 9220 19660 9276
rect 19660 9220 19716 9276
rect 19716 9220 19720 9276
rect 19656 9216 19720 9220
rect 19736 9276 19800 9280
rect 19736 9220 19740 9276
rect 19740 9220 19796 9276
rect 19796 9220 19800 9276
rect 19736 9216 19800 9220
rect 19816 9276 19880 9280
rect 19816 9220 19820 9276
rect 19820 9220 19876 9276
rect 19876 9220 19880 9276
rect 19816 9216 19880 9220
rect 4216 8732 4280 8736
rect 4216 8676 4220 8732
rect 4220 8676 4276 8732
rect 4276 8676 4280 8732
rect 4216 8672 4280 8676
rect 4296 8732 4360 8736
rect 4296 8676 4300 8732
rect 4300 8676 4356 8732
rect 4356 8676 4360 8732
rect 4296 8672 4360 8676
rect 4376 8732 4440 8736
rect 4376 8676 4380 8732
rect 4380 8676 4436 8732
rect 4436 8676 4440 8732
rect 4376 8672 4440 8676
rect 4456 8732 4520 8736
rect 4456 8676 4460 8732
rect 4460 8676 4516 8732
rect 4516 8676 4520 8732
rect 4456 8672 4520 8676
rect 34936 8732 35000 8736
rect 34936 8676 34940 8732
rect 34940 8676 34996 8732
rect 34996 8676 35000 8732
rect 34936 8672 35000 8676
rect 35016 8732 35080 8736
rect 35016 8676 35020 8732
rect 35020 8676 35076 8732
rect 35076 8676 35080 8732
rect 35016 8672 35080 8676
rect 35096 8732 35160 8736
rect 35096 8676 35100 8732
rect 35100 8676 35156 8732
rect 35156 8676 35160 8732
rect 35096 8672 35160 8676
rect 35176 8732 35240 8736
rect 35176 8676 35180 8732
rect 35180 8676 35236 8732
rect 35236 8676 35240 8732
rect 35176 8672 35240 8676
rect 19576 8188 19640 8192
rect 19576 8132 19580 8188
rect 19580 8132 19636 8188
rect 19636 8132 19640 8188
rect 19576 8128 19640 8132
rect 19656 8188 19720 8192
rect 19656 8132 19660 8188
rect 19660 8132 19716 8188
rect 19716 8132 19720 8188
rect 19656 8128 19720 8132
rect 19736 8188 19800 8192
rect 19736 8132 19740 8188
rect 19740 8132 19796 8188
rect 19796 8132 19800 8188
rect 19736 8128 19800 8132
rect 19816 8188 19880 8192
rect 19816 8132 19820 8188
rect 19820 8132 19876 8188
rect 19876 8132 19880 8188
rect 19816 8128 19880 8132
rect 4216 7644 4280 7648
rect 4216 7588 4220 7644
rect 4220 7588 4276 7644
rect 4276 7588 4280 7644
rect 4216 7584 4280 7588
rect 4296 7644 4360 7648
rect 4296 7588 4300 7644
rect 4300 7588 4356 7644
rect 4356 7588 4360 7644
rect 4296 7584 4360 7588
rect 4376 7644 4440 7648
rect 4376 7588 4380 7644
rect 4380 7588 4436 7644
rect 4436 7588 4440 7644
rect 4376 7584 4440 7588
rect 4456 7644 4520 7648
rect 4456 7588 4460 7644
rect 4460 7588 4516 7644
rect 4516 7588 4520 7644
rect 4456 7584 4520 7588
rect 34936 7644 35000 7648
rect 34936 7588 34940 7644
rect 34940 7588 34996 7644
rect 34996 7588 35000 7644
rect 34936 7584 35000 7588
rect 35016 7644 35080 7648
rect 35016 7588 35020 7644
rect 35020 7588 35076 7644
rect 35076 7588 35080 7644
rect 35016 7584 35080 7588
rect 35096 7644 35160 7648
rect 35096 7588 35100 7644
rect 35100 7588 35156 7644
rect 35156 7588 35160 7644
rect 35096 7584 35160 7588
rect 35176 7644 35240 7648
rect 35176 7588 35180 7644
rect 35180 7588 35236 7644
rect 35236 7588 35240 7644
rect 35176 7584 35240 7588
rect 20300 7516 20364 7580
rect 19576 7100 19640 7104
rect 19576 7044 19580 7100
rect 19580 7044 19636 7100
rect 19636 7044 19640 7100
rect 19576 7040 19640 7044
rect 19656 7100 19720 7104
rect 19656 7044 19660 7100
rect 19660 7044 19716 7100
rect 19716 7044 19720 7100
rect 19656 7040 19720 7044
rect 19736 7100 19800 7104
rect 19736 7044 19740 7100
rect 19740 7044 19796 7100
rect 19796 7044 19800 7100
rect 19736 7040 19800 7044
rect 19816 7100 19880 7104
rect 19816 7044 19820 7100
rect 19820 7044 19876 7100
rect 19876 7044 19880 7100
rect 19816 7040 19880 7044
rect 4216 6556 4280 6560
rect 4216 6500 4220 6556
rect 4220 6500 4276 6556
rect 4276 6500 4280 6556
rect 4216 6496 4280 6500
rect 4296 6556 4360 6560
rect 4296 6500 4300 6556
rect 4300 6500 4356 6556
rect 4356 6500 4360 6556
rect 4296 6496 4360 6500
rect 4376 6556 4440 6560
rect 4376 6500 4380 6556
rect 4380 6500 4436 6556
rect 4436 6500 4440 6556
rect 4376 6496 4440 6500
rect 4456 6556 4520 6560
rect 4456 6500 4460 6556
rect 4460 6500 4516 6556
rect 4516 6500 4520 6556
rect 4456 6496 4520 6500
rect 34936 6556 35000 6560
rect 34936 6500 34940 6556
rect 34940 6500 34996 6556
rect 34996 6500 35000 6556
rect 34936 6496 35000 6500
rect 35016 6556 35080 6560
rect 35016 6500 35020 6556
rect 35020 6500 35076 6556
rect 35076 6500 35080 6556
rect 35016 6496 35080 6500
rect 35096 6556 35160 6560
rect 35096 6500 35100 6556
rect 35100 6500 35156 6556
rect 35156 6500 35160 6556
rect 35096 6496 35160 6500
rect 35176 6556 35240 6560
rect 35176 6500 35180 6556
rect 35180 6500 35236 6556
rect 35236 6500 35240 6556
rect 35176 6496 35240 6500
rect 19576 6012 19640 6016
rect 19576 5956 19580 6012
rect 19580 5956 19636 6012
rect 19636 5956 19640 6012
rect 19576 5952 19640 5956
rect 19656 6012 19720 6016
rect 19656 5956 19660 6012
rect 19660 5956 19716 6012
rect 19716 5956 19720 6012
rect 19656 5952 19720 5956
rect 19736 6012 19800 6016
rect 19736 5956 19740 6012
rect 19740 5956 19796 6012
rect 19796 5956 19800 6012
rect 19736 5952 19800 5956
rect 19816 6012 19880 6016
rect 19816 5956 19820 6012
rect 19820 5956 19876 6012
rect 19876 5956 19880 6012
rect 19816 5952 19880 5956
rect 4216 5468 4280 5472
rect 4216 5412 4220 5468
rect 4220 5412 4276 5468
rect 4276 5412 4280 5468
rect 4216 5408 4280 5412
rect 4296 5468 4360 5472
rect 4296 5412 4300 5468
rect 4300 5412 4356 5468
rect 4356 5412 4360 5468
rect 4296 5408 4360 5412
rect 4376 5468 4440 5472
rect 4376 5412 4380 5468
rect 4380 5412 4436 5468
rect 4436 5412 4440 5468
rect 4376 5408 4440 5412
rect 4456 5468 4520 5472
rect 4456 5412 4460 5468
rect 4460 5412 4516 5468
rect 4516 5412 4520 5468
rect 4456 5408 4520 5412
rect 34936 5468 35000 5472
rect 34936 5412 34940 5468
rect 34940 5412 34996 5468
rect 34996 5412 35000 5468
rect 34936 5408 35000 5412
rect 35016 5468 35080 5472
rect 35016 5412 35020 5468
rect 35020 5412 35076 5468
rect 35076 5412 35080 5468
rect 35016 5408 35080 5412
rect 35096 5468 35160 5472
rect 35096 5412 35100 5468
rect 35100 5412 35156 5468
rect 35156 5412 35160 5468
rect 35096 5408 35160 5412
rect 35176 5468 35240 5472
rect 35176 5412 35180 5468
rect 35180 5412 35236 5468
rect 35236 5412 35240 5468
rect 35176 5408 35240 5412
rect 19576 4924 19640 4928
rect 19576 4868 19580 4924
rect 19580 4868 19636 4924
rect 19636 4868 19640 4924
rect 19576 4864 19640 4868
rect 19656 4924 19720 4928
rect 19656 4868 19660 4924
rect 19660 4868 19716 4924
rect 19716 4868 19720 4924
rect 19656 4864 19720 4868
rect 19736 4924 19800 4928
rect 19736 4868 19740 4924
rect 19740 4868 19796 4924
rect 19796 4868 19800 4924
rect 19736 4864 19800 4868
rect 19816 4924 19880 4928
rect 19816 4868 19820 4924
rect 19820 4868 19876 4924
rect 19876 4868 19880 4924
rect 19816 4864 19880 4868
rect 14044 4856 14108 4860
rect 14044 4800 14058 4856
rect 14058 4800 14108 4856
rect 14044 4796 14108 4800
rect 28948 4796 29012 4860
rect 9628 4524 9692 4588
rect 17908 4524 17972 4588
rect 4216 4380 4280 4384
rect 4216 4324 4220 4380
rect 4220 4324 4276 4380
rect 4276 4324 4280 4380
rect 4216 4320 4280 4324
rect 4296 4380 4360 4384
rect 4296 4324 4300 4380
rect 4300 4324 4356 4380
rect 4356 4324 4360 4380
rect 4296 4320 4360 4324
rect 4376 4380 4440 4384
rect 4376 4324 4380 4380
rect 4380 4324 4436 4380
rect 4436 4324 4440 4380
rect 4376 4320 4440 4324
rect 4456 4380 4520 4384
rect 4456 4324 4460 4380
rect 4460 4324 4516 4380
rect 4516 4324 4520 4380
rect 4456 4320 4520 4324
rect 34936 4380 35000 4384
rect 34936 4324 34940 4380
rect 34940 4324 34996 4380
rect 34996 4324 35000 4380
rect 34936 4320 35000 4324
rect 35016 4380 35080 4384
rect 35016 4324 35020 4380
rect 35020 4324 35076 4380
rect 35076 4324 35080 4380
rect 35016 4320 35080 4324
rect 35096 4380 35160 4384
rect 35096 4324 35100 4380
rect 35100 4324 35156 4380
rect 35156 4324 35160 4380
rect 35096 4320 35160 4324
rect 35176 4380 35240 4384
rect 35176 4324 35180 4380
rect 35180 4324 35236 4380
rect 35236 4324 35240 4380
rect 35176 4320 35240 4324
rect 9628 4312 9692 4316
rect 9628 4256 9642 4312
rect 9642 4256 9692 4312
rect 9628 4252 9692 4256
rect 17908 4252 17972 4316
rect 28948 4252 29012 4316
rect 14228 4040 14292 4044
rect 14228 3984 14278 4040
rect 14278 3984 14292 4040
rect 14228 3980 14292 3984
rect 19576 3836 19640 3840
rect 19576 3780 19580 3836
rect 19580 3780 19636 3836
rect 19636 3780 19640 3836
rect 19576 3776 19640 3780
rect 19656 3836 19720 3840
rect 19656 3780 19660 3836
rect 19660 3780 19716 3836
rect 19716 3780 19720 3836
rect 19656 3776 19720 3780
rect 19736 3836 19800 3840
rect 19736 3780 19740 3836
rect 19740 3780 19796 3836
rect 19796 3780 19800 3836
rect 19736 3776 19800 3780
rect 19816 3836 19880 3840
rect 19816 3780 19820 3836
rect 19820 3780 19876 3836
rect 19876 3780 19880 3836
rect 19816 3776 19880 3780
rect 4216 3292 4280 3296
rect 4216 3236 4220 3292
rect 4220 3236 4276 3292
rect 4276 3236 4280 3292
rect 4216 3232 4280 3236
rect 4296 3292 4360 3296
rect 4296 3236 4300 3292
rect 4300 3236 4356 3292
rect 4356 3236 4360 3292
rect 4296 3232 4360 3236
rect 4376 3292 4440 3296
rect 4376 3236 4380 3292
rect 4380 3236 4436 3292
rect 4436 3236 4440 3292
rect 4376 3232 4440 3236
rect 4456 3292 4520 3296
rect 4456 3236 4460 3292
rect 4460 3236 4516 3292
rect 4516 3236 4520 3292
rect 4456 3232 4520 3236
rect 34936 3292 35000 3296
rect 34936 3236 34940 3292
rect 34940 3236 34996 3292
rect 34996 3236 35000 3292
rect 34936 3232 35000 3236
rect 35016 3292 35080 3296
rect 35016 3236 35020 3292
rect 35020 3236 35076 3292
rect 35076 3236 35080 3292
rect 35016 3232 35080 3236
rect 35096 3292 35160 3296
rect 35096 3236 35100 3292
rect 35100 3236 35156 3292
rect 35156 3236 35160 3292
rect 35096 3232 35160 3236
rect 35176 3292 35240 3296
rect 35176 3236 35180 3292
rect 35180 3236 35236 3292
rect 35236 3236 35240 3292
rect 35176 3232 35240 3236
rect 19576 2748 19640 2752
rect 19576 2692 19580 2748
rect 19580 2692 19636 2748
rect 19636 2692 19640 2748
rect 19576 2688 19640 2692
rect 19656 2748 19720 2752
rect 19656 2692 19660 2748
rect 19660 2692 19716 2748
rect 19716 2692 19720 2748
rect 19656 2688 19720 2692
rect 19736 2748 19800 2752
rect 19736 2692 19740 2748
rect 19740 2692 19796 2748
rect 19796 2692 19800 2748
rect 19736 2688 19800 2692
rect 19816 2748 19880 2752
rect 19816 2692 19820 2748
rect 19820 2692 19876 2748
rect 19876 2692 19880 2748
rect 19816 2688 19880 2692
rect 28396 2680 28460 2684
rect 28396 2624 28446 2680
rect 28446 2624 28460 2680
rect 28396 2620 28460 2624
rect 4216 2204 4280 2208
rect 4216 2148 4220 2204
rect 4220 2148 4276 2204
rect 4276 2148 4280 2204
rect 4216 2144 4280 2148
rect 4296 2204 4360 2208
rect 4296 2148 4300 2204
rect 4300 2148 4356 2204
rect 4356 2148 4360 2204
rect 4296 2144 4360 2148
rect 4376 2204 4440 2208
rect 4376 2148 4380 2204
rect 4380 2148 4436 2204
rect 4436 2148 4440 2204
rect 4376 2144 4440 2148
rect 4456 2204 4520 2208
rect 4456 2148 4460 2204
rect 4460 2148 4516 2204
rect 4516 2148 4520 2204
rect 4456 2144 4520 2148
rect 34936 2204 35000 2208
rect 34936 2148 34940 2204
rect 34940 2148 34996 2204
rect 34996 2148 35000 2204
rect 34936 2144 35000 2148
rect 35016 2204 35080 2208
rect 35016 2148 35020 2204
rect 35020 2148 35076 2204
rect 35076 2148 35080 2204
rect 35016 2144 35080 2148
rect 35096 2204 35160 2208
rect 35096 2148 35100 2204
rect 35100 2148 35156 2204
rect 35156 2148 35160 2204
rect 35096 2144 35160 2148
rect 35176 2204 35240 2208
rect 35176 2148 35180 2204
rect 35180 2148 35236 2204
rect 35236 2148 35240 2204
rect 35176 2144 35240 2148
rect 30420 912 30484 916
rect 30420 856 30434 912
rect 30434 856 30484 912
rect 30420 852 30484 856
<< metal4 >>
rect 4208 77280 4528 77840
rect 4208 77216 4216 77280
rect 4280 77216 4296 77280
rect 4360 77216 4376 77280
rect 4440 77216 4456 77280
rect 4520 77216 4528 77280
rect 4208 76192 4528 77216
rect 4208 76128 4216 76192
rect 4280 76128 4296 76192
rect 4360 76128 4376 76192
rect 4440 76128 4456 76192
rect 4520 76128 4528 76192
rect 4208 75104 4528 76128
rect 4208 75040 4216 75104
rect 4280 75040 4296 75104
rect 4360 75040 4376 75104
rect 4440 75040 4456 75104
rect 4520 75040 4528 75104
rect 4208 74016 4528 75040
rect 4208 73952 4216 74016
rect 4280 73952 4296 74016
rect 4360 73952 4376 74016
rect 4440 73952 4456 74016
rect 4520 73952 4528 74016
rect 4208 72928 4528 73952
rect 4208 72864 4216 72928
rect 4280 72864 4296 72928
rect 4360 72864 4376 72928
rect 4440 72864 4456 72928
rect 4520 72864 4528 72928
rect 4208 71840 4528 72864
rect 4208 71776 4216 71840
rect 4280 71776 4296 71840
rect 4360 71776 4376 71840
rect 4440 71776 4456 71840
rect 4520 71776 4528 71840
rect 4208 70752 4528 71776
rect 4208 70688 4216 70752
rect 4280 70688 4296 70752
rect 4360 70688 4376 70752
rect 4440 70688 4456 70752
rect 4520 70688 4528 70752
rect 4208 69664 4528 70688
rect 4208 69600 4216 69664
rect 4280 69600 4296 69664
rect 4360 69600 4376 69664
rect 4440 69600 4456 69664
rect 4520 69600 4528 69664
rect 4208 68576 4528 69600
rect 4208 68512 4216 68576
rect 4280 68512 4296 68576
rect 4360 68512 4376 68576
rect 4440 68512 4456 68576
rect 4520 68512 4528 68576
rect 4208 67488 4528 68512
rect 4208 67424 4216 67488
rect 4280 67424 4296 67488
rect 4360 67424 4376 67488
rect 4440 67424 4456 67488
rect 4520 67424 4528 67488
rect 4208 66848 4528 67424
rect 4208 66612 4250 66848
rect 4486 66612 4528 66848
rect 4208 66400 4528 66612
rect 4208 66336 4216 66400
rect 4280 66336 4296 66400
rect 4360 66336 4376 66400
rect 4440 66336 4456 66400
rect 4520 66336 4528 66400
rect 4208 65312 4528 66336
rect 4208 65248 4216 65312
rect 4280 65248 4296 65312
rect 4360 65248 4376 65312
rect 4440 65248 4456 65312
rect 4520 65248 4528 65312
rect 4208 64224 4528 65248
rect 4208 64160 4216 64224
rect 4280 64160 4296 64224
rect 4360 64160 4376 64224
rect 4440 64160 4456 64224
rect 4520 64160 4528 64224
rect 4208 63136 4528 64160
rect 4208 63072 4216 63136
rect 4280 63072 4296 63136
rect 4360 63072 4376 63136
rect 4440 63072 4456 63136
rect 4520 63072 4528 63136
rect 4208 62048 4528 63072
rect 4208 61984 4216 62048
rect 4280 61984 4296 62048
rect 4360 61984 4376 62048
rect 4440 61984 4456 62048
rect 4520 61984 4528 62048
rect 4208 60960 4528 61984
rect 4208 60896 4216 60960
rect 4280 60896 4296 60960
rect 4360 60896 4376 60960
rect 4440 60896 4456 60960
rect 4520 60896 4528 60960
rect 4208 59872 4528 60896
rect 4208 59808 4216 59872
rect 4280 59808 4296 59872
rect 4360 59808 4376 59872
rect 4440 59808 4456 59872
rect 4520 59808 4528 59872
rect 4208 58784 4528 59808
rect 4208 58720 4216 58784
rect 4280 58720 4296 58784
rect 4360 58720 4376 58784
rect 4440 58720 4456 58784
rect 4520 58720 4528 58784
rect 4208 57696 4528 58720
rect 4208 57632 4216 57696
rect 4280 57632 4296 57696
rect 4360 57632 4376 57696
rect 4440 57632 4456 57696
rect 4520 57632 4528 57696
rect 4208 56608 4528 57632
rect 4208 56544 4216 56608
rect 4280 56544 4296 56608
rect 4360 56544 4376 56608
rect 4440 56544 4456 56608
rect 4520 56544 4528 56608
rect 4208 55520 4528 56544
rect 4208 55456 4216 55520
rect 4280 55456 4296 55520
rect 4360 55456 4376 55520
rect 4440 55456 4456 55520
rect 4520 55456 4528 55520
rect 4208 54432 4528 55456
rect 4208 54368 4216 54432
rect 4280 54368 4296 54432
rect 4360 54368 4376 54432
rect 4440 54368 4456 54432
rect 4520 54368 4528 54432
rect 4208 53344 4528 54368
rect 19568 77824 19888 77840
rect 19568 77760 19576 77824
rect 19640 77760 19656 77824
rect 19720 77760 19736 77824
rect 19800 77760 19816 77824
rect 19880 77760 19888 77824
rect 19568 76736 19888 77760
rect 19568 76672 19576 76736
rect 19640 76672 19656 76736
rect 19720 76672 19736 76736
rect 19800 76672 19816 76736
rect 19880 76672 19888 76736
rect 19568 75648 19888 76672
rect 19568 75584 19576 75648
rect 19640 75584 19656 75648
rect 19720 75584 19736 75648
rect 19800 75584 19816 75648
rect 19880 75584 19888 75648
rect 19568 74560 19888 75584
rect 19568 74496 19576 74560
rect 19640 74496 19656 74560
rect 19720 74496 19736 74560
rect 19800 74496 19816 74560
rect 19880 74496 19888 74560
rect 19568 73472 19888 74496
rect 19568 73408 19576 73472
rect 19640 73408 19656 73472
rect 19720 73408 19736 73472
rect 19800 73408 19816 73472
rect 19880 73408 19888 73472
rect 19568 72384 19888 73408
rect 34928 77280 35248 77840
rect 34928 77216 34936 77280
rect 35000 77216 35016 77280
rect 35080 77216 35096 77280
rect 35160 77216 35176 77280
rect 35240 77216 35248 77280
rect 34928 76192 35248 77216
rect 34928 76128 34936 76192
rect 35000 76128 35016 76192
rect 35080 76128 35096 76192
rect 35160 76128 35176 76192
rect 35240 76128 35248 76192
rect 34928 75104 35248 76128
rect 34928 75040 34936 75104
rect 35000 75040 35016 75104
rect 35080 75040 35096 75104
rect 35160 75040 35176 75104
rect 35240 75040 35248 75104
rect 34928 74016 35248 75040
rect 34928 73952 34936 74016
rect 35000 73952 35016 74016
rect 35080 73952 35096 74016
rect 35160 73952 35176 74016
rect 35240 73952 35248 74016
rect 28947 73268 29013 73269
rect 28947 73204 28948 73268
rect 29012 73204 29013 73268
rect 28947 73203 29013 73204
rect 28950 72997 29010 73203
rect 28947 72996 29013 72997
rect 28947 72932 28948 72996
rect 29012 72932 29013 72996
rect 28947 72931 29013 72932
rect 19568 72320 19576 72384
rect 19640 72320 19656 72384
rect 19720 72320 19736 72384
rect 19800 72320 19816 72384
rect 19880 72320 19888 72384
rect 19568 71296 19888 72320
rect 34928 72928 35248 73952
rect 34928 72864 34936 72928
rect 35000 72864 35016 72928
rect 35080 72864 35096 72928
rect 35160 72864 35176 72928
rect 35240 72864 35248 72928
rect 21035 71908 21101 71909
rect 21035 71844 21036 71908
rect 21100 71844 21101 71908
rect 21035 71843 21101 71844
rect 19568 71232 19576 71296
rect 19640 71232 19656 71296
rect 19720 71232 19736 71296
rect 19800 71232 19816 71296
rect 19880 71232 19888 71296
rect 19568 70208 19888 71232
rect 19568 70144 19576 70208
rect 19640 70144 19656 70208
rect 19720 70144 19736 70208
rect 19800 70144 19816 70208
rect 19880 70144 19888 70208
rect 19568 69120 19888 70144
rect 19568 69056 19576 69120
rect 19640 69056 19656 69120
rect 19720 69056 19736 69120
rect 19800 69056 19816 69120
rect 19880 69056 19888 69120
rect 19568 68032 19888 69056
rect 19568 67968 19576 68032
rect 19640 67968 19656 68032
rect 19720 67968 19736 68032
rect 19800 67968 19816 68032
rect 19880 67968 19888 68032
rect 19568 66944 19888 67968
rect 19568 66880 19576 66944
rect 19640 66880 19656 66944
rect 19720 66880 19736 66944
rect 19800 66880 19816 66944
rect 19880 66880 19888 66944
rect 19568 65856 19888 66880
rect 19568 65792 19576 65856
rect 19640 65792 19656 65856
rect 19720 65792 19736 65856
rect 19800 65792 19816 65856
rect 19880 65792 19888 65856
rect 19568 64768 19888 65792
rect 19568 64704 19576 64768
rect 19640 64704 19656 64768
rect 19720 64704 19736 64768
rect 19800 64704 19816 64768
rect 19880 64704 19888 64768
rect 19568 63680 19888 64704
rect 19568 63616 19576 63680
rect 19640 63616 19656 63680
rect 19720 63616 19736 63680
rect 19800 63616 19816 63680
rect 19880 63616 19888 63680
rect 19568 62592 19888 63616
rect 19568 62528 19576 62592
rect 19640 62528 19656 62592
rect 19720 62528 19736 62592
rect 19800 62528 19816 62592
rect 19880 62528 19888 62592
rect 19568 61504 19888 62528
rect 19568 61440 19576 61504
rect 19640 61440 19656 61504
rect 19720 61440 19736 61504
rect 19800 61440 19816 61504
rect 19880 61440 19888 61504
rect 19568 60416 19888 61440
rect 19568 60352 19576 60416
rect 19640 60352 19656 60416
rect 19720 60352 19736 60416
rect 19800 60352 19816 60416
rect 19880 60352 19888 60416
rect 19568 59328 19888 60352
rect 19568 59264 19576 59328
rect 19640 59264 19656 59328
rect 19720 59264 19736 59328
rect 19800 59264 19816 59328
rect 19880 59264 19888 59328
rect 19568 58240 19888 59264
rect 19568 58176 19576 58240
rect 19640 58176 19656 58240
rect 19720 58176 19736 58240
rect 19800 58176 19816 58240
rect 19880 58176 19888 58240
rect 19568 57152 19888 58176
rect 19568 57088 19576 57152
rect 19640 57088 19656 57152
rect 19720 57088 19736 57152
rect 19800 57088 19816 57152
rect 19880 57088 19888 57152
rect 19568 56064 19888 57088
rect 19568 56000 19576 56064
rect 19640 56000 19656 56064
rect 19720 56000 19736 56064
rect 19800 56000 19816 56064
rect 19880 56000 19888 56064
rect 19568 54976 19888 56000
rect 19568 54912 19576 54976
rect 19640 54912 19656 54976
rect 19720 54912 19736 54976
rect 19800 54912 19816 54976
rect 19880 54912 19888 54976
rect 14779 53956 14845 53957
rect 14779 53892 14780 53956
rect 14844 53892 14845 53956
rect 14779 53891 14845 53892
rect 4208 53280 4216 53344
rect 4280 53280 4296 53344
rect 4360 53280 4376 53344
rect 4440 53280 4456 53344
rect 4520 53280 4528 53344
rect 4208 52256 4528 53280
rect 4208 52192 4216 52256
rect 4280 52192 4296 52256
rect 4360 52192 4376 52256
rect 4440 52192 4456 52256
rect 4520 52192 4528 52256
rect 4208 51168 4528 52192
rect 4208 51104 4216 51168
rect 4280 51104 4296 51168
rect 4360 51104 4376 51168
rect 4440 51104 4456 51168
rect 4520 51104 4528 51168
rect 4208 50080 4528 51104
rect 4208 50016 4216 50080
rect 4280 50016 4296 50080
rect 4360 50016 4376 50080
rect 4440 50016 4456 50080
rect 4520 50016 4528 50080
rect 4208 48992 4528 50016
rect 4208 48928 4216 48992
rect 4280 48928 4296 48992
rect 4360 48928 4376 48992
rect 4440 48928 4456 48992
rect 4520 48928 4528 48992
rect 4208 47904 4528 48928
rect 4208 47840 4216 47904
rect 4280 47840 4296 47904
rect 4360 47840 4376 47904
rect 4440 47840 4456 47904
rect 4520 47840 4528 47904
rect 4208 46816 4528 47840
rect 4208 46752 4216 46816
rect 4280 46752 4296 46816
rect 4360 46752 4376 46816
rect 4440 46752 4456 46816
rect 4520 46752 4528 46816
rect 4208 45728 4528 46752
rect 4208 45664 4216 45728
rect 4280 45664 4296 45728
rect 4360 45664 4376 45728
rect 4440 45664 4456 45728
rect 4520 45664 4528 45728
rect 4208 44640 4528 45664
rect 4208 44576 4216 44640
rect 4280 44576 4296 44640
rect 4360 44576 4376 44640
rect 4440 44576 4456 44640
rect 4520 44576 4528 44640
rect 4208 43552 4528 44576
rect 4208 43488 4216 43552
rect 4280 43488 4296 43552
rect 4360 43488 4376 43552
rect 4440 43488 4456 43552
rect 4520 43488 4528 43552
rect 4208 42464 4528 43488
rect 4208 42400 4216 42464
rect 4280 42400 4296 42464
rect 4360 42400 4376 42464
rect 4440 42400 4456 42464
rect 4520 42400 4528 42464
rect 4208 41376 4528 42400
rect 14411 41852 14477 41853
rect 14411 41788 14412 41852
rect 14476 41788 14477 41852
rect 14411 41787 14477 41788
rect 4208 41312 4216 41376
rect 4280 41312 4296 41376
rect 4360 41312 4376 41376
rect 4440 41312 4456 41376
rect 4520 41312 4528 41376
rect 4208 40288 4528 41312
rect 13675 40492 13741 40493
rect 13675 40428 13676 40492
rect 13740 40428 13741 40492
rect 13675 40427 13741 40428
rect 4208 40224 4216 40288
rect 4280 40224 4296 40288
rect 4360 40224 4376 40288
rect 4440 40224 4456 40288
rect 4520 40224 4528 40288
rect 4208 39200 4528 40224
rect 4208 39136 4216 39200
rect 4280 39136 4296 39200
rect 4360 39136 4376 39200
rect 4440 39136 4456 39200
rect 4520 39136 4528 39200
rect 4208 38112 4528 39136
rect 4208 38048 4216 38112
rect 4280 38048 4296 38112
rect 4360 38048 4376 38112
rect 4440 38048 4456 38112
rect 4520 38048 4528 38112
rect 4208 37024 4528 38048
rect 4208 36960 4216 37024
rect 4280 36960 4296 37024
rect 4360 36960 4376 37024
rect 4440 36960 4456 37024
rect 4520 36960 4528 37024
rect 4208 36212 4528 36960
rect 4208 35976 4250 36212
rect 4486 35976 4528 36212
rect 9630 36141 9690 36942
rect 9627 36140 9693 36141
rect 9627 36076 9628 36140
rect 9692 36076 9693 36140
rect 9627 36075 9693 36076
rect 4208 35936 4528 35976
rect 4208 35872 4216 35936
rect 4280 35872 4296 35936
rect 4360 35872 4376 35936
rect 4440 35872 4456 35936
rect 4520 35872 4528 35936
rect 4208 34848 4528 35872
rect 4208 34784 4216 34848
rect 4280 34784 4296 34848
rect 4360 34784 4376 34848
rect 4440 34784 4456 34848
rect 4520 34784 4528 34848
rect 4208 33760 4528 34784
rect 13123 34644 13189 34645
rect 13123 34580 13124 34644
rect 13188 34580 13189 34644
rect 13123 34579 13189 34580
rect 8339 34508 8405 34509
rect 8339 34444 8340 34508
rect 8404 34444 8405 34508
rect 8339 34443 8405 34444
rect 4208 33696 4216 33760
rect 4280 33696 4296 33760
rect 4360 33696 4376 33760
rect 4440 33696 4456 33760
rect 4520 33696 4528 33760
rect 4208 32672 4528 33696
rect 4208 32608 4216 32672
rect 4280 32608 4296 32672
rect 4360 32608 4376 32672
rect 4440 32608 4456 32672
rect 4520 32608 4528 32672
rect 4208 31584 4528 32608
rect 4208 31520 4216 31584
rect 4280 31520 4296 31584
rect 4360 31520 4376 31584
rect 4440 31520 4456 31584
rect 4520 31520 4528 31584
rect 4208 30496 4528 31520
rect 4208 30432 4216 30496
rect 4280 30432 4296 30496
rect 4360 30432 4376 30496
rect 4440 30432 4456 30496
rect 4520 30432 4528 30496
rect 4208 29408 4528 30432
rect 4208 29344 4216 29408
rect 4280 29344 4296 29408
rect 4360 29344 4376 29408
rect 4440 29344 4456 29408
rect 4520 29344 4528 29408
rect 4208 28320 4528 29344
rect 8342 29205 8402 34443
rect 12571 34236 12637 34237
rect 12571 34172 12572 34236
rect 12636 34172 12637 34236
rect 12571 34171 12637 34172
rect 12574 30973 12634 34171
rect 13126 33146 13186 34579
rect 13491 33148 13557 33149
rect 13126 33086 13370 33146
rect 12571 30972 12637 30973
rect 12571 30908 12572 30972
rect 12636 30908 12637 30972
rect 12571 30907 12637 30908
rect 13123 30700 13189 30701
rect 13123 30636 13124 30700
rect 13188 30636 13189 30700
rect 13123 30635 13189 30636
rect 8339 29204 8405 29205
rect 8339 29140 8340 29204
rect 8404 29140 8405 29204
rect 8339 29139 8405 29140
rect 4208 28256 4216 28320
rect 4280 28256 4296 28320
rect 4360 28256 4376 28320
rect 4440 28256 4456 28320
rect 4520 28256 4528 28320
rect 4208 27232 4528 28256
rect 4208 27168 4216 27232
rect 4280 27168 4296 27232
rect 4360 27168 4376 27232
rect 4440 27168 4456 27232
rect 4520 27168 4528 27232
rect 4208 26144 4528 27168
rect 7235 26756 7301 26757
rect 7235 26692 7236 26756
rect 7300 26692 7301 26756
rect 7235 26691 7301 26692
rect 6683 26348 6749 26349
rect 6683 26298 6684 26348
rect 6748 26298 6749 26348
rect 4208 26080 4216 26144
rect 4280 26080 4296 26144
rect 4360 26080 4376 26144
rect 4440 26080 4456 26144
rect 4520 26080 4528 26144
rect 4208 25056 4528 26080
rect 4208 24992 4216 25056
rect 4280 24992 4296 25056
rect 4360 24992 4376 25056
rect 4440 24992 4456 25056
rect 4520 24992 4528 25056
rect 4208 23968 4528 24992
rect 4208 23904 4216 23968
rect 4280 23904 4296 23968
rect 4360 23904 4376 23968
rect 4440 23904 4456 23968
rect 4520 23904 4528 23968
rect 4208 22880 4528 23904
rect 4208 22816 4216 22880
rect 4280 22816 4296 22880
rect 4360 22816 4376 22880
rect 4440 22816 4456 22880
rect 4520 22816 4528 22880
rect 4208 21792 4528 22816
rect 4208 21728 4216 21792
rect 4280 21728 4296 21792
rect 4360 21728 4376 21792
rect 4440 21728 4456 21792
rect 4520 21728 4528 21792
rect 4208 20704 4528 21728
rect 7238 21538 7298 26691
rect 13126 26349 13186 30635
rect 13310 26485 13370 33086
rect 13491 33084 13492 33148
rect 13556 33084 13557 33148
rect 13491 33083 13557 33084
rect 13494 30701 13554 33083
rect 13491 30700 13557 30701
rect 13491 30636 13492 30700
rect 13556 30636 13557 30700
rect 13491 30635 13557 30636
rect 13307 26484 13373 26485
rect 13307 26420 13308 26484
rect 13372 26420 13373 26484
rect 13307 26419 13373 26420
rect 13123 26348 13189 26349
rect 13123 26284 13124 26348
rect 13188 26284 13189 26348
rect 13123 26283 13189 26284
rect 13678 24853 13738 40427
rect 14227 34780 14293 34781
rect 14227 34716 14228 34780
rect 14292 34716 14293 34780
rect 14227 34715 14293 34716
rect 13859 34644 13925 34645
rect 13859 34580 13860 34644
rect 13924 34580 13925 34644
rect 13859 34579 13925 34580
rect 13675 24852 13741 24853
rect 13675 24788 13676 24852
rect 13740 24788 13741 24852
rect 13675 24787 13741 24788
rect 4208 20640 4216 20704
rect 4280 20640 4296 20704
rect 4360 20640 4376 20704
rect 4440 20640 4456 20704
rect 4520 20640 4528 20704
rect 4208 19616 4528 20640
rect 4208 19552 4216 19616
rect 4280 19552 4296 19616
rect 4360 19552 4376 19616
rect 4440 19552 4456 19616
rect 4520 19552 4528 19616
rect 4208 18528 4528 19552
rect 4208 18464 4216 18528
rect 4280 18464 4296 18528
rect 4360 18464 4376 18528
rect 4440 18464 4456 18528
rect 4520 18464 4528 18528
rect 4208 17440 4528 18464
rect 4208 17376 4216 17440
rect 4280 17376 4296 17440
rect 4360 17376 4376 17440
rect 4440 17376 4456 17440
rect 4520 17376 4528 17440
rect 4208 16352 4528 17376
rect 4208 16288 4216 16352
rect 4280 16288 4296 16352
rect 4360 16288 4376 16352
rect 4440 16288 4456 16352
rect 4520 16288 4528 16352
rect 4208 15264 4528 16288
rect 4208 15200 4216 15264
rect 4280 15200 4296 15264
rect 4360 15200 4376 15264
rect 4440 15200 4456 15264
rect 4520 15200 4528 15264
rect 4208 14176 4528 15200
rect 13862 15061 13922 34579
rect 14230 31653 14290 34715
rect 14227 31652 14293 31653
rect 14227 31588 14228 31652
rect 14292 31588 14293 31652
rect 14227 31587 14293 31588
rect 14227 29204 14293 29205
rect 14227 29140 14228 29204
rect 14292 29140 14293 29204
rect 14227 29139 14293 29140
rect 14043 28252 14109 28253
rect 14043 28188 14044 28252
rect 14108 28188 14109 28252
rect 14043 28187 14109 28188
rect 14046 27301 14106 28187
rect 14043 27300 14109 27301
rect 14043 27236 14044 27300
rect 14108 27236 14109 27300
rect 14043 27235 14109 27236
rect 14230 27026 14290 29139
rect 14046 26966 14290 27026
rect 14046 23629 14106 26966
rect 14227 26892 14293 26893
rect 14227 26828 14228 26892
rect 14292 26828 14293 26892
rect 14227 26827 14293 26828
rect 14043 23628 14109 23629
rect 14043 23564 14044 23628
rect 14108 23564 14109 23628
rect 14043 23563 14109 23564
rect 13859 15060 13925 15061
rect 13859 14996 13860 15060
rect 13924 14996 13925 15060
rect 13859 14995 13925 14996
rect 4208 14112 4216 14176
rect 4280 14112 4296 14176
rect 4360 14112 4376 14176
rect 4440 14112 4456 14176
rect 4520 14112 4528 14176
rect 4208 13088 4528 14112
rect 4208 13024 4216 13088
rect 4280 13024 4296 13088
rect 4360 13024 4376 13088
rect 4440 13024 4456 13088
rect 4520 13024 4528 13088
rect 4208 12000 4528 13024
rect 9627 12476 9693 12477
rect 9627 12412 9628 12476
rect 9692 12412 9693 12476
rect 9627 12411 9693 12412
rect 4208 11936 4216 12000
rect 4280 11936 4296 12000
rect 4360 11936 4376 12000
rect 4440 11936 4456 12000
rect 4520 11936 4528 12000
rect 4208 10912 4528 11936
rect 9630 11797 9690 12411
rect 9627 11796 9693 11797
rect 9627 11732 9628 11796
rect 9692 11732 9693 11796
rect 9627 11731 9693 11732
rect 4208 10848 4216 10912
rect 4280 10848 4296 10912
rect 4360 10848 4376 10912
rect 4440 10848 4456 10912
rect 4520 10848 4528 10912
rect 4208 9824 4528 10848
rect 4208 9760 4216 9824
rect 4280 9760 4296 9824
rect 4360 9760 4376 9824
rect 4440 9760 4456 9824
rect 4520 9760 4528 9824
rect 4208 8736 4528 9760
rect 4208 8672 4216 8736
rect 4280 8672 4296 8736
rect 4360 8672 4376 8736
rect 4440 8672 4456 8736
rect 4520 8672 4528 8736
rect 4208 7648 4528 8672
rect 4208 7584 4216 7648
rect 4280 7584 4296 7648
rect 4360 7584 4376 7648
rect 4440 7584 4456 7648
rect 4520 7584 4528 7648
rect 4208 6560 4528 7584
rect 4208 6496 4216 6560
rect 4280 6496 4296 6560
rect 4360 6496 4376 6560
rect 4440 6496 4456 6560
rect 4520 6496 4528 6560
rect 4208 5576 4528 6496
rect 4208 5472 4250 5576
rect 4486 5472 4528 5576
rect 4208 5408 4216 5472
rect 4520 5408 4528 5472
rect 4208 5340 4250 5408
rect 4486 5340 4528 5408
rect 4208 4384 4528 5340
rect 14046 4861 14106 23563
rect 14043 4860 14109 4861
rect 14043 4796 14044 4860
rect 14108 4796 14109 4860
rect 14043 4795 14109 4796
rect 9627 4588 9693 4589
rect 9627 4524 9628 4588
rect 9692 4524 9693 4588
rect 9627 4523 9693 4524
rect 4208 4320 4216 4384
rect 4280 4320 4296 4384
rect 4360 4320 4376 4384
rect 4440 4320 4456 4384
rect 4520 4320 4528 4384
rect 4208 3296 4528 4320
rect 9630 4317 9690 4523
rect 9627 4316 9693 4317
rect 9627 4252 9628 4316
rect 9692 4252 9693 4316
rect 9627 4251 9693 4252
rect 14230 4045 14290 26827
rect 14414 13293 14474 41787
rect 14595 29204 14661 29205
rect 14595 29140 14596 29204
rect 14660 29140 14661 29204
rect 14595 29139 14661 29140
rect 14598 25125 14658 29139
rect 14595 25124 14661 25125
rect 14595 25060 14596 25124
rect 14660 25060 14661 25124
rect 14595 25059 14661 25060
rect 14782 13429 14842 53891
rect 19568 53888 19888 54912
rect 19568 53824 19576 53888
rect 19640 53824 19656 53888
rect 19720 53824 19736 53888
rect 19800 53824 19816 53888
rect 19880 53824 19888 53888
rect 19568 52800 19888 53824
rect 19568 52736 19576 52800
rect 19640 52736 19656 52800
rect 19720 52736 19736 52800
rect 19800 52736 19816 52800
rect 19880 52736 19888 52800
rect 19568 51712 19888 52736
rect 19568 51648 19576 51712
rect 19640 51648 19656 51712
rect 19720 51648 19736 51712
rect 19800 51648 19816 51712
rect 19880 51648 19888 51712
rect 19568 51530 19888 51648
rect 19568 51294 19610 51530
rect 19846 51294 19888 51530
rect 19568 50624 19888 51294
rect 19568 50560 19576 50624
rect 19640 50560 19656 50624
rect 19720 50560 19736 50624
rect 19800 50560 19816 50624
rect 19880 50560 19888 50624
rect 19568 49536 19888 50560
rect 19568 49472 19576 49536
rect 19640 49472 19656 49536
rect 19720 49472 19736 49536
rect 19800 49472 19816 49536
rect 19880 49472 19888 49536
rect 19568 48448 19888 49472
rect 19568 48384 19576 48448
rect 19640 48384 19656 48448
rect 19720 48384 19736 48448
rect 19800 48384 19816 48448
rect 19880 48384 19888 48448
rect 19568 47360 19888 48384
rect 19568 47296 19576 47360
rect 19640 47296 19656 47360
rect 19720 47296 19736 47360
rect 19800 47296 19816 47360
rect 19880 47296 19888 47360
rect 19568 46272 19888 47296
rect 20299 47020 20365 47021
rect 20299 46956 20300 47020
rect 20364 46956 20365 47020
rect 20299 46955 20365 46956
rect 19568 46208 19576 46272
rect 19640 46208 19656 46272
rect 19720 46208 19736 46272
rect 19800 46208 19816 46272
rect 19880 46208 19888 46272
rect 15699 46204 15765 46205
rect 15699 46140 15700 46204
rect 15764 46140 15765 46204
rect 15699 46139 15765 46140
rect 14963 35052 15029 35053
rect 14963 34988 14964 35052
rect 15028 34988 15029 35052
rect 14963 34987 15029 34988
rect 14966 34373 15026 34987
rect 14963 34372 15029 34373
rect 14963 34308 14964 34372
rect 15028 34308 15029 34372
rect 14963 34307 15029 34308
rect 15331 32468 15397 32469
rect 15331 32418 15332 32468
rect 15396 32418 15397 32468
rect 15334 31653 15394 32182
rect 14963 31652 15029 31653
rect 14963 31588 14964 31652
rect 15028 31588 15029 31652
rect 14963 31587 15029 31588
rect 15331 31652 15397 31653
rect 15331 31588 15332 31652
rect 15396 31588 15397 31652
rect 15331 31587 15397 31588
rect 14966 26893 15026 31587
rect 14963 26892 15029 26893
rect 14963 26828 14964 26892
rect 15028 26828 15029 26892
rect 14963 26827 15029 26828
rect 14779 13428 14845 13429
rect 14779 13364 14780 13428
rect 14844 13364 14845 13428
rect 14779 13363 14845 13364
rect 14411 13292 14477 13293
rect 14411 13228 14412 13292
rect 14476 13228 14477 13292
rect 14411 13227 14477 13228
rect 15702 12477 15762 46139
rect 19568 45184 19888 46208
rect 19568 45120 19576 45184
rect 19640 45120 19656 45184
rect 19720 45120 19736 45184
rect 19800 45120 19816 45184
rect 19880 45120 19888 45184
rect 19568 44096 19888 45120
rect 19568 44032 19576 44096
rect 19640 44032 19656 44096
rect 19720 44032 19736 44096
rect 19800 44032 19816 44096
rect 19880 44032 19888 44096
rect 19568 43008 19888 44032
rect 19568 42944 19576 43008
rect 19640 42944 19656 43008
rect 19720 42944 19736 43008
rect 19800 42944 19816 43008
rect 19880 42944 19888 43008
rect 19568 41920 19888 42944
rect 19568 41856 19576 41920
rect 19640 41856 19656 41920
rect 19720 41856 19736 41920
rect 19800 41856 19816 41920
rect 19880 41856 19888 41920
rect 19568 40832 19888 41856
rect 19568 40768 19576 40832
rect 19640 40768 19656 40832
rect 19720 40768 19736 40832
rect 19800 40768 19816 40832
rect 19880 40768 19888 40832
rect 19568 39744 19888 40768
rect 19568 39680 19576 39744
rect 19640 39680 19656 39744
rect 19720 39680 19736 39744
rect 19800 39680 19816 39744
rect 19880 39680 19888 39744
rect 15883 38724 15949 38725
rect 15883 38660 15884 38724
rect 15948 38660 15949 38724
rect 15883 38659 15949 38660
rect 15886 20773 15946 38659
rect 19568 38656 19888 39680
rect 19568 38592 19576 38656
rect 19640 38592 19656 38656
rect 19720 38592 19736 38656
rect 19800 38592 19816 38656
rect 19880 38592 19888 38656
rect 17171 37772 17237 37773
rect 17171 37708 17172 37772
rect 17236 37708 17237 37772
rect 17171 37707 17237 37708
rect 16803 34372 16869 34373
rect 16803 34308 16804 34372
rect 16868 34308 16869 34372
rect 16803 34307 16869 34308
rect 16067 33692 16133 33693
rect 16067 33628 16068 33692
rect 16132 33628 16133 33692
rect 16067 33627 16133 33628
rect 16070 31653 16130 33627
rect 16067 31652 16133 31653
rect 16067 31588 16068 31652
rect 16132 31588 16133 31652
rect 16067 31587 16133 31588
rect 16806 29205 16866 34307
rect 16803 29204 16869 29205
rect 16803 29140 16804 29204
rect 16868 29140 16869 29204
rect 16803 29139 16869 29140
rect 16619 28524 16685 28525
rect 16619 28460 16620 28524
rect 16684 28460 16685 28524
rect 16619 28459 16685 28460
rect 16622 23765 16682 28459
rect 17174 27165 17234 37707
rect 19568 37568 19888 38592
rect 19568 37504 19576 37568
rect 19640 37504 19656 37568
rect 19720 37504 19736 37568
rect 19800 37504 19816 37568
rect 19880 37504 19888 37568
rect 19568 36480 19888 37504
rect 19568 36416 19576 36480
rect 19640 36416 19656 36480
rect 19720 36416 19736 36480
rect 19800 36416 19816 36480
rect 19880 36416 19888 36480
rect 19568 35392 19888 36416
rect 19568 35328 19576 35392
rect 19640 35328 19656 35392
rect 19720 35328 19736 35392
rect 19800 35328 19816 35392
rect 19880 35328 19888 35392
rect 19568 34304 19888 35328
rect 19568 34240 19576 34304
rect 19640 34240 19656 34304
rect 19720 34240 19736 34304
rect 19800 34240 19816 34304
rect 19880 34240 19888 34304
rect 19568 33216 19888 34240
rect 20115 34236 20181 34237
rect 20115 34172 20116 34236
rect 20180 34172 20181 34236
rect 20115 34171 20181 34172
rect 19568 33152 19576 33216
rect 19640 33152 19656 33216
rect 19720 33152 19736 33216
rect 19800 33152 19816 33216
rect 19880 33152 19888 33216
rect 19568 32128 19888 33152
rect 19568 32064 19576 32128
rect 19640 32064 19656 32128
rect 19720 32064 19736 32128
rect 19800 32064 19816 32128
rect 19880 32064 19888 32128
rect 19568 31040 19888 32064
rect 19568 30976 19576 31040
rect 19640 30976 19656 31040
rect 19720 30976 19736 31040
rect 19800 30976 19816 31040
rect 19880 30976 19888 31040
rect 19568 29952 19888 30976
rect 19568 29888 19576 29952
rect 19640 29888 19656 29952
rect 19720 29888 19736 29952
rect 19800 29888 19816 29952
rect 19880 29888 19888 29952
rect 19568 28864 19888 29888
rect 19568 28800 19576 28864
rect 19640 28800 19656 28864
rect 19720 28800 19736 28864
rect 19800 28800 19816 28864
rect 19880 28800 19888 28864
rect 19568 27776 19888 28800
rect 20118 28661 20178 34171
rect 20115 28660 20181 28661
rect 20115 28596 20116 28660
rect 20180 28596 20181 28660
rect 20115 28595 20181 28596
rect 19568 27712 19576 27776
rect 19640 27712 19656 27776
rect 19720 27712 19736 27776
rect 19800 27712 19816 27776
rect 19880 27712 19888 27776
rect 17171 27164 17237 27165
rect 17171 27100 17172 27164
rect 17236 27100 17237 27164
rect 17171 27099 17237 27100
rect 19568 26688 19888 27712
rect 19568 26624 19576 26688
rect 19640 26624 19656 26688
rect 19720 26624 19736 26688
rect 19800 26624 19816 26688
rect 19880 26624 19888 26688
rect 19568 25600 19888 26624
rect 19568 25536 19576 25600
rect 19640 25536 19656 25600
rect 19720 25536 19736 25600
rect 19800 25536 19816 25600
rect 19880 25536 19888 25600
rect 19568 24512 19888 25536
rect 19568 24448 19576 24512
rect 19640 24448 19656 24512
rect 19720 24448 19736 24512
rect 19800 24448 19816 24512
rect 19880 24448 19888 24512
rect 16619 23764 16685 23765
rect 16619 23700 16620 23764
rect 16684 23700 16685 23764
rect 16619 23699 16685 23700
rect 16622 23578 16682 23699
rect 19568 23424 19888 24448
rect 19568 23360 19576 23424
rect 19640 23360 19656 23424
rect 19720 23360 19736 23424
rect 19800 23360 19816 23424
rect 19880 23360 19888 23424
rect 19568 22336 19888 23360
rect 19568 22272 19576 22336
rect 19640 22272 19656 22336
rect 19720 22272 19736 22336
rect 19800 22272 19816 22336
rect 19880 22272 19888 22336
rect 19568 21248 19888 22272
rect 19568 21184 19576 21248
rect 19640 21184 19656 21248
rect 19720 21184 19736 21248
rect 19800 21184 19816 21248
rect 19880 21184 19888 21248
rect 19568 20894 19888 21184
rect 15883 20772 15949 20773
rect 15883 20708 15884 20772
rect 15948 20708 15949 20772
rect 15883 20707 15949 20708
rect 19568 20658 19610 20894
rect 19846 20658 19888 20894
rect 19568 20160 19888 20658
rect 19568 20096 19576 20160
rect 19640 20096 19656 20160
rect 19720 20096 19736 20160
rect 19800 20096 19816 20160
rect 19880 20096 19888 20160
rect 19568 19072 19888 20096
rect 19568 19008 19576 19072
rect 19640 19008 19656 19072
rect 19720 19008 19736 19072
rect 19800 19008 19816 19072
rect 19880 19008 19888 19072
rect 19568 17984 19888 19008
rect 19568 17920 19576 17984
rect 19640 17920 19656 17984
rect 19720 17920 19736 17984
rect 19800 17920 19816 17984
rect 19880 17920 19888 17984
rect 19568 16896 19888 17920
rect 19568 16832 19576 16896
rect 19640 16832 19656 16896
rect 19720 16832 19736 16896
rect 19800 16832 19816 16896
rect 19880 16832 19888 16896
rect 19568 15808 19888 16832
rect 19568 15744 19576 15808
rect 19640 15744 19656 15808
rect 19720 15744 19736 15808
rect 19800 15744 19816 15808
rect 19880 15744 19888 15808
rect 19568 14720 19888 15744
rect 19568 14656 19576 14720
rect 19640 14656 19656 14720
rect 19720 14656 19736 14720
rect 19800 14656 19816 14720
rect 19880 14656 19888 14720
rect 19568 13632 19888 14656
rect 19568 13568 19576 13632
rect 19640 13568 19656 13632
rect 19720 13568 19736 13632
rect 19800 13568 19816 13632
rect 19880 13568 19888 13632
rect 19568 12544 19888 13568
rect 19568 12480 19576 12544
rect 19640 12480 19656 12544
rect 19720 12480 19736 12544
rect 19800 12480 19816 12544
rect 19880 12480 19888 12544
rect 15699 12476 15765 12477
rect 15699 12412 15700 12476
rect 15764 12412 15765 12476
rect 15699 12411 15765 12412
rect 19568 11456 19888 12480
rect 19568 11392 19576 11456
rect 19640 11392 19656 11456
rect 19720 11392 19736 11456
rect 19800 11392 19816 11456
rect 19880 11392 19888 11456
rect 19568 10368 19888 11392
rect 19568 10304 19576 10368
rect 19640 10304 19656 10368
rect 19720 10304 19736 10368
rect 19800 10304 19816 10368
rect 19880 10304 19888 10368
rect 19568 9280 19888 10304
rect 19568 9216 19576 9280
rect 19640 9216 19656 9280
rect 19720 9216 19736 9280
rect 19800 9216 19816 9280
rect 19880 9216 19888 9280
rect 19568 8192 19888 9216
rect 19568 8128 19576 8192
rect 19640 8128 19656 8192
rect 19720 8128 19736 8192
rect 19800 8128 19816 8192
rect 19880 8128 19888 8192
rect 19568 7104 19888 8128
rect 20302 7581 20362 46955
rect 20851 46476 20917 46477
rect 20851 46412 20852 46476
rect 20916 46412 20917 46476
rect 20851 46411 20917 46412
rect 20667 34372 20733 34373
rect 20667 34308 20668 34372
rect 20732 34308 20733 34372
rect 20667 34307 20733 34308
rect 20483 28252 20549 28253
rect 20483 28188 20484 28252
rect 20548 28188 20549 28252
rect 20483 28187 20549 28188
rect 20486 17917 20546 28187
rect 20670 27981 20730 34307
rect 20667 27980 20733 27981
rect 20667 27916 20668 27980
rect 20732 27916 20733 27980
rect 20667 27915 20733 27916
rect 20483 17916 20549 17917
rect 20483 17852 20484 17916
rect 20548 17852 20549 17916
rect 20483 17851 20549 17852
rect 20854 15605 20914 46411
rect 21038 17917 21098 71843
rect 34928 71840 35248 72864
rect 34928 71776 34936 71840
rect 35000 71776 35016 71840
rect 35080 71776 35096 71840
rect 35160 71776 35176 71840
rect 35240 71776 35248 71840
rect 34928 70752 35248 71776
rect 34928 70688 34936 70752
rect 35000 70688 35016 70752
rect 35080 70688 35096 70752
rect 35160 70688 35176 70752
rect 35240 70688 35248 70752
rect 34928 69664 35248 70688
rect 34928 69600 34936 69664
rect 35000 69600 35016 69664
rect 35080 69600 35096 69664
rect 35160 69600 35176 69664
rect 35240 69600 35248 69664
rect 30051 69052 30117 69053
rect 30051 68988 30052 69052
rect 30116 68988 30117 69052
rect 30051 68987 30117 68988
rect 28947 68372 29013 68373
rect 28947 68308 28948 68372
rect 29012 68308 29013 68372
rect 28947 68307 29013 68308
rect 28950 67965 29010 68307
rect 28947 67964 29013 67965
rect 28947 67900 28948 67964
rect 29012 67900 29013 67964
rect 28947 67899 29013 67900
rect 28395 67148 28461 67149
rect 28395 67084 28396 67148
rect 28460 67084 28461 67148
rect 28395 67083 28461 67084
rect 22507 62796 22573 62797
rect 22507 62732 22508 62796
rect 22572 62732 22573 62796
rect 22507 62731 22573 62732
rect 21771 54092 21837 54093
rect 21771 54028 21772 54092
rect 21836 54028 21837 54092
rect 21771 54027 21837 54028
rect 21774 50829 21834 54027
rect 21771 50828 21837 50829
rect 21771 50764 21772 50828
rect 21836 50764 21837 50828
rect 21771 50763 21837 50764
rect 21219 49740 21285 49741
rect 21219 49676 21220 49740
rect 21284 49676 21285 49740
rect 21219 49675 21285 49676
rect 21035 17916 21101 17917
rect 21035 17852 21036 17916
rect 21100 17852 21101 17916
rect 21035 17851 21101 17852
rect 21222 16557 21282 49675
rect 21587 31380 21653 31381
rect 21587 31316 21588 31380
rect 21652 31316 21653 31380
rect 21587 31315 21653 31316
rect 21403 27844 21469 27845
rect 21403 27780 21404 27844
rect 21468 27780 21469 27844
rect 21403 27779 21469 27780
rect 21406 24173 21466 27779
rect 21590 24581 21650 31315
rect 22142 30429 22202 30822
rect 21955 30428 22021 30429
rect 21955 30364 21956 30428
rect 22020 30364 22021 30428
rect 21955 30363 22021 30364
rect 22139 30428 22205 30429
rect 22139 30364 22140 30428
rect 22204 30364 22205 30428
rect 22139 30363 22205 30364
rect 21958 28930 22018 30363
rect 22323 29204 22389 29205
rect 22323 29140 22324 29204
rect 22388 29140 22389 29204
rect 22323 29139 22389 29140
rect 21958 28870 22202 28930
rect 21771 28524 21837 28525
rect 21771 28460 21772 28524
rect 21836 28460 21837 28524
rect 21771 28459 21837 28460
rect 21774 27570 21834 28459
rect 21958 28253 22018 28870
rect 22142 28797 22202 28870
rect 22139 28796 22205 28797
rect 22139 28732 22140 28796
rect 22204 28732 22205 28796
rect 22139 28731 22205 28732
rect 21955 28252 22021 28253
rect 21955 28188 21956 28252
rect 22020 28188 22021 28252
rect 21955 28187 22021 28188
rect 22326 27573 22386 29139
rect 22323 27572 22389 27573
rect 21774 27510 22202 27570
rect 21587 24580 21653 24581
rect 21587 24516 21588 24580
rect 21652 24516 21653 24580
rect 21587 24515 21653 24516
rect 21403 24172 21469 24173
rect 21403 24108 21404 24172
rect 21468 24108 21469 24172
rect 21403 24107 21469 24108
rect 21958 23629 22018 27510
rect 22142 27301 22202 27510
rect 22323 27508 22324 27572
rect 22388 27508 22389 27572
rect 22323 27507 22389 27508
rect 22139 27300 22205 27301
rect 22139 27236 22140 27300
rect 22204 27236 22205 27300
rect 22139 27235 22205 27236
rect 21955 23628 22021 23629
rect 21955 23564 21956 23628
rect 22020 23564 22021 23628
rect 21955 23563 22021 23564
rect 21219 16556 21285 16557
rect 21219 16492 21220 16556
rect 21284 16492 21285 16556
rect 21219 16491 21285 16492
rect 20851 15604 20917 15605
rect 20851 15540 20852 15604
rect 20916 15540 20917 15604
rect 20851 15539 20917 15540
rect 22510 15197 22570 62731
rect 28027 62252 28093 62253
rect 28027 62188 28028 62252
rect 28092 62188 28093 62252
rect 28027 62187 28093 62188
rect 24715 54228 24781 54229
rect 24715 54164 24716 54228
rect 24780 54164 24781 54228
rect 24715 54163 24781 54164
rect 24531 53956 24597 53957
rect 24531 53892 24532 53956
rect 24596 53892 24597 53956
rect 24531 53891 24597 53892
rect 24347 37364 24413 37365
rect 24347 37300 24348 37364
rect 24412 37300 24413 37364
rect 24347 37299 24413 37300
rect 23246 36277 23306 36942
rect 23243 36276 23309 36277
rect 23243 36212 23244 36276
rect 23308 36212 23309 36276
rect 23243 36211 23309 36212
rect 23795 32196 23861 32197
rect 23246 31653 23306 32182
rect 23795 32132 23796 32196
rect 23860 32132 23861 32196
rect 23795 32131 23861 32132
rect 23243 31652 23309 31653
rect 23243 31588 23244 31652
rect 23308 31588 23309 31652
rect 23243 31587 23309 31588
rect 22875 30020 22941 30021
rect 22875 29956 22876 30020
rect 22940 29956 22941 30020
rect 22875 29955 22941 29956
rect 22878 25397 22938 29955
rect 23798 28797 23858 32131
rect 23795 28796 23861 28797
rect 23795 28732 23796 28796
rect 23860 28732 23861 28796
rect 23795 28731 23861 28732
rect 23243 27164 23309 27165
rect 23243 27100 23244 27164
rect 23308 27100 23309 27164
rect 23243 27099 23309 27100
rect 22875 25396 22941 25397
rect 22875 25332 22876 25396
rect 22940 25332 22941 25396
rect 22875 25331 22941 25332
rect 23246 25125 23306 27099
rect 23243 25124 23309 25125
rect 23243 25060 23244 25124
rect 23308 25060 23309 25124
rect 23243 25059 23309 25060
rect 23246 23221 23306 23342
rect 23243 23220 23309 23221
rect 23243 23156 23244 23220
rect 23308 23156 23309 23220
rect 23243 23155 23309 23156
rect 22507 15196 22573 15197
rect 22507 15132 22508 15196
rect 22572 15132 22573 15196
rect 22507 15131 22573 15132
rect 24350 9757 24410 37299
rect 24534 15197 24594 53891
rect 24718 19957 24778 54163
rect 27843 51372 27909 51373
rect 27843 51308 27844 51372
rect 27908 51308 27909 51372
rect 27843 51307 27909 51308
rect 27846 42669 27906 51307
rect 27843 42668 27909 42669
rect 27843 42604 27844 42668
rect 27908 42604 27909 42668
rect 27843 42603 27909 42604
rect 28030 38453 28090 62187
rect 28211 47020 28277 47021
rect 28211 46956 28212 47020
rect 28276 46956 28277 47020
rect 28211 46955 28277 46956
rect 28214 41853 28274 46955
rect 28211 41852 28277 41853
rect 28211 41788 28212 41852
rect 28276 41788 28277 41852
rect 28211 41787 28277 41788
rect 28027 38452 28093 38453
rect 28027 38388 28028 38452
rect 28092 38388 28093 38452
rect 28027 38387 28093 38388
rect 27843 38044 27909 38045
rect 27843 37980 27844 38044
rect 27908 37980 27909 38044
rect 27843 37979 27909 37980
rect 27846 30157 27906 37979
rect 27843 30156 27909 30157
rect 27843 30092 27844 30156
rect 27908 30092 27909 30156
rect 27843 30091 27909 30092
rect 24715 19956 24781 19957
rect 24715 19892 24716 19956
rect 24780 19892 24781 19956
rect 24715 19891 24781 19892
rect 24531 15196 24597 15197
rect 24531 15132 24532 15196
rect 24596 15132 24597 15196
rect 24531 15131 24597 15132
rect 24347 9756 24413 9757
rect 24347 9692 24348 9756
rect 24412 9692 24413 9756
rect 24347 9691 24413 9692
rect 20299 7580 20365 7581
rect 20299 7516 20300 7580
rect 20364 7516 20365 7580
rect 20299 7515 20365 7516
rect 19568 7040 19576 7104
rect 19640 7040 19656 7104
rect 19720 7040 19736 7104
rect 19800 7040 19816 7104
rect 19880 7040 19888 7104
rect 19568 6016 19888 7040
rect 19568 5952 19576 6016
rect 19640 5952 19656 6016
rect 19720 5952 19736 6016
rect 19800 5952 19816 6016
rect 19880 5952 19888 6016
rect 19568 4928 19888 5952
rect 19568 4864 19576 4928
rect 19640 4864 19656 4928
rect 19720 4864 19736 4928
rect 19800 4864 19816 4928
rect 19880 4864 19888 4928
rect 17907 4588 17973 4589
rect 17907 4524 17908 4588
rect 17972 4524 17973 4588
rect 17907 4523 17973 4524
rect 17910 4317 17970 4523
rect 17907 4316 17973 4317
rect 17907 4252 17908 4316
rect 17972 4252 17973 4316
rect 17907 4251 17973 4252
rect 14227 4044 14293 4045
rect 14227 3980 14228 4044
rect 14292 3980 14293 4044
rect 14227 3979 14293 3980
rect 4208 3232 4216 3296
rect 4280 3232 4296 3296
rect 4360 3232 4376 3296
rect 4440 3232 4456 3296
rect 4520 3232 4528 3296
rect 4208 2208 4528 3232
rect 4208 2144 4216 2208
rect 4280 2144 4296 2208
rect 4360 2144 4376 2208
rect 4440 2144 4456 2208
rect 4520 2144 4528 2208
rect 4208 2128 4528 2144
rect 19568 3840 19888 4864
rect 19568 3776 19576 3840
rect 19640 3776 19656 3840
rect 19720 3776 19736 3840
rect 19800 3776 19816 3840
rect 19880 3776 19888 3840
rect 19568 2752 19888 3776
rect 19568 2688 19576 2752
rect 19640 2688 19656 2752
rect 19720 2688 19736 2752
rect 19800 2688 19816 2752
rect 19880 2688 19888 2752
rect 19568 2128 19888 2688
rect 28398 2685 28458 67083
rect 28579 51236 28645 51237
rect 28579 51172 28580 51236
rect 28644 51172 28645 51236
rect 28579 51171 28645 51172
rect 29131 51236 29197 51237
rect 29131 51172 29132 51236
rect 29196 51172 29197 51236
rect 29131 51171 29197 51172
rect 28582 43893 28642 51171
rect 29134 49469 29194 51171
rect 29131 49468 29197 49469
rect 29131 49404 29132 49468
rect 29196 49404 29197 49468
rect 29131 49403 29197 49404
rect 30054 48245 30114 68987
rect 34928 68576 35248 69600
rect 34928 68512 34936 68576
rect 35000 68512 35016 68576
rect 35080 68512 35096 68576
rect 35160 68512 35176 68576
rect 35240 68512 35248 68576
rect 34928 67488 35248 68512
rect 34928 67424 34936 67488
rect 35000 67424 35016 67488
rect 35080 67424 35096 67488
rect 35160 67424 35176 67488
rect 35240 67424 35248 67488
rect 34928 66848 35248 67424
rect 34928 66612 34970 66848
rect 35206 66612 35248 66848
rect 34928 66400 35248 66612
rect 34928 66336 34936 66400
rect 35000 66336 35016 66400
rect 35080 66336 35096 66400
rect 35160 66336 35176 66400
rect 35240 66336 35248 66400
rect 34928 65312 35248 66336
rect 34928 65248 34936 65312
rect 35000 65248 35016 65312
rect 35080 65248 35096 65312
rect 35160 65248 35176 65312
rect 35240 65248 35248 65312
rect 34928 64224 35248 65248
rect 34928 64160 34936 64224
rect 35000 64160 35016 64224
rect 35080 64160 35096 64224
rect 35160 64160 35176 64224
rect 35240 64160 35248 64224
rect 34928 63136 35248 64160
rect 34928 63072 34936 63136
rect 35000 63072 35016 63136
rect 35080 63072 35096 63136
rect 35160 63072 35176 63136
rect 35240 63072 35248 63136
rect 34928 62048 35248 63072
rect 34928 61984 34936 62048
rect 35000 61984 35016 62048
rect 35080 61984 35096 62048
rect 35160 61984 35176 62048
rect 35240 61984 35248 62048
rect 34928 60960 35248 61984
rect 34928 60896 34936 60960
rect 35000 60896 35016 60960
rect 35080 60896 35096 60960
rect 35160 60896 35176 60960
rect 35240 60896 35248 60960
rect 34928 59872 35248 60896
rect 34928 59808 34936 59872
rect 35000 59808 35016 59872
rect 35080 59808 35096 59872
rect 35160 59808 35176 59872
rect 35240 59808 35248 59872
rect 34928 58784 35248 59808
rect 34928 58720 34936 58784
rect 35000 58720 35016 58784
rect 35080 58720 35096 58784
rect 35160 58720 35176 58784
rect 35240 58720 35248 58784
rect 34928 57696 35248 58720
rect 34928 57632 34936 57696
rect 35000 57632 35016 57696
rect 35080 57632 35096 57696
rect 35160 57632 35176 57696
rect 35240 57632 35248 57696
rect 34928 56608 35248 57632
rect 34928 56544 34936 56608
rect 35000 56544 35016 56608
rect 35080 56544 35096 56608
rect 35160 56544 35176 56608
rect 35240 56544 35248 56608
rect 34928 55520 35248 56544
rect 34928 55456 34936 55520
rect 35000 55456 35016 55520
rect 35080 55456 35096 55520
rect 35160 55456 35176 55520
rect 35240 55456 35248 55520
rect 34928 54432 35248 55456
rect 34928 54368 34936 54432
rect 35000 54368 35016 54432
rect 35080 54368 35096 54432
rect 35160 54368 35176 54432
rect 35240 54368 35248 54432
rect 34928 53344 35248 54368
rect 34928 53280 34936 53344
rect 35000 53280 35016 53344
rect 35080 53280 35096 53344
rect 35160 53280 35176 53344
rect 35240 53280 35248 53344
rect 34928 52256 35248 53280
rect 34928 52192 34936 52256
rect 35000 52192 35016 52256
rect 35080 52192 35096 52256
rect 35160 52192 35176 52256
rect 35240 52192 35248 52256
rect 34928 51168 35248 52192
rect 34928 51104 34936 51168
rect 35000 51104 35016 51168
rect 35080 51104 35096 51168
rect 35160 51104 35176 51168
rect 35240 51104 35248 51168
rect 34928 50080 35248 51104
rect 34928 50016 34936 50080
rect 35000 50016 35016 50080
rect 35080 50016 35096 50080
rect 35160 50016 35176 50080
rect 35240 50016 35248 50080
rect 34928 48992 35248 50016
rect 34928 48928 34936 48992
rect 35000 48928 35016 48992
rect 35080 48928 35096 48992
rect 35160 48928 35176 48992
rect 35240 48928 35248 48992
rect 29683 48244 29749 48245
rect 29683 48180 29684 48244
rect 29748 48180 29749 48244
rect 29683 48179 29749 48180
rect 30051 48244 30117 48245
rect 30051 48180 30052 48244
rect 30116 48180 30117 48244
rect 30051 48179 30117 48180
rect 28947 46204 29013 46205
rect 28947 46140 28948 46204
rect 29012 46140 29013 46204
rect 28947 46139 29013 46140
rect 28950 45797 29010 46139
rect 28947 45796 29013 45797
rect 28947 45732 28948 45796
rect 29012 45732 29013 45796
rect 28947 45731 29013 45732
rect 28579 43892 28645 43893
rect 28579 43828 28580 43892
rect 28644 43828 28645 43892
rect 28579 43827 28645 43828
rect 29686 41309 29746 48179
rect 34928 47904 35248 48928
rect 34928 47840 34936 47904
rect 35000 47840 35016 47904
rect 35080 47840 35096 47904
rect 35160 47840 35176 47904
rect 35240 47840 35248 47904
rect 34928 46816 35248 47840
rect 34928 46752 34936 46816
rect 35000 46752 35016 46816
rect 35080 46752 35096 46816
rect 35160 46752 35176 46816
rect 35240 46752 35248 46816
rect 34928 45728 35248 46752
rect 34928 45664 34936 45728
rect 35000 45664 35016 45728
rect 35080 45664 35096 45728
rect 35160 45664 35176 45728
rect 35240 45664 35248 45728
rect 34928 44640 35248 45664
rect 34928 44576 34936 44640
rect 35000 44576 35016 44640
rect 35080 44576 35096 44640
rect 35160 44576 35176 44640
rect 35240 44576 35248 44640
rect 34928 43552 35248 44576
rect 34928 43488 34936 43552
rect 35000 43488 35016 43552
rect 35080 43488 35096 43552
rect 35160 43488 35176 43552
rect 35240 43488 35248 43552
rect 34928 42464 35248 43488
rect 34928 42400 34936 42464
rect 35000 42400 35016 42464
rect 35080 42400 35096 42464
rect 35160 42400 35176 42464
rect 35240 42400 35248 42464
rect 34928 41376 35248 42400
rect 34928 41312 34936 41376
rect 35000 41312 35016 41376
rect 35080 41312 35096 41376
rect 35160 41312 35176 41376
rect 35240 41312 35248 41376
rect 29683 41308 29749 41309
rect 29683 41244 29684 41308
rect 29748 41244 29749 41308
rect 29683 41243 29749 41244
rect 34928 40288 35248 41312
rect 34928 40224 34936 40288
rect 35000 40224 35016 40288
rect 35080 40224 35096 40288
rect 35160 40224 35176 40288
rect 35240 40224 35248 40288
rect 34928 39200 35248 40224
rect 34928 39136 34936 39200
rect 35000 39136 35016 39200
rect 35080 39136 35096 39200
rect 35160 39136 35176 39200
rect 35240 39136 35248 39200
rect 34928 38112 35248 39136
rect 34928 38048 34936 38112
rect 35000 38048 35016 38112
rect 35080 38048 35096 38112
rect 35160 38048 35176 38112
rect 35240 38048 35248 38112
rect 34928 37024 35248 38048
rect 34928 36960 34936 37024
rect 35000 36960 35016 37024
rect 35080 36960 35096 37024
rect 35160 36960 35176 37024
rect 35240 36960 35248 37024
rect 34928 36212 35248 36960
rect 34928 35976 34970 36212
rect 35206 35976 35248 36212
rect 34928 35936 35248 35976
rect 34928 35872 34936 35936
rect 35000 35872 35016 35936
rect 35080 35872 35096 35936
rect 35160 35872 35176 35936
rect 35240 35872 35248 35936
rect 34928 34848 35248 35872
rect 34928 34784 34936 34848
rect 35000 34784 35016 34848
rect 35080 34784 35096 34848
rect 35160 34784 35176 34848
rect 35240 34784 35248 34848
rect 34928 33760 35248 34784
rect 34928 33696 34936 33760
rect 35000 33696 35016 33760
rect 35080 33696 35096 33760
rect 35160 33696 35176 33760
rect 35240 33696 35248 33760
rect 34928 32672 35248 33696
rect 34928 32608 34936 32672
rect 35000 32608 35016 32672
rect 35080 32608 35096 32672
rect 35160 32608 35176 32672
rect 35240 32608 35248 32672
rect 34928 31584 35248 32608
rect 34928 31520 34936 31584
rect 35000 31520 35016 31584
rect 35080 31520 35096 31584
rect 35160 31520 35176 31584
rect 35240 31520 35248 31584
rect 34928 30496 35248 31520
rect 34928 30432 34936 30496
rect 35000 30432 35016 30496
rect 35080 30432 35096 30496
rect 35160 30432 35176 30496
rect 35240 30432 35248 30496
rect 34928 29408 35248 30432
rect 34928 29344 34936 29408
rect 35000 29344 35016 29408
rect 35080 29344 35096 29408
rect 35160 29344 35176 29408
rect 35240 29344 35248 29408
rect 34928 28320 35248 29344
rect 35571 29340 35637 29341
rect 35571 29276 35572 29340
rect 35636 29276 35637 29340
rect 35571 29275 35637 29276
rect 34928 28256 34936 28320
rect 35000 28256 35016 28320
rect 35080 28256 35096 28320
rect 35160 28256 35176 28320
rect 35240 28256 35248 28320
rect 34470 26621 34530 28102
rect 34928 27232 35248 28256
rect 34928 27168 34936 27232
rect 35000 27168 35016 27232
rect 35080 27168 35096 27232
rect 35160 27168 35176 27232
rect 35240 27168 35248 27232
rect 34467 26620 34533 26621
rect 34467 26556 34468 26620
rect 34532 26556 34533 26620
rect 34467 26555 34533 26556
rect 34928 26144 35248 27168
rect 34928 26080 34936 26144
rect 35000 26080 35016 26144
rect 35080 26080 35096 26144
rect 35160 26080 35176 26144
rect 35240 26080 35248 26144
rect 34470 25261 34530 26062
rect 34467 25260 34533 25261
rect 34467 25196 34468 25260
rect 34532 25196 34533 25260
rect 34467 25195 34533 25196
rect 34928 25056 35248 26080
rect 34928 24992 34936 25056
rect 35000 24992 35016 25056
rect 35080 24992 35096 25056
rect 35160 24992 35176 25056
rect 35240 24992 35248 25056
rect 34928 23968 35248 24992
rect 34928 23904 34936 23968
rect 35000 23904 35016 23968
rect 35080 23904 35096 23968
rect 35160 23904 35176 23968
rect 35240 23904 35248 23968
rect 34928 22880 35248 23904
rect 34928 22816 34936 22880
rect 35000 22816 35016 22880
rect 35080 22816 35096 22880
rect 35160 22816 35176 22880
rect 35240 22816 35248 22880
rect 34928 21792 35248 22816
rect 34928 21728 34936 21792
rect 35000 21728 35016 21792
rect 35080 21728 35096 21792
rect 35160 21728 35176 21792
rect 35240 21728 35248 21792
rect 34928 20704 35248 21728
rect 35574 21538 35634 29275
rect 34928 20640 34936 20704
rect 35000 20640 35016 20704
rect 35080 20640 35096 20704
rect 35160 20640 35176 20704
rect 35240 20640 35248 20704
rect 34928 19616 35248 20640
rect 34928 19552 34936 19616
rect 35000 19552 35016 19616
rect 35080 19552 35096 19616
rect 35160 19552 35176 19616
rect 35240 19552 35248 19616
rect 34928 18528 35248 19552
rect 34928 18464 34936 18528
rect 35000 18464 35016 18528
rect 35080 18464 35096 18528
rect 35160 18464 35176 18528
rect 35240 18464 35248 18528
rect 34928 17440 35248 18464
rect 34928 17376 34936 17440
rect 35000 17376 35016 17440
rect 35080 17376 35096 17440
rect 35160 17376 35176 17440
rect 35240 17376 35248 17440
rect 34928 16352 35248 17376
rect 34928 16288 34936 16352
rect 35000 16288 35016 16352
rect 35080 16288 35096 16352
rect 35160 16288 35176 16352
rect 35240 16288 35248 16352
rect 34928 15264 35248 16288
rect 34928 15200 34936 15264
rect 35000 15200 35016 15264
rect 35080 15200 35096 15264
rect 35160 15200 35176 15264
rect 35240 15200 35248 15264
rect 34928 14176 35248 15200
rect 34928 14112 34936 14176
rect 35000 14112 35016 14176
rect 35080 14112 35096 14176
rect 35160 14112 35176 14176
rect 35240 14112 35248 14176
rect 34928 13088 35248 14112
rect 34928 13024 34936 13088
rect 35000 13024 35016 13088
rect 35080 13024 35096 13088
rect 35160 13024 35176 13088
rect 35240 13024 35248 13088
rect 28947 12204 29013 12205
rect 28947 12140 28948 12204
rect 29012 12140 29013 12204
rect 28947 12139 29013 12140
rect 28950 11253 29010 12139
rect 34928 12000 35248 13024
rect 34928 11936 34936 12000
rect 35000 11936 35016 12000
rect 35080 11936 35096 12000
rect 35160 11936 35176 12000
rect 35240 11936 35248 12000
rect 28947 11252 29013 11253
rect 28947 11188 28948 11252
rect 29012 11188 29013 11252
rect 28947 11187 29013 11188
rect 34928 10912 35248 11936
rect 34928 10848 34936 10912
rect 35000 10848 35016 10912
rect 35080 10848 35096 10912
rect 35160 10848 35176 10912
rect 35240 10848 35248 10912
rect 34928 9824 35248 10848
rect 34928 9760 34936 9824
rect 35000 9760 35016 9824
rect 35080 9760 35096 9824
rect 35160 9760 35176 9824
rect 35240 9760 35248 9824
rect 30419 9620 30485 9621
rect 30419 9556 30420 9620
rect 30484 9556 30485 9620
rect 30419 9555 30485 9556
rect 28947 4860 29013 4861
rect 28947 4796 28948 4860
rect 29012 4796 29013 4860
rect 28947 4795 29013 4796
rect 28950 4317 29010 4795
rect 28947 4316 29013 4317
rect 28947 4252 28948 4316
rect 29012 4252 29013 4316
rect 28947 4251 29013 4252
rect 28395 2684 28461 2685
rect 28395 2620 28396 2684
rect 28460 2620 28461 2684
rect 28395 2619 28461 2620
rect 30422 917 30482 9555
rect 34928 8736 35248 9760
rect 34928 8672 34936 8736
rect 35000 8672 35016 8736
rect 35080 8672 35096 8736
rect 35160 8672 35176 8736
rect 35240 8672 35248 8736
rect 34928 7648 35248 8672
rect 34928 7584 34936 7648
rect 35000 7584 35016 7648
rect 35080 7584 35096 7648
rect 35160 7584 35176 7648
rect 35240 7584 35248 7648
rect 34928 6560 35248 7584
rect 34928 6496 34936 6560
rect 35000 6496 35016 6560
rect 35080 6496 35096 6560
rect 35160 6496 35176 6560
rect 35240 6496 35248 6560
rect 34928 5576 35248 6496
rect 34928 5472 34970 5576
rect 35206 5472 35248 5576
rect 34928 5408 34936 5472
rect 35240 5408 35248 5472
rect 34928 5340 34970 5408
rect 35206 5340 35248 5408
rect 34928 4384 35248 5340
rect 34928 4320 34936 4384
rect 35000 4320 35016 4384
rect 35080 4320 35096 4384
rect 35160 4320 35176 4384
rect 35240 4320 35248 4384
rect 34928 3296 35248 4320
rect 34928 3232 34936 3296
rect 35000 3232 35016 3296
rect 35080 3232 35096 3296
rect 35160 3232 35176 3296
rect 35240 3232 35248 3296
rect 34928 2208 35248 3232
rect 34928 2144 34936 2208
rect 35000 2144 35016 2208
rect 35080 2144 35096 2208
rect 35160 2144 35176 2208
rect 35240 2144 35248 2208
rect 34928 2128 35248 2144
rect 30419 916 30485 917
rect 30419 852 30420 916
rect 30484 852 30485 916
rect 30419 851 30485 852
<< via4 >>
rect 4250 66612 4486 66848
rect 9542 36942 9778 37178
rect 4250 35976 4486 36212
rect 12670 30292 12906 30378
rect 12670 30228 12756 30292
rect 12756 30228 12820 30292
rect 12820 30228 12906 30292
rect 12670 30142 12906 30228
rect 6598 26284 6684 26298
rect 6684 26284 6748 26298
rect 6748 26284 6834 26298
rect 6598 26062 6834 26284
rect 7150 21302 7386 21538
rect 4250 5472 4486 5576
rect 4250 5408 4280 5472
rect 4280 5408 4296 5472
rect 4296 5408 4360 5472
rect 4360 5408 4376 5472
rect 4376 5408 4440 5472
rect 4440 5408 4456 5472
rect 4456 5408 4486 5472
rect 4250 5340 4486 5408
rect 19610 51294 19846 51530
rect 15246 32404 15332 32418
rect 15332 32404 15396 32418
rect 15396 32404 15482 32418
rect 15246 32182 15482 32404
rect 16534 23342 16770 23578
rect 19610 20658 19846 20894
rect 22054 30822 22290 31058
rect 23158 36942 23394 37178
rect 23158 32332 23394 32418
rect 23158 32268 23244 32332
rect 23244 32268 23308 32332
rect 23308 32268 23394 32332
rect 23158 32182 23394 32268
rect 23894 28252 24130 28338
rect 23894 28188 23980 28252
rect 23980 28188 24044 28252
rect 24044 28188 24130 28252
rect 23894 28102 24130 28188
rect 23158 23342 23394 23578
rect 34970 66612 35206 66848
rect 34970 35976 35206 36212
rect 34382 28102 34618 28338
rect 34382 26062 34618 26298
rect 35486 21302 35722 21538
rect 34970 5472 35206 5576
rect 34970 5408 35000 5472
rect 35000 5408 35016 5472
rect 35016 5408 35080 5472
rect 35080 5408 35096 5472
rect 35096 5408 35160 5472
rect 35160 5408 35176 5472
rect 35176 5408 35206 5472
rect 34970 5340 35206 5408
<< metal5 >>
rect 1104 66848 38824 66890
rect 1104 66612 4250 66848
rect 4486 66612 34970 66848
rect 35206 66612 38824 66848
rect 1104 66570 38824 66612
rect 1104 51530 38824 51572
rect 1104 51294 19610 51530
rect 19846 51294 38824 51530
rect 1104 51252 38824 51294
rect 9500 37178 23436 37220
rect 9500 36942 9542 37178
rect 9778 36942 23158 37178
rect 23394 36942 23436 37178
rect 9500 36900 23436 36942
rect 1104 36212 38824 36254
rect 1104 35976 4250 36212
rect 4486 35976 34970 36212
rect 35206 35976 38824 36212
rect 1104 35934 38824 35976
rect 15204 32418 23436 32460
rect 15204 32182 15246 32418
rect 15482 32182 23158 32418
rect 23394 32182 23436 32418
rect 15204 32140 23436 32182
rect 15020 31058 22332 31100
rect 15020 30822 22054 31058
rect 22290 30822 22332 31058
rect 15020 30780 22332 30822
rect 15020 30420 15340 30780
rect 12628 30378 15340 30420
rect 12628 30142 12670 30378
rect 12906 30142 15340 30378
rect 12628 30100 15340 30142
rect 23852 28338 34660 28380
rect 23852 28102 23894 28338
rect 24130 28102 34382 28338
rect 34618 28102 34660 28338
rect 23852 28060 34660 28102
rect 6556 26298 34660 26340
rect 6556 26062 6598 26298
rect 6834 26062 34382 26298
rect 34618 26062 34660 26298
rect 6556 26020 34660 26062
rect 16492 23578 23436 23620
rect 16492 23342 16534 23578
rect 16770 23342 23158 23578
rect 23394 23342 23436 23578
rect 16492 23300 23436 23342
rect 7108 21538 35764 21580
rect 7108 21302 7150 21538
rect 7386 21302 35486 21538
rect 35722 21302 35764 21538
rect 7108 21260 35764 21302
rect 1104 20894 38824 20936
rect 1104 20658 19610 20894
rect 19846 20658 38824 20894
rect 1104 20616 38824 20658
rect 1104 5576 38824 5618
rect 1104 5340 4250 5576
rect 4486 5340 34970 5576
rect 35206 5340 38824 5576
rect 1104 5298 38824 5340
use sky130_fd_sc_hd__decap_3  PHY_0 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 1104 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606120350
transform 1 0 1104 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 1380 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1606120350
transform 1 0 2484 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1606120350
transform 1 0 1380 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_15
timestamp 1606120350
transform 1 0 2484 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 3956 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 3588 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1606120350
transform 1 0 4048 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1606120350
transform 1 0 5152 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1606120350
transform 1 0 3588 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1606120350
transform 1 0 4692 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1606120350
transform 1 0 6808 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1606120350
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 6256 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1606120350
transform 1 0 6900 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 5796 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 6532 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1606120350
transform 1 0 6808 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1606120350
transform 1 0 8004 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1606120350
transform 1 0 9108 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_74
timestamp 1606120350
transform 1 0 7912 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_86
timestamp 1606120350
transform 1 0 9016 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1606120350
transform 1 0 9660 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1606120350
transform 1 0 9752 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1606120350
transform 1 0 10856 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_98
timestamp 1606120350
transform 1 0 10120 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_110
timestamp 1606120350
transform 1 0 11224 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_123
timestamp 1606120350
transform 1 0 12420 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_1_118
timestamp 1606120350
transform 1 0 11960 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_120
timestamp 1606120350
transform 1 0 12144 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__CLK /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 12144 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__CLK
timestamp 1606120350
transform 1 0 11960 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1125__D
timestamp 1606120350
transform 1 0 12328 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1606120350
transform 1 0 12328 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1606120350
transform 1 0 12512 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_132 /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 13248 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_128
timestamp 1606120350
transform 1 0 12880 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__D
timestamp 1606120350
transform 1 0 13340 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1131__D
timestamp 1606120350
transform 1 0 12696 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1143_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 13524 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1125_
timestamp 1606120350
transform 1 0 12604 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1606120350
transform 1 0 15364 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_144
timestamp 1606120350
transform 1 0 14352 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_152
timestamp 1606120350
transform 1 0 15088 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1606120350
transform 1 0 15456 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_154
timestamp 1606120350
transform 1 0 15272 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__CLK
timestamp 1606120350
transform 1 0 17664 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1606120350
transform 1 0 16560 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_182
timestamp 1606120350
transform 1 0 17848 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_166
timestamp 1606120350
transform 1 0 16376 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_178
timestamp 1606120350
transform 1 0 17480 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_182
timestamp 1606120350
transform 1 0 17848 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1215_
timestamp 1606120350
transform 1 0 18584 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1606120350
transform 1 0 18216 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1606120350
transform 1 0 17940 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1215__D
timestamp 1606120350
transform 1 0 18032 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_187
timestamp 1606120350
transform 1 0 18308 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1606120350
transform 1 0 18032 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1606120350
transform 1 0 19136 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1227_
timestamp 1606120350
transform 1 0 20700 0 1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1606120350
transform 1 0 21068 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__D
timestamp 1606120350
transform 1 0 20516 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1227__CLK
timestamp 1606120350
transform 1 0 20700 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_209
timestamp 1606120350
transform 1 0 20332 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_215
timestamp 1606120350
transform 1 0 20884 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1606120350
transform 1 0 21160 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_208
timestamp 1606120350
transform 1 0 20240 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1606120350
transform 1 0 23920 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1606120350
transform 1 0 23552 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__D
timestamp 1606120350
transform 1 0 23736 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1204__CLK
timestamp 1606120350
transform 1 0 23368 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_230
timestamp 1606120350
transform 1 0 22264 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_244
timestamp 1606120350
transform 1 0 23552 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1606120350
transform 1 0 24012 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_232
timestamp 1606120350
transform 1 0 22448 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245
timestamp 1606120350
transform 1 0 23644 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1204_
timestamp 1606120350
transform 1 0 24288 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__CLK
timestamp 1606120350
transform 1 0 26220 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_271
timestamp 1606120350
transform 1 0 26036 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_257
timestamp 1606120350
transform 1 0 24748 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_269
timestamp 1606120350
transform 1 0 25852 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1198_
timestamp 1606120350
transform 1 0 26864 0 -1 2720
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1606120350
transform 1 0 26772 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1198__D
timestamp 1606120350
transform 1 0 26588 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_275
timestamp 1606120350
transform 1 0 26404 0 -1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1606120350
transform 1 0 26956 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1606120350
transform 1 0 28060 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1606120350
transform 1 0 29624 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1606120350
transform 1 0 29164 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_299
timestamp 1606120350
transform 1 0 28612 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_307
timestamp 1606120350
transform 1 0 29348 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_311
timestamp 1606120350
transform 1 0 29716 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_306
timestamp 1606120350
transform 1 0 29256 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_318
timestamp 1606120350
transform 1 0 30360 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1606120350
transform 1 0 32476 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_323
timestamp 1606120350
transform 1 0 30820 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_335
timestamp 1606120350
transform 1 0 31924 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_342
timestamp 1606120350
transform 1 0 32568 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_330
timestamp 1606120350
transform 1 0 31464 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_342
timestamp 1606120350
transform 1 0 32568 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_354
timestamp 1606120350
transform 1 0 33672 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_354
timestamp 1606120350
transform 1 0 33672 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1606120350
transform 1 0 35328 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1606120350
transform 1 0 34776 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_366
timestamp 1606120350
transform 1 0 34776 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_373
timestamp 1606120350
transform 1 0 35420 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_385
timestamp 1606120350
transform 1 0 36524 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_367
timestamp 1606120350
transform 1 0 34868 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_379
timestamp 1606120350
transform 1 0 35972 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606120350
transform -1 0 38824 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606120350
transform -1 0 38824 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1606120350
transform 1 0 38180 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_397
timestamp 1606120350
transform 1 0 37628 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_404
timestamp 1606120350
transform 1 0 38272 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_391
timestamp 1606120350
transform 1 0 37076 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_403
timestamp 1606120350
transform 1 0 38180 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606120350
transform 1 0 1104 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_3
timestamp 1606120350
transform 1 0 1380 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_15
timestamp 1606120350
transform 1 0 2484 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1606120350
transform 1 0 3956 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_27
timestamp 1606120350
transform 1 0 3588 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1606120350
transform 1 0 4048 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1606120350
transform 1 0 5152 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1606120350
transform 1 0 6256 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1606120350
transform 1 0 7360 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1606120350
transform 1 0 8464 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1606120350
transform 1 0 9568 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1606120350
transform 1 0 9660 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1606120350
transform 1 0 10764 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1131_
timestamp 1606120350
transform 1 0 12696 0 -1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_2_117
timestamp 1606120350
transform 1 0 11868 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_125
timestamp 1606120350
transform 1 0 12604 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1606120350
transform 1 0 15180 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_145
timestamp 1606120350
transform 1 0 14444 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1606120350
transform 1 0 15272 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1606120350
transform 1 0 16376 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1606120350
transform 1 0 17480 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__CLK
timestamp 1606120350
transform 1 0 19504 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_190
timestamp 1606120350
transform 1 0 18584 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_198
timestamp 1606120350
transform 1 0 19320 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1606120350
transform 1 0 19688 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1606120350
transform 1 0 20792 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1606120350
transform 1 0 20884 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1606120350
transform 1 0 21988 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1606120350
transform 1 0 23092 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_251
timestamp 1606120350
transform 1 0 24196 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_263
timestamp 1606120350
transform 1 0 25300 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1606120350
transform 1 0 26404 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_276
timestamp 1606120350
transform 1 0 26496 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_288
timestamp 1606120350
transform 1 0 27600 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_300
timestamp 1606120350
transform 1 0 28704 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_312
timestamp 1606120350
transform 1 0 29808 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1606120350
transform 1 0 32016 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_324
timestamp 1606120350
transform 1 0 30912 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_337
timestamp 1606120350
transform 1 0 32108 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_349
timestamp 1606120350
transform 1 0 33212 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_361
timestamp 1606120350
transform 1 0 34316 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_373
timestamp 1606120350
transform 1 0 35420 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_385
timestamp 1606120350
transform 1 0 36524 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606120350
transform -1 0 38824 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1606120350
transform 1 0 37628 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_398
timestamp 1606120350
transform 1 0 37720 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_406
timestamp 1606120350
transform 1 0 38456 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606120350
transform 1 0 1104 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1606120350
transform 1 0 1380 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1606120350
transform 1 0 2484 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1606120350
transform 1 0 3588 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1606120350
transform 1 0 4692 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1606120350
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1606120350
transform 1 0 5796 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1606120350
transform 1 0 6532 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1606120350
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1606120350
transform 1 0 7912 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_86
timestamp 1606120350
transform 1 0 9016 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_98
timestamp 1606120350
transform 1 0 10120 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_110
timestamp 1606120350
transform 1 0 11224 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1606120350
transform 1 0 12328 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__D
timestamp 1606120350
transform 1 0 12604 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1119__CLK
timestamp 1606120350
transform 1 0 12972 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1143__CLK
timestamp 1606120350
transform 1 0 13524 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_123
timestamp 1606120350
transform 1 0 12420 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_3_127
timestamp 1606120350
transform 1 0 12788 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_131
timestamp 1606120350
transform 1 0 13156 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_137
timestamp 1606120350
transform 1 0 13708 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_149
timestamp 1606120350
transform 1 0 14812 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_161
timestamp 1606120350
transform 1 0 15916 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_173
timestamp 1606120350
transform 1 0 17020 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_181
timestamp 1606120350
transform 1 0 17756 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1210_
timestamp 1606120350
transform 1 0 19504 0 1 3808
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1606120350
transform 1 0 17940 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1210__D
timestamp 1606120350
transform 1 0 19320 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1606120350
transform 1 0 18032 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_196
timestamp 1606120350
transform 1 0 19136 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_219
timestamp 1606120350
transform 1 0 21252 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1606120350
transform 1 0 23552 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_231
timestamp 1606120350
transform 1 0 22356 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_243
timestamp 1606120350
transform 1 0 23460 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_245
timestamp 1606120350
transform 1 0 23644 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_257
timestamp 1606120350
transform 1 0 24748 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_269
timestamp 1606120350
transform 1 0 25852 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1606120350
transform 1 0 26956 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1606120350
transform 1 0 28060 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1606120350
transform 1 0 29164 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_306
timestamp 1606120350
transform 1 0 29256 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_318
timestamp 1606120350
transform 1 0 30360 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_330
timestamp 1606120350
transform 1 0 31464 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_342
timestamp 1606120350
transform 1 0 32568 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_354
timestamp 1606120350
transform 1 0 33672 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1606120350
transform 1 0 34776 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_367
timestamp 1606120350
transform 1 0 34868 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_379
timestamp 1606120350
transform 1 0 35972 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606120350
transform -1 0 38824 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_391
timestamp 1606120350
transform 1 0 37076 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_403
timestamp 1606120350
transform 1 0 38180 0 1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606120350
transform 1 0 1104 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1606120350
transform 1 0 1380 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1606120350
transform 1 0 2484 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1606120350
transform 1 0 3956 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1606120350
transform 1 0 3588 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1606120350
transform 1 0 4048 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1606120350
transform 1 0 5152 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1606120350
transform 1 0 6256 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1606120350
transform 1 0 7360 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1606120350
transform 1 0 8464 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1606120350
transform 1 0 9568 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1606120350
transform 1 0 9660 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1606120350
transform 1 0 10764 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1119_
timestamp 1606120350
transform 1 0 12420 0 -1 4896
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_4_117
timestamp 1606120350
transform 1 0 11868 0 -1 4896
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1606120350
transform 1 0 15180 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_142
timestamp 1606120350
transform 1 0 14168 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_150
timestamp 1606120350
transform 1 0 14904 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1606120350
transform 1 0 15272 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1606120350
transform 1 0 16376 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1606120350
transform 1 0 17480 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1606120350
transform 1 0 18584 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1606120350
transform 1 0 19688 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1606120350
transform 1 0 20792 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1606120350
transform 1 0 20884 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1606120350
transform 1 0 21988 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_239
timestamp 1606120350
transform 1 0 23092 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_251
timestamp 1606120350
transform 1 0 24196 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_263
timestamp 1606120350
transform 1 0 25300 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1606120350
transform 1 0 26404 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_276
timestamp 1606120350
transform 1 0 26496 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_288
timestamp 1606120350
transform 1 0 27600 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_300
timestamp 1606120350
transform 1 0 28704 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_312
timestamp 1606120350
transform 1 0 29808 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1606120350
transform 1 0 32016 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_324
timestamp 1606120350
transform 1 0 30912 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_337
timestamp 1606120350
transform 1 0 32108 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_349
timestamp 1606120350
transform 1 0 33212 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_361
timestamp 1606120350
transform 1 0 34316 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_373
timestamp 1606120350
transform 1 0 35420 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_385
timestamp 1606120350
transform 1 0 36524 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606120350
transform -1 0 38824 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1606120350
transform 1 0 37628 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_398
timestamp 1606120350
transform 1 0 37720 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_406
timestamp 1606120350
transform 1 0 38456 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606120350
transform 1 0 1104 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1606120350
transform 1 0 1380 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1606120350
transform 1 0 2484 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1606120350
transform 1 0 3588 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1606120350
transform 1 0 4692 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1606120350
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1606120350
transform 1 0 5796 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1606120350
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1606120350
transform 1 0 6808 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_74
timestamp 1606120350
transform 1 0 7912 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_86
timestamp 1606120350
transform 1 0 9016 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_98
timestamp 1606120350
transform 1 0 10120 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_110
timestamp 1606120350
transform 1 0 11224 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1606120350
transform 1 0 12328 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1606120350
transform 1 0 12420 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1606120350
transform 1 0 13524 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1606120350
transform 1 0 14628 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1606120350
transform 1 0 15732 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1606120350
transform 1 0 16836 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1606120350
transform 1 0 17940 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1606120350
transform 1 0 18032 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1606120350
transform 1 0 19136 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1606120350
transform 1 0 20240 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_220
timestamp 1606120350
transform 1 0 21344 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1606120350
transform 1 0 23552 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_232
timestamp 1606120350
transform 1 0 22448 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1606120350
transform 1 0 23644 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_257
timestamp 1606120350
transform 1 0 24748 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_269
timestamp 1606120350
transform 1 0 25852 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1606120350
transform 1 0 26956 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1606120350
transform 1 0 28060 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1606120350
transform 1 0 29164 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_306
timestamp 1606120350
transform 1 0 29256 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_318
timestamp 1606120350
transform 1 0 30360 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_330
timestamp 1606120350
transform 1 0 31464 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_342
timestamp 1606120350
transform 1 0 32568 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_354
timestamp 1606120350
transform 1 0 33672 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1606120350
transform 1 0 34776 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_367
timestamp 1606120350
transform 1 0 34868 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_379
timestamp 1606120350
transform 1 0 35972 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606120350
transform -1 0 38824 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_391
timestamp 1606120350
transform 1 0 37076 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_403
timestamp 1606120350
transform 1 0 38180 0 1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606120350
transform 1 0 1104 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606120350
transform 1 0 1104 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1606120350
transform 1 0 1380 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1606120350
transform 1 0 2484 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1606120350
transform 1 0 1380 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1606120350
transform 1 0 2484 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1606120350
transform 1 0 3956 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1606120350
transform 1 0 3588 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1606120350
transform 1 0 4048 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_44
timestamp 1606120350
transform 1 0 5152 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1606120350
transform 1 0 3588 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1606120350
transform 1 0 4692 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1606120350
transform 1 0 6716 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_56
timestamp 1606120350
transform 1 0 6256 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_68
timestamp 1606120350
transform 1 0 7360 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1606120350
transform 1 0 5796 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1606120350
transform 1 0 6532 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1606120350
transform 1 0 6808 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_80
timestamp 1606120350
transform 1 0 8464 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_74
timestamp 1606120350
transform 1 0 7912 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1606120350
transform 1 0 9016 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1606120350
transform 1 0 9568 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_93
timestamp 1606120350
transform 1 0 9660 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_105
timestamp 1606120350
transform 1 0 10764 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1606120350
transform 1 0 10120 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1606120350
transform 1 0 11224 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1606120350
transform 1 0 12328 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_117
timestamp 1606120350
transform 1 0 11868 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_129
timestamp 1606120350
transform 1 0 12972 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1606120350
transform 1 0 12420 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1606120350
transform 1 0 13524 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1606120350
transform 1 0 15180 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1606120350
transform 1 0 14076 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1606120350
transform 1 0 15272 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1606120350
transform 1 0 14628 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1606120350
transform 1 0 15732 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1606120350
transform 1 0 16376 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1606120350
transform 1 0 17480 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1606120350
transform 1 0 16836 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1606120350
transform 1 0 17940 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1606120350
transform 1 0 18584 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_202
timestamp 1606120350
transform 1 0 19688 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1606120350
transform 1 0 18032 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1606120350
transform 1 0 19136 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1606120350
transform 1 0 20792 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_215
timestamp 1606120350
transform 1 0 20884 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_227
timestamp 1606120350
transform 1 0 21988 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1606120350
transform 1 0 20240 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_220
timestamp 1606120350
transform 1 0 21344 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1606120350
transform 1 0 23552 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_239
timestamp 1606120350
transform 1 0 23092 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_251
timestamp 1606120350
transform 1 0 24196 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_232
timestamp 1606120350
transform 1 0 22448 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1606120350
transform 1 0 23644 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_263
timestamp 1606120350
transform 1 0 25300 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1606120350
transform 1 0 24748 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_269
timestamp 1606120350
transform 1 0 25852 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1606120350
transform 1 0 26404 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_276
timestamp 1606120350
transform 1 0 26496 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_288
timestamp 1606120350
transform 1 0 27600 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1606120350
transform 1 0 26956 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1606120350
transform 1 0 28060 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1606120350
transform 1 0 29164 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_300
timestamp 1606120350
transform 1 0 28704 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_312
timestamp 1606120350
transform 1 0 29808 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_306
timestamp 1606120350
transform 1 0 29256 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_318
timestamp 1606120350
transform 1 0 30360 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1606120350
transform 1 0 32016 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_324
timestamp 1606120350
transform 1 0 30912 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_337
timestamp 1606120350
transform 1 0 32108 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_330
timestamp 1606120350
transform 1 0 31464 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_342
timestamp 1606120350
transform 1 0 32568 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_349
timestamp 1606120350
transform 1 0 33212 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_361
timestamp 1606120350
transform 1 0 34316 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_354
timestamp 1606120350
transform 1 0 33672 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1166_
timestamp 1606120350
transform 1 0 35972 0 1 5984
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1606120350
transform 1 0 34776 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__D
timestamp 1606120350
transform 1 0 35788 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1166__CLK
timestamp 1606120350
transform 1 0 35972 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_373
timestamp 1606120350
transform 1 0 35420 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_6_381
timestamp 1606120350
transform 1 0 36156 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_367
timestamp 1606120350
transform 1 0 34868 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_375
timestamp 1606120350
transform 1 0 35604 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606120350
transform -1 0 38824 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606120350
transform -1 0 38824 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1606120350
transform 1 0 37628 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_393
timestamp 1606120350
transform 1 0 37260 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_398
timestamp 1606120350
transform 1 0 37720 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_406
timestamp 1606120350
transform 1 0 38456 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_398
timestamp 1606120350
transform 1 0 37720 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_406
timestamp 1606120350
transform 1 0 38456 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606120350
transform 1 0 1104 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1606120350
transform 1 0 1380 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1606120350
transform 1 0 2484 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1606120350
transform 1 0 3956 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1606120350
transform 1 0 3588 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1606120350
transform 1 0 4048 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1606120350
transform 1 0 5152 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1606120350
transform 1 0 6256 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_68
timestamp 1606120350
transform 1 0 7360 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1606120350
transform 1 0 8464 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1606120350
transform 1 0 9568 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1606120350
transform 1 0 9660 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1606120350
transform 1 0 10764 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1606120350
transform 1 0 11868 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1606120350
transform 1 0 12972 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1606120350
transform 1 0 15180 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1606120350
transform 1 0 14076 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1606120350
transform 1 0 15272 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1606120350
transform 1 0 16376 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1606120350
transform 1 0 17480 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_190
timestamp 1606120350
transform 1 0 18584 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_202
timestamp 1606120350
transform 1 0 19688 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1606120350
transform 1 0 20792 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1606120350
transform 1 0 20884 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_227
timestamp 1606120350
transform 1 0 21988 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_239
timestamp 1606120350
transform 1 0 23092 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_251
timestamp 1606120350
transform 1 0 24196 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_263
timestamp 1606120350
transform 1 0 25300 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1606120350
transform 1 0 26404 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_276
timestamp 1606120350
transform 1 0 26496 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_288
timestamp 1606120350
transform 1 0 27600 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_300
timestamp 1606120350
transform 1 0 28704 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_312
timestamp 1606120350
transform 1 0 29808 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1606120350
transform 1 0 32016 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_324
timestamp 1606120350
transform 1 0 30912 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_337
timestamp 1606120350
transform 1 0 32108 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_349
timestamp 1606120350
transform 1 0 33212 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_361
timestamp 1606120350
transform 1 0 34316 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_373
timestamp 1606120350
transform 1 0 35420 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_385
timestamp 1606120350
transform 1 0 36524 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606120350
transform -1 0 38824 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1606120350
transform 1 0 37628 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_398
timestamp 1606120350
transform 1 0 37720 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_406
timestamp 1606120350
transform 1 0 38456 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606120350
transform 1 0 1104 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1606120350
transform 1 0 1380 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1606120350
transform 1 0 2484 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1606120350
transform 1 0 3588 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1606120350
transform 1 0 4692 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1606120350
transform 1 0 6716 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1606120350
transform 1 0 5796 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1606120350
transform 1 0 6532 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1606120350
transform 1 0 6808 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_74
timestamp 1606120350
transform 1 0 7912 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_86
timestamp 1606120350
transform 1 0 9016 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_98
timestamp 1606120350
transform 1 0 10120 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_110
timestamp 1606120350
transform 1 0 11224 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1606120350
transform 1 0 12328 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1606120350
transform 1 0 12420 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1606120350
transform 1 0 13524 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_147
timestamp 1606120350
transform 1 0 14628 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_159
timestamp 1606120350
transform 1 0 15732 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_171
timestamp 1606120350
transform 1 0 16836 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1606120350
transform 1 0 17940 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1606120350
transform 1 0 18032 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1606120350
transform 1 0 19136 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1606120350
transform 1 0 20240 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_220
timestamp 1606120350
transform 1 0 21344 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1606120350
transform 1 0 23552 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_232
timestamp 1606120350
transform 1 0 22448 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1606120350
transform 1 0 23644 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1606120350
transform 1 0 24748 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_269
timestamp 1606120350
transform 1 0 25852 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1606120350
transform 1 0 26956 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1606120350
transform 1 0 28060 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1606120350
transform 1 0 29164 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_306
timestamp 1606120350
transform 1 0 29256 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_318
timestamp 1606120350
transform 1 0 30360 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_330
timestamp 1606120350
transform 1 0 31464 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_342
timestamp 1606120350
transform 1 0 32568 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_354
timestamp 1606120350
transform 1 0 33672 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1606120350
transform 1 0 34776 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_367
timestamp 1606120350
transform 1 0 34868 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_379
timestamp 1606120350
transform 1 0 35972 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606120350
transform -1 0 38824 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_391
timestamp 1606120350
transform 1 0 37076 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_403
timestamp 1606120350
transform 1 0 38180 0 1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606120350
transform 1 0 1104 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1606120350
transform 1 0 1380 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1606120350
transform 1 0 2484 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1606120350
transform 1 0 3956 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1606120350
transform 1 0 3588 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1606120350
transform 1 0 4048 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1606120350
transform 1 0 5152 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1606120350
transform 1 0 6256 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1606120350
transform 1 0 7360 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_80
timestamp 1606120350
transform 1 0 8464 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1606120350
transform 1 0 9568 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1606120350
transform 1 0 9660 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_105
timestamp 1606120350
transform 1 0 10764 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_117
timestamp 1606120350
transform 1 0 11868 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_129
timestamp 1606120350
transform 1 0 12972 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1606120350
transform 1 0 15180 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1606120350
transform 1 0 14076 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1606120350
transform 1 0 15272 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_166
timestamp 1606120350
transform 1 0 16376 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_178
timestamp 1606120350
transform 1 0 17480 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_190
timestamp 1606120350
transform 1 0 18584 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_202
timestamp 1606120350
transform 1 0 19688 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1606120350
transform 1 0 20792 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1606120350
transform 1 0 20884 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1606120350
transform 1 0 21988 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1606120350
transform 1 0 23092 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_251
timestamp 1606120350
transform 1 0 24196 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_263
timestamp 1606120350
transform 1 0 25300 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1606120350
transform 1 0 26404 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_276
timestamp 1606120350
transform 1 0 26496 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_288
timestamp 1606120350
transform 1 0 27600 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_300
timestamp 1606120350
transform 1 0 28704 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_312
timestamp 1606120350
transform 1 0 29808 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1606120350
transform 1 0 32016 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_324
timestamp 1606120350
transform 1 0 30912 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_337
timestamp 1606120350
transform 1 0 32108 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_349
timestamp 1606120350
transform 1 0 33212 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_361
timestamp 1606120350
transform 1 0 34316 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_373
timestamp 1606120350
transform 1 0 35420 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_385
timestamp 1606120350
transform 1 0 36524 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606120350
transform -1 0 38824 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1606120350
transform 1 0 37628 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_398
timestamp 1606120350
transform 1 0 37720 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_406
timestamp 1606120350
transform 1 0 38456 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606120350
transform 1 0 1104 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1606120350
transform 1 0 1380 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1606120350
transform 1 0 2484 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1606120350
transform 1 0 3588 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1606120350
transform 1 0 4692 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1606120350
transform 1 0 6716 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1606120350
transform 1 0 5796 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1606120350
transform 1 0 6532 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1606120350
transform 1 0 6808 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_74
timestamp 1606120350
transform 1 0 7912 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_86
timestamp 1606120350
transform 1 0 9016 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_98
timestamp 1606120350
transform 1 0 10120 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_110
timestamp 1606120350
transform 1 0 11224 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1606120350
transform 1 0 12328 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1606120350
transform 1 0 12420 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1606120350
transform 1 0 13524 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_147
timestamp 1606120350
transform 1 0 14628 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_159
timestamp 1606120350
transform 1 0 15732 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_171
timestamp 1606120350
transform 1 0 16836 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1606120350
transform 1 0 17940 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1606120350
transform 1 0 18032 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1606120350
transform 1 0 19136 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1606120350
transform 1 0 20240 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_220
timestamp 1606120350
transform 1 0 21344 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1606120350
transform 1 0 23552 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_232
timestamp 1606120350
transform 1 0 22448 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_245
timestamp 1606120350
transform 1 0 23644 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_257
timestamp 1606120350
transform 1 0 24748 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_269
timestamp 1606120350
transform 1 0 25852 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1606120350
transform 1 0 26956 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1606120350
transform 1 0 28060 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1606120350
transform 1 0 29164 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_306
timestamp 1606120350
transform 1 0 29256 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_318
timestamp 1606120350
transform 1 0 30360 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_330
timestamp 1606120350
transform 1 0 31464 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_342
timestamp 1606120350
transform 1 0 32568 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_354
timestamp 1606120350
transform 1 0 33672 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1606120350
transform 1 0 34776 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_367
timestamp 1606120350
transform 1 0 34868 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_379
timestamp 1606120350
transform 1 0 35972 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606120350
transform -1 0 38824 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_391
timestamp 1606120350
transform 1 0 37076 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_403
timestamp 1606120350
transform 1 0 38180 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606120350
transform 1 0 1104 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1606120350
transform 1 0 1380 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1606120350
transform 1 0 2484 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1606120350
transform 1 0 3956 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1606120350
transform 1 0 3588 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1606120350
transform 1 0 4048 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1606120350
transform 1 0 5152 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1606120350
transform 1 0 6256 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1606120350
transform 1 0 7360 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1606120350
transform 1 0 8464 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1606120350
transform 1 0 9568 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1606120350
transform 1 0 9660 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_105
timestamp 1606120350
transform 1 0 10764 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_117
timestamp 1606120350
transform 1 0 11868 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_129
timestamp 1606120350
transform 1 0 12972 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1606120350
transform 1 0 15180 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1606120350
transform 1 0 14076 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1606120350
transform 1 0 15272 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1606120350
transform 1 0 16376 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1606120350
transform 1 0 17480 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_190
timestamp 1606120350
transform 1 0 18584 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_202
timestamp 1606120350
transform 1 0 19688 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1606120350
transform 1 0 20792 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1606120350
transform 1 0 20884 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1606120350
transform 1 0 21988 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1606120350
transform 1 0 23092 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_251
timestamp 1606120350
transform 1 0 24196 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_263
timestamp 1606120350
transform 1 0 25300 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1606120350
transform 1 0 26404 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_276
timestamp 1606120350
transform 1 0 26496 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_288
timestamp 1606120350
transform 1 0 27600 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_300
timestamp 1606120350
transform 1 0 28704 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_312
timestamp 1606120350
transform 1 0 29808 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1606120350
transform 1 0 32016 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_324
timestamp 1606120350
transform 1 0 30912 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_337
timestamp 1606120350
transform 1 0 32108 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_349
timestamp 1606120350
transform 1 0 33212 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_361
timestamp 1606120350
transform 1 0 34316 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_373
timestamp 1606120350
transform 1 0 35420 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_385
timestamp 1606120350
transform 1 0 36524 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606120350
transform -1 0 38824 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1606120350
transform 1 0 37628 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_398
timestamp 1606120350
transform 1 0 37720 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_406
timestamp 1606120350
transform 1 0 38456 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1218_
timestamp 1606120350
transform 1 0 1472 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606120350
transform 1 0 1104 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606120350
transform 1 0 1104 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__D
timestamp 1606120350
transform 1 0 1564 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1218__CLK
timestamp 1606120350
transform 1 0 1932 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_3
timestamp 1606120350
transform 1 0 1380 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_13_7
timestamp 1606120350
transform 1 0 1748 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_11
timestamp 1606120350
transform 1 0 2116 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_3
timestamp 1606120350
transform 1 0 1380 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1606120350
transform 1 0 3956 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_23
timestamp 1606120350
transform 1 0 3220 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_35
timestamp 1606120350
transform 1 0 4324 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_23
timestamp 1606120350
transform 1 0 3220 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1606120350
transform 1 0 4048 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1606120350
transform 1 0 5152 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1202_
timestamp 1606120350
transform 1 0 7084 0 -1 10336
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1606120350
transform 1 0 6716 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__D
timestamp 1606120350
transform 1 0 7084 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_47
timestamp 1606120350
transform 1 0 5428 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1606120350
transform 1 0 6532 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_13_62
timestamp 1606120350
transform 1 0 6808 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_13_67
timestamp 1606120350
transform 1 0 7268 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_14_56
timestamp 1606120350
transform 1 0 6256 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_64
timestamp 1606120350
transform 1 0 6992 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1202__CLK
timestamp 1606120350
transform 1 0 7452 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_71
timestamp 1606120350
transform 1 0 7636 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_83
timestamp 1606120350
transform 1 0 8740 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_84
timestamp 1606120350
transform 1 0 8832 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1606120350
transform 1 0 9568 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_95
timestamp 1606120350
transform 1 0 9844 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_107
timestamp 1606120350
transform 1 0 10948 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1606120350
transform 1 0 9660 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_105
timestamp 1606120350
transform 1 0 10764 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1606120350
transform 1 0 12328 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_119
timestamp 1606120350
transform 1 0 12052 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1606120350
transform 1 0 12420 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_135
timestamp 1606120350
transform 1 0 13524 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_117
timestamp 1606120350
transform 1 0 11868 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_129
timestamp 1606120350
transform 1 0 12972 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1606120350
transform 1 0 15180 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_147
timestamp 1606120350
transform 1 0 14628 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_159
timestamp 1606120350
transform 1 0 15732 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1606120350
transform 1 0 14076 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_154
timestamp 1606120350
transform 1 0 15272 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_171
timestamp 1606120350
transform 1 0 16836 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_166
timestamp 1606120350
transform 1 0 16376 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_178
timestamp 1606120350
transform 1 0 17480 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1606120350
transform 1 0 17940 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1606120350
transform 1 0 18032 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1606120350
transform 1 0 19136 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_190
timestamp 1606120350
transform 1 0 18584 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_202
timestamp 1606120350
transform 1 0 19688 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1606120350
transform 1 0 20792 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1606120350
transform 1 0 20240 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_220
timestamp 1606120350
transform 1 0 21344 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_215
timestamp 1606120350
transform 1 0 20884 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_227
timestamp 1606120350
transform 1 0 21988 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1606120350
transform 1 0 23552 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_232
timestamp 1606120350
transform 1 0 22448 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_245
timestamp 1606120350
transform 1 0 23644 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_239
timestamp 1606120350
transform 1 0 23092 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_251
timestamp 1606120350
transform 1 0 24196 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_257
timestamp 1606120350
transform 1 0 24748 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_269
timestamp 1606120350
transform 1 0 25852 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_263
timestamp 1606120350
transform 1 0 25300 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1606120350
transform 1 0 26404 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1606120350
transform 1 0 26956 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1606120350
transform 1 0 28060 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_276
timestamp 1606120350
transform 1 0 26496 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_288
timestamp 1606120350
transform 1 0 27600 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1606120350
transform 1 0 29164 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_306
timestamp 1606120350
transform 1 0 29256 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_318
timestamp 1606120350
transform 1 0 30360 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_300
timestamp 1606120350
transform 1 0 28704 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_312
timestamp 1606120350
transform 1 0 29808 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1606120350
transform 1 0 32016 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_330
timestamp 1606120350
transform 1 0 31464 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_342
timestamp 1606120350
transform 1 0 32568 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_324
timestamp 1606120350
transform 1 0 30912 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_337
timestamp 1606120350
transform 1 0 32108 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_354
timestamp 1606120350
transform 1 0 33672 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_349
timestamp 1606120350
transform 1 0 33212 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_361
timestamp 1606120350
transform 1 0 34316 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1606120350
transform 1 0 34776 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_367
timestamp 1606120350
transform 1 0 34868 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_379
timestamp 1606120350
transform 1 0 35972 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_373
timestamp 1606120350
transform 1 0 35420 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_385
timestamp 1606120350
transform 1 0 36524 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606120350
transform -1 0 38824 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606120350
transform -1 0 38824 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1606120350
transform 1 0 37628 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_391
timestamp 1606120350
transform 1 0 37076 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_403
timestamp 1606120350
transform 1 0 38180 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_398
timestamp 1606120350
transform 1 0 37720 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_406
timestamp 1606120350
transform 1 0 38456 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606120350
transform 1 0 1104 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1606120350
transform 1 0 1380 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1606120350
transform 1 0 2484 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1606120350
transform 1 0 3588 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1606120350
transform 1 0 4692 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1606120350
transform 1 0 6716 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1606120350
transform 1 0 5796 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1606120350
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1606120350
transform 1 0 6808 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_74
timestamp 1606120350
transform 1 0 7912 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_86
timestamp 1606120350
transform 1 0 9016 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_98
timestamp 1606120350
transform 1 0 10120 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_110
timestamp 1606120350
transform 1 0 11224 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1606120350
transform 1 0 12328 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1606120350
transform 1 0 12420 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_135
timestamp 1606120350
transform 1 0 13524 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__A1
timestamp 1606120350
transform 1 0 15548 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__A2
timestamp 1606120350
transform 1 0 15180 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_147
timestamp 1606120350
transform 1 0 14628 0 1 10336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_15_155
timestamp 1606120350
transform 1 0 15364 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_159
timestamp 1606120350
transform 1 0 15732 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__B1
timestamp 1606120350
transform 1 0 15916 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0794__B2
timestamp 1606120350
transform 1 0 16284 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__D
timestamp 1606120350
transform 1 0 17572 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_163
timestamp 1606120350
transform 1 0 16100 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_167
timestamp 1606120350
transform 1 0 16468 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_181
timestamp 1606120350
transform 1 0 17756 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1606120350
transform 1 0 17940 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1097__CLK
timestamp 1606120350
transform 1 0 18216 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_15_184
timestamp 1606120350
transform 1 0 18032 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_188
timestamp 1606120350
transform 1 0 18400 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_200
timestamp 1606120350
transform 1 0 19504 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_212
timestamp 1606120350
transform 1 0 20608 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_224
timestamp 1606120350
transform 1 0 21712 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1606120350
transform 1 0 23552 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_236
timestamp 1606120350
transform 1 0 22816 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_245
timestamp 1606120350
transform 1 0 23644 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_257
timestamp 1606120350
transform 1 0 24748 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_269
timestamp 1606120350
transform 1 0 25852 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1606120350
transform 1 0 26956 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1606120350
transform 1 0 28060 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1606120350
transform 1 0 29164 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_306
timestamp 1606120350
transform 1 0 29256 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_318
timestamp 1606120350
transform 1 0 30360 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_330
timestamp 1606120350
transform 1 0 31464 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_342
timestamp 1606120350
transform 1 0 32568 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_354
timestamp 1606120350
transform 1 0 33672 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1606120350
transform 1 0 34776 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_367
timestamp 1606120350
transform 1 0 34868 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_379
timestamp 1606120350
transform 1 0 35972 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606120350
transform -1 0 38824 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_391
timestamp 1606120350
transform 1 0 37076 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_403
timestamp 1606120350
transform 1 0 38180 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606120350
transform 1 0 1104 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1606120350
transform 1 0 1380 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1606120350
transform 1 0 2484 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1606120350
transform 1 0 3956 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1606120350
transform 1 0 3588 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1606120350
transform 1 0 4048 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1606120350
transform 1 0 5152 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1606120350
transform 1 0 6256 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1606120350
transform 1 0 7360 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1606120350
transform 1 0 8464 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1606120350
transform 1 0 9568 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1606120350
transform 1 0 9660 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_105
timestamp 1606120350
transform 1 0 10764 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_117
timestamp 1606120350
transform 1 0 11868 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_129
timestamp 1606120350
transform 1 0 12972 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _0794_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 15548 0 -1 11424
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1606120350
transform 1 0 15180 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1606120350
transform 1 0 14076 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_154
timestamp 1606120350
transform 1 0 15272 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1097_
timestamp 1606120350
transform 1 0 17572 0 -1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_16_171
timestamp 1606120350
transform 1 0 16836 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__CLK
timestamp 1606120350
transform 1 0 19504 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_16_198
timestamp 1606120350
transform 1 0 19320 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_202
timestamp 1606120350
transform 1 0 19688 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1606120350
transform 1 0 20792 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1606120350
transform 1 0 20884 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_227
timestamp 1606120350
transform 1 0 21988 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_239
timestamp 1606120350
transform 1 0 23092 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_251
timestamp 1606120350
transform 1 0 24196 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_263
timestamp 1606120350
transform 1 0 25300 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1606120350
transform 1 0 26404 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_276
timestamp 1606120350
transform 1 0 26496 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_288
timestamp 1606120350
transform 1 0 27600 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_300
timestamp 1606120350
transform 1 0 28704 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_312
timestamp 1606120350
transform 1 0 29808 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1606120350
transform 1 0 32016 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_324
timestamp 1606120350
transform 1 0 30912 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_337
timestamp 1606120350
transform 1 0 32108 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_349
timestamp 1606120350
transform 1 0 33212 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_361
timestamp 1606120350
transform 1 0 34316 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_373
timestamp 1606120350
transform 1 0 35420 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_385
timestamp 1606120350
transform 1 0 36524 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606120350
transform -1 0 38824 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1606120350
transform 1 0 37628 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_398
timestamp 1606120350
transform 1 0 37720 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_406
timestamp 1606120350
transform 1 0 38456 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606120350
transform 1 0 1104 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1606120350
transform 1 0 1380 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1606120350
transform 1 0 2484 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1606120350
transform 1 0 3588 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1606120350
transform 1 0 4692 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1606120350
transform 1 0 6716 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1606120350
transform 1 0 5796 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1606120350
transform 1 0 6532 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1606120350
transform 1 0 6808 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_74
timestamp 1606120350
transform 1 0 7912 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_86
timestamp 1606120350
transform 1 0 9016 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_98
timestamp 1606120350
transform 1 0 10120 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_110
timestamp 1606120350
transform 1 0 11224 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1606120350
transform 1 0 12328 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__A1
timestamp 1606120350
transform 1 0 13156 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__B1
timestamp 1606120350
transform 1 0 13524 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__A2
timestamp 1606120350
transform 1 0 12788 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_123
timestamp 1606120350
transform 1 0 12420 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_17_129
timestamp 1606120350
transform 1 0 12972 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_133
timestamp 1606120350
transform 1 0 13340 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_137
timestamp 1606120350
transform 1 0 13708 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1096_
timestamp 1606120350
transform 1 0 15456 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0786__B2
timestamp 1606120350
transform 1 0 13892 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__D
timestamp 1606120350
transform 1 0 15272 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__CLK
timestamp 1606120350
transform 1 0 14904 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_141
timestamp 1606120350
transform 1 0 14076 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_149
timestamp 1606120350
transform 1 0 14812 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_152
timestamp 1606120350
transform 1 0 15088 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__B2
timestamp 1606120350
transform 1 0 17756 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1094__CLK
timestamp 1606120350
transform 1 0 17388 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_175
timestamp 1606120350
transform 1 0 17204 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_179
timestamp 1606120350
transform 1 0 17572 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1139_
timestamp 1606120350
transform 1 0 19412 0 1 11424
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1606120350
transform 1 0 17940 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1139__D
timestamp 1606120350
transform 1 0 19228 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__A1
timestamp 1606120350
transform 1 0 18584 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__B1
timestamp 1606120350
transform 1 0 18216 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_184
timestamp 1606120350
transform 1 0 18032 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_17_188
timestamp 1606120350
transform 1 0 18400 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_192
timestamp 1606120350
transform 1 0 18768 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_196
timestamp 1606120350
transform 1 0 19136 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_218
timestamp 1606120350
transform 1 0 21160 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1606120350
transform 1 0 23552 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_230
timestamp 1606120350
transform 1 0 22264 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_242
timestamp 1606120350
transform 1 0 23368 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_245
timestamp 1606120350
transform 1 0 23644 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_257
timestamp 1606120350
transform 1 0 24748 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_269
timestamp 1606120350
transform 1 0 25852 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1606120350
transform 1 0 26956 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1606120350
transform 1 0 28060 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1606120350
transform 1 0 29164 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_306
timestamp 1606120350
transform 1 0 29256 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_318
timestamp 1606120350
transform 1 0 30360 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_330
timestamp 1606120350
transform 1 0 31464 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_342
timestamp 1606120350
transform 1 0 32568 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_354
timestamp 1606120350
transform 1 0 33672 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1606120350
transform 1 0 34776 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_367
timestamp 1606120350
transform 1 0 34868 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_379
timestamp 1606120350
transform 1 0 35972 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606120350
transform -1 0 38824 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_391
timestamp 1606120350
transform 1 0 37076 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_403
timestamp 1606120350
transform 1 0 38180 0 1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606120350
transform 1 0 1104 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1606120350
transform 1 0 1380 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1606120350
transform 1 0 2484 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1606120350
transform 1 0 3956 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1606120350
transform 1 0 3588 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1606120350
transform 1 0 4048 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1606120350
transform 1 0 5152 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1606120350
transform 1 0 6256 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1606120350
transform 1 0 7360 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_80
timestamp 1606120350
transform 1 0 8464 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1606120350
transform 1 0 9568 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1606120350
transform 1 0 9660 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1606120350
transform 1 0 10764 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _0786_
timestamp 1606120350
transform 1 0 13156 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_18_117
timestamp 1606120350
transform 1 0 11868 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_129
timestamp 1606120350
transform 1 0 12972 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1606120350
transform 1 0 15180 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1096__D
timestamp 1606120350
transform 1 0 15456 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_145
timestamp 1606120350
transform 1 0 14444 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_154
timestamp 1606120350
transform 1 0 15272 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_158
timestamp 1606120350
transform 1 0 15640 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1094_
timestamp 1606120350
transform 1 0 16100 0 -1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_18_162
timestamp 1606120350
transform 1 0 16008 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_18_182
timestamp 1606120350
transform 1 0 17848 0 -1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_4  _0796_
timestamp 1606120350
transform 1 0 18584 0 -1 12512
box -38 -48 1326 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0796__A2
timestamp 1606120350
transform 1 0 18400 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_18_204
timestamp 1606120350
transform 1 0 19872 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1606120350
transform 1 0 20792 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_18_212
timestamp 1606120350
transform 1 0 20608 0 -1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_18_215
timestamp 1606120350
transform 1 0 20884 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_227
timestamp 1606120350
transform 1 0 21988 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_239
timestamp 1606120350
transform 1 0 23092 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_251
timestamp 1606120350
transform 1 0 24196 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_263
timestamp 1606120350
transform 1 0 25300 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1606120350
transform 1 0 26404 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_276
timestamp 1606120350
transform 1 0 26496 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_288
timestamp 1606120350
transform 1 0 27600 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_300
timestamp 1606120350
transform 1 0 28704 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_312
timestamp 1606120350
transform 1 0 29808 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1606120350
transform 1 0 32016 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_324
timestamp 1606120350
transform 1 0 30912 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_337
timestamp 1606120350
transform 1 0 32108 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_349
timestamp 1606120350
transform 1 0 33212 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_361
timestamp 1606120350
transform 1 0 34316 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_373
timestamp 1606120350
transform 1 0 35420 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_385
timestamp 1606120350
transform 1 0 36524 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606120350
transform -1 0 38824 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1606120350
transform 1 0 37628 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_398
timestamp 1606120350
transform 1 0 37720 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_406
timestamp 1606120350
transform 1 0 38456 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606120350
transform 1 0 1104 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606120350
transform 1 0 1104 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1606120350
transform 1 0 1380 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1606120350
transform 1 0 2484 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1606120350
transform 1 0 1380 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1606120350
transform 1 0 2484 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1606120350
transform 1 0 3956 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1606120350
transform 1 0 3588 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1606120350
transform 1 0 4692 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1606120350
transform 1 0 3588 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1606120350
transform 1 0 4048 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1606120350
transform 1 0 5152 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1606120350
transform 1 0 6716 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1606120350
transform 1 0 5796 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1606120350
transform 1 0 6532 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1606120350
transform 1 0 6808 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_56
timestamp 1606120350
transform 1 0 6256 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_68
timestamp 1606120350
transform 1 0 7360 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_74
timestamp 1606120350
transform 1 0 7912 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_86
timestamp 1606120350
transform 1 0 9016 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_80
timestamp 1606120350
transform 1 0 8464 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1606120350
transform 1 0 9568 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_98
timestamp 1606120350
transform 1 0 10120 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_110
timestamp 1606120350
transform 1 0 11224 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1606120350
transform 1 0 9660 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1606120350
transform 1 0 10764 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1093_
timestamp 1606120350
transform 1 0 13616 0 1 12512
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1606120350
transform 1 0 12328 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__D
timestamp 1606120350
transform 1 0 13432 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1093__CLK
timestamp 1606120350
transform 1 0 13616 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_123
timestamp 1606120350
transform 1 0 12420 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_131
timestamp 1606120350
transform 1 0 13156 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1606120350
transform 1 0 11868 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_129
timestamp 1606120350
transform 1 0 12972 0 -1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_135
timestamp 1606120350
transform 1 0 13524 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1606120350
transform 1 0 15180 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_155
timestamp 1606120350
transform 1 0 15364 0 1 12512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_138
timestamp 1606120350
transform 1 0 13800 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_150
timestamp 1606120350
transform 1 0 14904 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_154
timestamp 1606120350
transform 1 0 15272 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_162
timestamp 1606120350
transform 1 0 16008 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_19_171
timestamp 1606120350
transform 1 0 16836 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_167
timestamp 1606120350
transform 1 0 16468 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_19_163
timestamp 1606120350
transform 1 0 16100 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__A2
timestamp 1606120350
transform 1 0 15916 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__B1
timestamp 1606120350
transform 1 0 16652 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__A1
timestamp 1606120350
transform 1 0 16284 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_175
timestamp 1606120350
transform 1 0 17204 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0789__B2
timestamp 1606120350
transform 1 0 17020 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_179
timestamp 1606120350
transform 1 0 17572 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _0789_
timestamp 1606120350
transform 1 0 16284 0 -1 13600
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1606120350
transform 1 0 17940 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1606120350
transform 1 0 18032 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1606120350
transform 1 0 19136 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_191
timestamp 1606120350
transform 1 0 18676 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_203
timestamp 1606120350
transform 1 0 19780 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_215
timestamp 1606120350
transform 1 0 20884 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_211
timestamp 1606120350
transform 1 0 20516 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1606120350
transform 1 0 20792 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_20_223
timestamp 1606120350
transform 1 0 21620 0 -1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_19_224
timestamp 1606120350
transform 1 0 21712 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_220
timestamp 1606120350
transform 1 0 21344 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_4_0_clk_A
timestamp 1606120350
transform 1 0 21804 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_4_0_clk /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 21804 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_228
timestamp 1606120350
transform 1 0 22080 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_227
timestamp 1606120350
transform 1 0 21988 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1606120350
transform 1 0 20240 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1606120350
transform 1 0 23552 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_239
timestamp 1606120350
transform 1 0 23092 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_243
timestamp 1606120350
transform 1 0 23460 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_245
timestamp 1606120350
transform 1 0 23644 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_240
timestamp 1606120350
transform 1 0 23184 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_257
timestamp 1606120350
transform 1 0 24748 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_269
timestamp 1606120350
transform 1 0 25852 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_252
timestamp 1606120350
transform 1 0 24288 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_264
timestamp 1606120350
transform 1 0 25392 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_272
timestamp 1606120350
transform 1 0 26128 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1606120350
transform 1 0 26404 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1606120350
transform 1 0 26956 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1606120350
transform 1 0 28060 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_276
timestamp 1606120350
transform 1 0 26496 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_288
timestamp 1606120350
transform 1 0 27600 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1606120350
transform 1 0 29164 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_306
timestamp 1606120350
transform 1 0 29256 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_318
timestamp 1606120350
transform 1 0 30360 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_300
timestamp 1606120350
transform 1 0 28704 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_312
timestamp 1606120350
transform 1 0 29808 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1606120350
transform 1 0 32016 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_330
timestamp 1606120350
transform 1 0 31464 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_342
timestamp 1606120350
transform 1 0 32568 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_324
timestamp 1606120350
transform 1 0 30912 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_337
timestamp 1606120350
transform 1 0 32108 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_354
timestamp 1606120350
transform 1 0 33672 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_349
timestamp 1606120350
transform 1 0 33212 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_361
timestamp 1606120350
transform 1 0 34316 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1606120350
transform 1 0 34776 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_367
timestamp 1606120350
transform 1 0 34868 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_379
timestamp 1606120350
transform 1 0 35972 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_373
timestamp 1606120350
transform 1 0 35420 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_385
timestamp 1606120350
transform 1 0 36524 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606120350
transform -1 0 38824 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606120350
transform -1 0 38824 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1606120350
transform 1 0 37628 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_391
timestamp 1606120350
transform 1 0 37076 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_403
timestamp 1606120350
transform 1 0 38180 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_398
timestamp 1606120350
transform 1 0 37720 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_406
timestamp 1606120350
transform 1 0 38456 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606120350
transform 1 0 1104 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1606120350
transform 1 0 1380 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1606120350
transform 1 0 2484 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1606120350
transform 1 0 3588 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1606120350
transform 1 0 4692 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1606120350
transform 1 0 6716 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1606120350
transform 1 0 5796 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1606120350
transform 1 0 6532 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1606120350
transform 1 0 6808 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_74
timestamp 1606120350
transform 1 0 7912 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_86
timestamp 1606120350
transform 1 0 9016 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_1_0_clk_A
timestamp 1606120350
transform 1 0 11408 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_98
timestamp 1606120350
transform 1 0 10120 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_110
timestamp 1606120350
transform 1 0 11224 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_114
timestamp 1606120350
transform 1 0 11592 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1606120350
transform 1 0 12328 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_123
timestamp 1606120350
transform 1 0 12420 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_135
timestamp 1606120350
transform 1 0 13524 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__A
timestamp 1606120350
transform 1 0 15272 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0714__B
timestamp 1606120350
transform 1 0 15640 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_147
timestamp 1606120350
transform 1 0 14628 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_153
timestamp 1606120350
transform 1 0 15180 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_156
timestamp 1606120350
transform 1 0 15456 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__D
timestamp 1606120350
transform 1 0 17572 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_160
timestamp 1606120350
transform 1 0 15824 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_172
timestamp 1606120350
transform 1 0 16928 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_178
timestamp 1606120350
transform 1 0 17480 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_181
timestamp 1606120350
transform 1 0 17756 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1606120350
transform 1 0 17940 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1095__CLK
timestamp 1606120350
transform 1 0 18216 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_184
timestamp 1606120350
transform 1 0 18032 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_188
timestamp 1606120350
transform 1 0 18400 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_200
timestamp 1606120350
transform 1 0 19504 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_212
timestamp 1606120350
transform 1 0 20608 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_224
timestamp 1606120350
transform 1 0 21712 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1606120350
transform 1 0 23552 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_2_0_clk_A
timestamp 1606120350
transform 1 0 23092 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_21_236
timestamp 1606120350
transform 1 0 22816 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_21_241
timestamp 1606120350
transform 1 0 23276 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_245
timestamp 1606120350
transform 1 0 23644 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_5_0_clk
timestamp 1606120350
transform 1 0 24932 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_5_0_clk_A
timestamp 1606120350
transform 1 0 25392 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_257
timestamp 1606120350
transform 1 0 24748 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_21_262
timestamp 1606120350
transform 1 0 25208 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_266
timestamp 1606120350
transform 1 0 25576 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_278
timestamp 1606120350
transform 1 0 26680 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_290
timestamp 1606120350
transform 1 0 27784 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1606120350
transform 1 0 29164 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_302
timestamp 1606120350
transform 1 0 28888 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_306
timestamp 1606120350
transform 1 0 29256 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_318
timestamp 1606120350
transform 1 0 30360 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_330
timestamp 1606120350
transform 1 0 31464 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_342
timestamp 1606120350
transform 1 0 32568 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_354
timestamp 1606120350
transform 1 0 33672 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1606120350
transform 1 0 34776 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_367
timestamp 1606120350
transform 1 0 34868 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_379
timestamp 1606120350
transform 1 0 35972 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606120350
transform -1 0 38824 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_391
timestamp 1606120350
transform 1 0 37076 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_403
timestamp 1606120350
transform 1 0 38180 0 1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606120350
transform 1 0 1104 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1606120350
transform 1 0 1380 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1606120350
transform 1 0 2484 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1606120350
transform 1 0 3956 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1606120350
transform 1 0 3588 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1606120350
transform 1 0 4048 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1606120350
transform 1 0 5152 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1606120350
transform 1 0 6256 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1606120350
transform 1 0 7360 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_80
timestamp 1606120350
transform 1 0 8464 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1606120350
transform 1 0 9568 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_1_0_clk
timestamp 1606120350
transform 1 0 11408 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1606120350
transform 1 0 9660 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_105
timestamp 1606120350
transform 1 0 10764 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_111
timestamp 1606120350
transform 1 0 11316 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__CLK
timestamp 1606120350
transform 1 0 13524 0 -1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_115
timestamp 1606120350
transform 1 0 11684 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_127
timestamp 1606120350
transform 1 0 12788 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_22_137
timestamp 1606120350
transform 1 0 13708 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _0714_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 15272 0 -1 14688
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1606120350
transform 1 0 15180 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_149
timestamp 1606120350
transform 1 0 14812 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1095_
timestamp 1606120350
transform 1 0 17572 0 -1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_22_161
timestamp 1606120350
transform 1 0 15916 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_173
timestamp 1606120350
transform 1 0 17020 0 -1 14688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_198
timestamp 1606120350
transform 1 0 19320 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1606120350
transform 1 0 20792 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_210
timestamp 1606120350
transform 1 0 20424 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_215
timestamp 1606120350
transform 1 0 20884 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_227
timestamp 1606120350
transform 1 0 21988 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_2_0_clk
timestamp 1606120350
transform 1 0 23092 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_242
timestamp 1606120350
transform 1 0 23368 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_254
timestamp 1606120350
transform 1 0 24472 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_266
timestamp 1606120350
transform 1 0 25576 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_274
timestamp 1606120350
transform 1 0 26312 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1606120350
transform 1 0 26404 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_276
timestamp 1606120350
transform 1 0 26496 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_288
timestamp 1606120350
transform 1 0 27600 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_300
timestamp 1606120350
transform 1 0 28704 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_312
timestamp 1606120350
transform 1 0 29808 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1606120350
transform 1 0 32016 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_324
timestamp 1606120350
transform 1 0 30912 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_337
timestamp 1606120350
transform 1 0 32108 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_349
timestamp 1606120350
transform 1 0 33212 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_361
timestamp 1606120350
transform 1 0 34316 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_373
timestamp 1606120350
transform 1 0 35420 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_385
timestamp 1606120350
transform 1 0 36524 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606120350
transform -1 0 38824 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1606120350
transform 1 0 37628 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_398
timestamp 1606120350
transform 1 0 37720 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_406
timestamp 1606120350
transform 1 0 38456 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606120350
transform 1 0 1104 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1606120350
transform 1 0 1380 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1606120350
transform 1 0 2484 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1606120350
transform 1 0 3588 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1606120350
transform 1 0 4692 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1606120350
transform 1 0 6716 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1606120350
transform 1 0 5796 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1606120350
transform 1 0 6532 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1606120350
transform 1 0 6808 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_74
timestamp 1606120350
transform 1 0 7912 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1606120350
transform 1 0 9016 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1606120350
transform 1 0 10120 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1606120350
transform 1 0 11224 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1084_
timestamp 1606120350
transform 1 0 13524 0 1 14688
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1606120350
transform 1 0 12328 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1084__D
timestamp 1606120350
transform 1 0 13340 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_123
timestamp 1606120350
transform 1 0 12420 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_131
timestamp 1606120350
transform 1 0 13156 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__A2
timestamp 1606120350
transform 1 0 15456 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_154
timestamp 1606120350
transform 1 0 15272 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_158
timestamp 1606120350
transform 1 0 15640 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0715_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 16008 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__A1
timestamp 1606120350
transform 1 0 15824 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__A1
timestamp 1606120350
transform 1 0 17756 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__B2
timestamp 1606120350
transform 1 0 17388 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_23_174
timestamp 1606120350
transform 1 0 17112 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_179
timestamp 1606120350
transform 1 0 17572 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0791_
timestamp 1606120350
transform 1 0 18032 0 1 14688
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1606120350
transform 1 0 17940 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_198
timestamp 1606120350
transform 1 0 19320 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__D
timestamp 1606120350
transform 1 0 20884 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1214__CLK
timestamp 1606120350
transform 1 0 21252 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_210
timestamp 1606120350
transform 1 0 20424 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_214
timestamp 1606120350
transform 1 0 20792 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_217
timestamp 1606120350
transform 1 0 21068 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_221
timestamp 1606120350
transform 1 0 21436 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1606120350
transform 1 0 23552 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_233
timestamp 1606120350
transform 1 0 22540 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_241
timestamp 1606120350
transform 1 0 23276 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_245
timestamp 1606120350
transform 1 0 23644 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_257
timestamp 1606120350
transform 1 0 24748 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_269
timestamp 1606120350
transform 1 0 25852 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_281
timestamp 1606120350
transform 1 0 26956 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_293
timestamp 1606120350
transform 1 0 28060 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1606120350
transform 1 0 29164 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_306
timestamp 1606120350
transform 1 0 29256 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_318
timestamp 1606120350
transform 1 0 30360 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_330
timestamp 1606120350
transform 1 0 31464 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_342
timestamp 1606120350
transform 1 0 32568 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_354
timestamp 1606120350
transform 1 0 33672 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1606120350
transform 1 0 34776 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_367
timestamp 1606120350
transform 1 0 34868 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_379
timestamp 1606120350
transform 1 0 35972 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606120350
transform -1 0 38824 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_391
timestamp 1606120350
transform 1 0 37076 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_403
timestamp 1606120350
transform 1 0 38180 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606120350
transform 1 0 1104 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__D
timestamp 1606120350
transform 1 0 1564 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_3
timestamp 1606120350
transform 1 0 1380 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_7
timestamp 1606120350
transform 1 0 1748 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_19
timestamp 1606120350
transform 1 0 2852 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1606120350
transform 1 0 3956 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1606120350
transform 1 0 4048 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1606120350
transform 1 0 5152 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_56
timestamp 1606120350
transform 1 0 6256 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_68
timestamp 1606120350
transform 1 0 7360 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_80
timestamp 1606120350
transform 1 0 8464 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1606120350
transform 1 0 9568 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1606120350
transform 1 0 9660 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1606120350
transform 1 0 10764 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1606120350
transform 1 0 11868 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1606120350
transform 1 0 12972 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1606120350
transform 1 0 15180 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1606120350
transform 1 0 14076 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_154
timestamp 1606120350
transform 1 0 15272 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0715__B1
timestamp 1606120350
transform 1 0 16008 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_164
timestamp 1606120350
transform 1 0 16192 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_176
timestamp 1606120350
transform 1 0 17296 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__B1
timestamp 1606120350
transform 1 0 18032 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0791__A2
timestamp 1606120350
transform 1 0 18400 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_186
timestamp 1606120350
transform 1 0 18216 0 -1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1606120350
transform 1 0 18584 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1606120350
transform 1 0 19688 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1214_
timestamp 1606120350
transform 1 0 20884 0 -1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1606120350
transform 1 0 20792 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_234
timestamp 1606120350
transform 1 0 22632 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_246
timestamp 1606120350
transform 1 0 23736 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_258
timestamp 1606120350
transform 1 0 24840 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_270
timestamp 1606120350
transform 1 0 25944 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_274
timestamp 1606120350
transform 1 0 26312 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1606120350
transform 1 0 26404 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_276
timestamp 1606120350
transform 1 0 26496 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_288
timestamp 1606120350
transform 1 0 27600 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_300
timestamp 1606120350
transform 1 0 28704 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_312
timestamp 1606120350
transform 1 0 29808 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1606120350
transform 1 0 32016 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_324
timestamp 1606120350
transform 1 0 30912 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_337
timestamp 1606120350
transform 1 0 32108 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_349
timestamp 1606120350
transform 1 0 33212 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_361
timestamp 1606120350
transform 1 0 34316 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_373
timestamp 1606120350
transform 1 0 35420 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_385
timestamp 1606120350
transform 1 0 36524 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606120350
transform -1 0 38824 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1606120350
transform 1 0 37628 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_398
timestamp 1606120350
transform 1 0 37720 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_406
timestamp 1606120350
transform 1 0 38456 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1219_
timestamp 1606120350
transform 1 0 1380 0 1 15776
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606120350
transform 1 0 1104 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_22
timestamp 1606120350
transform 1 0 3128 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_34
timestamp 1606120350
transform 1 0 4232 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1606120350
transform 1 0 6716 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_46
timestamp 1606120350
transform 1 0 5336 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_58
timestamp 1606120350
transform 1 0 6440 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1606120350
transform 1 0 6808 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_74
timestamp 1606120350
transform 1 0 7912 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_86
timestamp 1606120350
transform 1 0 9016 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_0_0_clk
timestamp 1606120350
transform 1 0 10028 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_0_0_clk_A
timestamp 1606120350
transform 1 0 10488 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_94
timestamp 1606120350
transform 1 0 9752 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_25_100
timestamp 1606120350
transform 1 0 10304 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_104
timestamp 1606120350
transform 1 0 10672 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1606120350
transform 1 0 12328 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__A1
timestamp 1606120350
transform 1 0 13340 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__B1
timestamp 1606120350
transform 1 0 13708 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_116
timestamp 1606120350
transform 1 0 11776 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_123
timestamp 1606120350
transform 1 0 12420 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_131
timestamp 1606120350
transform 1 0 13156 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_135
timestamp 1606120350
transform 1 0 13524 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0785_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 15180 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0785__A
timestamp 1606120350
transform 1 0 15640 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0666__A2
timestamp 1606120350
transform 1 0 14076 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_139
timestamp 1606120350
transform 1 0 13892 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_143
timestamp 1606120350
transform 1 0 14260 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_151
timestamp 1606120350
transform 1 0 14996 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_156
timestamp 1606120350
transform 1 0 15456 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__A1_N
timestamp 1606120350
transform 1 0 16744 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__B2
timestamp 1606120350
transform 1 0 17112 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__A2_N
timestamp 1606120350
transform 1 0 17480 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0790__B1
timestamp 1606120350
transform 1 0 16376 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_160
timestamp 1606120350
transform 1 0 15824 0 1 15776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_25_168
timestamp 1606120350
transform 1 0 16560 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_172
timestamp 1606120350
transform 1 0 16928 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_176
timestamp 1606120350
transform 1 0 17296 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_25_180
timestamp 1606120350
transform 1 0 17664 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1606120350
transform 1 0 17940 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1606120350
transform 1 0 18032 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1606120350
transform 1 0 19136 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1606120350
transform 1 0 20240 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_220
timestamp 1606120350
transform 1 0 21344 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1606120350
transform 1 0 23552 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__D
timestamp 1606120350
transform 1 0 23828 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1167__CLK
timestamp 1606120350
transform 1 0 24196 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_232
timestamp 1606120350
transform 1 0 22448 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_245
timestamp 1606120350
transform 1 0 23644 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_249
timestamp 1606120350
transform 1 0 24012 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_25_253
timestamp 1606120350
transform 1 0 24380 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_265
timestamp 1606120350
transform 1 0 25484 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_277
timestamp 1606120350
transform 1 0 26588 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_289
timestamp 1606120350
transform 1 0 27692 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1606120350
transform 1 0 29164 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_301
timestamp 1606120350
transform 1 0 28796 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_306
timestamp 1606120350
transform 1 0 29256 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_318
timestamp 1606120350
transform 1 0 30360 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_330
timestamp 1606120350
transform 1 0 31464 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_342
timestamp 1606120350
transform 1 0 32568 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_354
timestamp 1606120350
transform 1 0 33672 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1606120350
transform 1 0 34776 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_367
timestamp 1606120350
transform 1 0 34868 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_379
timestamp 1606120350
transform 1 0 35972 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606120350
transform -1 0 38824 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_391
timestamp 1606120350
transform 1 0 37076 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_403
timestamp 1606120350
transform 1 0 38180 0 1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606120350
transform 1 0 1104 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606120350
transform 1 0 1104 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1219__CLK
timestamp 1606120350
transform 1 0 1564 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_3
timestamp 1606120350
transform 1 0 1380 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_7
timestamp 1606120350
transform 1 0 1748 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_19
timestamp 1606120350
transform 1 0 2852 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1606120350
transform 1 0 1380 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1606120350
transform 1 0 2484 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1606120350
transform 1 0 3956 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1606120350
transform 1 0 4048 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1606120350
transform 1 0 5152 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_27
timestamp 1606120350
transform 1 0 3588 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_39
timestamp 1606120350
transform 1 0 4692 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1606120350
transform 1 0 6716 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1606120350
transform 1 0 6256 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1606120350
transform 1 0 7360 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_51
timestamp 1606120350
transform 1 0 5796 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_59
timestamp 1606120350
transform 1 0 6532 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1606120350
transform 1 0 6808 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_0_0_clk
timestamp 1606120350
transform 1 0 8372 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_0_0_clk_A
timestamp 1606120350
transform 1 0 8832 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1606120350
transform 1 0 8464 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_74
timestamp 1606120350
transform 1 0 7912 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_78
timestamp 1606120350
transform 1 0 8280 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_82
timestamp 1606120350
transform 1 0 8648 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_86
timestamp 1606120350
transform 1 0 9016 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1606120350
transform 1 0 9568 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__B2
timestamp 1606120350
transform 1 0 11592 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1606120350
transform 1 0 9660 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1606120350
transform 1 0 10764 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_98
timestamp 1606120350
transform 1 0 10120 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_110
timestamp 1606120350
transform 1 0 11224 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_123
timestamp 1606120350
transform 1 0 12420 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_120
timestamp 1606120350
transform 1 0 12144 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_116
timestamp 1606120350
transform 1 0 11776 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_120
timestamp 1606120350
transform 1 0 12144 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_117
timestamp 1606120350
transform 1 0 11868 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__A2
timestamp 1606120350
transform 1 0 11960 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__A1
timestamp 1606120350
transform 1 0 12604 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0817__B1
timestamp 1606120350
transform 1 0 11960 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1606120350
transform 1 0 12328 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_127
timestamp 1606120350
transform 1 0 12788 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_130
timestamp 1606120350
transform 1 0 13064 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__D
timestamp 1606120350
transform 1 0 12880 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1083_
timestamp 1606120350
transform 1 0 12880 0 1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__a21o_4  _0666_
timestamp 1606120350
transform 1 0 13340 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_147
timestamp 1606120350
transform 1 0 14628 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_145
timestamp 1606120350
transform 1 0 14444 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_155
timestamp 1606120350
transform 1 0 15364 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_151
timestamp 1606120350
transform 1 0 14996 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_26_158
timestamp 1606120350
transform 1 0 15640 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_154
timestamp 1606120350
transform 1 0 15272 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0665__A
timestamp 1606120350
transform 1 0 14812 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__B1
timestamp 1606120350
transform 1 0 15732 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0665__B
timestamp 1606120350
transform 1 0 15180 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__A1_N
timestamp 1606120350
transform 1 0 15548 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1606120350
transform 1 0 15180 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0788_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 15732 0 1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__a2bb2o_4  _0790_
timestamp 1606120350
transform 1 0 16744 0 -1 16864
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__A1_N
timestamp 1606120350
transform 1 0 17388 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__B2
timestamp 1606120350
transform 1 0 17756 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__B2
timestamp 1606120350
transform 1 0 16100 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_26_161
timestamp 1606120350
transform 1 0 15916 0 -1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_165
timestamp 1606120350
transform 1 0 16284 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_169
timestamp 1606120350
transform 1 0 16652 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_175
timestamp 1606120350
transform 1 0 17204 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_179
timestamp 1606120350
transform 1 0 17572 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_27_192
timestamp 1606120350
transform 1 0 18768 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_27_188
timestamp 1606120350
transform 1 0 18400 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_184
timestamp 1606120350
transform 1 0 18032 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__B1
timestamp 1606120350
transform 1 0 18584 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0795__A2_N
timestamp 1606120350
transform 1 0 18216 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1606120350
transform 1 0 17940 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0575__A
timestamp 1606120350
transform 1 0 19044 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_197
timestamp 1606120350
transform 1 0 19228 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_198
timestamp 1606120350
transform 1 0 19320 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_186
timestamp 1606120350
transform 1 0 18216 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1606120350
transform 1 0 20792 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_210
timestamp 1606120350
transform 1 0 20424 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1606120350
transform 1 0 20884 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_227
timestamp 1606120350
transform 1 0 21988 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_209
timestamp 1606120350
transform 1 0 20332 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_221
timestamp 1606120350
transform 1 0 21436 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1167_
timestamp 1606120350
transform 1 0 23644 0 -1 16864
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1606120350
transform 1 0 23552 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_239
timestamp 1606120350
transform 1 0 23092 0 -1 16864
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_233
timestamp 1606120350
transform 1 0 22540 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_241
timestamp 1606120350
transform 1 0 23276 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_245
timestamp 1606120350
transform 1 0 23644 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_264
timestamp 1606120350
transform 1 0 25392 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_272
timestamp 1606120350
transform 1 0 26128 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_257
timestamp 1606120350
transform 1 0 24748 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_269
timestamp 1606120350
transform 1 0 25852 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1606120350
transform 1 0 26404 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_276
timestamp 1606120350
transform 1 0 26496 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_288
timestamp 1606120350
transform 1 0 27600 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1606120350
transform 1 0 26956 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1606120350
transform 1 0 28060 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1606120350
transform 1 0 29164 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_300
timestamp 1606120350
transform 1 0 28704 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_312
timestamp 1606120350
transform 1 0 29808 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_306
timestamp 1606120350
transform 1 0 29256 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_318
timestamp 1606120350
transform 1 0 30360 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1606120350
transform 1 0 32016 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_324
timestamp 1606120350
transform 1 0 30912 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_337
timestamp 1606120350
transform 1 0 32108 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_330
timestamp 1606120350
transform 1 0 31464 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_342
timestamp 1606120350
transform 1 0 32568 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_349
timestamp 1606120350
transform 1 0 33212 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_361
timestamp 1606120350
transform 1 0 34316 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_354
timestamp 1606120350
transform 1 0 33672 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1606120350
transform 1 0 34776 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_373
timestamp 1606120350
transform 1 0 35420 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_385
timestamp 1606120350
transform 1 0 36524 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_367
timestamp 1606120350
transform 1 0 34868 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_379
timestamp 1606120350
transform 1 0 35972 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606120350
transform -1 0 38824 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606120350
transform -1 0 38824 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1606120350
transform 1 0 37628 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_398
timestamp 1606120350
transform 1 0 37720 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_406
timestamp 1606120350
transform 1 0 38456 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_391
timestamp 1606120350
transform 1 0 37076 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_403
timestamp 1606120350
transform 1 0 38180 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1606120350
transform 1 0 1104 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1606120350
transform 1 0 1380 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1606120350
transform 1 0 2484 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1606120350
transform 1 0 3956 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1606120350
transform 1 0 3588 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1606120350
transform 1 0 4048 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1606120350
transform 1 0 5152 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1606120350
transform 1 0 6256 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1606120350
transform 1 0 7360 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1606120350
transform 1 0 8464 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1606120350
transform 1 0 9568 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__A2
timestamp 1606120350
transform 1 0 11408 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__CLK
timestamp 1606120350
transform 1 0 9844 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_93
timestamp 1606120350
transform 1 0 9660 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_97
timestamp 1606120350
transform 1 0 10028 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_109
timestamp 1606120350
transform 1 0 11132 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_114
timestamp 1606120350
transform 1 0 11592 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0817_
timestamp 1606120350
transform 1 0 11960 0 -1 17952
box -38 -48 1326 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__A1
timestamp 1606120350
transform 1 0 11776 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1083__CLK
timestamp 1606120350
transform 1 0 13432 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_132
timestamp 1606120350
transform 1 0 13248 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_136
timestamp 1606120350
transform 1 0 13616 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _0665_
timestamp 1606120350
transform 1 0 15272 0 -1 17952
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1606120350
transform 1 0 15180 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__A2
timestamp 1606120350
transform 1 0 14904 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_148
timestamp 1606120350
transform 1 0 14720 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_152
timestamp 1606120350
transform 1 0 15088 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _0795_
timestamp 1606120350
transform 1 0 16836 0 -1 17952
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0788__A2_N
timestamp 1606120350
transform 1 0 16100 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_161
timestamp 1606120350
transform 1 0 15916 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_28_165
timestamp 1606120350
transform 1 0 16284 0 -1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__inv_8  _0575_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 19044 0 -1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0568__A1
timestamp 1606120350
transform 1 0 18492 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0568__B1
timestamp 1606120350
transform 1 0 18860 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_187
timestamp 1606120350
transform 1 0 18308 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_28_191
timestamp 1606120350
transform 1 0 18676 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_204
timestamp 1606120350
transform 1 0 19872 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1606120350
transform 1 0 20792 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_212
timestamp 1606120350
transform 1 0 20608 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1606120350
transform 1 0 20884 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1606120350
transform 1 0 21988 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1606120350
transform 1 0 23092 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_251
timestamp 1606120350
transform 1 0 24196 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_263
timestamp 1606120350
transform 1 0 25300 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1606120350
transform 1 0 26404 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_276
timestamp 1606120350
transform 1 0 26496 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_288
timestamp 1606120350
transform 1 0 27600 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_300
timestamp 1606120350
transform 1 0 28704 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_312
timestamp 1606120350
transform 1 0 29808 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1606120350
transform 1 0 32016 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_324
timestamp 1606120350
transform 1 0 30912 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_337
timestamp 1606120350
transform 1 0 32108 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_349
timestamp 1606120350
transform 1 0 33212 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_361
timestamp 1606120350
transform 1 0 34316 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_373
timestamp 1606120350
transform 1 0 35420 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_385
timestamp 1606120350
transform 1 0 36524 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1606120350
transform -1 0 38824 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1606120350
transform 1 0 37628 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_398
timestamp 1606120350
transform 1 0 37720 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_406
timestamp 1606120350
transform 1 0 38456 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1606120350
transform 1 0 1104 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1606120350
transform 1 0 1380 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1606120350
transform 1 0 2484 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1606120350
transform 1 0 3588 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1606120350
transform 1 0 4692 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1606120350
transform 1 0 6716 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1606120350
transform 1 0 5796 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1606120350
transform 1 0 6532 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1606120350
transform 1 0 6808 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_74
timestamp 1606120350
transform 1 0 7912 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_86
timestamp 1606120350
transform 1 0 9016 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _1129_
timestamp 1606120350
transform 1 0 9844 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1129__D
timestamp 1606120350
transform 1 0 9660 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_29_92
timestamp 1606120350
transform 1 0 9568 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_29_114
timestamp 1606120350
transform 1 0 11592 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1110_
timestamp 1606120350
transform 1 0 12420 0 1 17952
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1606120350
transform 1 0 12328 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__B1
timestamp 1606120350
transform 1 0 11868 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_119
timestamp 1606120350
transform 1 0 12052 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_4  _0784_
timestamp 1606120350
transform 1 0 14904 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__A1
timestamp 1606120350
transform 1 0 14720 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0691__A
timestamp 1606120350
transform 1 0 14352 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_142
timestamp 1606120350
transform 1 0 14168 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_146
timestamp 1606120350
transform 1 0 14536 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_162
timestamp 1606120350
transform 1 0 16008 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_166
timestamp 1606120350
transform 1 0 16376 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__A1
timestamp 1606120350
transform 1 0 16192 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_170
timestamp 1606120350
transform 1 0 16744 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__A2
timestamp 1606120350
transform 1 0 16560 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_174
timestamp 1606120350
transform 1 0 17112 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0793__B1
timestamp 1606120350
transform 1 0 16928 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_29_178
timestamp 1606120350
transform 1 0 17480 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0787__A
timestamp 1606120350
transform 1 0 17296 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0568__A2
timestamp 1606120350
transform 1 0 17756 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0604_
timestamp 1606120350
transform 1 0 18676 0 1 17952
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1606120350
transform 1 0 17940 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0604__A
timestamp 1606120350
transform 1 0 18492 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_184
timestamp 1606120350
transform 1 0 18032 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_188
timestamp 1606120350
transform 1 0 18400 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_200
timestamp 1606120350
transform 1 0 19504 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_212
timestamp 1606120350
transform 1 0 20608 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_224
timestamp 1606120350
transform 1 0 21712 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1606120350
transform 1 0 23552 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__D
timestamp 1606120350
transform 1 0 22448 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1142__CLK
timestamp 1606120350
transform 1 0 22816 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_234
timestamp 1606120350
transform 1 0 22632 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_238
timestamp 1606120350
transform 1 0 23000 0 1 17952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_245
timestamp 1606120350
transform 1 0 23644 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_257
timestamp 1606120350
transform 1 0 24748 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_269
timestamp 1606120350
transform 1 0 25852 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1606120350
transform 1 0 26956 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_293
timestamp 1606120350
transform 1 0 28060 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1606120350
transform 1 0 29164 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_306
timestamp 1606120350
transform 1 0 29256 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_318
timestamp 1606120350
transform 1 0 30360 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_330
timestamp 1606120350
transform 1 0 31464 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_342
timestamp 1606120350
transform 1 0 32568 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_354
timestamp 1606120350
transform 1 0 33672 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1606120350
transform 1 0 34776 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_367
timestamp 1606120350
transform 1 0 34868 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_379
timestamp 1606120350
transform 1 0 35972 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1606120350
transform -1 0 38824 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_391
timestamp 1606120350
transform 1 0 37076 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_403
timestamp 1606120350
transform 1 0 38180 0 1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1606120350
transform 1 0 1104 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1606120350
transform 1 0 1380 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1606120350
transform 1 0 2484 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1606120350
transform 1 0 3956 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1606120350
transform 1 0 3588 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1606120350
transform 1 0 4048 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1606120350
transform 1 0 5152 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1606120350
transform 1 0 6256 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1606120350
transform 1 0 7360 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1606120350
transform 1 0 8464 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1606120350
transform 1 0 9568 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1606120350
transform 1 0 9660 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_105
timestamp 1606120350
transform 1 0 10764 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_113
timestamp 1606120350
transform 1 0 11500 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0816_
timestamp 1606120350
transform 1 0 11868 0 -1 19040
box -38 -48 1326 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0816__B2
timestamp 1606120350
transform 1 0 11684 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__D
timestamp 1606120350
transform 1 0 13340 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1110__CLK
timestamp 1606120350
transform 1 0 13708 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_131
timestamp 1606120350
transform 1 0 13156 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_135
timestamp 1606120350
transform 1 0 13524 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0691_
timestamp 1606120350
transform 1 0 13984 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_4  _0793_
timestamp 1606120350
transform 1 0 15456 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1606120350
transform 1 0 15180 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0784__B1
timestamp 1606120350
transform 1 0 14904 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1606120350
transform 1 0 13892 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_143
timestamp 1606120350
transform 1 0 14260 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_149
timestamp 1606120350
transform 1 0 14812 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_30_152
timestamp 1606120350
transform 1 0 15088 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_154
timestamp 1606120350
transform 1 0 15272 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0787_
timestamp 1606120350
transform 1 0 17296 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0560__A
timestamp 1606120350
transform 1 0 16744 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0559__B1
timestamp 1606120350
transform 1 0 17756 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_30_168
timestamp 1606120350
transform 1 0 16560 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_172
timestamp 1606120350
transform 1 0 16928 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_30_179
timestamp 1606120350
transform 1 0 17572 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _0568_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 18492 0 -1 19040
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__B1
timestamp 1606120350
transform 1 0 18308 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_183
timestamp 1606120350
transform 1 0 17940 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_202
timestamp 1606120350
transform 1 0 19688 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1606120350
transform 1 0 20792 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1606120350
transform 1 0 20884 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_227
timestamp 1606120350
transform 1 0 21988 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1142_
timestamp 1606120350
transform 1 0 22448 0 -1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_30_231
timestamp 1606120350
transform 1 0 22356 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_251
timestamp 1606120350
transform 1 0 24196 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_263
timestamp 1606120350
transform 1 0 25300 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1606120350
transform 1 0 26404 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_276
timestamp 1606120350
transform 1 0 26496 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_288
timestamp 1606120350
transform 1 0 27600 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__CLK
timestamp 1606120350
transform 1 0 30084 0 -1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_300
timestamp 1606120350
transform 1 0 28704 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_312
timestamp 1606120350
transform 1 0 29808 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_317
timestamp 1606120350
transform 1 0 30268 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1606120350
transform 1 0 32016 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_329
timestamp 1606120350
transform 1 0 31372 0 -1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_335
timestamp 1606120350
transform 1 0 31924 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_337
timestamp 1606120350
transform 1 0 32108 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_349
timestamp 1606120350
transform 1 0 33212 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_361
timestamp 1606120350
transform 1 0 34316 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_373
timestamp 1606120350
transform 1 0 35420 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_385
timestamp 1606120350
transform 1 0 36524 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1606120350
transform -1 0 38824 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1606120350
transform 1 0 37628 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_398
timestamp 1606120350
transform 1 0 37720 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_406
timestamp 1606120350
transform 1 0 38456 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1606120350
transform 1 0 1104 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1606120350
transform 1 0 1380 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1606120350
transform 1 0 2484 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__D
timestamp 1606120350
transform 1 0 4416 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1137__CLK
timestamp 1606120350
transform 1 0 4784 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_27
timestamp 1606120350
transform 1 0 3588 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_35
timestamp 1606120350
transform 1 0 4324 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_38
timestamp 1606120350
transform 1 0 4600 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_42
timestamp 1606120350
transform 1 0 4968 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1606120350
transform 1 0 6716 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_54
timestamp 1606120350
transform 1 0 6072 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_60
timestamp 1606120350
transform 1 0 6624 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1606120350
transform 1 0 6808 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_74
timestamp 1606120350
transform 1 0 7912 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_86
timestamp 1606120350
transform 1 0 9016 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_98
timestamp 1606120350
transform 1 0 10120 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_110
timestamp 1606120350
transform 1 0 11224 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1109_
timestamp 1606120350
transform 1 0 12420 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1606120350
transform 1 0 12328 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__D
timestamp 1606120350
transform 1 0 12144 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_118
timestamp 1606120350
transform 1 0 11960 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0783_
timestamp 1606120350
transform 1 0 14904 0 1 19040
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__B
timestamp 1606120350
transform 1 0 14720 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0637__A
timestamp 1606120350
transform 1 0 14352 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_142
timestamp 1606120350
transform 1 0 14168 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_146
timestamp 1606120350
transform 1 0 14536 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_157
timestamp 1606120350
transform 1 0 15548 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  _0560_
timestamp 1606120350
transform 1 0 16376 0 1 19040
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__B
timestamp 1606120350
transform 1 0 15916 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0559__A1_N
timestamp 1606120350
transform 1 0 17388 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0559__A2_N
timestamp 1606120350
transform 1 0 17756 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_163
timestamp 1606120350
transform 1 0 16100 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_31_175
timestamp 1606120350
transform 1 0 17204 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_179
timestamp 1606120350
transform 1 0 17572 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0605_
timestamp 1606120350
transform 1 0 18860 0 1 19040
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1606120350
transform 1 0 17940 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0559__B2
timestamp 1606120350
transform 1 0 18216 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__A2_N
timestamp 1606120350
transform 1 0 18676 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_184
timestamp 1606120350
transform 1 0 18032 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_31_188
timestamp 1606120350
transform 1 0 18400 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0557__A
timestamp 1606120350
transform 1 0 20884 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__B2
timestamp 1606120350
transform 1 0 20516 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_209
timestamp 1606120350
transform 1 0 20332 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_31_213
timestamp 1606120350
transform 1 0 20700 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_217
timestamp 1606120350
transform 1 0 21068 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1606120350
transform 1 0 23552 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_229
timestamp 1606120350
transform 1 0 22172 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_241
timestamp 1606120350
transform 1 0 23276 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_245
timestamp 1606120350
transform 1 0 23644 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_257
timestamp 1606120350
transform 1 0 24748 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_269
timestamp 1606120350
transform 1 0 25852 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1606120350
transform 1 0 26956 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_293
timestamp 1606120350
transform 1 0 28060 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1144_
timestamp 1606120350
transform 1 0 30084 0 1 19040
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1606120350
transform 1 0 29164 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1144__D
timestamp 1606120350
transform 1 0 29900 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_306
timestamp 1606120350
transform 1 0 29256 0 1 19040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_312
timestamp 1606120350
transform 1 0 29808 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_334
timestamp 1606120350
transform 1 0 31832 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_346
timestamp 1606120350
transform 1 0 32936 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_358
timestamp 1606120350
transform 1 0 34040 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1606120350
transform 1 0 34776 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_367
timestamp 1606120350
transform 1 0 34868 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_379
timestamp 1606120350
transform 1 0 35972 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1606120350
transform -1 0 38824 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_391
timestamp 1606120350
transform 1 0 37076 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_403
timestamp 1606120350
transform 1 0 38180 0 1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1606120350
transform 1 0 1104 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1606120350
transform 1 0 1380 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1606120350
transform 1 0 2484 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1137_
timestamp 1606120350
transform 1 0 4416 0 -1 20128
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1606120350
transform 1 0 3956 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1606120350
transform 1 0 3588 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_32
timestamp 1606120350
transform 1 0 4048 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_55
timestamp 1606120350
transform 1 0 6164 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_67
timestamp 1606120350
transform 1 0 7268 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_79
timestamp 1606120350
transform 1 0 8372 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_91
timestamp 1606120350
transform 1 0 9476 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1606120350
transform 1 0 9568 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1606120350
transform 1 0 9660 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1606120350
transform 1 0 10764 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0637_
timestamp 1606120350
transform 1 0 13708 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1109__CLK
timestamp 1606120350
transform 1 0 12420 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_117
timestamp 1606120350
transform 1 0 11868 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_32_125
timestamp 1606120350
transform 1 0 12604 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1606120350
transform 1 0 15180 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0783__A
timestamp 1606120350
transform 1 0 14904 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_140
timestamp 1606120350
transform 1 0 13984 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_148
timestamp 1606120350
transform 1 0 14720 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_152
timestamp 1606120350
transform 1 0 15088 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_154
timestamp 1606120350
transform 1 0 15272 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_4  _0559_
timestamp 1606120350
transform 1 0 17388 0 -1 20128
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_4  _0792_
timestamp 1606120350
transform 1 0 15916 0 -1 20128
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0792__A
timestamp 1606120350
transform 1 0 16744 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0603__A
timestamp 1606120350
transform 1 0 17204 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_160
timestamp 1606120350
transform 1 0 15824 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_168
timestamp 1606120350
transform 1 0 16560 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_32_172
timestamp 1606120350
transform 1 0 16928 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0577__A2_N
timestamp 1606120350
transform 1 0 19044 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0605__A1_N
timestamp 1606120350
transform 1 0 19412 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_193
timestamp 1606120350
transform 1 0 18860 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_197
timestamp 1606120350
transform 1 0 19228 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_32_201
timestamp 1606120350
transform 1 0 19596 0 -1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0557_
timestamp 1606120350
transform 1 0 20884 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1606120350
transform 1 0 20792 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0562__A
timestamp 1606120350
transform 1 0 21344 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0578__B
timestamp 1606120350
transform 1 0 20148 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0578__D
timestamp 1606120350
transform 1 0 20516 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_32_209
timestamp 1606120350
transform 1 0 20332 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_213
timestamp 1606120350
transform 1 0 20700 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_218
timestamp 1606120350
transform 1 0 21160 0 -1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_222
timestamp 1606120350
transform 1 0 21528 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_234
timestamp 1606120350
transform 1 0 22632 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_246
timestamp 1606120350
transform 1 0 23736 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_258
timestamp 1606120350
transform 1 0 24840 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_270
timestamp 1606120350
transform 1 0 25944 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_274
timestamp 1606120350
transform 1 0 26312 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1606120350
transform 1 0 26404 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_276
timestamp 1606120350
transform 1 0 26496 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_288
timestamp 1606120350
transform 1 0 27600 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_300
timestamp 1606120350
transform 1 0 28704 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_312
timestamp 1606120350
transform 1 0 29808 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1606120350
transform 1 0 32016 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_324
timestamp 1606120350
transform 1 0 30912 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_337
timestamp 1606120350
transform 1 0 32108 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_349
timestamp 1606120350
transform 1 0 33212 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_361
timestamp 1606120350
transform 1 0 34316 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_373
timestamp 1606120350
transform 1 0 35420 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_385
timestamp 1606120350
transform 1 0 36524 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1606120350
transform -1 0 38824 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1606120350
transform 1 0 37628 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_398
timestamp 1606120350
transform 1 0 37720 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_406
timestamp 1606120350
transform 1 0 38456 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1606120350
transform 1 0 1104 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1606120350
transform 1 0 1104 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1606120350
transform 1 0 1380 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1606120350
transform 1 0 2484 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1606120350
transform 1 0 1380 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1606120350
transform 1 0 2484 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1606120350
transform 1 0 3956 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1606120350
transform 1 0 3588 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1606120350
transform 1 0 4692 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1606120350
transform 1 0 3588 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1606120350
transform 1 0 4048 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1606120350
transform 1 0 5152 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1606120350
transform 1 0 6716 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_51
timestamp 1606120350
transform 1 0 5796 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_59
timestamp 1606120350
transform 1 0 6532 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1606120350
transform 1 0 6808 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1606120350
transform 1 0 6256 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1606120350
transform 1 0 7360 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_74
timestamp 1606120350
transform 1 0 7912 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_86
timestamp 1606120350
transform 1 0 9016 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1606120350
transform 1 0 8464 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1606120350
transform 1 0 9568 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_98
timestamp 1606120350
transform 1 0 10120 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_110
timestamp 1606120350
transform 1 0 11224 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_114
timestamp 1606120350
transform 1 0 11592 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1606120350
transform 1 0 9660 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_105
timestamp 1606120350
transform 1 0 10764 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_113
timestamp 1606120350
transform 1 0 11500 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_123
timestamp 1606120350
transform 1 0 12420 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_121
timestamp 1606120350
transform 1 0 12236 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_117
timestamp 1606120350
transform 1 0 11868 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__CLK
timestamp 1606120350
transform 1 0 12052 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1112__D
timestamp 1606120350
transform 1 0 11684 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1606120350
transform 1 0 12328 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_136
timestamp 1606120350
transform 1 0 13616 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_131
timestamp 1606120350
transform 1 0 13156 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0678_
timestamp 1606120350
transform 1 0 13340 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_134
timestamp 1606120350
transform 1 0 13432 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1112_
timestamp 1606120350
transform 1 0 11684 0 -1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__buf_1  _0667_
timestamp 1606120350
transform 1 0 15364 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1606120350
transform 1 0 15180 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0678__A
timestamp 1606120350
transform 1 0 13800 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_140
timestamp 1606120350
transform 1 0 13984 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_152
timestamp 1606120350
transform 1 0 15088 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_33_158
timestamp 1606120350
transform 1 0 15640 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_34_146
timestamp 1606120350
transform 1 0 14536 0 -1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_152
timestamp 1606120350
transform 1 0 15088 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1606120350
transform 1 0 15272 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_168
timestamp 1606120350
transform 1 0 16560 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_162
timestamp 1606120350
transform 1 0 16008 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0614__A
timestamp 1606120350
transform 1 0 16192 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__A
timestamp 1606120350
transform 1 0 16376 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0667__A
timestamp 1606120350
transform 1 0 15824 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0614_
timestamp 1606120350
transform 1 0 16376 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_34_172
timestamp 1606120350
transform 1 0 16928 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_179
timestamp 1606120350
transform 1 0 17572 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_175
timestamp 1606120350
transform 1 0 17204 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0554__A
timestamp 1606120350
transform 1 0 17388 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__B1
timestamp 1606120350
transform 1 0 16744 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0554_
timestamp 1606120350
transform 1 0 17020 0 -1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_34_182
timestamp 1606120350
transform 1 0 17848 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0577__A1_N
timestamp 1606120350
transform 1 0 17756 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_186
timestamp 1606120350
transform 1 0 18216 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_33_193
timestamp 1606120350
transform 1 0 18860 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__A1
timestamp 1606120350
transform 1 0 18400 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0633__A
timestamp 1606120350
transform 1 0 18032 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1606120350
transform 1 0 17940 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0603_
timestamp 1606120350
transform 1 0 18032 0 1 20128
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_33_201
timestamp 1606120350
transform 1 0 19596 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_33_197
timestamp 1606120350
transform 1 0 19228 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0578__A
timestamp 1606120350
transform 1 0 19964 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0577__B2
timestamp 1606120350
transform 1 0 19412 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0577__B1
timestamp 1606120350
transform 1 0 19044 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0577_
timestamp 1606120350
transform 1 0 18584 0 -1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_34_210
timestamp 1606120350
transform 1 0 20424 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_34_206
timestamp 1606120350
transform 1 0 20056 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0615__A1_N
timestamp 1606120350
transform 1 0 20608 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0578__C
timestamp 1606120350
transform 1 0 20240 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1606120350
transform 1 0 20792 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0562_
timestamp 1606120350
transform 1 0 20884 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_34_218
timestamp 1606120350
transform 1 0 21160 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0607__A
timestamp 1606120350
transform 1 0 21344 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_222
timestamp 1606120350
transform 1 0 21528 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_224
timestamp 1606120350
transform 1 0 21712 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__nor4_4  _0578_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 20148 0 1 20128
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1606120350
transform 1 0 23552 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_236
timestamp 1606120350
transform 1 0 22816 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_245
timestamp 1606120350
transform 1 0 23644 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_234
timestamp 1606120350
transform 1 0 22632 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_246
timestamp 1606120350
transform 1 0 23736 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__CLK
timestamp 1606120350
transform 1 0 24840 0 -1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_257
timestamp 1606120350
transform 1 0 24748 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_269
timestamp 1606120350
transform 1 0 25852 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_260
timestamp 1606120350
transform 1 0 25024 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_272
timestamp 1606120350
transform 1 0 26128 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1606120350
transform 1 0 26404 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1606120350
transform 1 0 26956 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_293
timestamp 1606120350
transform 1 0 28060 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_276
timestamp 1606120350
transform 1 0 26496 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_288
timestamp 1606120350
transform 1 0 27600 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1606120350
transform 1 0 29164 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_306
timestamp 1606120350
transform 1 0 29256 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_318
timestamp 1606120350
transform 1 0 30360 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_300
timestamp 1606120350
transform 1 0 28704 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_312
timestamp 1606120350
transform 1 0 29808 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1606120350
transform 1 0 32016 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_330
timestamp 1606120350
transform 1 0 31464 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_342
timestamp 1606120350
transform 1 0 32568 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_324
timestamp 1606120350
transform 1 0 30912 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_337
timestamp 1606120350
transform 1 0 32108 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_354
timestamp 1606120350
transform 1 0 33672 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_349
timestamp 1606120350
transform 1 0 33212 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_361
timestamp 1606120350
transform 1 0 34316 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1606120350
transform 1 0 34776 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_367
timestamp 1606120350
transform 1 0 34868 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_379
timestamp 1606120350
transform 1 0 35972 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_373
timestamp 1606120350
transform 1 0 35420 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_385
timestamp 1606120350
transform 1 0 36524 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1606120350
transform -1 0 38824 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1606120350
transform -1 0 38824 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1606120350
transform 1 0 37628 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_391
timestamp 1606120350
transform 1 0 37076 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_403
timestamp 1606120350
transform 1 0 38180 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_398
timestamp 1606120350
transform 1 0 37720 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_406
timestamp 1606120350
transform 1 0 38456 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1606120350
transform 1 0 1104 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1606120350
transform 1 0 1380 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1606120350
transform 1 0 2484 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1606120350
transform 1 0 3588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1606120350
transform 1 0 4692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1606120350
transform 1 0 6716 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_51
timestamp 1606120350
transform 1 0 5796 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1606120350
transform 1 0 6532 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1606120350
transform 1 0 6808 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_74
timestamp 1606120350
transform 1 0 7912 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_86
timestamp 1606120350
transform 1 0 9016 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__B1
timestamp 1606120350
transform 1 0 11592 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__B2
timestamp 1606120350
transform 1 0 11224 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__A2
timestamp 1606120350
transform 1 0 10856 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_98
timestamp 1606120350
transform 1 0 10120 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_108
timestamp 1606120350
transform 1 0 11040 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_112
timestamp 1606120350
transform 1 0 11408 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1606120350
transform 1 0 12328 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0819__A1
timestamp 1606120350
transform 1 0 11960 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__CLK
timestamp 1606120350
transform 1 0 13616 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_116
timestamp 1606120350
transform 1 0 11776 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_120
timestamp 1606120350
transform 1 0 12144 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_123
timestamp 1606120350
transform 1 0 12420 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_135
timestamp 1606120350
transform 1 0 13524 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0801__A
timestamp 1606120350
transform 1 0 14168 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0692__A
timestamp 1606120350
transform 1 0 15640 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_138
timestamp 1606120350
transform 1 0 13800 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_144
timestamp 1606120350
transform 1 0 14352 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_156
timestamp 1606120350
transform 1 0 15456 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0639_
timestamp 1606120350
transform 1 0 16560 0 1 21216
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0692__B
timestamp 1606120350
transform 1 0 16008 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0627__A
timestamp 1606120350
transform 1 0 17756 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0633__B
timestamp 1606120350
transform 1 0 17388 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0639__B
timestamp 1606120350
transform 1 0 16376 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_160
timestamp 1606120350
transform 1 0 15824 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_164
timestamp 1606120350
transform 1 0 16192 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_175
timestamp 1606120350
transform 1 0 17204 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_179
timestamp 1606120350
transform 1 0 17572 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0615_
timestamp 1606120350
transform 1 0 19688 0 1 21216
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_8  _0627_
timestamp 1606120350
transform 1 0 18124 0 1 21216
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1606120350
transform 1 0 17940 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0607__B
timestamp 1606120350
transform 1 0 19136 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0615__B2
timestamp 1606120350
transform 1 0 19504 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_184
timestamp 1606120350
transform 1 0 18032 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_194
timestamp 1606120350
transform 1 0 18952 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_198
timestamp 1606120350
transform 1 0 19320 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0608__B
timestamp 1606120350
transform 1 0 21344 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0608__A
timestamp 1606120350
transform 1 0 21712 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0615__B1
timestamp 1606120350
transform 1 0 22080 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_218
timestamp 1606120350
transform 1 0 21160 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_222
timestamp 1606120350
transform 1 0 21528 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_35_226
timestamp 1606120350
transform 1 0 21896 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1606120350
transform 1 0 23552 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__D
timestamp 1606120350
transform 1 0 23092 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1135__CLK
timestamp 1606120350
transform 1 0 23828 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_230
timestamp 1606120350
transform 1 0 22264 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_238
timestamp 1606120350
transform 1 0 23000 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_241
timestamp 1606120350
transform 1 0 23276 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_35_245
timestamp 1606120350
transform 1 0 23644 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_35_249
timestamp 1606120350
transform 1 0 24012 0 1 21216
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _1175_
timestamp 1606120350
transform 1 0 24840 0 1 21216
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1175__D
timestamp 1606120350
transform 1 0 24656 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_35_255
timestamp 1606120350
transform 1 0 24564 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_277
timestamp 1606120350
transform 1 0 26588 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_289
timestamp 1606120350
transform 1 0 27692 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1606120350
transform 1 0 29164 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_301
timestamp 1606120350
transform 1 0 28796 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_306
timestamp 1606120350
transform 1 0 29256 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_318
timestamp 1606120350
transform 1 0 30360 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_330
timestamp 1606120350
transform 1 0 31464 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_342
timestamp 1606120350
transform 1 0 32568 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_354
timestamp 1606120350
transform 1 0 33672 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1606120350
transform 1 0 34776 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_367
timestamp 1606120350
transform 1 0 34868 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_379
timestamp 1606120350
transform 1 0 35972 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1606120350
transform -1 0 38824 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_391
timestamp 1606120350
transform 1 0 37076 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_403
timestamp 1606120350
transform 1 0 38180 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1606120350
transform 1 0 1104 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__D
timestamp 1606120350
transform 1 0 1564 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_3
timestamp 1606120350
transform 1 0 1380 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_7
timestamp 1606120350
transform 1 0 1748 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_19
timestamp 1606120350
transform 1 0 2852 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1606120350
transform 1 0 3956 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1606120350
transform 1 0 4048 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1606120350
transform 1 0 5152 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_56
timestamp 1606120350
transform 1 0 6256 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_68
timestamp 1606120350
transform 1 0 7360 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_80
timestamp 1606120350
transform 1 0 8464 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _0819_
timestamp 1606120350
transform 1 0 11592 0 -1 22304
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1606120350
transform 1 0 9568 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_93
timestamp 1606120350
transform 1 0 9660 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_105
timestamp 1606120350
transform 1 0 10764 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_113
timestamp 1606120350
transform 1 0 11500 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__A1
timestamp 1606120350
transform 1 0 13156 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__A2
timestamp 1606120350
transform 1 0 13524 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_128
timestamp 1606120350
transform 1 0 12880 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_133
timestamp 1606120350
transform 1 0 13340 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_137
timestamp 1606120350
transform 1 0 13708 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1103__D
timestamp 1606120350
transform 1 0 13892 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_36_141
timestamp 1606120350
transform 1 0 14076 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0801_
timestamp 1606120350
transform 1 0 14168 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_145
timestamp 1606120350
transform 1 0 14444 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__D
timestamp 1606120350
transform 1 0 14628 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_149
timestamp 1606120350
transform 1 0 14812 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__A
timestamp 1606120350
transform 1 0 14996 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_154
timestamp 1606120350
transform 1 0 15272 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__A
timestamp 1606120350
transform 1 0 15456 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1606120350
transform 1 0 15180 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_36_158
timestamp 1606120350
transform 1 0 15640 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0633_
timestamp 1606120350
transform 1 0 17388 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _0692_
timestamp 1606120350
transform 1 0 16008 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__B1
timestamp 1606120350
transform 1 0 17204 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__A2
timestamp 1606120350
transform 1 0 16836 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0693__A1
timestamp 1606120350
transform 1 0 15824 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_169
timestamp 1606120350
transform 1 0 16652 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_173
timestamp 1606120350
transform 1 0 17020 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0607_
timestamp 1606120350
transform 1 0 18768 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0574__B
timestamp 1606120350
transform 1 0 19688 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__B2
timestamp 1606120350
transform 1 0 18584 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__A
timestamp 1606120350
transform 1 0 18216 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_184
timestamp 1606120350
transform 1 0 18032 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_188
timestamp 1606120350
transform 1 0 18400 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_36_199
timestamp 1606120350
transform 1 0 19412 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_204
timestamp 1606120350
transform 1 0 19872 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_212
timestamp 1606120350
transform 1 0 20608 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_208
timestamp 1606120350
transform 1 0 20240 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0615__A2_N
timestamp 1606120350
transform 1 0 20424 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0574__C
timestamp 1606120350
transform 1 0 20056 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1606120350
transform 1 0 20792 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0608_
timestamp 1606120350
transform 1 0 20884 0 -1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_36_226
timestamp 1606120350
transform 1 0 21896 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_222
timestamp 1606120350
transform 1 0 21528 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__D
timestamp 1606120350
transform 1 0 22080 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0572__A
timestamp 1606120350
transform 1 0 21712 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1135_
timestamp 1606120350
transform 1 0 23092 0 -1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0570__B
timestamp 1606120350
transform 1 0 22448 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_36_230
timestamp 1606120350
transform 1 0 22264 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_234
timestamp 1606120350
transform 1 0 22632 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_238
timestamp 1606120350
transform 1 0 23000 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_258
timestamp 1606120350
transform 1 0 24840 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_270
timestamp 1606120350
transform 1 0 25944 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_274
timestamp 1606120350
transform 1 0 26312 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1606120350
transform 1 0 26404 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_276
timestamp 1606120350
transform 1 0 26496 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_288
timestamp 1606120350
transform 1 0 27600 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_300
timestamp 1606120350
transform 1 0 28704 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_312
timestamp 1606120350
transform 1 0 29808 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1606120350
transform 1 0 32016 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_324
timestamp 1606120350
transform 1 0 30912 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_337
timestamp 1606120350
transform 1 0 32108 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_349
timestamp 1606120350
transform 1 0 33212 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_361
timestamp 1606120350
transform 1 0 34316 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_373
timestamp 1606120350
transform 1 0 35420 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_385
timestamp 1606120350
transform 1 0 36524 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1606120350
transform -1 0 38824 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1606120350
transform 1 0 37628 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_398
timestamp 1606120350
transform 1 0 37720 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_406
timestamp 1606120350
transform 1 0 38456 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1140_
timestamp 1606120350
transform 1 0 1564 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1606120350
transform 1 0 1104 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1606120350
transform 1 0 1380 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_24
timestamp 1606120350
transform 1 0 3312 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_36
timestamp 1606120350
transform 1 0 4416 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1606120350
transform 1 0 6716 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_48
timestamp 1606120350
transform 1 0 5520 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_60
timestamp 1606120350
transform 1 0 6624 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_62
timestamp 1606120350
transform 1 0 6808 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_74
timestamp 1606120350
transform 1 0 7912 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_86
timestamp 1606120350
transform 1 0 9016 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__B1
timestamp 1606120350
transform 1 0 10488 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__B2
timestamp 1606120350
transform 1 0 10856 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__A1
timestamp 1606120350
transform 1 0 11224 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0814__A2
timestamp 1606120350
transform 1 0 10120 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_100
timestamp 1606120350
transform 1 0 10304 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_104
timestamp 1606120350
transform 1 0 10672 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_108
timestamp 1606120350
transform 1 0 11040 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_112
timestamp 1606120350
transform 1 0 11408 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_118
timestamp 1606120350
transform 1 0 11960 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0670__A
timestamp 1606120350
transform 1 0 11776 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__B1
timestamp 1606120350
transform 1 0 12144 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1606120350
transform 1 0 12328 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0670_
timestamp 1606120350
transform 1 0 12420 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_37_133
timestamp 1606120350
transform 1 0 13340 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_37_130
timestamp 1606120350
transform 1 0 13064 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_126
timestamp 1606120350
transform 1 0 12696 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0807__B2
timestamp 1606120350
transform 1 0 13156 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1103_
timestamp 1606120350
transform 1 0 13616 0 1 22304
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0687__B
timestamp 1606120350
transform 1 0 15548 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_155
timestamp 1606120350
transform 1 0 15364 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_37_159
timestamp 1606120350
transform 1 0 15732 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _0638_
timestamp 1606120350
transform 1 0 16560 0 1 22304
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0638__B
timestamp 1606120350
transform 1 0 17388 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__B
timestamp 1606120350
transform 1 0 17756 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__A1
timestamp 1606120350
transform 1 0 16376 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0638__A
timestamp 1606120350
transform 1 0 16008 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_164
timestamp 1606120350
transform 1 0 16192 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_175
timestamp 1606120350
transform 1 0 17204 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_179
timestamp 1606120350
transform 1 0 17572 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__nor3_4  _0574_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 19688 0 1 22304
box -38 -48 1234 592
use sky130_fd_sc_hd__and4_4  _0602_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 18124 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1606120350
transform 1 0 17940 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0574__A
timestamp 1606120350
transform 1 0 19504 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0625__A2
timestamp 1606120350
transform 1 0 19136 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_184
timestamp 1606120350
transform 1 0 18032 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_194
timestamp 1606120350
transform 1 0 18952 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_198
timestamp 1606120350
transform 1 0 19320 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0572_
timestamp 1606120350
transform 1 0 21620 0 1 22304
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__A
timestamp 1606120350
transform 1 0 21068 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__C
timestamp 1606120350
transform 1 0 21436 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_215
timestamp 1606120350
transform 1 0 20884 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_219
timestamp 1606120350
transform 1 0 21252 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1606120350
transform 1 0 23552 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0553__A
timestamp 1606120350
transform 1 0 22632 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0598__A
timestamp 1606120350
transform 1 0 23828 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__B1
timestamp 1606120350
transform 1 0 23000 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_232
timestamp 1606120350
transform 1 0 22448 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_37_236
timestamp 1606120350
transform 1 0 22816 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_240
timestamp 1606120350
transform 1 0 23184 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_37_245
timestamp 1606120350
transform 1 0 23644 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_249
timestamp 1606120350
transform 1 0 24012 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_1_0_clk_A
timestamp 1606120350
transform 1 0 24472 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_37_253
timestamp 1606120350
transform 1 0 24380 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_256
timestamp 1606120350
transform 1 0 24656 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_268
timestamp 1606120350
transform 1 0 25760 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_280
timestamp 1606120350
transform 1 0 26864 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_292
timestamp 1606120350
transform 1 0 27968 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1606120350
transform 1 0 29164 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_37_304
timestamp 1606120350
transform 1 0 29072 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_306
timestamp 1606120350
transform 1 0 29256 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_318
timestamp 1606120350
transform 1 0 30360 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_330
timestamp 1606120350
transform 1 0 31464 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_342
timestamp 1606120350
transform 1 0 32568 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_354
timestamp 1606120350
transform 1 0 33672 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1606120350
transform 1 0 34776 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_367
timestamp 1606120350
transform 1 0 34868 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_379
timestamp 1606120350
transform 1 0 35972 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1606120350
transform -1 0 38824 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_391
timestamp 1606120350
transform 1 0 37076 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_403
timestamp 1606120350
transform 1 0 38180 0 1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1606120350
transform 1 0 1104 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1140__CLK
timestamp 1606120350
transform 1 0 1564 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__CLK
timestamp 1606120350
transform 1 0 2024 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_3
timestamp 1606120350
transform 1 0 1380 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_7
timestamp 1606120350
transform 1 0 1748 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_12
timestamp 1606120350
transform 1 0 2208 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1606120350
transform 1 0 3956 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_24
timestamp 1606120350
transform 1 0 3312 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_30
timestamp 1606120350
transform 1 0 3864 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1606120350
transform 1 0 4048 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1606120350
transform 1 0 5152 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_56
timestamp 1606120350
transform 1 0 6256 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_68
timestamp 1606120350
transform 1 0 7360 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_80
timestamp 1606120350
transform 1 0 8464 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _0814_
timestamp 1606120350
transform 1 0 10488 0 -1 23392
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1606120350
transform 1 0 9568 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_93
timestamp 1606120350
transform 1 0 9660 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_101
timestamp 1606120350
transform 1 0 10396 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0807_
timestamp 1606120350
transform 1 0 13156 0 -1 23392
box -38 -48 1326 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0495__A
timestamp 1606120350
transform 1 0 12788 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__D
timestamp 1606120350
transform 1 0 12420 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0543__A
timestamp 1606120350
transform 1 0 11960 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_116
timestamp 1606120350
transform 1 0 11776 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_38_120
timestamp 1606120350
transform 1 0 12144 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_125
timestamp 1606120350
transform 1 0 12604 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_129
timestamp 1606120350
transform 1 0 12972 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0687_
timestamp 1606120350
transform 1 0 15364 0 -1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1606120350
transform 1 0 15180 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__B1
timestamp 1606120350
transform 1 0 14996 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__B2
timestamp 1606120350
transform 1 0 14628 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_145
timestamp 1606120350
transform 1 0 14444 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_149
timestamp 1606120350
transform 1 0 14812 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_38_154
timestamp 1606120350
transform 1 0 15272 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _0693_
timestamp 1606120350
transform 1 0 16744 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0634__B
timestamp 1606120350
transform 1 0 16468 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_162
timestamp 1606120350
transform 1 0 16008 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_166
timestamp 1606120350
transform 1 0 16376 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_169
timestamp 1606120350
transform 1 0 16652 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_182
timestamp 1606120350
transform 1 0 17848 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_4  _0625_
timestamp 1606120350
transform 1 0 18768 0 -1 23392
box -38 -48 1326 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0612__A
timestamp 1606120350
transform 1 0 18216 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0602__C
timestamp 1606120350
transform 1 0 18584 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_188
timestamp 1606120350
transform 1 0 18400 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0599_
timestamp 1606120350
transform 1 0 20884 0 -1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1606120350
transform 1 0 20792 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__B2
timestamp 1606120350
transform 1 0 20516 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0599__B
timestamp 1606120350
transform 1 0 21896 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_206
timestamp 1606120350
transform 1 0 20056 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_210
timestamp 1606120350
transform 1 0 20424 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_38_213
timestamp 1606120350
transform 1 0 20700 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_224
timestamp 1606120350
transform 1 0 21712 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_228
timestamp 1606120350
transform 1 0 22080 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__C
timestamp 1606120350
transform 1 0 22264 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0553_
timestamp 1606120350
transform 1 0 22448 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_38_235
timestamp 1606120350
transform 1 0 22724 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__D
timestamp 1606120350
transform 1 0 22908 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_239
timestamp 1606120350
transform 1 0 23092 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__A1
timestamp 1606120350
transform 1 0 23276 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_38_246
timestamp 1606120350
transform 1 0 23736 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0598_
timestamp 1606120350
transform 1 0 23460 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_250
timestamp 1606120350
transform 1 0 24104 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0525__A
timestamp 1606120350
transform 1 0 23920 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_1_0_clk
timestamp 1606120350
transform 1 0 24472 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0593__A
timestamp 1606120350
transform 1 0 25208 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__CLK
timestamp 1606120350
transform 1 0 25576 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_257
timestamp 1606120350
transform 1 0 24748 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_261
timestamp 1606120350
transform 1 0 25116 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_38_264
timestamp 1606120350
transform 1 0 25392 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_38_268
timestamp 1606120350
transform 1 0 25760 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_274
timestamp 1606120350
transform 1 0 26312 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1606120350
transform 1 0 26404 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_276
timestamp 1606120350
transform 1 0 26496 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_288
timestamp 1606120350
transform 1 0 27600 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_300
timestamp 1606120350
transform 1 0 28704 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_312
timestamp 1606120350
transform 1 0 29808 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1606120350
transform 1 0 32016 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_324
timestamp 1606120350
transform 1 0 30912 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_337
timestamp 1606120350
transform 1 0 32108 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_349
timestamp 1606120350
transform 1 0 33212 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_361
timestamp 1606120350
transform 1 0 34316 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_373
timestamp 1606120350
transform 1 0 35420 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_385
timestamp 1606120350
transform 1 0 36524 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1606120350
transform -1 0 38824 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1606120350
transform 1 0 37628 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_398
timestamp 1606120350
transform 1 0 37720 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_406
timestamp 1606120350
transform 1 0 38456 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1136_
timestamp 1606120350
transform 1 0 2024 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1606120350
transform 1 0 1104 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1606120350
transform 1 0 1104 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1136__D
timestamp 1606120350
transform 1 0 1840 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1606120350
transform 1 0 1380 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_7
timestamp 1606120350
transform 1 0 1748 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1606120350
transform 1 0 1380 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1606120350
transform 1 0 2484 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1606120350
transform 1 0 3956 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_29
timestamp 1606120350
transform 1 0 3772 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_41
timestamp 1606120350
transform 1 0 4876 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1606120350
transform 1 0 3588 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1606120350
transform 1 0 4048 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1606120350
transform 1 0 5152 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1606120350
transform 1 0 6716 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_53
timestamp 1606120350
transform 1 0 5980 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_62
timestamp 1606120350
transform 1 0 6808 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_56
timestamp 1606120350
transform 1 0 6256 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_68
timestamp 1606120350
transform 1 0 7360 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_0_0_clk
timestamp 1606120350
transform 1 0 7912 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__B1
timestamp 1606120350
transform 1 0 9384 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_0_0_clk_A
timestamp 1606120350
transform 1 0 7912 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__CLK
timestamp 1606120350
transform 1 0 9200 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_76
timestamp 1606120350
transform 1 0 8096 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_90
timestamp 1606120350
transform 1 0 9384 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_77
timestamp 1606120350
transform 1 0 8188 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_89
timestamp 1606120350
transform 1 0 9292 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_101
timestamp 1606120350
transform 1 0 10396 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_97
timestamp 1606120350
transform 1 0 10028 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_93
timestamp 1606120350
transform 1 0 9660 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1108__D
timestamp 1606120350
transform 1 0 9568 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__B2
timestamp 1606120350
transform 1 0 10212 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A1
timestamp 1606120350
transform 1 0 9844 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1606120350
transform 1 0 9568 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_40_112
timestamp 1606120350
transform 1 0 11408 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_108
timestamp 1606120350
transform 1 0 11040 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_113
timestamp 1606120350
transform 1 0 11500 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__CLK
timestamp 1606120350
transform 1 0 10580 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1107__CLK
timestamp 1606120350
transform 1 0 11224 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__A2
timestamp 1606120350
transform 1 0 11592 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0808_
timestamp 1606120350
transform 1 0 10764 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1108_
timestamp 1606120350
transform 1 0 9752 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_40_123
timestamp 1606120350
transform 1 0 12420 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_119
timestamp 1606120350
transform 1 0 12052 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_39_117
timestamp 1606120350
transform 1 0 11868 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0609__A
timestamp 1606120350
transform 1 0 12144 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__A1
timestamp 1606120350
transform 1 0 12512 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0808__A
timestamp 1606120350
transform 1 0 11684 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1606120350
transform 1 0 12328 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0543_
timestamp 1606120350
transform 1 0 11776 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_134
timestamp 1606120350
transform 1 0 13432 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_130
timestamp 1606120350
transform 1 0 13064 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_40_126
timestamp 1606120350
transform 1 0 12696 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__A1
timestamp 1606120350
transform 1 0 13248 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__B1
timestamp 1606120350
transform 1 0 13616 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0495_
timestamp 1606120350
transform 1 0 12788 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1107_
timestamp 1606120350
transform 1 0 12420 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_40_145
timestamp 1606120350
transform 1 0 14444 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_146
timestamp 1606120350
transform 1 0 14536 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_142
timestamp 1606120350
transform 1 0 14168 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0609__B
timestamp 1606120350
transform 1 0 14352 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0609_
timestamp 1606120350
transform 1 0 13800 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_40_154
timestamp 1606120350
transform 1 0 15272 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_40_149
timestamp 1606120350
transform 1 0 14812 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__A4
timestamp 1606120350
transform 1 0 14628 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0635__B
timestamp 1606120350
transform 1 0 14996 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0494__A
timestamp 1606120350
transform 1 0 14720 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1606120350
transform 1 0 15180 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0494_
timestamp 1606120350
transform 1 0 14904 0 1 23392
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_39_159
timestamp 1606120350
transform 1 0 15732 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__A2
timestamp 1606120350
transform 1 0 15640 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_163
timestamp 1606120350
transform 1 0 16100 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__A1_N
timestamp 1606120350
transform 1 0 16284 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0765__A2_N
timestamp 1606120350
transform 1 0 15916 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0634_
timestamp 1606120350
transform 1 0 16468 0 1 23392
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_40_180
timestamp 1606120350
transform 1 0 17664 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_176
timestamp 1606120350
transform 1 0 17296 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_179
timestamp 1606120350
transform 1 0 17572 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_174
timestamp 1606120350
transform 1 0 17112 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0612__D
timestamp 1606120350
transform 1 0 17480 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0612__C
timestamp 1606120350
transform 1 0 17848 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0612__B
timestamp 1606120350
transform 1 0 17388 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0626__A
timestamp 1606120350
transform 1 0 17756 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0765_
timestamp 1606120350
transform 1 0 15824 0 -1 24480
box -38 -48 1510 592
use sky130_fd_sc_hd__fill_2  FILLER_39_184
timestamp 1606120350
transform 1 0 18032 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1606120350
transform 1 0 17940 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_40_205
timestamp 1606120350
transform 1 0 19964 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_40_201
timestamp 1606120350
transform 1 0 19596 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_197
timestamp 1606120350
transform 1 0 19228 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_203
timestamp 1606120350
transform 1 0 19780 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0626__B
timestamp 1606120350
transform 1 0 19780 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0611__C
timestamp 1606120350
transform 1 0 19412 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__C
timestamp 1606120350
transform 1 0 19964 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__nor3_4  _0626_
timestamp 1606120350
transform 1 0 18032 0 -1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__nor4_4  _0612_
timestamp 1606120350
transform 1 0 18216 0 1 23392
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_40_210
timestamp 1606120350
transform 1 0 20424 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_39_207
timestamp 1606120350
transform 1 0 20148 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__A
timestamp 1606120350
transform 1 0 20240 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0613__B
timestamp 1606120350
transform 1 0 20608 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0573__A2
timestamp 1606120350
transform 1 0 20332 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1606120350
transform 1 0 20792 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _0613_
timestamp 1606120350
transform 1 0 20884 0 -1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_40_228
timestamp 1606120350
transform 1 0 22080 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_224
timestamp 1606120350
transform 1 0 21712 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_228
timestamp 1606120350
transform 1 0 22080 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__D
timestamp 1606120350
transform 1 0 21896 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__a22oi_4  _0573_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 20516 0 1 23392
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_39_234
timestamp 1606120350
transform 1 0 22632 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__D
timestamp 1606120350
transform 1 0 22816 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__A
timestamp 1606120350
transform 1 0 22264 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0570__A
timestamp 1606120350
transform 1 0 22448 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0570_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 22448 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_40_243
timestamp 1606120350
transform 1 0 23460 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_239
timestamp 1606120350
transform 1 0 23092 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_238
timestamp 1606120350
transform 1 0 23000 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__D
timestamp 1606120350
transform 1 0 23276 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0528__A
timestamp 1606120350
transform 1 0 23368 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1606120350
transform 1 0 23552 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_248
timestamp 1606120350
transform 1 0 23920 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__D
timestamp 1606120350
transform 1 0 23644 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0525__B
timestamp 1606120350
transform 1 0 24104 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0528_
timestamp 1606120350
transform 1 0 23644 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _0525_
timestamp 1606120350
transform 1 0 23828 0 -1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_40_258
timestamp 1606120350
transform 1 0 24840 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_40_254
timestamp 1606120350
transform 1 0 24472 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_39_252
timestamp 1606120350
transform 1 0 24288 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0489__A
timestamp 1606120350
transform 1 0 25024 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__A2
timestamp 1606120350
transform 1 0 24656 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1133__D
timestamp 1606120350
transform 1 0 24564 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0593_
timestamp 1606120350
transform 1 0 25208 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_40_269
timestamp 1606120350
transform 1 0 25852 0 -1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_40_265
timestamp 1606120350
transform 1 0 25484 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1101__CLK
timestamp 1606120350
transform 1 0 25668 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1133_
timestamp 1606120350
transform 1 0 24748 0 1 23392
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1606120350
transform 1 0 26404 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_276
timestamp 1606120350
transform 1 0 26496 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_288
timestamp 1606120350
transform 1 0 27600 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_276
timestamp 1606120350
transform 1 0 26496 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_288
timestamp 1606120350
transform 1 0 27600 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1606120350
transform 1 0 29164 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_300
timestamp 1606120350
transform 1 0 28704 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_304
timestamp 1606120350
transform 1 0 29072 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_306
timestamp 1606120350
transform 1 0 29256 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_318
timestamp 1606120350
transform 1 0 30360 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_300
timestamp 1606120350
transform 1 0 28704 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_312
timestamp 1606120350
transform 1 0 29808 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1606120350
transform 1 0 32016 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_330
timestamp 1606120350
transform 1 0 31464 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_342
timestamp 1606120350
transform 1 0 32568 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_324
timestamp 1606120350
transform 1 0 30912 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_337
timestamp 1606120350
transform 1 0 32108 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_354
timestamp 1606120350
transform 1 0 33672 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_349
timestamp 1606120350
transform 1 0 33212 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_361
timestamp 1606120350
transform 1 0 34316 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1606120350
transform 1 0 34776 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_367
timestamp 1606120350
transform 1 0 34868 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_379
timestamp 1606120350
transform 1 0 35972 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_373
timestamp 1606120350
transform 1 0 35420 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_385
timestamp 1606120350
transform 1 0 36524 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1606120350
transform -1 0 38824 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1606120350
transform -1 0 38824 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1606120350
transform 1 0 37628 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_391
timestamp 1606120350
transform 1 0 37076 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_403
timestamp 1606120350
transform 1 0 38180 0 1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_398
timestamp 1606120350
transform 1 0 37720 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_406
timestamp 1606120350
transform 1 0 38456 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1606120350
transform 1 0 1104 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1606120350
transform 1 0 1380 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1606120350
transform 1 0 2484 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1606120350
transform 1 0 3588 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1606120350
transform 1 0 4692 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1606120350
transform 1 0 6716 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_51
timestamp 1606120350
transform 1 0 5796 0 1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_59
timestamp 1606120350
transform 1 0 6532 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_41_62
timestamp 1606120350
transform 1 0 6808 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1124_
timestamp 1606120350
transform 1 0 9108 0 1 24480
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__D
timestamp 1606120350
transform 1 0 8924 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1124__CLK
timestamp 1606120350
transform 1 0 8556 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_74
timestamp 1606120350
transform 1 0 7912 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_80
timestamp 1606120350
transform 1 0 8464 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_83
timestamp 1606120350
transform 1 0 8740 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__B2
timestamp 1606120350
transform 1 0 11408 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0811__A2
timestamp 1606120350
transform 1 0 11040 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_106
timestamp 1606120350
transform 1 0 10856 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_110
timestamp 1606120350
transform 1 0 11224 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_114
timestamp 1606120350
transform 1 0 11592 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0812_
timestamp 1606120350
transform 1 0 12512 0 1 24480
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1606120350
transform 1 0 12328 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__B1
timestamp 1606120350
transform 1 0 12144 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0799__A
timestamp 1606120350
transform 1 0 11776 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_118
timestamp 1606120350
transform 1 0 11960 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_123
timestamp 1606120350
transform 1 0 12420 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_138
timestamp 1606120350
transform 1 0 13800 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0751__B1
timestamp 1606120350
transform 1 0 13984 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_142
timestamp 1606120350
transform 1 0 14168 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__A3
timestamp 1606120350
transform 1 0 14352 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0497_
timestamp 1606120350
transform 1 0 14536 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_149
timestamp 1606120350
transform 1 0 14812 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0497__A
timestamp 1606120350
transform 1 0 14996 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_153
timestamp 1606120350
transform 1 0 15180 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0519__A
timestamp 1606120350
transform 1 0 15364 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_41_157
timestamp 1606120350
transform 1 0 15548 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_4  _0635_
timestamp 1606120350
transform 1 0 15824 0 1 24480
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__A1
timestamp 1606120350
transform 1 0 17756 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0626__C
timestamp 1606120350
transform 1 0 17388 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_173
timestamp 1606120350
transform 1 0 17020 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_179
timestamp 1606120350
transform 1 0 17572 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _0632_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 18032 0 1 24480
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1606120350
transform 1 0 17940 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0611__B
timestamp 1606120350
transform 1 0 19504 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0611__A
timestamp 1606120350
transform 1 0 19872 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_198
timestamp 1606120350
transform 1 0 19320 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_202
timestamp 1606120350
transform 1 0 19688 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0529_
timestamp 1606120350
transform 1 0 21620 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0647_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 20056 0 1 24480
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0529__A
timestamp 1606120350
transform 1 0 21436 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__A
timestamp 1606120350
transform 1 0 21068 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_215
timestamp 1606120350
transform 1 0 20884 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_219
timestamp 1606120350
transform 1 0 21252 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0524_
timestamp 1606120350
transform 1 0 23644 0 1 24480
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1606120350
transform 1 0 23552 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0524__A
timestamp 1606120350
transform 1 0 23368 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__C
timestamp 1606120350
transform 1 0 22632 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__B
timestamp 1606120350
transform 1 0 23000 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_232
timestamp 1606120350
transform 1 0 22448 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_236
timestamp 1606120350
transform 1 0 22816 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_240
timestamp 1606120350
transform 1 0 23184 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_256
timestamp 1606120350
transform 1 0 24656 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_252
timestamp 1606120350
transform 1 0 24288 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0524__B
timestamp 1606120350
transform 1 0 24472 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__A1
timestamp 1606120350
transform 1 0 24840 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0526_
timestamp 1606120350
transform 1 0 25024 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_41_263
timestamp 1606120350
transform 1 0 25300 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0526__A
timestamp 1606120350
transform 1 0 25484 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_41_267
timestamp 1606120350
transform 1 0 25668 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0522__A
timestamp 1606120350
transform 1 0 25852 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_271
timestamp 1606120350
transform 1 0 26036 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0592__A
timestamp 1606120350
transform 1 0 26496 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_41_275
timestamp 1606120350
transform 1 0 26404 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_278
timestamp 1606120350
transform 1 0 26680 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_290
timestamp 1606120350
transform 1 0 27784 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1606120350
transform 1 0 29164 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_41_302
timestamp 1606120350
transform 1 0 28888 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_306
timestamp 1606120350
transform 1 0 29256 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_318
timestamp 1606120350
transform 1 0 30360 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_330
timestamp 1606120350
transform 1 0 31464 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_342
timestamp 1606120350
transform 1 0 32568 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_354
timestamp 1606120350
transform 1 0 33672 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1606120350
transform 1 0 34776 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_367
timestamp 1606120350
transform 1 0 34868 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_379
timestamp 1606120350
transform 1 0 35972 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1606120350
transform -1 0 38824 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_391
timestamp 1606120350
transform 1 0 37076 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_403
timestamp 1606120350
transform 1 0 38180 0 1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1606120350
transform 1 0 1104 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1606120350
transform 1 0 1380 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1606120350
transform 1 0 2484 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1606120350
transform 1 0 3956 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1606120350
transform 1 0 3588 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1606120350
transform 1 0 4048 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1606120350
transform 1 0 5152 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_56
timestamp 1606120350
transform 1 0 6256 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_68
timestamp 1606120350
transform 1 0 7360 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__D
timestamp 1606120350
transform 1 0 9016 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1111__D
timestamp 1606120350
transform 1 0 9384 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_42_80
timestamp 1606120350
transform 1 0 8464 0 -1 25568
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_42_88
timestamp 1606120350
transform 1 0 9200 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0811_
timestamp 1606120350
transform 1 0 9660 0 -1 25568
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1606120350
transform 1 0 9568 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__A2
timestamp 1606120350
transform 1 0 11316 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_107
timestamp 1606120350
transform 1 0 10948 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_42_113
timestamp 1606120350
transform 1 0 11500 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0751_
timestamp 1606120350
transform 1 0 13340 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0799_
timestamp 1606120350
transform 1 0 12236 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__B1
timestamp 1606120350
transform 1 0 13156 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__B1
timestamp 1606120350
transform 1 0 12788 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__A2
timestamp 1606120350
transform 1 0 12052 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0812__A2
timestamp 1606120350
transform 1 0 11684 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_117
timestamp 1606120350
transform 1 0 11868 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_42_124
timestamp 1606120350
transform 1 0 12512 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_42_129
timestamp 1606120350
transform 1 0 12972 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0519_
timestamp 1606120350
transform 1 0 15364 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1606120350
transform 1 0 15180 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__C
timestamp 1606120350
transform 1 0 14628 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0635__C
timestamp 1606120350
transform 1 0 14996 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_145
timestamp 1606120350
transform 1 0 14444 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_149
timestamp 1606120350
transform 1 0 14812 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_154
timestamp 1606120350
transform 1 0 15272 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_158
timestamp 1606120350
transform 1 0 15640 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__o41a_4  _0649_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 16376 0 -1 25568
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0635__A
timestamp 1606120350
transform 1 0 15824 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0649__A1
timestamp 1606120350
transform 1 0 16192 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_162
timestamp 1606120350
transform 1 0 16008 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__nor3_4  _0611_
timestamp 1606120350
transform 1 0 18676 0 -1 25568
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__B1
timestamp 1606120350
transform 1 0 18124 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__A2
timestamp 1606120350
transform 1 0 18492 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_183
timestamp 1606120350
transform 1 0 17940 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_187
timestamp 1606120350
transform 1 0 18308 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_204
timestamp 1606120350
transform 1 0 19872 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_215
timestamp 1606120350
transform 1 0 20884 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_212
timestamp 1606120350
transform 1 0 20608 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_208
timestamp 1606120350
transform 1 0 20240 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__C1
timestamp 1606120350
transform 1 0 20424 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0632__B1
timestamp 1606120350
transform 1 0 20056 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1606120350
transform 1 0 20792 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_42_223
timestamp 1606120350
transform 1 0 21620 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_219
timestamp 1606120350
transform 1 0 21252 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0647__B
timestamp 1606120350
transform 1 0 21436 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__A
timestamp 1606120350
transform 1 0 21068 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0489_
timestamp 1606120350
transform 1 0 21712 0 -1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_4  _1101_
timestamp 1606120350
transform 1 0 23368 0 -1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__B
timestamp 1606120350
transform 1 0 22724 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__C
timestamp 1606120350
transform 1 0 23092 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_233
timestamp 1606120350
transform 1 0 22540 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_237
timestamp 1606120350
transform 1 0 22908 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_42_241
timestamp 1606120350
transform 1 0 23276 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0703__B
timestamp 1606120350
transform 1 0 25300 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__B2
timestamp 1606120350
transform 1 0 25668 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0804__B1
timestamp 1606120350
transform 1 0 26036 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_261
timestamp 1606120350
transform 1 0 25116 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_265
timestamp 1606120350
transform 1 0 25484 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_269
timestamp 1606120350
transform 1 0 25852 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_273
timestamp 1606120350
transform 1 0 26220 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0592_
timestamp 1606120350
transform 1 0 26496 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1606120350
transform 1 0 26404 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0556__C
timestamp 1606120350
transform 1 0 26956 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_42_279
timestamp 1606120350
transform 1 0 26772 0 -1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_283
timestamp 1606120350
transform 1 0 27140 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_295
timestamp 1606120350
transform 1 0 28244 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_307
timestamp 1606120350
transform 1 0 29348 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_319
timestamp 1606120350
transform 1 0 30452 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1606120350
transform 1 0 32016 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_331
timestamp 1606120350
transform 1 0 31556 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_335
timestamp 1606120350
transform 1 0 31924 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_337
timestamp 1606120350
transform 1 0 32108 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_349
timestamp 1606120350
transform 1 0 33212 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_361
timestamp 1606120350
transform 1 0 34316 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_373
timestamp 1606120350
transform 1 0 35420 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_385
timestamp 1606120350
transform 1 0 36524 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1606120350
transform -1 0 38824 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1606120350
transform 1 0 37628 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_398
timestamp 1606120350
transform 1 0 37720 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_406
timestamp 1606120350
transform 1 0 38456 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1606120350
transform 1 0 1104 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1606120350
transform 1 0 1380 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1606120350
transform 1 0 2484 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1606120350
transform 1 0 3588 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1606120350
transform 1 0 4692 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1606120350
transform 1 0 6716 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__D
timestamp 1606120350
transform 1 0 6072 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1120__CLK
timestamp 1606120350
transform 1 0 6440 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_51
timestamp 1606120350
transform 1 0 5796 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_56
timestamp 1606120350
transform 1 0 6256 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_43_60
timestamp 1606120350
transform 1 0 6624 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_62
timestamp 1606120350
transform 1 0 6808 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1106_
timestamp 1606120350
transform 1 0 9016 0 1 25568
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0813__A
timestamp 1606120350
transform 1 0 8556 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1106__CLK
timestamp 1606120350
transform 1 0 8188 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_74
timestamp 1606120350
transform 1 0 7912 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_79
timestamp 1606120350
transform 1 0 8372 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_83
timestamp 1606120350
transform 1 0 8740 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__D
timestamp 1606120350
transform 1 0 11408 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__D
timestamp 1606120350
transform 1 0 11040 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_105
timestamp 1606120350
transform 1 0 10764 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_110
timestamp 1606120350
transform 1 0 11224 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_114
timestamp 1606120350
transform 1 0 11592 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0688_
timestamp 1606120350
transform 1 0 12420 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_565
timestamp 1606120350
transform 1 0 12328 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__A1
timestamp 1606120350
transform 1 0 13340 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__A
timestamp 1606120350
transform 1 0 12144 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0752__A2
timestamp 1606120350
transform 1 0 11776 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_118
timestamp 1606120350
transform 1 0 11960 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_130
timestamp 1606120350
transform 1 0 13064 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_43_135
timestamp 1606120350
transform 1 0 13524 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _0631_
timestamp 1606120350
transform 1 0 13800 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _0766_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 15364 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__A
timestamp 1606120350
transform 1 0 14812 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0541__A
timestamp 1606120350
transform 1 0 15180 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_147
timestamp 1606120350
transform 1 0 14628 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_151
timestamp 1606120350
transform 1 0 14996 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__A
timestamp 1606120350
transform 1 0 16652 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__A2
timestamp 1606120350
transform 1 0 17756 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__C1
timestamp 1606120350
transform 1 0 17388 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__B
timestamp 1606120350
transform 1 0 17020 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_167
timestamp 1606120350
transform 1 0 16468 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_171
timestamp 1606120350
transform 1 0 16836 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_175
timestamp 1606120350
transform 1 0 17204 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_179
timestamp 1606120350
transform 1 0 17572 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__a2111oi_4  _0610_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 18032 0 1 25568
box -38 -48 2062 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_566
timestamp 1606120350
transform 1 0 17940 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0703_
timestamp 1606120350
transform 1 0 20792 0 1 25568
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__A
timestamp 1606120350
transform 1 0 20240 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0571__A
timestamp 1606120350
transform 1 0 21804 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__B
timestamp 1606120350
transform 1 0 20608 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_206
timestamp 1606120350
transform 1 0 20056 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_210
timestamp 1606120350
transform 1 0 20424 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_223
timestamp 1606120350
transform 1 0 21620 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_227
timestamp 1606120350
transform 1 0 21988 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_238
timestamp 1606120350
transform 1 0 23000 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_234
timestamp 1606120350
transform 1 0 22632 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0556__D
timestamp 1606120350
transform 1 0 22172 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0556__B
timestamp 1606120350
transform 1 0 22816 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0571_
timestamp 1606120350
transform 1 0 22356 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_43_245
timestamp 1606120350
transform 1 0 23644 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_242
timestamp 1606120350
transform 1 0 23368 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0556__A
timestamp 1606120350
transform 1 0 23184 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_567
timestamp 1606120350
transform 1 0 23552 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _0804_
timestamp 1606120350
transform 1 0 23828 0 1 25568
box -38 -48 1326 592
use sky130_fd_sc_hd__or2_4  _0527_
timestamp 1606120350
transform 1 0 25852 0 1 25568
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0527__A
timestamp 1606120350
transform 1 0 25668 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__C
timestamp 1606120350
transform 1 0 25300 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_261
timestamp 1606120350
transform 1 0 25116 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_265
timestamp 1606120350
transform 1 0 25484 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0527__B
timestamp 1606120350
transform 1 0 26680 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0523__A
timestamp 1606120350
transform 1 0 27048 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0601__A
timestamp 1606120350
transform 1 0 27508 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_276
timestamp 1606120350
transform 1 0 26496 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_43_280
timestamp 1606120350
transform 1 0 26864 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_43_284
timestamp 1606120350
transform 1 0 27232 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_289
timestamp 1606120350
transform 1 0 27692 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_568
timestamp 1606120350
transform 1 0 29164 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_301
timestamp 1606120350
transform 1 0 28796 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_306
timestamp 1606120350
transform 1 0 29256 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_318
timestamp 1606120350
transform 1 0 30360 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_330
timestamp 1606120350
transform 1 0 31464 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_342
timestamp 1606120350
transform 1 0 32568 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_354
timestamp 1606120350
transform 1 0 33672 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_569
timestamp 1606120350
transform 1 0 34776 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_367
timestamp 1606120350
transform 1 0 34868 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_379
timestamp 1606120350
transform 1 0 35972 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1606120350
transform -1 0 38824 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_391
timestamp 1606120350
transform 1 0 37076 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_403
timestamp 1606120350
transform 1 0 38180 0 1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1606120350
transform 1 0 1104 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__D
timestamp 1606120350
transform 1 0 1564 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1216__CLK
timestamp 1606120350
transform 1 0 1932 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1606120350
transform 1 0 1380 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_7
timestamp 1606120350
transform 1 0 1748 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_11
timestamp 1606120350
transform 1 0 2116 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_570
timestamp 1606120350
transform 1 0 3956 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_23
timestamp 1606120350
transform 1 0 3220 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_32
timestamp 1606120350
transform 1 0 4048 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_44
timestamp 1606120350
transform 1 0 5152 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1120_
timestamp 1606120350
transform 1 0 6072 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_44_52
timestamp 1606120350
transform 1 0 5888 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0813_
timestamp 1606120350
transform 1 0 8556 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__B1
timestamp 1606120350
transform 1 0 9384 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0532__A
timestamp 1606120350
transform 1 0 9016 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_73
timestamp 1606120350
transform 1 0 7820 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_84
timestamp 1606120350
transform 1 0 8832 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_88
timestamp 1606120350
transform 1 0 9200 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1111_
timestamp 1606120350
transform 1 0 10488 0 -1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_571
timestamp 1606120350
transform 1 0 9568 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A1
timestamp 1606120350
transform 1 0 10304 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__B2
timestamp 1606120350
transform 1 0 9936 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_93
timestamp 1606120350
transform 1 0 9660 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_98
timestamp 1606120350
transform 1 0 10120 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _0752_
timestamp 1606120350
transform 1 0 13340 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0688__B
timestamp 1606120350
transform 1 0 12420 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__B1
timestamp 1606120350
transform 1 0 12972 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_121
timestamp 1606120350
transform 1 0 12236 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_125
timestamp 1606120350
transform 1 0 12604 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_131
timestamp 1606120350
transform 1 0 13156 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0541_
timestamp 1606120350
transform 1 0 15548 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_572
timestamp 1606120350
transform 1 0 15180 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0631__B
timestamp 1606120350
transform 1 0 14628 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__D
timestamp 1606120350
transform 1 0 14996 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_145
timestamp 1606120350
transform 1 0 14444 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_149
timestamp 1606120350
transform 1 0 14812 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_44_154
timestamp 1606120350
transform 1 0 15272 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_4  _0636_
timestamp 1606120350
transform 1 0 16560 0 -1 26656
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0766__A1
timestamp 1606120350
transform 1 0 16008 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__C
timestamp 1606120350
transform 1 0 16376 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_160
timestamp 1606120350
transform 1 0 15824 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_164
timestamp 1606120350
transform 1 0 16192 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_181
timestamp 1606120350
transform 1 0 17756 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0696_
timestamp 1606120350
transform 1 0 18860 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__A
timestamp 1606120350
transform 1 0 19872 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__C
timestamp 1606120350
transform 1 0 17940 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0696__C
timestamp 1606120350
transform 1 0 18676 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0610__D1
timestamp 1606120350
transform 1 0 18308 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_185
timestamp 1606120350
transform 1 0 18124 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_189
timestamp 1606120350
transform 1 0 18492 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_202
timestamp 1606120350
transform 1 0 19688 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0704_
timestamp 1606120350
transform 1 0 20884 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_573
timestamp 1606120350
transform 1 0 20792 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__D
timestamp 1606120350
transform 1 0 20240 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__B
timestamp 1606120350
transform 1 0 21896 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__A
timestamp 1606120350
transform 1 0 20608 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_206
timestamp 1606120350
transform 1 0 20056 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_210
timestamp 1606120350
transform 1 0 20424 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_224
timestamp 1606120350
transform 1 0 21712 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_228
timestamp 1606120350
transform 1 0 22080 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0522_
timestamp 1606120350
transform 1 0 24012 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0556_
timestamp 1606120350
transform 1 0 22448 0 -1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0561__B
timestamp 1606120350
transform 1 0 23644 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__B
timestamp 1606120350
transform 1 0 22264 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_241
timestamp 1606120350
transform 1 0 23276 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_44_247
timestamp 1606120350
transform 1 0 23828 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__B
timestamp 1606120350
transform 1 0 25024 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0704__D
timestamp 1606120350
transform 1 0 25392 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__D
timestamp 1606120350
transform 1 0 25760 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__D
timestamp 1606120350
transform 1 0 26128 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_258
timestamp 1606120350
transform 1 0 24840 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_262
timestamp 1606120350
transform 1 0 25208 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_266
timestamp 1606120350
transform 1 0 25576 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_270
timestamp 1606120350
transform 1 0 25944 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_44_274
timestamp 1606120350
transform 1 0 26312 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_44_283
timestamp 1606120350
transform 1 0 27140 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_44_279
timestamp 1606120350
transform 1 0 26772 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__D
timestamp 1606120350
transform 1 0 27324 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__D
timestamp 1606120350
transform 1 0 26956 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_574
timestamp 1606120350
transform 1 0 26404 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0523_
timestamp 1606120350
transform 1 0 26496 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_290
timestamp 1606120350
transform 1 0 27784 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0561__C
timestamp 1606120350
transform 1 0 27968 0 -1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0601_
timestamp 1606120350
transform 1 0 27508 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_294
timestamp 1606120350
transform 1 0 28152 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_306
timestamp 1606120350
transform 1 0 29256 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_318
timestamp 1606120350
transform 1 0 30360 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_575
timestamp 1606120350
transform 1 0 32016 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_330
timestamp 1606120350
transform 1 0 31464 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_337
timestamp 1606120350
transform 1 0 32108 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_349
timestamp 1606120350
transform 1 0 33212 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_361
timestamp 1606120350
transform 1 0 34316 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_373
timestamp 1606120350
transform 1 0 35420 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_385
timestamp 1606120350
transform 1 0 36524 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1606120350
transform -1 0 38824 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_576
timestamp 1606120350
transform 1 0 37628 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_398
timestamp 1606120350
transform 1 0 37720 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_406
timestamp 1606120350
transform 1 0 38456 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1216_
timestamp 1606120350
transform 1 0 1564 0 1 26656
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1606120350
transform 1 0 1104 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_3
timestamp 1606120350
transform 1 0 1380 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_24
timestamp 1606120350
transform 1 0 3312 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_36
timestamp 1606120350
transform 1 0 4416 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_577
timestamp 1606120350
transform 1 0 6716 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__D
timestamp 1606120350
transform 1 0 6992 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1200__CLK
timestamp 1606120350
transform 1 0 7360 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_48
timestamp 1606120350
transform 1 0 5520 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_60
timestamp 1606120350
transform 1 0 6624 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_62
timestamp 1606120350
transform 1 0 6808 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_66
timestamp 1606120350
transform 1 0 7176 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0630_
timestamp 1606120350
transform 1 0 9292 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0662_
timestamp 1606120350
transform 1 0 8280 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0662__A
timestamp 1606120350
transform 1 0 8740 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0818__A2
timestamp 1606120350
transform 1 0 9108 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_70
timestamp 1606120350
transform 1 0 7544 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_81
timestamp 1606120350
transform 1 0 8556 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_85
timestamp 1606120350
transform 1 0 8924 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0818_
timestamp 1606120350
transform 1 0 10304 0 1 26656
box -38 -48 1326 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0630__A
timestamp 1606120350
transform 1 0 9752 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0806__A
timestamp 1606120350
transform 1 0 10120 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_92
timestamp 1606120350
transform 1 0 9568 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_96
timestamp 1606120350
transform 1 0 9936 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_114
timestamp 1606120350
transform 1 0 11592 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _0759_
timestamp 1606120350
transform 1 0 12880 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_578
timestamp 1606120350
transform 1 0 12328 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A2
timestamp 1606120350
transform 1 0 12696 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__B
timestamp 1606120350
transform 1 0 11776 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0757__A
timestamp 1606120350
transform 1 0 12144 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_118
timestamp 1606120350
transform 1 0 11960 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_123
timestamp 1606120350
transform 1 0 12420 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_4  _0758_
timestamp 1606120350
transform 1 0 14720 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__B
timestamp 1606120350
transform 1 0 14536 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__B1
timestamp 1606120350
transform 1 0 14168 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_140
timestamp 1606120350
transform 1 0 13984 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_144
timestamp 1606120350
transform 1 0 14352 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0532_
timestamp 1606120350
transform 1 0 16560 0 1 26656
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0532__B
timestamp 1606120350
transform 1 0 17388 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0694__A
timestamp 1606120350
transform 1 0 17756 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__A
timestamp 1606120350
transform 1 0 16008 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0690__B
timestamp 1606120350
transform 1 0 16376 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_160
timestamp 1606120350
transform 1 0 15824 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_164
timestamp 1606120350
transform 1 0 16192 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_175
timestamp 1606120350
transform 1 0 17204 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_179
timestamp 1606120350
transform 1 0 17572 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0563_
timestamp 1606120350
transform 1 0 18216 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__nand4_4  _0567_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 19228 0 1 26656
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_579
timestamp 1606120350
transform 1 0 17940 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0563__A
timestamp 1606120350
transform 1 0 18676 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__C
timestamp 1606120350
transform 1 0 19044 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_184
timestamp 1606120350
transform 1 0 18032 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_189
timestamp 1606120350
transform 1 0 18492 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_193
timestamp 1606120350
transform 1 0 18860 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0641_
timestamp 1606120350
transform 1 0 21528 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__A
timestamp 1606120350
transform 1 0 21344 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0641__C
timestamp 1606120350
transform 1 0 20976 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_214
timestamp 1606120350
transform 1 0 20792 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_218
timestamp 1606120350
transform 1 0 21160 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0561_
timestamp 1606120350
transform 1 0 23644 0 1 26656
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_580
timestamp 1606120350
transform 1 0 23552 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0561__A
timestamp 1606120350
transform 1 0 23368 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__A
timestamp 1606120350
transform 1 0 22540 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__C
timestamp 1606120350
transform 1 0 22908 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_231
timestamp 1606120350
transform 1 0 22356 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_235
timestamp 1606120350
transform 1 0 22724 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_45_239
timestamp 1606120350
transform 1 0 23092 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_254
timestamp 1606120350
transform 1 0 24472 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_258
timestamp 1606120350
transform 1 0 24840 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__C
timestamp 1606120350
transform 1 0 24656 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__A
timestamp 1606120350
transform 1 0 25024 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0565_
timestamp 1606120350
transform 1 0 25208 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_265
timestamp 1606120350
transform 1 0 25484 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_269
timestamp 1606120350
transform 1 0 25852 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0565__A
timestamp 1606120350
transform 1 0 25668 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__D
timestamp 1606120350
transform 1 0 26036 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0490_
timestamp 1606120350
transform 1 0 26220 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_276
timestamp 1606120350
transform 1 0 26496 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_280
timestamp 1606120350
transform 1 0 26864 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0490__A
timestamp 1606120350
transform 1 0 26680 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0517__A
timestamp 1606120350
transform 1 0 27048 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0518_
timestamp 1606120350
transform 1 0 27232 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_45_287
timestamp 1606120350
transform 1 0 27508 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0518__A
timestamp 1606120350
transform 1 0 27692 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_291
timestamp 1606120350
transform 1 0 27876 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0640__A
timestamp 1606120350
transform 1 0 28060 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_45_295
timestamp 1606120350
transform 1 0 28244 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_581
timestamp 1606120350
transform 1 0 29164 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0561__D
timestamp 1606120350
transform 1 0 28428 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_299
timestamp 1606120350
transform 1 0 28612 0 1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_306
timestamp 1606120350
transform 1 0 29256 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_318
timestamp 1606120350
transform 1 0 30360 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_330
timestamp 1606120350
transform 1 0 31464 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_342
timestamp 1606120350
transform 1 0 32568 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_354
timestamp 1606120350
transform 1 0 33672 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_582
timestamp 1606120350
transform 1 0 34776 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_367
timestamp 1606120350
transform 1 0 34868 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_379
timestamp 1606120350
transform 1 0 35972 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1606120350
transform -1 0 38824 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_391
timestamp 1606120350
transform 1 0 37076 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_403
timestamp 1606120350
transform 1 0 38180 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_10
timestamp 1606120350
transform 1 0 2024 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_3
timestamp 1606120350
transform 1 0 1380 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0486__A
timestamp 1606120350
transform 1 0 1564 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1606120350
transform 1 0 1104 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1606120350
transform 1 0 1104 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _0486_
timestamp 1606120350
transform 1 0 1380 0 1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0486__B
timestamp 1606120350
transform 1 0 2208 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_14
timestamp 1606120350
transform 1 0 2392 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_19
timestamp 1606120350
transform 1 0 2852 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_7
timestamp 1606120350
transform 1 0 1748 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_583
timestamp 1606120350
transform 1 0 3956 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_32
timestamp 1606120350
transform 1 0 4048 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_44
timestamp 1606120350
transform 1 0 5152 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_26
timestamp 1606120350
transform 1 0 3496 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_38
timestamp 1606120350
transform 1 0 4600 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1200_
timestamp 1606120350
transform 1 0 6716 0 -1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_590
timestamp 1606120350
transform 1 0 6716 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__B1
timestamp 1606120350
transform 1 0 7176 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_56
timestamp 1606120350
transform 1 0 6256 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_60
timestamp 1606120350
transform 1 0 6624 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_50
timestamp 1606120350
transform 1 0 5704 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_58
timestamp 1606120350
transform 1 0 6440 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_62
timestamp 1606120350
transform 1 0 6808 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_47_68
timestamp 1606120350
transform 1 0 7360 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_72
timestamp 1606120350
transform 1 0 7728 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__A1
timestamp 1606120350
transform 1 0 7544 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_76
timestamp 1606120350
transform 1 0 8096 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__B2
timestamp 1606120350
transform 1 0 7912 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_80
timestamp 1606120350
transform 1 0 8464 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_80
timestamp 1606120350
transform 1 0 8464 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0810__A2
timestamp 1606120350
transform 1 0 8280 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__A1
timestamp 1606120350
transform 1 0 8648 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__A1
timestamp 1606120350
transform 1 0 8740 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_85
timestamp 1606120350
transform 1 0 8924 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_84
timestamp 1606120350
transform 1 0 8832 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0760__A1
timestamp 1606120350
transform 1 0 9016 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A1
timestamp 1606120350
transform 1 0 9108 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_88
timestamp 1606120350
transform 1 0 9200 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__A1
timestamp 1606120350
transform 1 0 9384 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0624_
timestamp 1606120350
transform 1 0 9292 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_96
timestamp 1606120350
transform 1 0 9936 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_92
timestamp 1606120350
transform 1 0 9568 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_99
timestamp 1606120350
transform 1 0 10212 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_93
timestamp 1606120350
transform 1 0 9660 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__B2
timestamp 1606120350
transform 1 0 10028 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__B1
timestamp 1606120350
transform 1 0 10120 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0624__A
timestamp 1606120350
transform 1 0 9752 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_584
timestamp 1606120350
transform 1 0 9568 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_107
timestamp 1606120350
transform 1 0 10948 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_103
timestamp 1606120350
transform 1 0 10580 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_106
timestamp 1606120350
transform 1 0 10856 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__B2
timestamp 1606120350
transform 1 0 10396 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0661__A
timestamp 1606120350
transform 1 0 10764 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0806_
timestamp 1606120350
transform 1 0 10580 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0654_
timestamp 1606120350
transform 1 0 10304 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_114
timestamp 1606120350
transform 1 0 11592 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_110
timestamp 1606120350
transform 1 0 11224 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__A2
timestamp 1606120350
transform 1 0 11040 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__A1
timestamp 1606120350
transform 1 0 11408 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0654__A
timestamp 1606120350
transform 1 0 11132 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0757_
timestamp 1606120350
transform 1 0 11592 0 -1 27744
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _0711_
timestamp 1606120350
transform 1 0 11316 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_123
timestamp 1606120350
transform 1 0 12420 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_118
timestamp 1606120350
transform 1 0 11960 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_125
timestamp 1606120350
transform 1 0 12604 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_121
timestamp 1606120350
transform 1 0 12236 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0761__A2
timestamp 1606120350
transform 1 0 12420 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__A2
timestamp 1606120350
transform 1 0 12144 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0711__A
timestamp 1606120350
transform 1 0 11776 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_591
timestamp 1606120350
transform 1 0 12328 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_133
timestamp 1606120350
transform 1 0 13340 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_129
timestamp 1606120350
transform 1 0 12972 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0759__B1
timestamp 1606120350
transform 1 0 12788 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__B1
timestamp 1606120350
transform 1 0 13524 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0535__A
timestamp 1606120350
transform 1 0 13156 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0535_
timestamp 1606120350
transform 1 0 12696 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _0768_
timestamp 1606120350
transform 1 0 13708 0 1 27744
box -38 -48 1326 592
use sky130_fd_sc_hd__o21a_4  _0760_
timestamp 1606120350
transform 1 0 12972 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_146
timestamp 1606120350
transform 1 0 14536 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_141
timestamp 1606120350
transform 1 0 14076 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__A
timestamp 1606120350
transform 1 0 14352 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0758__A1
timestamp 1606120350
transform 1 0 14720 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_156
timestamp 1606120350
transform 1 0 15456 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_47_151
timestamp 1606120350
transform 1 0 14996 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_154
timestamp 1606120350
transform 1 0 15272 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_46_150
timestamp 1606120350
transform 1 0 14904 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__B
timestamp 1606120350
transform 1 0 15640 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0767__A2
timestamp 1606120350
transform 1 0 15272 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_585
timestamp 1606120350
transform 1 0 15180 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _0537_
timestamp 1606120350
transform 1 0 15732 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_169
timestamp 1606120350
transform 1 0 16652 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0690_
timestamp 1606120350
transform 1 0 15824 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_179
timestamp 1606120350
transform 1 0 17572 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_175
timestamp 1606120350
transform 1 0 17204 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_171
timestamp 1606120350
transform 1 0 16836 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_173
timestamp 1606120350
transform 1 0 17020 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__B
timestamp 1606120350
transform 1 0 17204 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0636__C
timestamp 1606120350
transform 1 0 16836 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0537__B1
timestamp 1606120350
transform 1 0 17388 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0537__A1
timestamp 1606120350
transform 1 0 17020 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0694_
timestamp 1606120350
transform 1 0 17388 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0566__A
timestamp 1606120350
transform 1 0 17756 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0538_
timestamp 1606120350
transform 1 0 18308 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_592
timestamp 1606120350
transform 1 0 17940 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__C
timestamp 1606120350
transform 1 0 18400 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_186
timestamp 1606120350
transform 1 0 18216 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_47_184
timestamp 1606120350
transform 1 0 18032 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0538__A
timestamp 1606120350
transform 1 0 18768 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__A
timestamp 1606120350
transform 1 0 18768 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_190
timestamp 1606120350
transform 1 0 18584 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_190
timestamp 1606120350
transform 1 0 18584 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_194
timestamp 1606120350
transform 1 0 18952 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0699_
timestamp 1606120350
transform 1 0 18952 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_46_203
timestamp 1606120350
transform 1 0 19780 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0567__B
timestamp 1606120350
transform 1 0 19964 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__A
timestamp 1606120350
transform 1 0 19136 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__nor4_4  _0618_
timestamp 1606120350
transform 1 0 19320 0 1 27744
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_47_215
timestamp 1606120350
transform 1 0 20884 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_46_211
timestamp 1606120350
transform 1 0 20516 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_207
timestamp 1606120350
transform 1 0 20148 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__A
timestamp 1606120350
transform 1 0 20608 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_586
timestamp 1606120350
transform 1 0 20792 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0646_
timestamp 1606120350
transform 1 0 20884 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_219
timestamp 1606120350
transform 1 0 21252 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_224
timestamp 1606120350
transform 1 0 21712 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__C
timestamp 1606120350
transform 1 0 21068 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__A
timestamp 1606120350
transform 1 0 21436 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0642_
timestamp 1606120350
transform 1 0 21620 0 1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_46_228
timestamp 1606120350
transform 1 0 22080 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__B
timestamp 1606120350
transform 1 0 21896 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_236
timestamp 1606120350
transform 1 0 22816 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_232
timestamp 1606120350
transform 1 0 22448 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__C
timestamp 1606120350
transform 1 0 22264 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__C
timestamp 1606120350
transform 1 0 23000 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__A
timestamp 1606120350
transform 1 0 22632 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0705_
timestamp 1606120350
transform 1 0 22448 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_47_240
timestamp 1606120350
transform 1 0 23184 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_245
timestamp 1606120350
transform 1 0 23644 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_241
timestamp 1606120350
transform 1 0 23276 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0646__D
timestamp 1606120350
transform 1 0 23460 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0702__B
timestamp 1606120350
transform 1 0 23828 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0643__B
timestamp 1606120350
transform 1 0 23368 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_593
timestamp 1606120350
transform 1 0 23552 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _0702_
timestamp 1606120350
transform 1 0 24012 0 -1 27744
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_4  _0805_
timestamp 1606120350
transform 1 0 23644 0 1 27744
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_46_258
timestamp 1606120350
transform 1 0 24840 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_259
timestamp 1606120350
transform 1 0 24932 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_262
timestamp 1606120350
transform 1 0 25208 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0699__C
timestamp 1606120350
transform 1 0 25024 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__B1
timestamp 1606120350
transform 1 0 25116 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_263
timestamp 1606120350
transform 1 0 25300 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_266
timestamp 1606120350
transform 1 0 25576 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0705__D
timestamp 1606120350
transform 1 0 25392 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0564__A
timestamp 1606120350
transform 1 0 25484 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_270
timestamp 1606120350
transform 1 0 25944 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_46_270
timestamp 1606120350
transform 1 0 25944 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__A2
timestamp 1606120350
transform 1 0 25760 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0564_
timestamp 1606120350
transform 1 0 25668 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_274
timestamp 1606120350
transform 1 0 26312 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0576__B
timestamp 1606120350
transform 1 0 26220 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0576__D
timestamp 1606120350
transform 1 0 26128 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_283
timestamp 1606120350
transform 1 0 27140 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_279
timestamp 1606120350
transform 1 0 26772 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0576__C
timestamp 1606120350
transform 1 0 27324 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0576__A
timestamp 1606120350
transform 1 0 26956 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__D
timestamp 1606120350
transform 1 0 26496 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_587
timestamp 1606120350
transform 1 0 26404 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0517_
timestamp 1606120350
transform 1 0 26496 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_46_294
timestamp 1606120350
transform 1 0 28152 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_290
timestamp 1606120350
transform 1 0 27784 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0698__D
timestamp 1606120350
transform 1 0 28336 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0642__D
timestamp 1606120350
transform 1 0 27968 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0640_
timestamp 1606120350
transform 1 0 27508 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1188_
timestamp 1606120350
transform 1 0 26680 0 1 27744
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_47_301
timestamp 1606120350
transform 1 0 28796 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_47_297
timestamp 1606120350
transform 1 0 28428 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_46_298
timestamp 1606120350
transform 1 0 28520 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1188__CLK
timestamp 1606120350
transform 1 0 28704 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__D
timestamp 1606120350
transform 1 0 28980 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0530__A
timestamp 1606120350
transform 1 0 28612 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_594
timestamp 1606120350
transform 1 0 29164 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0600_
timestamp 1606120350
transform 1 0 29256 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_309
timestamp 1606120350
transform 1 0 29532 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0600__A
timestamp 1606120350
transform 1 0 29716 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_313
timestamp 1606120350
transform 1 0 29900 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_314
timestamp 1606120350
transform 1 0 29992 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_302
timestamp 1606120350
transform 1 0 28888 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_588
timestamp 1606120350
transform 1 0 32016 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__D
timestamp 1606120350
transform 1 0 32384 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_326
timestamp 1606120350
transform 1 0 31096 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_334
timestamp 1606120350
transform 1 0 31832 0 -1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_337
timestamp 1606120350
transform 1 0 32108 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_325
timestamp 1606120350
transform 1 0 31004 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_47_337
timestamp 1606120350
transform 1 0 32108 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_47_342
timestamp 1606120350
transform 1 0 32568 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1141__CLK
timestamp 1606120350
transform 1 0 32752 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_349
timestamp 1606120350
transform 1 0 33212 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_361
timestamp 1606120350
transform 1 0 34316 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_346
timestamp 1606120350
transform 1 0 32936 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_358
timestamp 1606120350
transform 1 0 34040 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_595
timestamp 1606120350
transform 1 0 34776 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_373
timestamp 1606120350
transform 1 0 35420 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_385
timestamp 1606120350
transform 1 0 36524 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_367
timestamp 1606120350
transform 1 0 34868 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_379
timestamp 1606120350
transform 1 0 35972 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1606120350
transform -1 0 38824 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1606120350
transform -1 0 38824 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_589
timestamp 1606120350
transform 1 0 37628 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_398
timestamp 1606120350
transform 1 0 37720 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_406
timestamp 1606120350
transform 1 0 38456 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_391
timestamp 1606120350
transform 1 0 37076 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_403
timestamp 1606120350
transform 1 0 38180 0 1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1606120350
transform 1 0 1104 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1606120350
transform 1 0 1380 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1606120350
transform 1 0 2484 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_596
timestamp 1606120350
transform 1 0 3956 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_27
timestamp 1606120350
transform 1 0 3588 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_32
timestamp 1606120350
transform 1 0 4048 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_44
timestamp 1606120350
transform 1 0 5152 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__D
timestamp 1606120350
transform 1 0 7268 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1105__CLK
timestamp 1606120350
transform 1 0 6900 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_56
timestamp 1606120350
transform 1 0 6256 0 -1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_62
timestamp 1606120350
transform 1 0 6808 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_65
timestamp 1606120350
transform 1 0 7084 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0810_
timestamp 1606120350
transform 1 0 7544 0 -1 28832
box -38 -48 1326 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__D
timestamp 1606120350
transform 1 0 9384 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__A1
timestamp 1606120350
transform 1 0 9016 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_69
timestamp 1606120350
transform 1 0 7452 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_84
timestamp 1606120350
transform 1 0 8832 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_88
timestamp 1606120350
transform 1 0 9200 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0661_
timestamp 1606120350
transform 1 0 10672 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_597
timestamp 1606120350
transform 1 0 9568 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__B2
timestamp 1606120350
transform 1 0 10488 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0768__B1
timestamp 1606120350
transform 1 0 10120 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_93
timestamp 1606120350
transform 1 0 9660 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_97
timestamp 1606120350
transform 1 0 10028 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_100
timestamp 1606120350
transform 1 0 10304 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_113
timestamp 1606120350
transform 1 0 11500 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _0761_
timestamp 1606120350
transform 1 0 12236 0 -1 28832
box -38 -48 1326 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0542__C
timestamp 1606120350
transform 1 0 11776 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__B1
timestamp 1606120350
transform 1 0 13708 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_118
timestamp 1606120350
transform 1 0 11960 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_135
timestamp 1606120350
transform 1 0 13524 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _0767_
timestamp 1606120350
transform 1 0 15272 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_598
timestamp 1606120350
transform 1 0 15180 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__B
timestamp 1606120350
transform 1 0 14996 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__B
timestamp 1606120350
transform 1 0 14628 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__C
timestamp 1606120350
transform 1 0 14260 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_139
timestamp 1606120350
transform 1 0 13892 0 -1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_145
timestamp 1606120350
transform 1 0 14444 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_149
timestamp 1606120350
transform 1 0 14812 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0566_
timestamp 1606120350
transform 1 0 17388 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0537__A2
timestamp 1606120350
transform 1 0 16560 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__A
timestamp 1606120350
transform 1 0 16928 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__C
timestamp 1606120350
transform 1 0 17848 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_166
timestamp 1606120350
transform 1 0 16376 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_170
timestamp 1606120350
transform 1 0 16744 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_174
timestamp 1606120350
transform 1 0 17112 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_48_180
timestamp 1606120350
transform 1 0 17664 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0698_
timestamp 1606120350
transform 1 0 18400 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__A
timestamp 1606120350
transform 1 0 19412 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__C
timestamp 1606120350
transform 1 0 19872 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0618__B
timestamp 1606120350
transform 1 0 18216 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_184
timestamp 1606120350
transform 1 0 18032 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1606120350
transform 1 0 19228 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_48_201
timestamp 1606120350
transform 1 0 19596 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _0645_
timestamp 1606120350
transform 1 0 20884 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_599
timestamp 1606120350
transform 1 0 20792 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__A
timestamp 1606120350
transform 1 0 21896 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0645__B
timestamp 1606120350
transform 1 0 20608 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0644__C
timestamp 1606120350
transform 1 0 20240 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_206
timestamp 1606120350
transform 1 0 20056 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_210
timestamp 1606120350
transform 1 0 20424 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_224
timestamp 1606120350
transform 1 0 21712 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_228
timestamp 1606120350
transform 1 0 22080 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0516_
timestamp 1606120350
transform 1 0 24012 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _0643_
timestamp 1606120350
transform 1 0 22448 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__B
timestamp 1606120350
transform 1 0 23828 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__B
timestamp 1606120350
transform 1 0 22264 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__A
timestamp 1606120350
transform 1 0 23460 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_241
timestamp 1606120350
transform 1 0 23276 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_245
timestamp 1606120350
transform 1 0 23644 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__A1
timestamp 1606120350
transform 1 0 25024 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0805__B2
timestamp 1606120350
transform 1 0 25392 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__B1_N
timestamp 1606120350
transform 1 0 26128 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__A1
timestamp 1606120350
transform 1 0 25760 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_258
timestamp 1606120350
transform 1 0 24840 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_262
timestamp 1606120350
transform 1 0 25208 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_266
timestamp 1606120350
transform 1 0 25576 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_270
timestamp 1606120350
transform 1 0 25944 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_48_274
timestamp 1606120350
transform 1 0 26312 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0530_
timestamp 1606120350
transform 1 0 28060 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _0576_
timestamp 1606120350
transform 1 0 26496 0 -1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_600
timestamp 1606120350
transform 1 0 26404 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0644__D
timestamp 1606120350
transform 1 0 27508 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1102__D
timestamp 1606120350
transform 1 0 27876 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_285
timestamp 1606120350
transform 1 0 27324 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_289
timestamp 1606120350
transform 1 0 27692 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_296
timestamp 1606120350
transform 1 0 28336 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0516__A
timestamp 1606120350
transform 1 0 28520 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1102__CLK
timestamp 1606120350
transform 1 0 28888 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_48_300
timestamp 1606120350
transform 1 0 28704 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_304
timestamp 1606120350
transform 1 0 29072 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_316
timestamp 1606120350
transform 1 0 30176 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1141_
timestamp 1606120350
transform 1 0 32384 0 -1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_601
timestamp 1606120350
transform 1 0 32016 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_328
timestamp 1606120350
transform 1 0 31280 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_337
timestamp 1606120350
transform 1 0 32108 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_359
timestamp 1606120350
transform 1 0 34132 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_371
timestamp 1606120350
transform 1 0 35236 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_383
timestamp 1606120350
transform 1 0 36340 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1606120350
transform -1 0 38824 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_602
timestamp 1606120350
transform 1 0 37628 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_48_395
timestamp 1606120350
transform 1 0 37444 0 -1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_398
timestamp 1606120350
transform 1 0 37720 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_406
timestamp 1606120350
transform 1 0 38456 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1606120350
transform 1 0 1104 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__D
timestamp 1606120350
transform 1 0 1564 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1165__CLK
timestamp 1606120350
transform 1 0 1932 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_3
timestamp 1606120350
transform 1 0 1380 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_7
timestamp 1606120350
transform 1 0 1748 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_11
timestamp 1606120350
transform 1 0 2116 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_23
timestamp 1606120350
transform 1 0 3220 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_35
timestamp 1606120350
transform 1 0 4324 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1105_
timestamp 1606120350
transform 1 0 7268 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_603
timestamp 1606120350
transform 1 0 6716 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__D
timestamp 1606120350
transform 1 0 6992 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1104__CLK
timestamp 1606120350
transform 1 0 6532 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_47
timestamp 1606120350
transform 1 0 5428 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_62
timestamp 1606120350
transform 1 0 6808 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_66
timestamp 1606120350
transform 1 0 7176 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__D
timestamp 1606120350
transform 1 0 9384 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_86
timestamp 1606120350
transform 1 0 9016 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_92
timestamp 1606120350
transform 1 0 9568 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0713__A
timestamp 1606120350
transform 1 0 9752 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_96
timestamp 1606120350
transform 1 0 9936 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__A2
timestamp 1606120350
transform 1 0 10120 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0520_
timestamp 1606120350
transform 1 0 10304 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_103
timestamp 1606120350
transform 1 0 10580 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0520__A
timestamp 1606120350
transform 1 0 10764 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_107
timestamp 1606120350
transform 1 0 10948 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0536__A
timestamp 1606120350
transform 1 0 11132 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_114
timestamp 1606120350
transform 1 0 11592 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0534_
timestamp 1606120350
transform 1 0 11316 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _0754_
timestamp 1606120350
transform 1 0 13340 0 1 28832
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_604
timestamp 1606120350
transform 1 0 12328 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0753__A2
timestamp 1606120350
transform 1 0 13156 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0542__B
timestamp 1606120350
transform 1 0 11776 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0534__A
timestamp 1606120350
transform 1 0 12144 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0542__A
timestamp 1606120350
transform 1 0 12604 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_118
timestamp 1606120350
transform 1 0 11960 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_123
timestamp 1606120350
transform 1 0 12420 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_127
timestamp 1606120350
transform 1 0 12788 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0514_
timestamp 1606120350
transform 1 0 15364 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__B
timestamp 1606120350
transform 1 0 15180 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0686__C
timestamp 1606120350
transform 1 0 14812 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_147
timestamp 1606120350
transform 1 0 14628 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_151
timestamp 1606120350
transform 1 0 14996 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_158
timestamp 1606120350
transform 1 0 15640 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0689_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 16376 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0514__A
timestamp 1606120350
transform 1 0 15824 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0689__A
timestamp 1606120350
transform 1 0 16192 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__C
timestamp 1606120350
transform 1 0 17756 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0700__A
timestamp 1606120350
transform 1 0 17388 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_162
timestamp 1606120350
transform 1 0 16008 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_175
timestamp 1606120350
transform 1 0 17204 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_179
timestamp 1606120350
transform 1 0 17572 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0697_
timestamp 1606120350
transform 1 0 18584 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_605
timestamp 1606120350
transform 1 0 17940 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0581__A
timestamp 1606120350
transform 1 0 19596 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__C
timestamp 1606120350
transform 1 0 18400 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_184
timestamp 1606120350
transform 1 0 18032 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_199
timestamp 1606120350
transform 1 0 19412 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_203
timestamp 1606120350
transform 1 0 19780 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _0558_
timestamp 1606120350
transform 1 0 21896 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _0644_
timestamp 1606120350
transform 1 0 20332 0 1 28832
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__D
timestamp 1606120350
transform 1 0 21712 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0644__A
timestamp 1606120350
transform 1 0 20148 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__C
timestamp 1606120350
transform 1 0 21344 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_218
timestamp 1606120350
transform 1 0 21160 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_222
timestamp 1606120350
transform 1 0 21528 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1102_
timestamp 1606120350
transform 1 0 23644 0 1 28832
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_606
timestamp 1606120350
transform 1 0 23552 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__A
timestamp 1606120350
transform 1 0 23368 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0597__C
timestamp 1606120350
transform 1 0 23000 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_49_235
timestamp 1606120350
transform 1 0 22724 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_49_240
timestamp 1606120350
transform 1 0 23184 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__a21bo_4  _0929_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 26128 0 1 28832
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__A
timestamp 1606120350
transform 1 0 25944 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__B
timestamp 1606120350
transform 1 0 25576 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_264
timestamp 1606120350
transform 1 0 25392 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_268
timestamp 1606120350
transform 1 0 25760 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0606_
timestamp 1606120350
transform 1 0 28060 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__C
timestamp 1606120350
transform 1 0 27508 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0929__A2
timestamp 1606120350
transform 1 0 27876 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_285
timestamp 1606120350
transform 1 0 27324 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_289
timestamp 1606120350
transform 1 0 27692 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_296
timestamp 1606120350
transform 1 0 28336 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_607
timestamp 1606120350
transform 1 0 29164 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0606__A
timestamp 1606120350
transform 1 0 28520 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0581__B
timestamp 1606120350
transform 1 0 28888 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0555__A
timestamp 1606120350
transform 1 0 29440 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_49_300
timestamp 1606120350
transform 1 0 28704 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_49_304
timestamp 1606120350
transform 1 0 29072 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_49_306
timestamp 1606120350
transform 1 0 29256 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_310
timestamp 1606120350
transform 1 0 29624 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_322
timestamp 1606120350
transform 1 0 30728 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_334
timestamp 1606120350
transform 1 0 31832 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_346
timestamp 1606120350
transform 1 0 32936 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_358
timestamp 1606120350
transform 1 0 34040 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_608
timestamp 1606120350
transform 1 0 34776 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_367
timestamp 1606120350
transform 1 0 34868 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_379
timestamp 1606120350
transform 1 0 35972 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1606120350
transform -1 0 38824 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_391
timestamp 1606120350
transform 1 0 37076 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_403
timestamp 1606120350
transform 1 0 38180 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1165_
timestamp 1606120350
transform 1 0 1380 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1606120350
transform 1 0 1104 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_50_22
timestamp 1606120350
transform 1 0 3128 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_609
timestamp 1606120350
transform 1 0 3956 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_50_30
timestamp 1606120350
transform 1 0 3864 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_32
timestamp 1606120350
transform 1 0 4048 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_44
timestamp 1606120350
transform 1 0 5152 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1104_
timestamp 1606120350
transform 1 0 6808 0 -1 29920
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__D
timestamp 1606120350
transform 1 0 6624 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_56
timestamp 1606120350
transform 1 0 6256 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__B2
timestamp 1606120350
transform 1 0 9384 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0542__D
timestamp 1606120350
transform 1 0 9016 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_81
timestamp 1606120350
transform 1 0 8556 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_85
timestamp 1606120350
transform 1 0 8924 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_50_88
timestamp 1606120350
transform 1 0 9200 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_50_93
timestamp 1606120350
transform 1 0 9660 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_610
timestamp 1606120350
transform 1 0 9568 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0713_
timestamp 1606120350
transform 1 0 9752 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_97
timestamp 1606120350
transform 1 0 10028 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0539__A
timestamp 1606120350
transform 1 0 10212 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_101
timestamp 1606120350
transform 1 0 10396 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0754__B1
timestamp 1606120350
transform 1 0 10580 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0536_
timestamp 1606120350
transform 1 0 10764 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_108
timestamp 1606120350
transform 1 0 11040 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0540__A
timestamp 1606120350
transform 1 0 11224 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_112
timestamp 1606120350
transform 1 0 11408 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__A1
timestamp 1606120350
transform 1 0 11592 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0542_
timestamp 1606120350
transform 1 0 11776 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _0753_
timestamp 1606120350
transform 1 0 13340 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__C
timestamp 1606120350
transform 1 0 13156 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__D
timestamp 1606120350
transform 1 0 12788 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_125
timestamp 1606120350
transform 1 0 12604 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_129
timestamp 1606120350
transform 1 0 12972 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_611
timestamp 1606120350
transform 1 0 15180 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0515__A
timestamp 1606120350
transform 1 0 15456 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__A
timestamp 1606120350
transform 1 0 14720 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_145
timestamp 1606120350
transform 1 0 14444 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_50_150
timestamp 1606120350
transform 1 0 14904 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_154
timestamp 1606120350
transform 1 0 15272 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_158
timestamp 1606120350
transform 1 0 15640 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _0686_
timestamp 1606120350
transform 1 0 16192 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _0700_
timestamp 1606120350
transform 1 0 17756 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__C
timestamp 1606120350
transform 1 0 17204 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__A
timestamp 1606120350
transform 1 0 16008 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__A
timestamp 1606120350
transform 1 0 17572 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_173
timestamp 1606120350
transform 1 0 17020 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_177
timestamp 1606120350
transform 1 0 17388 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0581_
timestamp 1606120350
transform 1 0 19412 0 -1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__B1
timestamp 1606120350
transform 1 0 19228 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__D1
timestamp 1606120350
transform 1 0 18860 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_190
timestamp 1606120350
transform 1 0 18584 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_50_195
timestamp 1606120350
transform 1 0 19044 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0701_
timestamp 1606120350
transform 1 0 20884 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_612
timestamp 1606120350
transform 1 0 20792 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__A2
timestamp 1606120350
transform 1 0 20240 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__C
timestamp 1606120350
transform 1 0 21896 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0644__B
timestamp 1606120350
transform 1 0 20608 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_206
timestamp 1606120350
transform 1 0 20056 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_210
timestamp 1606120350
transform 1 0 20424 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_224
timestamp 1606120350
transform 1 0 21712 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_228
timestamp 1606120350
transform 1 0 22080 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0555_
timestamp 1606120350
transform 1 0 22448 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__or3_4  _0597_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 24012 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0545__C
timestamp 1606120350
transform 1 0 22264 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__B
timestamp 1606120350
transform 1 0 23828 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__C
timestamp 1606120350
transform 1 0 23460 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_241
timestamp 1606120350
transform 1 0 23276 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_245
timestamp 1606120350
transform 1 0 23644 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0586__B
timestamp 1606120350
transform 1 0 25208 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__D
timestamp 1606120350
transform 1 0 25576 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__C
timestamp 1606120350
transform 1 0 25944 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_258
timestamp 1606120350
transform 1 0 24840 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_50_264
timestamp 1606120350
transform 1 0 25392 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_268
timestamp 1606120350
transform 1 0 25760 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_50_272
timestamp 1606120350
transform 1 0 26128 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _0584_
timestamp 1606120350
transform 1 0 26496 0 -1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_613
timestamp 1606120350
transform 1 0 26404 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0701__D
timestamp 1606120350
transform 1 0 27508 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0584__D
timestamp 1606120350
transform 1 0 27876 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0697__D
timestamp 1606120350
transform 1 0 28244 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_285
timestamp 1606120350
transform 1 0 27324 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_289
timestamp 1606120350
transform 1 0 27692 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_293
timestamp 1606120350
transform 1 0 28060 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0558__B
timestamp 1606120350
transform 1 0 28612 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_50_297
timestamp 1606120350
transform 1 0 28428 0 -1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_301
timestamp 1606120350
transform 1 0 28796 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_313
timestamp 1606120350
transform 1 0 29900 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_614
timestamp 1606120350
transform 1 0 32016 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_325
timestamp 1606120350
transform 1 0 31004 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_333
timestamp 1606120350
transform 1 0 31740 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_337
timestamp 1606120350
transform 1 0 32108 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_349
timestamp 1606120350
transform 1 0 33212 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_361
timestamp 1606120350
transform 1 0 34316 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_373
timestamp 1606120350
transform 1 0 35420 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_385
timestamp 1606120350
transform 1 0 36524 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1606120350
transform -1 0 38824 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_615
timestamp 1606120350
transform 1 0 37628 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_398
timestamp 1606120350
transform 1 0 37720 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_406
timestamp 1606120350
transform 1 0 38456 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1606120350
transform 1 0 1104 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1606120350
transform 1 0 1380 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1606120350
transform 1 0 2484 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1606120350
transform 1 0 3588 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1606120350
transform 1 0 4692 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_616
timestamp 1606120350
transform 1 0 6716 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__A1
timestamp 1606120350
transform 1 0 7084 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__D
timestamp 1606120350
transform 1 0 6532 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0540__D
timestamp 1606120350
transform 1 0 6164 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1606120350
transform 1 0 5796 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_57
timestamp 1606120350
transform 1 0 6348 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_62
timestamp 1606120350
transform 1 0 6808 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_67
timestamp 1606120350
transform 1 0 7268 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0809_
timestamp 1606120350
transform 1 0 7636 0 1 29920
box -38 -48 1326 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0652__A
timestamp 1606120350
transform 1 0 9108 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0680__A
timestamp 1606120350
transform 1 0 7452 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_85
timestamp 1606120350
transform 1 0 8924 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_89
timestamp 1606120350
transform 1 0 9292 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0531_
timestamp 1606120350
transform 1 0 9752 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _0540_
timestamp 1606120350
transform 1 0 10764 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0540__B
timestamp 1606120350
transform 1 0 10580 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0540__C
timestamp 1606120350
transform 1 0 10212 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0531__A
timestamp 1606120350
transform 1 0 9568 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_97
timestamp 1606120350
transform 1 0 10028 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_101
timestamp 1606120350
transform 1 0 10396 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_114
timestamp 1606120350
transform 1 0 11592 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0721_
timestamp 1606120350
transform 1 0 13156 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_617
timestamp 1606120350
transform 1 0 12328 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__B
timestamp 1606120350
transform 1 0 12972 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__A
timestamp 1606120350
transform 1 0 12604 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__B
timestamp 1606120350
transform 1 0 12144 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__C
timestamp 1606120350
transform 1 0 11776 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_118
timestamp 1606120350
transform 1 0 11960 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_123
timestamp 1606120350
transform 1 0 12420 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_127
timestamp 1606120350
transform 1 0 12788 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0675_
timestamp 1606120350
transform 1 0 14720 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0723__B
timestamp 1606120350
transform 1 0 14168 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__C
timestamp 1606120350
transform 1 0 14536 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_140
timestamp 1606120350
transform 1 0 13984 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_144
timestamp 1606120350
transform 1 0 14352 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_157
timestamp 1606120350
transform 1 0 15548 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _0738_
timestamp 1606120350
transform 1 0 16376 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__B
timestamp 1606120350
transform 1 0 17756 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__A
timestamp 1606120350
transform 1 0 17388 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__A
timestamp 1606120350
transform 1 0 16192 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0738__B
timestamp 1606120350
transform 1 0 15824 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_162
timestamp 1606120350
transform 1 0 16008 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_175
timestamp 1606120350
transform 1 0 17204 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_179
timestamp 1606120350
transform 1 0 17572 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__a2111oi_4  _0596_
timestamp 1606120350
transform 1 0 19688 0 1 29920
box -38 -48 2062 592
use sky130_fd_sc_hd__and4_4  _0741_
timestamp 1606120350
transform 1 0 18032 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_618
timestamp 1606120350
transform 1 0 17940 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__B
timestamp 1606120350
transform 1 0 19044 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__C1
timestamp 1606120350
transform 1 0 19504 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_193
timestamp 1606120350
transform 1 0 18860 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_197
timestamp 1606120350
transform 1 0 19228 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__A
timestamp 1606120350
transform 1 0 21896 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_224
timestamp 1606120350
transform 1 0 21712 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_228
timestamp 1606120350
transform 1 0 22080 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0569_
timestamp 1606120350
transform 1 0 22448 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _0619_
timestamp 1606120350
transform 1 0 23644 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_619
timestamp 1606120350
transform 1 0 23552 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__B
timestamp 1606120350
transform 1 0 22264 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0545__A
timestamp 1606120350
transform 1 0 22908 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0545__B
timestamp 1606120350
transform 1 0 23276 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_235
timestamp 1606120350
transform 1 0 22724 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_239
timestamp 1606120350
transform 1 0 23092 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_243
timestamp 1606120350
transform 1 0 23460 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _0586_
timestamp 1606120350
transform 1 0 25208 0 1 29920
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0586__A
timestamp 1606120350
transform 1 0 25024 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0588__A
timestamp 1606120350
transform 1 0 24656 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0619__A
timestamp 1606120350
transform 1 0 26220 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_254
timestamp 1606120350
transform 1 0 24472 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_258
timestamp 1606120350
transform 1 0 24840 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_271
timestamp 1606120350
transform 1 0 26036 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0617_
timestamp 1606120350
transform 1 0 26772 0 1 29920
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0617__A
timestamp 1606120350
transform 1 0 27600 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0617__B
timestamp 1606120350
transform 1 0 26588 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0586__D
timestamp 1606120350
transform 1 0 27968 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0569__A
timestamp 1606120350
transform 1 0 28336 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_275
timestamp 1606120350
transform 1 0 26404 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_286
timestamp 1606120350
transform 1 0 27416 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_290
timestamp 1606120350
transform 1 0 27784 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_294
timestamp 1606120350
transform 1 0 28152 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_620
timestamp 1606120350
transform 1 0 29164 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__D
timestamp 1606120350
transform 1 0 28704 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1152__CLK
timestamp 1606120350
transform 1 0 29440 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_51_298
timestamp 1606120350
transform 1 0 28520 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_51_302
timestamp 1606120350
transform 1 0 28888 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_306
timestamp 1606120350
transform 1 0 29256 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_310
timestamp 1606120350
transform 1 0 29624 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_322
timestamp 1606120350
transform 1 0 30728 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_334
timestamp 1606120350
transform 1 0 31832 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_346
timestamp 1606120350
transform 1 0 32936 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_358
timestamp 1606120350
transform 1 0 34040 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_621
timestamp 1606120350
transform 1 0 34776 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_367
timestamp 1606120350
transform 1 0 34868 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_379
timestamp 1606120350
transform 1 0 35972 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1606120350
transform -1 0 38824 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_391
timestamp 1606120350
transform 1 0 37076 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_403
timestamp 1606120350
transform 1 0 38180 0 1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1606120350
transform 1 0 1104 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1606120350
transform 1 0 1104 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1606120350
transform 1 0 1380 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1606120350
transform 1 0 2484 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1606120350
transform 1 0 1380 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1606120350
transform 1 0 2484 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_622
timestamp 1606120350
transform 1 0 3956 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_27
timestamp 1606120350
transform 1 0 3588 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_32
timestamp 1606120350
transform 1 0 4048 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_44
timestamp 1606120350
transform 1 0 5152 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1606120350
transform 1 0 3588 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1606120350
transform 1 0 4692 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_51
timestamp 1606120350
transform 1 0 5796 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_62
timestamp 1606120350
transform 1 0 6808 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_62
timestamp 1606120350
transform 1 0 6808 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_56
timestamp 1606120350
transform 1 0 6256 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__CLK
timestamp 1606120350
transform 1 0 6532 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__A2
timestamp 1606120350
transform 1 0 6624 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_629
timestamp 1606120350
transform 1 0 6716 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_66
timestamp 1606120350
transform 1 0 7176 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_66
timestamp 1606120350
transform 1 0 7176 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1098__D
timestamp 1606120350
transform 1 0 6992 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__D
timestamp 1606120350
transform 1 0 6992 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__B1
timestamp 1606120350
transform 1 0 7360 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0669__A
timestamp 1606120350
transform 1 0 7360 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_77
timestamp 1606120350
transform 1 0 8188 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_73
timestamp 1606120350
transform 1 0 7820 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__A2
timestamp 1606120350
transform 1 0 8372 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0809__B2
timestamp 1606120350
transform 1 0 8004 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0680_
timestamp 1606120350
transform 1 0 7544 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_89
timestamp 1606120350
transform 1 0 9292 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_88
timestamp 1606120350
transform 1 0 9200 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_84
timestamp 1606120350
transform 1 0 8832 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0675__D
timestamp 1606120350
transform 1 0 9016 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__D
timestamp 1606120350
transform 1 0 9384 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0653__A
timestamp 1606120350
transform 1 0 9476 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0652_
timestamp 1606120350
transform 1 0 8556 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1150_
timestamp 1606120350
transform 1 0 7544 0 1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_623
timestamp 1606120350
transform 1 0 9568 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__A2
timestamp 1606120350
transform 1 0 9844 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0800__B1
timestamp 1606120350
transform 1 0 9936 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_93
timestamp 1606120350
transform 1 0 9660 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_93
timestamp 1606120350
transform 1 0 9660 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0539_
timestamp 1606120350
transform 1 0 10120 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0521__C
timestamp 1606120350
transform 1 0 10212 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_101
timestamp 1606120350
transform 1 0 10396 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_53_97
timestamp 1606120350
transform 1 0 10028 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_101
timestamp 1606120350
transform 1 0 10396 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_114
timestamp 1606120350
transform 1 0 11592 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_107
timestamp 1606120350
transform 1 0 10948 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0521__B
timestamp 1606120350
transform 1 0 10764 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0521__A
timestamp 1606120350
transform 1 0 10580 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0521_
timestamp 1606120350
transform 1 0 10764 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_4  _0800_
timestamp 1606120350
transform 1 0 11132 0 -1 31008
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_53_118
timestamp 1606120350
transform 1 0 11960 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_123
timestamp 1606120350
transform 1 0 12420 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__D
timestamp 1606120350
transform 1 0 11776 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__A
timestamp 1606120350
transform 1 0 12144 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_630
timestamp 1606120350
transform 1 0 12328 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_135
timestamp 1606120350
transform 1 0 13524 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_132
timestamp 1606120350
transform 1 0 13248 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_128
timestamp 1606120350
transform 1 0 12880 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__D
timestamp 1606120350
transform 1 0 12696 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0721__A
timestamp 1606120350
transform 1 0 13064 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__C
timestamp 1606120350
transform 1 0 13432 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__B
timestamp 1606120350
transform 1 0 13708 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0723_
timestamp 1606120350
transform 1 0 13616 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_4  _0798_
timestamp 1606120350
transform 1 0 12420 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_143
timestamp 1606120350
transform 1 0 14260 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_139
timestamp 1606120350
transform 1 0 13892 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_145
timestamp 1606120350
transform 1 0 14444 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__C
timestamp 1606120350
transform 1 0 14536 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0676__A
timestamp 1606120350
transform 1 0 14076 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_149
timestamp 1606120350
transform 1 0 14812 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0546__D
timestamp 1606120350
transform 1 0 14628 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0546__B
timestamp 1606120350
transform 1 0 14996 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_624
timestamp 1606120350
transform 1 0 15180 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _0677_
timestamp 1606120350
transform 1 0 14720 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0515_
timestamp 1606120350
transform 1 0 15272 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_157
timestamp 1606120350
transform 1 0 15548 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_157
timestamp 1606120350
transform 1 0 15548 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__C
timestamp 1606120350
transform 1 0 15732 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0546__A
timestamp 1606120350
transform 1 0 15732 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_161
timestamp 1606120350
transform 1 0 15916 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_161
timestamp 1606120350
transform 1 0 15916 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__B
timestamp 1606120350
transform 1 0 16100 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__A
timestamp 1606120350
transform 1 0 16192 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0682_
timestamp 1606120350
transform 1 0 16376 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _0679_
timestamp 1606120350
transform 1 0 16284 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_179
timestamp 1606120350
transform 1 0 17572 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_175
timestamp 1606120350
transform 1 0 17204 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_178
timestamp 1606120350
transform 1 0 17480 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_52_174
timestamp 1606120350
transform 1 0 17112 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0679__C
timestamp 1606120350
transform 1 0 17296 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__B
timestamp 1606120350
transform 1 0 17388 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_52_182
timestamp 1606120350
transform 1 0 17848 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__A
timestamp 1606120350
transform 1 0 17756 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__C
timestamp 1606120350
transform 1 0 17940 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_631
timestamp 1606120350
transform 1 0 17940 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _0743_
timestamp 1606120350
transform 1 0 18124 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _0726_
timestamp 1606120350
transform 1 0 18032 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_197
timestamp 1606120350
transform 1 0 19228 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_193
timestamp 1606120350
transform 1 0 18860 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_198
timestamp 1606120350
transform 1 0 19320 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1606120350
transform 1 0 18952 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__B2
timestamp 1606120350
transform 1 0 19136 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__D
timestamp 1606120350
transform 1 0 19044 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__C
timestamp 1606120350
transform 1 0 19596 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__B
timestamp 1606120350
transform 1 0 19412 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0742_
timestamp 1606120350
transform 1 0 19596 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0582_
timestamp 1606120350
transform 1 0 19780 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_214
timestamp 1606120350
transform 1 0 20792 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_210
timestamp 1606120350
transform 1 0 20424 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_210
timestamp 1606120350
transform 1 0 20424 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_206
timestamp 1606120350
transform 1 0 20056 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0589__C
timestamp 1606120350
transform 1 0 20608 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0582__A
timestamp 1606120350
transform 1 0 20240 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__C
timestamp 1606120350
transform 1 0 20608 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_625
timestamp 1606120350
transform 1 0 20792 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _0724_
timestamp 1606120350
transform 1 0 20884 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_52_224
timestamp 1606120350
transform 1 0 21712 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__B
timestamp 1606120350
transform 1 0 20976 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0725_
timestamp 1606120350
transform 1 0 21160 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_227
timestamp 1606120350
transform 1 0 21988 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_228
timestamp 1606120350
transform 1 0 22080 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0589__A
timestamp 1606120350
transform 1 0 21896 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_53_235
timestamp 1606120350
transform 1 0 22724 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_231
timestamp 1606120350
transform 1 0 22356 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0589__D
timestamp 1606120350
transform 1 0 22264 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0589__B
timestamp 1606120350
transform 1 0 22540 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__B
timestamp 1606120350
transform 1 0 23000 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__A
timestamp 1606120350
transform 1 0 22172 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _0545_
timestamp 1606120350
transform 1 0 22448 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_240
timestamp 1606120350
transform 1 0 23184 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_247
timestamp 1606120350
transform 1 0 23828 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_241
timestamp 1606120350
transform 1 0 23276 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__A
timestamp 1606120350
transform 1 0 23644 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__A
timestamp 1606120350
transform 1 0 23368 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_632
timestamp 1606120350
transform 1 0 23552 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _0587_
timestamp 1606120350
transform 1 0 23644 0 1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0588_
timestamp 1606120350
transform 1 0 24012 0 -1 31008
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_53_254
timestamp 1606120350
transform 1 0 24472 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__C
timestamp 1606120350
transform 1 0 24656 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_258
timestamp 1606120350
transform 1 0 24840 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_258
timestamp 1606120350
transform 1 0 24840 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__C
timestamp 1606120350
transform 1 0 25024 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_265
timestamp 1606120350
transform 1 0 25484 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_264
timestamp 1606120350
transform 1 0 25392 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0586__C
timestamp 1606120350
transform 1 0 25208 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0510_
timestamp 1606120350
transform 1 0 25208 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_269
timestamp 1606120350
transform 1 0 25852 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_52_268
timestamp 1606120350
transform 1 0 25760 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__D
timestamp 1606120350
transform 1 0 25668 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0743__D
timestamp 1606120350
transform 1 0 25944 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0619__C
timestamp 1606120350
transform 1 0 25576 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_272
timestamp 1606120350
transform 1 0 26128 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0741__D
timestamp 1606120350
transform 1 0 26036 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0503_
timestamp 1606120350
transform 1 0 26220 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_280
timestamp 1606120350
transform 1 0 26864 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_276
timestamp 1606120350
transform 1 0 26496 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_52_280
timestamp 1606120350
transform 1 0 26864 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_52_276
timestamp 1606120350
transform 1 0 26496 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0585__D
timestamp 1606120350
transform 1 0 27048 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0596__A1
timestamp 1606120350
transform 1 0 26680 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1160__D
timestamp 1606120350
transform 1 0 26680 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_626
timestamp 1606120350
transform 1 0 26404 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0533_
timestamp 1606120350
transform 1 0 27232 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_295
timestamp 1606120350
transform 1 0 28244 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_291
timestamp 1606120350
transform 1 0 27876 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_287
timestamp 1606120350
transform 1 0 27508 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0726__C
timestamp 1606120350
transform 1 0 28060 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0533__A
timestamp 1606120350
transform 1 0 27692 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1152_
timestamp 1606120350
transform 1 0 27140 0 -1 31008
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_53_306
timestamp 1606120350
transform 1 0 29256 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_303
timestamp 1606120350
transform 1 0 28980 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_53_299
timestamp 1606120350
transform 1 0 28612 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0587__B
timestamp 1606120350
transform 1 0 28796 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0510__A
timestamp 1606120350
transform 1 0 28428 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__D
timestamp 1606120350
transform 1 0 29440 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_633
timestamp 1606120350
transform 1 0 29164 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_310
timestamp 1606120350
transform 1 0 29624 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1134__CLK
timestamp 1606120350
transform 1 0 29808 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_314
timestamp 1606120350
transform 1 0 29992 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_314
timestamp 1606120350
transform 1 0 29992 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_302
timestamp 1606120350
transform 1 0 28888 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_627
timestamp 1606120350
transform 1 0 32016 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_326
timestamp 1606120350
transform 1 0 31096 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_334
timestamp 1606120350
transform 1 0 31832 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_337
timestamp 1606120350
transform 1 0 32108 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_326
timestamp 1606120350
transform 1 0 31096 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_338
timestamp 1606120350
transform 1 0 32200 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_349
timestamp 1606120350
transform 1 0 33212 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_361
timestamp 1606120350
transform 1 0 34316 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_350
timestamp 1606120350
transform 1 0 33304 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_362
timestamp 1606120350
transform 1 0 34408 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_634
timestamp 1606120350
transform 1 0 34776 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_373
timestamp 1606120350
transform 1 0 35420 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_385
timestamp 1606120350
transform 1 0 36524 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_367
timestamp 1606120350
transform 1 0 34868 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_379
timestamp 1606120350
transform 1 0 35972 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1606120350
transform -1 0 38824 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1606120350
transform -1 0 38824 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_628
timestamp 1606120350
transform 1 0 37628 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_398
timestamp 1606120350
transform 1 0 37720 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_406
timestamp 1606120350
transform 1 0 38456 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_391
timestamp 1606120350
transform 1 0 37076 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_403
timestamp 1606120350
transform 1 0 38180 0 1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1606120350
transform 1 0 1104 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1606120350
transform 1 0 1380 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1606120350
transform 1 0 2484 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_635
timestamp 1606120350
transform 1 0 3956 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_27
timestamp 1606120350
transform 1 0 3588 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_32
timestamp 1606120350
transform 1 0 4048 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_44
timestamp 1606120350
transform 1 0 5152 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__D
timestamp 1606120350
transform 1 0 7360 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1150__CLK
timestamp 1606120350
transform 1 0 6992 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_54_56
timestamp 1606120350
transform 1 0 6256 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_66
timestamp 1606120350
transform 1 0 7176 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0669_
timestamp 1606120350
transform 1 0 7544 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_73
timestamp 1606120350
transform 1 0 7820 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__D
timestamp 1606120350
transform 1 0 8004 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_77
timestamp 1606120350
transform 1 0 8188 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__A
timestamp 1606120350
transform 1 0 8372 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0653_
timestamp 1606120350
transform 1 0 8556 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_84
timestamp 1606120350
transform 1 0 8832 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__B2
timestamp 1606120350
transform 1 0 9016 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_88
timestamp 1606120350
transform 1 0 9200 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__A1
timestamp 1606120350
transform 1 0 9384 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1098_
timestamp 1606120350
transform 1 0 10488 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_636
timestamp 1606120350
transform 1 0 9568 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0798__B1
timestamp 1606120350
transform 1 0 10304 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0521__D
timestamp 1606120350
transform 1 0 9936 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_54_93
timestamp 1606120350
transform 1 0 9660 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_98
timestamp 1606120350
transform 1 0 10120 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0676_
timestamp 1606120350
transform 1 0 13616 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__B1
timestamp 1606120350
transform 1 0 13432 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__A1
timestamp 1606120350
transform 1 0 13064 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__C1
timestamp 1606120350
transform 1 0 12696 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_121
timestamp 1606120350
transform 1 0 12236 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_125
timestamp 1606120350
transform 1 0 12604 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_128
timestamp 1606120350
transform 1 0 12880 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_132
timestamp 1606120350
transform 1 0 13248 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__nor4_4  _0546_
timestamp 1606120350
transform 1 0 15272 0 -1 32096
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_637
timestamp 1606120350
transform 1 0 15180 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0546__C
timestamp 1606120350
transform 1 0 14996 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__A
timestamp 1606120350
transform 1 0 14628 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_145
timestamp 1606120350
transform 1 0 14444 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_149
timestamp 1606120350
transform 1 0 14812 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__nor4_4  _0684_
timestamp 1606120350
transform 1 0 17572 0 -1 32096
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0682__B
timestamp 1606120350
transform 1 0 17020 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__A2
timestamp 1606120350
transform 1 0 17388 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_171
timestamp 1606120350
transform 1 0 16836 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_175
timestamp 1606120350
transform 1 0 17204 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__A
timestamp 1606120350
transform 1 0 19596 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__B1
timestamp 1606120350
transform 1 0 19964 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_196
timestamp 1606120350
transform 1 0 19136 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_200
timestamp 1606120350
transform 1 0 19504 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_203
timestamp 1606120350
transform 1 0 19780 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__nor4_4  _0589_
timestamp 1606120350
transform 1 0 21068 0 -1 32096
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_638
timestamp 1606120350
transform 1 0 20792 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__B
timestamp 1606120350
transform 1 0 20608 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_207
timestamp 1606120350
transform 1 0 20148 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_211
timestamp 1606120350
transform 1 0 20516 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_215
timestamp 1606120350
transform 1 0 20884 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0585_
timestamp 1606120350
transform 1 0 23368 0 -1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__B
timestamp 1606120350
transform 1 0 22816 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0742__D
timestamp 1606120350
transform 1 0 23184 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_234
timestamp 1606120350
transform 1 0 22632 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_238
timestamp 1606120350
transform 1 0 23000 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_251
timestamp 1606120350
transform 1 0 24196 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_255
timestamp 1606120350
transform 1 0 24564 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0619__B
timestamp 1606120350
transform 1 0 24380 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__C
timestamp 1606120350
transform 1 0 24748 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_262
timestamp 1606120350
transform 1 0 25208 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0504_
timestamp 1606120350
transform 1 0 24932 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_54_266
timestamp 1606120350
transform 1 0 25576 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0724__D
timestamp 1606120350
transform 1 0 25392 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_54_270
timestamp 1606120350
transform 1 0 25944 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0595__A
timestamp 1606120350
transform 1 0 25760 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_54_274
timestamp 1606120350
transform 1 0 26312 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0725__D
timestamp 1606120350
transform 1 0 26128 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1160_
timestamp 1606120350
transform 1 0 26680 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_639
timestamp 1606120350
transform 1 0 26404 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_276
timestamp 1606120350
transform 1 0 26496 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1134_
timestamp 1606120350
transform 1 0 29164 0 -1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_54_297
timestamp 1606120350
transform 1 0 28428 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_640
timestamp 1606120350
transform 1 0 32016 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_324
timestamp 1606120350
transform 1 0 30912 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_337
timestamp 1606120350
transform 1 0 32108 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_349
timestamp 1606120350
transform 1 0 33212 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_361
timestamp 1606120350
transform 1 0 34316 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_373
timestamp 1606120350
transform 1 0 35420 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_385
timestamp 1606120350
transform 1 0 36524 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1606120350
transform -1 0 38824 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_641
timestamp 1606120350
transform 1 0 37628 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_398
timestamp 1606120350
transform 1 0 37720 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_406
timestamp 1606120350
transform 1 0 38456 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1606120350
transform 1 0 1104 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1606120350
transform 1 0 1380 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1606120350
transform 1 0 2484 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_2_0_clk
timestamp 1606120350
transform 1 0 4876 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1606120350
transform 1 0 3588 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_39
timestamp 1606120350
transform 1 0 4692 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_44
timestamp 1606120350
transform 1 0 5152 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_642
timestamp 1606120350
transform 1 0 6716 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_2_0_clk_A
timestamp 1606120350
transform 1 0 5336 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__CLK
timestamp 1606120350
transform 1 0 7268 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_48
timestamp 1606120350
transform 1 0 5520 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_60
timestamp 1606120350
transform 1 0 6624 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_62
timestamp 1606120350
transform 1 0 6808 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_66
timestamp 1606120350
transform 1 0 7176 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0717_
timestamp 1606120350
transform 1 0 8188 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0797__B
timestamp 1606120350
transform 1 0 9384 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__B
timestamp 1606120350
transform 1 0 9016 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0717__A
timestamp 1606120350
transform 1 0 8004 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0668__A
timestamp 1606120350
transform 1 0 7636 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_69
timestamp 1606120350
transform 1 0 7452 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_73
timestamp 1606120350
transform 1 0 7820 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_84
timestamp 1606120350
transform 1 0 8832 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_88
timestamp 1606120350
transform 1 0 9200 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0655_
timestamp 1606120350
transform 1 0 10948 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _0797_
timestamp 1606120350
transform 1 0 9568 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1123__D
timestamp 1606120350
transform 1 0 10396 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__D
timestamp 1606120350
transform 1 0 10764 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_99
timestamp 1606120350
transform 1 0 10212 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_103
timestamp 1606120350
transform 1 0 10580 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_114
timestamp 1606120350
transform 1 0 11592 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_123
timestamp 1606120350
transform 1 0 12420 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_118
timestamp 1606120350
transform 1 0 11960 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0655__B
timestamp 1606120350
transform 1 0 11776 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0491__A
timestamp 1606120350
transform 1 0 12144 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_643
timestamp 1606120350
transform 1 0 12328 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0511_
timestamp 1606120350
transform 1 0 12512 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_131
timestamp 1606120350
transform 1 0 13156 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_127
timestamp 1606120350
transform 1 0 12788 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__A1
timestamp 1606120350
transform 1 0 13340 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0511__A
timestamp 1606120350
transform 1 0 12972 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _0772_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 13524 0 1 32096
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__B
timestamp 1606120350
transform 1 0 15732 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0512__A
timestamp 1606120350
transform 1 0 15272 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_152
timestamp 1606120350
transform 1 0 15088 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_55_156
timestamp 1606120350
transform 1 0 15456 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _0683_
timestamp 1606120350
transform 1 0 15916 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_clk
timestamp 1606120350
transform 1 0 17480 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__D
timestamp 1606120350
transform 1 0 16928 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__A1
timestamp 1606120350
transform 1 0 17296 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_170
timestamp 1606120350
transform 1 0 16744 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_174
timestamp 1606120350
transform 1 0 17112 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_181
timestamp 1606120350
transform 1 0 17756 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _0590_
timestamp 1606120350
transform 1 0 18308 0 1 32096
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_644
timestamp 1606120350
transform 1 0 17940 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_55_184
timestamp 1606120350
transform 1 0 18032 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_204
timestamp 1606120350
transform 1 0 19872 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0727_
timestamp 1606120350
transform 1 0 20608 0 1 32096
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0513__A
timestamp 1606120350
transform 1 0 20056 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__A
timestamp 1606120350
transform 1 0 20424 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__A
timestamp 1606120350
transform 1 0 21620 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0628__A
timestamp 1606120350
transform 1 0 21988 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_208
timestamp 1606120350
transform 1 0 20240 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_221
timestamp 1606120350
transform 1 0 21436 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1606120350
transform 1 0 21804 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0595_
timestamp 1606120350
transform 1 0 22172 0 1 32096
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_4  _1099_
timestamp 1606120350
transform 1 0 23644 0 1 32096
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_645
timestamp 1606120350
transform 1 0 23552 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0628__B
timestamp 1606120350
transform 1 0 23000 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__C
timestamp 1606120350
transform 1 0 23368 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_236
timestamp 1606120350
transform 1 0 22816 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_240
timestamp 1606120350
transform 1 0 23184 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0695_
timestamp 1606120350
transform 1 0 26128 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__D
timestamp 1606120350
transform 1 0 25576 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__D
timestamp 1606120350
transform 1 0 25944 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_264
timestamp 1606120350
transform 1 0 25392 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_268
timestamp 1606120350
transform 1 0 25760 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_275
timestamp 1606120350
transform 1 0 26404 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0695__A
timestamp 1606120350
transform 1 0 26588 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_279
timestamp 1606120350
transform 1 0 26772 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0503__A
timestamp 1606120350
transform 1 0 26956 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_3_0_clk
timestamp 1606120350
transform 1 0 27140 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_55_286
timestamp 1606120350
transform 1 0 27416 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_3_0_clk_A
timestamp 1606120350
transform 1 0 27600 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_290
timestamp 1606120350
transform 1 0 27784 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_294
timestamp 1606120350
transform 1 0 28152 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_7_0_clk_A
timestamp 1606120350
transform 1 0 28244 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_646
timestamp 1606120350
transform 1 0 29164 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_7_0_clk
timestamp 1606120350
transform 1 0 28428 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__D
timestamp 1606120350
transform 1 0 28888 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1121__CLK
timestamp 1606120350
transform 1 0 29440 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_55_300
timestamp 1606120350
transform 1 0 28704 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_304
timestamp 1606120350
transform 1 0 29072 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_306
timestamp 1606120350
transform 1 0 29256 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_310
timestamp 1606120350
transform 1 0 29624 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_322
timestamp 1606120350
transform 1 0 30728 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_334
timestamp 1606120350
transform 1 0 31832 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_346
timestamp 1606120350
transform 1 0 32936 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_358
timestamp 1606120350
transform 1 0 34040 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_647
timestamp 1606120350
transform 1 0 34776 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_367
timestamp 1606120350
transform 1 0 34868 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_379
timestamp 1606120350
transform 1 0 35972 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1606120350
transform -1 0 38824 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_391
timestamp 1606120350
transform 1 0 37076 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_403
timestamp 1606120350
transform 1 0 38180 0 1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1606120350
transform 1 0 1104 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1606120350
transform 1 0 1380 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1606120350
transform 1 0 2484 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_648
timestamp 1606120350
transform 1 0 3956 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_27
timestamp 1606120350
transform 1 0 3588 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_32
timestamp 1606120350
transform 1 0 4048 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_44
timestamp 1606120350
transform 1 0 5152 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_56
timestamp 1606120350
transform 1 0 6256 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_68
timestamp 1606120350
transform 1 0 7360 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0668_
timestamp 1606120350
transform 1 0 8556 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__B1
timestamp 1606120350
transform 1 0 9384 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0655__A
timestamp 1606120350
transform 1 0 9016 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__A3
timestamp 1606120350
transform 1 0 8372 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__A2
timestamp 1606120350
transform 1 0 8004 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_74
timestamp 1606120350
transform 1 0 7912 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_77
timestamp 1606120350
transform 1 0 8188 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_84
timestamp 1606120350
transform 1 0 8832 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_88
timestamp 1606120350
transform 1 0 9200 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1123_
timestamp 1606120350
transform 1 0 9660 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_649
timestamp 1606120350
transform 1 0 9568 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__C
timestamp 1606120350
transform 1 0 11592 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_112
timestamp 1606120350
transform 1 0 11408 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0491_
timestamp 1606120350
transform 1 0 12144 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_4  _0657_
timestamp 1606120350
transform 1 0 13156 0 -1 33184
box -38 -48 1326 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0657__B1
timestamp 1606120350
transform 1 0 12972 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0772__A2
timestamp 1606120350
transform 1 0 12604 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__B
timestamp 1606120350
transform 1 0 11960 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_116
timestamp 1606120350
transform 1 0 11776 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_123
timestamp 1606120350
transform 1 0 12420 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_127
timestamp 1606120350
transform 1 0 12788 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0512_
timestamp 1606120350
transform 1 0 15272 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_650
timestamp 1606120350
transform 1 0 15180 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__A2
timestamp 1606120350
transform 1 0 14628 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0677__B
timestamp 1606120350
transform 1 0 14996 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_145
timestamp 1606120350
transform 1 0 14444 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_149
timestamp 1606120350
transform 1 0 14812 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_157
timestamp 1606120350
transform 1 0 15548 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _0681_
timestamp 1606120350
transform 1 0 16376 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0683__A
timestamp 1606120350
transform 1 0 15916 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__A
timestamp 1606120350
transform 1 0 17572 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_56_163
timestamp 1606120350
transform 1 0 16100 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_175
timestamp 1606120350
transform 1 0 17204 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_56_181
timestamp 1606120350
transform 1 0 17756 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0513_
timestamp 1606120350
transform 1 0 19504 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _0744_
timestamp 1606120350
transform 1 0 17940 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0590__A3
timestamp 1606120350
transform 1 0 18952 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__C
timestamp 1606120350
transform 1 0 19320 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__D
timestamp 1606120350
transform 1 0 19964 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_192
timestamp 1606120350
transform 1 0 18768 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_196
timestamp 1606120350
transform 1 0 19136 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_203
timestamp 1606120350
transform 1 0 19780 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0583_
timestamp 1606120350
transform 1 0 20884 0 -1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_651
timestamp 1606120350
transform 1 0 20792 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__A
timestamp 1606120350
transform 1 0 21896 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__C
timestamp 1606120350
transform 1 0 20608 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_207
timestamp 1606120350
transform 1 0 20148 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_211
timestamp 1606120350
transform 1 0 20516 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_56_224
timestamp 1606120350
transform 1 0 21712 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_228
timestamp 1606120350
transform 1 0 22080 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0628_
timestamp 1606120350
transform 1 0 22448 0 -1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__dfxtp_4  _1151_
timestamp 1606120350
transform 1 0 23920 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0595__B
timestamp 1606120350
transform 1 0 22264 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__B
timestamp 1606120350
transform 1 0 23276 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__B
timestamp 1606120350
transform 1 0 23644 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_239
timestamp 1606120350
transform 1 0 23092 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_243
timestamp 1606120350
transform 1 0 23460 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_56_247
timestamp 1606120350
transform 1 0 23828 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0583__D
timestamp 1606120350
transform 1 0 25852 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0504__A
timestamp 1606120350
transform 1 0 26220 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_267
timestamp 1606120350
transform 1 0 25668 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_271
timestamp 1606120350
transform 1 0 26036 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_652
timestamp 1606120350
transform 1 0 26404 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1099__CLK
timestamp 1606120350
transform 1 0 26680 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1160__CLK
timestamp 1606120350
transform 1 0 27048 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_276
timestamp 1606120350
transform 1 0 26496 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_56_280
timestamp 1606120350
transform 1 0 26864 0 -1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_284
timestamp 1606120350
transform 1 0 27232 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_296
timestamp 1606120350
transform 1 0 28336 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1121_
timestamp 1606120350
transform 1 0 28612 0 -1 33184
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_56_318
timestamp 1606120350
transform 1 0 30360 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_653
timestamp 1606120350
transform 1 0 32016 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_330
timestamp 1606120350
transform 1 0 31464 0 -1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_56_337
timestamp 1606120350
transform 1 0 32108 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_349
timestamp 1606120350
transform 1 0 33212 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_361
timestamp 1606120350
transform 1 0 34316 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_373
timestamp 1606120350
transform 1 0 35420 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_385
timestamp 1606120350
transform 1 0 36524 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1606120350
transform -1 0 38824 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_654
timestamp 1606120350
transform 1 0 37628 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_398
timestamp 1606120350
transform 1 0 37720 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_406
timestamp 1606120350
transform 1 0 38456 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1606120350
transform 1 0 1104 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1606120350
transform 1 0 1380 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1606120350
transform 1 0 2484 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1606120350
transform 1 0 3588 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1606120350
transform 1 0 4692 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_655
timestamp 1606120350
transform 1 0 6716 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_1_0_clk
timestamp 1606120350
transform 1 0 6440 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_1_0_clk_A
timestamp 1606120350
transform 1 0 6992 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_51
timestamp 1606120350
transform 1 0 5796 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_57
timestamp 1606120350
transform 1 0 6348 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_62
timestamp 1606120350
transform 1 0 6808 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_57_66
timestamp 1606120350
transform 1 0 7176 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_57_71
timestamp 1606120350
transform 1 0 7636 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_3_0_clk_A
timestamp 1606120350
transform 1 0 7452 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_75
timestamp 1606120350
transform 1 0 8004 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__D
timestamp 1606120350
transform 1 0 7820 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_79
timestamp 1606120350
transform 1 0 8372 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__A
timestamp 1606120350
transform 1 0 8188 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_83
timestamp 1606120350
transform 1 0 8740 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__A1
timestamp 1606120350
transform 1 0 8556 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_87
timestamp 1606120350
transform 1 0 9108 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__A2
timestamp 1606120350
transform 1 0 8924 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__A1
timestamp 1606120350
transform 1 0 9292 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0750_
timestamp 1606120350
transform 1 0 9476 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _0773_
timestamp 1606120350
transform 1 0 10488 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0750__A
timestamp 1606120350
transform 1 0 9936 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__B1
timestamp 1606120350
transform 1 0 10304 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_94
timestamp 1606120350
transform 1 0 9752 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_98
timestamp 1606120350
transform 1 0 10120 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_114
timestamp 1606120350
transform 1 0 11592 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _0774_
timestamp 1606120350
transform 1 0 12420 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_656
timestamp 1606120350
transform 1 0 12328 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__A2
timestamp 1606120350
transform 1 0 12144 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__A1
timestamp 1606120350
transform 1 0 13708 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__C
timestamp 1606120350
transform 1 0 11776 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_118
timestamp 1606120350
transform 1 0 11960 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_135
timestamp 1606120350
transform 1 0 13524 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _0735_
timestamp 1606120350
transform 1 0 14260 0 1 33184
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__A1
timestamp 1606120350
transform 1 0 14076 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_139
timestamp 1606120350
transform 1 0 13892 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0771_
timestamp 1606120350
transform 1 0 16560 0 1 33184
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__B
timestamp 1606120350
transform 1 0 17756 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__B
timestamp 1606120350
transform 1 0 17388 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__B
timestamp 1606120350
transform 1 0 16008 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__A
timestamp 1606120350
transform 1 0 16376 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_160
timestamp 1606120350
transform 1 0 15824 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_164
timestamp 1606120350
transform 1 0 16192 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_175
timestamp 1606120350
transform 1 0 17204 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_179
timestamp 1606120350
transform 1 0 17572 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0616_
timestamp 1606120350
transform 1 0 19596 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _0739_
timestamp 1606120350
transform 1 0 18032 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_657
timestamp 1606120350
transform 1 0 17940 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__B
timestamp 1606120350
transform 1 0 19412 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__A
timestamp 1606120350
transform 1 0 19044 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_193
timestamp 1606120350
transform 1 0 18860 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_197
timestamp 1606120350
transform 1 0 19228 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0579_
timestamp 1606120350
transform 1 0 21160 0 1 33184
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0505__A
timestamp 1606120350
transform 1 0 20884 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_210
timestamp 1606120350
transform 1 0 20424 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_214
timestamp 1606120350
transform 1 0 20792 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_217
timestamp 1606120350
transform 1 0 21068 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_227
timestamp 1606120350
transform 1 0 21988 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0802_
timestamp 1606120350
transform 1 0 23644 0 1 33184
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_658
timestamp 1606120350
transform 1 0 23552 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_6_0_clk
timestamp 1606120350
transform 1 0 23276 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__D
timestamp 1606120350
transform 1 0 22724 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0505__B
timestamp 1606120350
transform 1 0 22172 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__D
timestamp 1606120350
transform 1 0 23092 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_231
timestamp 1606120350
transform 1 0 22356 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_57_237
timestamp 1606120350
transform 1 0 22908 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__A1
timestamp 1606120350
transform 1 0 25116 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__D
timestamp 1606120350
transform 1 0 25484 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__A
timestamp 1606120350
transform 1 0 25852 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__CLK
timestamp 1606120350
transform 1 0 26220 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_259
timestamp 1606120350
transform 1 0 24932 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_263
timestamp 1606120350
transform 1 0 25300 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_267
timestamp 1606120350
transform 1 0 25668 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_271
timestamp 1606120350
transform 1 0 26036 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__D
timestamp 1606120350
transform 1 0 27324 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1223__CLK
timestamp 1606120350
transform 1 0 27692 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_57_275
timestamp 1606120350
transform 1 0 26404 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_283
timestamp 1606120350
transform 1 0 27140 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_57_287
timestamp 1606120350
transform 1 0 27508 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_291
timestamp 1606120350
transform 1 0 27876 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_659
timestamp 1606120350
transform 1 0 29164 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_303
timestamp 1606120350
transform 1 0 28980 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_306
timestamp 1606120350
transform 1 0 29256 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_318
timestamp 1606120350
transform 1 0 30360 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__D
timestamp 1606120350
transform 1 0 32108 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1118__CLK
timestamp 1606120350
transform 1 0 32476 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_330
timestamp 1606120350
transform 1 0 31464 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_336
timestamp 1606120350
transform 1 0 32016 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_339
timestamp 1606120350
transform 1 0 32292 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_343
timestamp 1606120350
transform 1 0 32660 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_355
timestamp 1606120350
transform 1 0 33764 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_363
timestamp 1606120350
transform 1 0 34500 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_660
timestamp 1606120350
transform 1 0 34776 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_367
timestamp 1606120350
transform 1 0 34868 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_379
timestamp 1606120350
transform 1 0 35972 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1606120350
transform -1 0 38824 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_391
timestamp 1606120350
transform 1 0 37076 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_403
timestamp 1606120350
transform 1 0 38180 0 1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1606120350
transform 1 0 1104 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__D
timestamp 1606120350
transform 1 0 1656 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_3
timestamp 1606120350
transform 1 0 1380 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_8
timestamp 1606120350
transform 1 0 1840 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_20
timestamp 1606120350
transform 1 0 2944 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_661
timestamp 1606120350
transform 1 0 3956 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_28
timestamp 1606120350
transform 1 0 3680 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_32
timestamp 1606120350
transform 1 0 4048 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_44
timestamp 1606120350
transform 1 0 5152 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_56
timestamp 1606120350
transform 1 0 6256 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_68
timestamp 1606120350
transform 1 0 7360 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_3_0_clk
timestamp 1606120350
transform 1 0 8648 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__B2
timestamp 1606120350
transform 1 0 9384 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__A1
timestamp 1606120350
transform 1 0 8464 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0502__A
timestamp 1606120350
transform 1 0 8096 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_78
timestamp 1606120350
transform 1 0 8280 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_85
timestamp 1606120350
transform 1 0 8924 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_89
timestamp 1606120350
transform 1 0 9292 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0502_
timestamp 1606120350
transform 1 0 10764 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_662
timestamp 1606120350
transform 1 0 9568 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0774__B1
timestamp 1606120350
transform 1 0 10580 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0773__B1
timestamp 1606120350
transform 1 0 10212 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0775__A2
timestamp 1606120350
transform 1 0 9844 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_93
timestamp 1606120350
transform 1 0 9660 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_97
timestamp 1606120350
transform 1 0 10028 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_101
timestamp 1606120350
transform 1 0 10396 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_114
timestamp 1606120350
transform 1 0 11592 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0775_
timestamp 1606120350
transform 1 0 12328 0 -1 34272
box -38 -48 1326 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__A3
timestamp 1606120350
transform 1 0 12144 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__A3
timestamp 1606120350
transform 1 0 11776 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_118
timestamp 1606120350
transform 1 0 11960 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_136
timestamp 1606120350
transform 1 0 13616 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_140
timestamp 1606120350
transform 1 0 13984 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__A1
timestamp 1606120350
transform 1 0 13800 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0735__B2
timestamp 1606120350
transform 1 0 14260 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_145
timestamp 1606120350
transform 1 0 14444 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__B2
timestamp 1606120350
transform 1 0 14628 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_149
timestamp 1606120350
transform 1 0 14812 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__A1
timestamp 1606120350
transform 1 0 14996 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_154
timestamp 1606120350
transform 1 0 15272 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0740__A
timestamp 1606120350
transform 1 0 15456 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_663
timestamp 1606120350
transform 1 0 15180 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_58_158
timestamp 1606120350
transform 1 0 15640 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0722_
timestamp 1606120350
transform 1 0 17572 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _0740_
timestamp 1606120350
transform 1 0 16008 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0544__A
timestamp 1606120350
transform 1 0 17296 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__D
timestamp 1606120350
transform 1 0 15824 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_171
timestamp 1606120350
transform 1 0 16836 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_175
timestamp 1606120350
transform 1 0 17204 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_58_178
timestamp 1606120350
transform 1 0 17480 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _0580_
timestamp 1606120350
transform 1 0 19228 0 -1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__A
timestamp 1606120350
transform 1 0 19044 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__B
timestamp 1606120350
transform 1 0 18676 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_58_188
timestamp 1606120350
transform 1 0 18400 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_58_193
timestamp 1606120350
transform 1 0 18860 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_210
timestamp 1606120350
transform 1 0 20424 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_206
timestamp 1606120350
transform 1 0 20056 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__D
timestamp 1606120350
transform 1 0 20608 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0684__C
timestamp 1606120350
transform 1 0 20240 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_664
timestamp 1606120350
transform 1 0 20792 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0505_
timestamp 1606120350
transform 1 0 20884 0 -1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_58_226
timestamp 1606120350
transform 1 0 21896 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_222
timestamp 1606120350
transform 1 0 21528 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0727__C
timestamp 1606120350
transform 1 0 22080 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0579__B
timestamp 1606120350
transform 1 0 21712 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1180_
timestamp 1606120350
transform 1 0 22724 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0744__A
timestamp 1606120350
transform 1 0 22448 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_230
timestamp 1606120350
transform 1 0 22264 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_234
timestamp 1606120350
transform 1 0 22632 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__A2
timestamp 1606120350
transform 1 0 24656 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0616__C
timestamp 1606120350
transform 1 0 25024 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_6_0_clk_A
timestamp 1606120350
transform 1 0 25392 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__CLK
timestamp 1606120350
transform 1 0 26220 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_254
timestamp 1606120350
transform 1 0 24472 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_258
timestamp 1606120350
transform 1 0 24840 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_262
timestamp 1606120350
transform 1 0 25208 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_58_266
timestamp 1606120350
transform 1 0 25576 0 -1 34272
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_272
timestamp 1606120350
transform 1 0 26128 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1223_
timestamp 1606120350
transform 1 0 27324 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_665
timestamp 1606120350
transform 1 0 26404 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_276
timestamp 1606120350
transform 1 0 26496 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_284
timestamp 1606120350
transform 1 0 27232 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__CLK
timestamp 1606120350
transform 1 0 29256 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_58_304
timestamp 1606120350
transform 1 0 29072 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_58_308
timestamp 1606120350
transform 1 0 29440 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1118_
timestamp 1606120350
transform 1 0 32108 0 -1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_666
timestamp 1606120350
transform 1 0 32016 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_320
timestamp 1606120350
transform 1 0 30544 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_332
timestamp 1606120350
transform 1 0 31648 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_356
timestamp 1606120350
transform 1 0 33856 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_368
timestamp 1606120350
transform 1 0 34960 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_380
timestamp 1606120350
transform 1 0 36064 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1606120350
transform -1 0 38824 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_667
timestamp 1606120350
transform 1 0 37628 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_392
timestamp 1606120350
transform 1 0 37168 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_396
timestamp 1606120350
transform 1 0 37536 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_398
timestamp 1606120350
transform 1 0 37720 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_406
timestamp 1606120350
transform 1 0 38456 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1205_
timestamp 1606120350
transform 1 0 1656 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1606120350
transform 1 0 1104 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1606120350
transform 1 0 1104 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1205__CLK
timestamp 1606120350
transform 1 0 1656 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_3
timestamp 1606120350
transform 1 0 1380 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_60_3
timestamp 1606120350
transform 1 0 1380 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_8
timestamp 1606120350
transform 1 0 1840 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_20
timestamp 1606120350
transform 1 0 2944 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_674
timestamp 1606120350
transform 1 0 3956 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_25
timestamp 1606120350
transform 1 0 3404 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_37
timestamp 1606120350
transform 1 0 4508 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_28
timestamp 1606120350
transform 1 0 3680 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_32
timestamp 1606120350
transform 1 0 4048 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_44
timestamp 1606120350
transform 1 0 5152 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_668
timestamp 1606120350
transform 1 0 6716 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_49
timestamp 1606120350
transform 1 0 5612 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_62
timestamp 1606120350
transform 1 0 6808 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_56
timestamp 1606120350
transform 1 0 6256 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_68
timestamp 1606120350
transform 1 0 7360 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1122_
timestamp 1606120350
transform 1 0 9384 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__D
timestamp 1606120350
transform 1 0 9200 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__A2
timestamp 1606120350
transform 1 0 8832 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1122__CLK
timestamp 1606120350
transform 1 0 9384 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_74
timestamp 1606120350
transform 1 0 7912 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_82
timestamp 1606120350
transform 1 0 8648 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_86
timestamp 1606120350
transform 1 0 9016 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_60_80
timestamp 1606120350
transform 1 0 8464 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_88
timestamp 1606120350
transform 1 0 9200 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_93
timestamp 1606120350
transform 1 0 9660 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_675
timestamp 1606120350
transform 1 0 9568 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_60_100
timestamp 1606120350
transform 1 0 10304 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_60_97
timestamp 1606120350
transform 1 0 10028 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__B
timestamp 1606120350
transform 1 0 10120 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_104
timestamp 1606120350
transform 1 0 10672 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__C1
timestamp 1606120350
transform 1 0 10488 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_108
timestamp 1606120350
transform 1 0 11040 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_109
timestamp 1606120350
transform 1 0 11132 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__D
timestamp 1606120350
transform 1 0 10856 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__B2
timestamp 1606120350
transform 1 0 11224 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_112
timestamp 1606120350
transform 1 0 11408 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_114
timestamp 1606120350
transform 1 0 11592 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__A3
timestamp 1606120350
transform 1 0 11592 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0716__A
timestamp 1606120350
transform 1 0 11408 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_123
timestamp 1606120350
transform 1 0 12420 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_118
timestamp 1606120350
transform 1 0 11960 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0656__A
timestamp 1606120350
transform 1 0 11776 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0656__B
timestamp 1606120350
transform 1 0 12144 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__A1_N
timestamp 1606120350
transform 1 0 12604 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_669
timestamp 1606120350
transform 1 0 12328 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0716_
timestamp 1606120350
transform 1 0 11776 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _0656_
timestamp 1606120350
transform 1 0 12420 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_60_127
timestamp 1606120350
transform 1 0 12788 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_134
timestamp 1606120350
transform 1 0 13432 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_130
timestamp 1606120350
transform 1 0 13064 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0659__B
timestamp 1606120350
transform 1 0 12972 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0736__B1
timestamp 1606120350
transform 1 0 13248 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__B1
timestamp 1606120350
transform 1 0 13616 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _0736_
timestamp 1606120350
transform 1 0 13156 0 -1 35360
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_60_145
timestamp 1606120350
transform 1 0 14444 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0671__A2
timestamp 1606120350
transform 1 0 14628 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_149
timestamp 1606120350
transform 1 0 14812 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_159
timestamp 1606120350
transform 1 0 15732 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_155
timestamp 1606120350
transform 1 0 15364 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__A1
timestamp 1606120350
transform 1 0 14996 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__B1
timestamp 1606120350
transform 1 0 15548 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_676
timestamp 1606120350
transform 1 0 15180 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__a211o_4  _0672_
timestamp 1606120350
transform 1 0 15272 0 -1 35360
box -38 -48 1326 592
use sky130_fd_sc_hd__a32o_4  _0671_
timestamp 1606120350
transform 1 0 13800 0 1 34272
box -38 -48 1602 592
use sky130_fd_sc_hd__fill_2  FILLER_60_168
timestamp 1606120350
transform 1 0 16560 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0771__B
timestamp 1606120350
transform 1 0 15916 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0728_
timestamp 1606120350
transform 1 0 16100 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_60_172
timestamp 1606120350
transform 1 0 16928 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_178
timestamp 1606120350
transform 1 0 17480 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_172
timestamp 1606120350
transform 1 0 16928 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__C1
timestamp 1606120350
transform 1 0 16744 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0544__C
timestamp 1606120350
transform 1 0 17112 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0544__B
timestamp 1606120350
transform 1 0 17296 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0544_
timestamp 1606120350
transform 1 0 17296 0 -1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0507__A
timestamp 1606120350
transform 1 0 17756 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_189
timestamp 1606120350
transform 1 0 18492 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_185
timestamp 1606120350
transform 1 0 18124 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0739__C
timestamp 1606120350
transform 1 0 18676 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__A
timestamp 1606120350
transform 1 0 18308 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_670
timestamp 1606120350
transform 1 0 17940 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0507_
timestamp 1606120350
transform 1 0 18032 0 1 34272
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_60_200
timestamp 1606120350
transform 1 0 19504 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_197
timestamp 1606120350
transform 1 0 19228 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_193
timestamp 1606120350
transform 1 0 18860 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__B
timestamp 1606120350
transform 1 0 19688 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0722__C
timestamp 1606120350
transform 1 0 19412 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__B
timestamp 1606120350
transform 1 0 19044 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0720_
timestamp 1606120350
transform 1 0 18860 0 -1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _0594_
timestamp 1606120350
transform 1 0 19596 0 1 34272
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_60_204
timestamp 1606120350
transform 1 0 19872 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__A
timestamp 1606120350
transform 1 0 20056 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_208
timestamp 1606120350
transform 1 0 20240 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_208
timestamp 1606120350
transform 1 0 20240 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0594__B
timestamp 1606120350
transform 1 0 20424 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__C
timestamp 1606120350
transform 1 0 20424 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_212
timestamp 1606120350
transform 1 0 20608 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_212
timestamp 1606120350
transform 1 0 20608 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0508_
timestamp 1606120350
transform 1 0 20976 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_677
timestamp 1606120350
transform 1 0 20792 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0728__B
timestamp 1606120350
transform 1 0 20792 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_223
timestamp 1606120350
transform 1 0 21620 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_219
timestamp 1606120350
transform 1 0 21252 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0508__A
timestamp 1606120350
transform 1 0 21804 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__B1
timestamp 1606120350
transform 1 0 21436 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0629_
timestamp 1606120350
transform 1 0 21988 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _0803_
timestamp 1606120350
transform 1 0 20884 0 -1 35360
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_60_229
timestamp 1606120350
transform 1 0 22172 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_230
timestamp 1606120350
transform 1 0 22264 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__B2
timestamp 1606120350
transform 1 0 22356 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_233
timestamp 1606120350
transform 1 0 22540 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_234
timestamp 1606120350
transform 1 0 22632 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0629__A
timestamp 1606120350
transform 1 0 22448 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0720__A
timestamp 1606120350
transform 1 0 22724 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__A1
timestamp 1606120350
transform 1 0 22816 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_237
timestamp 1606120350
transform 1 0 22908 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_238
timestamp 1606120350
transform 1 0 23000 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0594__A
timestamp 1606120350
transform 1 0 23092 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_241
timestamp 1606120350
transform 1 0 23276 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_242
timestamp 1606120350
transform 1 0 23368 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0803__A2
timestamp 1606120350
transform 1 0 23184 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_245
timestamp 1606120350
transform 1 0 23644 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_245
timestamp 1606120350
transform 1 0 23644 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0580__D
timestamp 1606120350
transform 1 0 23460 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_671
timestamp 1606120350
transform 1 0 23552 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_0_0_clk_A
timestamp 1606120350
transform 1 0 23828 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__B2
timestamp 1606120350
transform 1 0 23828 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_60_249
timestamp 1606120350
transform 1 0 24012 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_249
timestamp 1606120350
transform 1 0 24012 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1180__CLK
timestamp 1606120350
transform 1 0 24196 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0802__B1
timestamp 1606120350
transform 1 0 24196 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1196_
timestamp 1606120350
transform 1 0 26220 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1196__D
timestamp 1606120350
transform 1 0 26036 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1151__D
timestamp 1606120350
transform 1 0 24564 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_253
timestamp 1606120350
transform 1 0 24380 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_257
timestamp 1606120350
transform 1 0 24748 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_269
timestamp 1606120350
transform 1 0 25852 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_253
timestamp 1606120350
transform 1 0 24380 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_265
timestamp 1606120350
transform 1 0 25484 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_273
timestamp 1606120350
transform 1 0 26220 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_678
timestamp 1606120350
transform 1 0 26404 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_292
timestamp 1606120350
transform 1 0 27968 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_276
timestamp 1606120350
transform 1 0 26496 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_288
timestamp 1606120350
transform 1 0 27600 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1130_
timestamp 1606120350
transform 1 0 29256 0 1 34272
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_672
timestamp 1606120350
transform 1 0 29164 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1130__D
timestamp 1606120350
transform 1 0 28980 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_59_300
timestamp 1606120350
transform 1 0 28704 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_300
timestamp 1606120350
transform 1 0 28704 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_312
timestamp 1606120350
transform 1 0 29808 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_679
timestamp 1606120350
transform 1 0 32016 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_325
timestamp 1606120350
transform 1 0 31004 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_337
timestamp 1606120350
transform 1 0 32108 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_324
timestamp 1606120350
transform 1 0 30912 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_337
timestamp 1606120350
transform 1 0 32108 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_349
timestamp 1606120350
transform 1 0 33212 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_361
timestamp 1606120350
transform 1 0 34316 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_365
timestamp 1606120350
transform 1 0 34684 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_349
timestamp 1606120350
transform 1 0 33212 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_361
timestamp 1606120350
transform 1 0 34316 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_673
timestamp 1606120350
transform 1 0 34776 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_367
timestamp 1606120350
transform 1 0 34868 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_379
timestamp 1606120350
transform 1 0 35972 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_373
timestamp 1606120350
transform 1 0 35420 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_385
timestamp 1606120350
transform 1 0 36524 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1606120350
transform -1 0 38824 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1606120350
transform -1 0 38824 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_680
timestamp 1606120350
transform 1 0 37628 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_391
timestamp 1606120350
transform 1 0 37076 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_403
timestamp 1606120350
transform 1 0 38180 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_398
timestamp 1606120350
transform 1 0 37720 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_406
timestamp 1606120350
transform 1 0 38456 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1606120350
transform 1 0 1104 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1606120350
transform 1 0 1380 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1606120350
transform 1 0 2484 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1606120350
transform 1 0 3588 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1606120350
transform 1 0 4692 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_681
timestamp 1606120350
transform 1 0 6716 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_51
timestamp 1606120350
transform 1 0 5796 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_59
timestamp 1606120350
transform 1 0 6532 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_62
timestamp 1606120350
transform 1 0 6808 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_74
timestamp 1606120350
transform 1 0 7912 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_86
timestamp 1606120350
transform 1 0 9016 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_94
timestamp 1606120350
transform 1 0 9752 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0672__A2
timestamp 1606120350
transform 1 0 9936 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_98
timestamp 1606120350
transform 1 0 10120 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__B1
timestamp 1606120350
transform 1 0 10304 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_102
timestamp 1606120350
transform 1 0 10488 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__A2
timestamp 1606120350
transform 1 0 10672 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_110
timestamp 1606120350
transform 1 0 11224 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_61_106
timestamp 1606120350
transform 1 0 10856 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0496__A
timestamp 1606120350
transform 1 0 11040 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_114
timestamp 1606120350
transform 1 0 11592 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_121
timestamp 1606120350
transform 1 0 12236 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_117
timestamp 1606120350
transform 1 0 11868 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__A2_N
timestamp 1606120350
transform 1 0 11684 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__B2
timestamp 1606120350
transform 1 0 12052 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_682
timestamp 1606120350
transform 1 0 12328 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_123
timestamp 1606120350
transform 1 0 12420 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0659_
timestamp 1606120350
transform 1 0 12512 0 1 35360
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_61_135
timestamp 1606120350
transform 1 0 13524 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_131
timestamp 1606120350
transform 1 0 13156 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0659__A
timestamp 1606120350
transform 1 0 13340 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__B1
timestamp 1606120350
transform 1 0 13708 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _0712_
timestamp 1606120350
transform 1 0 13892 0 1 35360
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__A
timestamp 1606120350
transform 1 0 15640 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_156
timestamp 1606120350
transform 1 0 15456 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0718_
timestamp 1606120350
transform 1 0 16192 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__C
timestamp 1606120350
transform 1 0 16008 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0544__D
timestamp 1606120350
transform 1 0 17296 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__A
timestamp 1606120350
transform 1 0 17664 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_160
timestamp 1606120350
transform 1 0 15824 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_173
timestamp 1606120350
transform 1 0 17020 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_178
timestamp 1606120350
transform 1 0 17480 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_61_182
timestamp 1606120350
transform 1 0 17848 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0506_
timestamp 1606120350
transform 1 0 19596 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _0729_
timestamp 1606120350
transform 1 0 18032 0 1 35360
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_683
timestamp 1606120350
transform 1 0 17940 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__B
timestamp 1606120350
transform 1 0 19136 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_193
timestamp 1606120350
transform 1 0 18860 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_61_198
timestamp 1606120350
transform 1 0 19320 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_204
timestamp 1606120350
transform 1 0 19872 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1100_
timestamp 1606120350
transform 1 0 20884 0 1 35360
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0506__A
timestamp 1606120350
transform 1 0 20056 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0718__D
timestamp 1606120350
transform 1 0 20424 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_208
timestamp 1606120350
transform 1 0 20240 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_61_212
timestamp 1606120350
transform 1 0 20608 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_684
timestamp 1606120350
transform 1 0 23552 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__D
timestamp 1606120350
transform 1 0 23092 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1179__CLK
timestamp 1606120350
transform 1 0 23828 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_234
timestamp 1606120350
transform 1 0 22632 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_238
timestamp 1606120350
transform 1 0 23000 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_61_241
timestamp 1606120350
transform 1 0 23276 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_61_245
timestamp 1606120350
transform 1 0 23644 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_249
timestamp 1606120350
transform 1 0 24012 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_261
timestamp 1606120350
transform 1 0 25116 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_273
timestamp 1606120350
transform 1 0 26220 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1168__D
timestamp 1606120350
transform 1 0 28152 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_285
timestamp 1606120350
transform 1 0 27324 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_293
timestamp 1606120350
transform 1 0 28060 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_296
timestamp 1606120350
transform 1 0 28336 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_685
timestamp 1606120350
transform 1 0 29164 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1168__CLK
timestamp 1606120350
transform 1 0 28520 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_300
timestamp 1606120350
transform 1 0 28704 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_304
timestamp 1606120350
transform 1 0 29072 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_306
timestamp 1606120350
transform 1 0 29256 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_318
timestamp 1606120350
transform 1 0 30360 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_330
timestamp 1606120350
transform 1 0 31464 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_342
timestamp 1606120350
transform 1 0 32568 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_354
timestamp 1606120350
transform 1 0 33672 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_686
timestamp 1606120350
transform 1 0 34776 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_367
timestamp 1606120350
transform 1 0 34868 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_379
timestamp 1606120350
transform 1 0 35972 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1606120350
transform -1 0 38824 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_391
timestamp 1606120350
transform 1 0 37076 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_403
timestamp 1606120350
transform 1 0 38180 0 1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1606120350
transform 1 0 1104 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1606120350
transform 1 0 1380 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1606120350
transform 1 0 2484 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_687
timestamp 1606120350
transform 1 0 3956 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_27
timestamp 1606120350
transform 1 0 3588 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_32
timestamp 1606120350
transform 1 0 4048 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_44
timestamp 1606120350
transform 1 0 5152 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_56
timestamp 1606120350
transform 1 0 6256 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_68
timestamp 1606120350
transform 1 0 7360 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_80
timestamp 1606120350
transform 1 0 8464 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0496_
timestamp 1606120350
transform 1 0 11040 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_688
timestamp 1606120350
transform 1 0 9568 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__A2
timestamp 1606120350
transform 1 0 11500 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__A3
timestamp 1606120350
transform 1 0 10856 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_62_93
timestamp 1606120350
transform 1 0 9660 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_105
timestamp 1606120350
transform 1 0 10764 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_62_111
timestamp 1606120350
transform 1 0 11316 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _0778_
timestamp 1606120350
transform 1 0 12052 0 -1 36448
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0778__B1
timestamp 1606120350
transform 1 0 11868 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_115
timestamp 1606120350
transform 1 0 11684 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_135
timestamp 1606120350
transform 1 0 13524 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_4  _0731_
timestamp 1606120350
transform 1 0 15272 0 -1 36448
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_689
timestamp 1606120350
transform 1 0 15180 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__A1
timestamp 1606120350
transform 1 0 14444 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__A1
timestamp 1606120350
transform 1 0 13892 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__A1
timestamp 1606120350
transform 1 0 14812 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_141
timestamp 1606120350
transform 1 0 14076 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_62_147
timestamp 1606120350
transform 1 0 14628 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_151
timestamp 1606120350
transform 1 0 14996 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0745_
timestamp 1606120350
transform 1 0 17572 0 -1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0681__C
timestamp 1606120350
transform 1 0 17020 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__A2
timestamp 1606120350
transform 1 0 17388 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_171
timestamp 1606120350
transform 1 0 16836 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_175
timestamp 1606120350
transform 1 0 17204 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0737_
timestamp 1606120350
transform 1 0 19136 0 -1 36448
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0648__B1
timestamp 1606120350
transform 1 0 18584 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__A1
timestamp 1606120350
transform 1 0 18952 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__B
timestamp 1606120350
transform 1 0 19964 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_188
timestamp 1606120350
transform 1 0 18400 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_192
timestamp 1606120350
transform 1 0 18768 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_203
timestamp 1606120350
transform 1 0 19780 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_207
timestamp 1606120350
transform 1 0 20148 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0729__C
timestamp 1606120350
transform 1 0 20332 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_62_211
timestamp 1606120350
transform 1 0 20516 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_690
timestamp 1606120350
transform 1 0 20792 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0487_
timestamp 1606120350
transform 1 0 20884 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_62_218
timestamp 1606120350
transform 1 0 21160 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__B
timestamp 1606120350
transform 1 0 21344 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_222
timestamp 1606120350
transform 1 0 21528 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0737__A
timestamp 1606120350
transform 1 0 21712 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_226
timestamp 1606120350
transform 1 0 21896 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0487__A
timestamp 1606120350
transform 1 0 22080 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1179_
timestamp 1606120350
transform 1 0 23092 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__CLK
timestamp 1606120350
transform 1 0 22448 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_62_230
timestamp 1606120350
transform 1 0 22264 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_234
timestamp 1606120350
transform 1 0 22632 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_238
timestamp 1606120350
transform 1 0 23000 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__CLK
timestamp 1606120350
transform 1 0 25392 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_62_258
timestamp 1606120350
transform 1 0 24840 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_62_266
timestamp 1606120350
transform 1 0 25576 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_274
timestamp 1606120350
transform 1 0 26312 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1168_
timestamp 1606120350
transform 1 0 28152 0 -1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_691
timestamp 1606120350
transform 1 0 26404 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_276
timestamp 1606120350
transform 1 0 26496 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_288
timestamp 1606120350
transform 1 0 27600 0 -1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_62_313
timestamp 1606120350
transform 1 0 29900 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_692
timestamp 1606120350
transform 1 0 32016 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_325
timestamp 1606120350
transform 1 0 31004 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_333
timestamp 1606120350
transform 1 0 31740 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_337
timestamp 1606120350
transform 1 0 32108 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_349
timestamp 1606120350
transform 1 0 33212 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_361
timestamp 1606120350
transform 1 0 34316 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_373
timestamp 1606120350
transform 1 0 35420 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_385
timestamp 1606120350
transform 1 0 36524 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1606120350
transform -1 0 38824 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_693
timestamp 1606120350
transform 1 0 37628 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_398
timestamp 1606120350
transform 1 0 37720 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_406
timestamp 1606120350
transform 1 0 38456 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1606120350
transform 1 0 1104 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1606120350
transform 1 0 1380 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1606120350
transform 1 0 2484 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1606120350
transform 1 0 3588 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1606120350
transform 1 0 4692 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_694
timestamp 1606120350
transform 1 0 6716 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_51
timestamp 1606120350
transform 1 0 5796 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_59
timestamp 1606120350
transform 1 0 6532 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_62
timestamp 1606120350
transform 1 0 6808 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_74
timestamp 1606120350
transform 1 0 7912 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_86
timestamp 1606120350
transform 1 0 9016 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  _0673_
timestamp 1606120350
transform 1 0 10764 0 1 36448
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0710__B1
timestamp 1606120350
transform 1 0 10580 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0673__A
timestamp 1606120350
transform 1 0 10212 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__D
timestamp 1606120350
transform 1 0 9844 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_94
timestamp 1606120350
transform 1 0 9752 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_97
timestamp 1606120350
transform 1 0 10028 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_101
timestamp 1606120350
transform 1 0 10396 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_114
timestamp 1606120350
transform 1 0 11592 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__a21bo_4  _0660_
timestamp 1606120350
transform 1 0 12512 0 1 36448
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_695
timestamp 1606120350
transform 1 0 12328 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__A1
timestamp 1606120350
transform 1 0 12144 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__B1_N
timestamp 1606120350
transform 1 0 11776 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_118
timestamp 1606120350
transform 1 0 11960 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_123
timestamp 1606120350
transform 1 0 12420 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_137
timestamp 1606120350
transform 1 0 13708 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _0747_
timestamp 1606120350
transform 1 0 14444 0 1 36448
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__B2
timestamp 1606120350
transform 1 0 14260 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0712__A2
timestamp 1606120350
transform 1 0 13892 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_141
timestamp 1606120350
transform 1 0 14076 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_162
timestamp 1606120350
transform 1 0 16008 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_166
timestamp 1606120350
transform 1 0 16376 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0709__A
timestamp 1606120350
transform 1 0 16192 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_170
timestamp 1606120350
transform 1 0 16744 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__A2
timestamp 1606120350
transform 1 0 16560 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_175
timestamp 1606120350
transform 1 0 17204 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0550_
timestamp 1606120350
transform 1 0 16928 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_179
timestamp 1606120350
transform 1 0 17572 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0550__A
timestamp 1606120350
transform 1 0 17388 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0648__A1
timestamp 1606120350
transform 1 0 17756 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_4  _0648_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 18032 0 1 36448
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_696
timestamp 1606120350
transform 1 0 17940 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__A2
timestamp 1606120350
transform 1 0 19412 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0648__A2
timestamp 1606120350
transform 1 0 19780 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_197
timestamp 1606120350
transform 1 0 19228 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_201
timestamp 1606120350
transform 1 0 19596 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_205
timestamp 1606120350
transform 1 0 19964 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_213
timestamp 1606120350
transform 1 0 20700 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_209
timestamp 1606120350
transform 1 0 20332 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0745__C
timestamp 1606120350
transform 1 0 20884 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__B1
timestamp 1606120350
transform 1 0 20516 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0708__B1
timestamp 1606120350
transform 1 0 20148 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_221
timestamp 1606120350
transform 1 0 21436 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_217
timestamp 1606120350
transform 1 0 21068 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__A1
timestamp 1606120350
transform 1 0 21620 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1100__D
timestamp 1606120350
transform 1 0 21252 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_225
timestamp 1606120350
transform 1 0 21804 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_697
timestamp 1606120350
transform 1 0 23552 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__D
timestamp 1606120350
transform 1 0 23092 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1132__CLK
timestamp 1606120350
transform 1 0 23828 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_237
timestamp 1606120350
transform 1 0 22908 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_63_241
timestamp 1606120350
transform 1 0 23276 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_245
timestamp 1606120350
transform 1 0 23644 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_249
timestamp 1606120350
transform 1 0 24012 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1116_
timestamp 1606120350
transform 1 0 25392 0 1 36448
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1116__D
timestamp 1606120350
transform 1 0 25208 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_63_261
timestamp 1606120350
transform 1 0 25116 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0830__A
timestamp 1606120350
transform 1 0 27324 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_63_283
timestamp 1606120350
transform 1 0 27140 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_287
timestamp 1606120350
transform 1 0 27508 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_698
timestamp 1606120350
transform 1 0 29164 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_299
timestamp 1606120350
transform 1 0 28612 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_306
timestamp 1606120350
transform 1 0 29256 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_318
timestamp 1606120350
transform 1 0 30360 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__D
timestamp 1606120350
transform 1 0 32108 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1201__CLK
timestamp 1606120350
transform 1 0 32476 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_330
timestamp 1606120350
transform 1 0 31464 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_336
timestamp 1606120350
transform 1 0 32016 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_339
timestamp 1606120350
transform 1 0 32292 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_343
timestamp 1606120350
transform 1 0 32660 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_355
timestamp 1606120350
transform 1 0 33764 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_363
timestamp 1606120350
transform 1 0 34500 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_699
timestamp 1606120350
transform 1 0 34776 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_367
timestamp 1606120350
transform 1 0 34868 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_379
timestamp 1606120350
transform 1 0 35972 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1606120350
transform -1 0 38824 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_391
timestamp 1606120350
transform 1 0 37076 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_403
timestamp 1606120350
transform 1 0 38180 0 1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1606120350
transform 1 0 1104 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1606120350
transform 1 0 1380 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1606120350
transform 1 0 2484 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_700
timestamp 1606120350
transform 1 0 3956 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_27
timestamp 1606120350
transform 1 0 3588 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_32
timestamp 1606120350
transform 1 0 4048 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_44
timestamp 1606120350
transform 1 0 5152 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_56
timestamp 1606120350
transform 1 0 6256 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_68
timestamp 1606120350
transform 1 0 7360 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_80
timestamp 1606120350
transform 1 0 8464 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1091_
timestamp 1606120350
transform 1 0 10764 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_701
timestamp 1606120350
transform 1 0 9568 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1091__CLK
timestamp 1606120350
transform 1 0 10580 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_93
timestamp 1606120350
transform 1 0 9660 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_101
timestamp 1606120350
transform 1 0 10396 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _0710_
timestamp 1606120350
transform 1 0 13248 0 -1 37536
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0660__A2
timestamp 1606120350
transform 1 0 12696 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__A1_N
timestamp 1606120350
transform 1 0 13064 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_124
timestamp 1606120350
transform 1 0 12512 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_128
timestamp 1606120350
transform 1 0 12880 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0709_
timestamp 1606120350
transform 1 0 15272 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_702
timestamp 1606120350
transform 1 0 15180 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__A2
timestamp 1606120350
transform 1 0 14628 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__B1
timestamp 1606120350
transform 1 0 14996 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_145
timestamp 1606120350
transform 1 0 14444 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_149
timestamp 1606120350
transform 1 0 14812 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_157
timestamp 1606120350
transform 1 0 15548 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _0730_
timestamp 1606120350
transform 1 0 16284 0 -1 37536
box -38 -48 1326 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0551__A2
timestamp 1606120350
transform 1 0 16008 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__B1
timestamp 1606120350
transform 1 0 17756 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_64_161
timestamp 1606120350
transform 1 0 15916 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_164
timestamp 1606120350
transform 1 0 16192 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_64_179
timestamp 1606120350
transform 1 0 17572 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_4  _0708_
timestamp 1606120350
transform 1 0 18308 0 -1 37536
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0621__B1
timestamp 1606120350
transform 1 0 18124 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__A2
timestamp 1606120350
transform 1 0 19964 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_183
timestamp 1606120350
transform 1 0 17940 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_200
timestamp 1606120350
transform 1 0 19504 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_204
timestamp 1606120350
transform 1 0 19872 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_703
timestamp 1606120350
transform 1 0 20792 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__A1
timestamp 1606120350
transform 1 0 20332 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_207
timestamp 1606120350
transform 1 0 20148 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_211
timestamp 1606120350
transform 1 0 20516 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_215
timestamp 1606120350
transform 1 0 20884 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_227
timestamp 1606120350
transform 1 0 21988 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1132_
timestamp 1606120350
transform 1 0 23092 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__B1
timestamp 1606120350
transform 1 0 25024 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_258
timestamp 1606120350
transform 1 0 24840 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_262
timestamp 1606120350
transform 1 0 25208 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_274
timestamp 1606120350
transform 1 0 26312 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0830_
timestamp 1606120350
transform 1 0 26864 0 -1 37536
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_704
timestamp 1606120350
transform 1 0 26404 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_276
timestamp 1606120350
transform 1 0 26496 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_289
timestamp 1606120350
transform 1 0 27692 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_301
timestamp 1606120350
transform 1 0 28796 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_313
timestamp 1606120350
transform 1 0 29900 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1201_
timestamp 1606120350
transform 1 0 32108 0 -1 37536
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_705
timestamp 1606120350
transform 1 0 32016 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_325
timestamp 1606120350
transform 1 0 31004 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_333
timestamp 1606120350
transform 1 0 31740 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_356
timestamp 1606120350
transform 1 0 33856 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_368
timestamp 1606120350
transform 1 0 34960 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_380
timestamp 1606120350
transform 1 0 36064 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1606120350
transform -1 0 38824 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_706
timestamp 1606120350
transform 1 0 37628 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_392
timestamp 1606120350
transform 1 0 37168 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_396
timestamp 1606120350
transform 1 0 37536 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_398
timestamp 1606120350
transform 1 0 37720 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_406
timestamp 1606120350
transform 1 0 38456 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1606120350
transform 1 0 1104 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1606120350
transform 1 0 1380 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1606120350
transform 1 0 2484 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1606120350
transform 1 0 3588 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1606120350
transform 1 0 4692 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_707
timestamp 1606120350
transform 1 0 6716 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_65_51
timestamp 1606120350
transform 1 0 5796 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_59
timestamp 1606120350
transform 1 0 6532 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_65_62
timestamp 1606120350
transform 1 0 6808 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_74
timestamp 1606120350
transform 1 0 7912 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_86
timestamp 1606120350
transform 1 0 9016 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__B1
timestamp 1606120350
transform 1 0 11316 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__A1
timestamp 1606120350
transform 1 0 10948 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__B2
timestamp 1606120350
transform 1 0 10580 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_98
timestamp 1606120350
transform 1 0 10120 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_102
timestamp 1606120350
transform 1 0 10488 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_105
timestamp 1606120350
transform 1 0 10764 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_109
timestamp 1606120350
transform 1 0 11132 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_65_113
timestamp 1606120350
transform 1 0 11500 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _0781_
timestamp 1606120350
transform 1 0 12420 0 1 37536
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_708
timestamp 1606120350
transform 1 0 12328 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__B2
timestamp 1606120350
transform 1 0 12144 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__A2_N
timestamp 1606120350
transform 1 0 11776 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_118
timestamp 1606120350
transform 1 0 11960 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_139
timestamp 1606120350
transform 1 0 13892 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__B1
timestamp 1606120350
transform 1 0 14076 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_143
timestamp 1606120350
transform 1 0 14260 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_147
timestamp 1606120350
transform 1 0 14628 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0719__A
timestamp 1606120350
transform 1 0 14720 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0719_
timestamp 1606120350
transform 1 0 14904 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_153
timestamp 1606120350
transform 1 0 15180 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__A2
timestamp 1606120350
transform 1 0 15364 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_157
timestamp 1606120350
transform 1 0 15548 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0551__A1
timestamp 1606120350
transform 1 0 15732 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _0746_
timestamp 1606120350
transform 1 0 15916 0 1 37536
box -38 -48 1326 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0551__B1
timestamp 1606120350
transform 1 0 17388 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0621__A1
timestamp 1606120350
transform 1 0 17756 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_175
timestamp 1606120350
transform 1 0 17204 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_179
timestamp 1606120350
transform 1 0 17572 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a21oi_4  _0706_
timestamp 1606120350
transform 1 0 18032 0 1 37536
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_4  _0707_
timestamp 1606120350
transform 1 0 19964 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_709
timestamp 1606120350
transform 1 0 17940 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0707__B1
timestamp 1606120350
transform 1 0 19780 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0621__A2
timestamp 1606120350
transform 1 0 19412 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_197
timestamp 1606120350
transform 1 0 19228 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_201
timestamp 1606120350
transform 1 0 19596 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0591__A
timestamp 1606120350
transform 1 0 21252 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0591__B
timestamp 1606120350
transform 1 0 21620 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_217
timestamp 1606120350
transform 1 0 21068 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_221
timestamp 1606120350
transform 1 0 21436 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_65_225
timestamp 1606120350
transform 1 0 21804 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_710
timestamp 1606120350
transform 1 0 23552 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A2
timestamp 1606120350
transform 1 0 23920 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__B1_N
timestamp 1606120350
transform 1 0 23368 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_237
timestamp 1606120350
transform 1 0 22908 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_241
timestamp 1606120350
transform 1 0 23276 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_65_245
timestamp 1606120350
transform 1 0 23644 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_250
timestamp 1606120350
transform 1 0 24104 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _0850_
timestamp 1606120350
transform 1 0 24840 0 1 37536
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__A1
timestamp 1606120350
transform 1 0 24656 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0850__A2
timestamp 1606120350
transform 1 0 24288 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A2
timestamp 1606120350
transform 1 0 26220 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_254
timestamp 1606120350
transform 1 0 24472 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_271
timestamp 1606120350
transform 1 0 26036 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__a21bo_4  _0924_
timestamp 1606120350
transform 1 0 26772 0 1 37536
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__D
timestamp 1606120350
transform 1 0 28152 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__B1_N
timestamp 1606120350
transform 1 0 26588 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_275
timestamp 1606120350
transform 1 0 26404 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_292
timestamp 1606120350
transform 1 0 27968 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_65_296
timestamp 1606120350
transform 1 0 28336 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_711
timestamp 1606120350
transform 1 0 29164 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1184__CLK
timestamp 1606120350
transform 1 0 28520 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_65_300
timestamp 1606120350
transform 1 0 28704 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_304
timestamp 1606120350
transform 1 0 29072 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_306
timestamp 1606120350
transform 1 0 29256 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_318
timestamp 1606120350
transform 1 0 30360 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_330
timestamp 1606120350
transform 1 0 31464 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_342
timestamp 1606120350
transform 1 0 32568 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_354
timestamp 1606120350
transform 1 0 33672 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_712
timestamp 1606120350
transform 1 0 34776 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_367
timestamp 1606120350
transform 1 0 34868 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_379
timestamp 1606120350
transform 1 0 35972 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1606120350
transform -1 0 38824 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_391
timestamp 1606120350
transform 1 0 37076 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_403
timestamp 1606120350
transform 1 0 38180 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1164_
timestamp 1606120350
transform 1 0 1380 0 1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1606120350
transform 1 0 1104 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1606120350
transform 1 0 1104 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__D
timestamp 1606120350
transform 1 0 1564 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1164__CLK
timestamp 1606120350
transform 1 0 1932 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_3
timestamp 1606120350
transform 1 0 1380 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_7
timestamp 1606120350
transform 1 0 1748 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_11
timestamp 1606120350
transform 1 0 2116 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_22
timestamp 1606120350
transform 1 0 3128 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_713
timestamp 1606120350
transform 1 0 3956 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_23
timestamp 1606120350
transform 1 0 3220 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_32
timestamp 1606120350
transform 1 0 4048 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_44
timestamp 1606120350
transform 1 0 5152 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_34
timestamp 1606120350
transform 1 0 4232 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_720
timestamp 1606120350
transform 1 0 6716 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_56
timestamp 1606120350
transform 1 0 6256 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_68
timestamp 1606120350
transform 1 0 7360 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_46
timestamp 1606120350
transform 1 0 5336 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_58
timestamp 1606120350
transform 1 0 6440 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_62
timestamp 1606120350
transform 1 0 6808 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__D
timestamp 1606120350
transform 1 0 9384 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1126__CLK
timestamp 1606120350
transform 1 0 9016 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_80
timestamp 1606120350
transform 1 0 8464 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_74
timestamp 1606120350
transform 1 0 7912 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_88
timestamp 1606120350
transform 1 0 9200 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _0780_
timestamp 1606120350
transform 1 0 11316 0 -1 38624
box -38 -48 1326 592
use sky130_fd_sc_hd__dfxtp_4  _1126_
timestamp 1606120350
transform 1 0 9568 0 1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_714
timestamp 1606120350
transform 1 0 9568 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0780__A2
timestamp 1606120350
transform 1 0 11132 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_93
timestamp 1606120350
transform 1 0 9660 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_105
timestamp 1606120350
transform 1 0 10764 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_67_111
timestamp 1606120350
transform 1 0 11316 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_67_123
timestamp 1606120350
transform 1 0 12420 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_119
timestamp 1606120350
transform 1 0 12052 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_66_125
timestamp 1606120350
transform 1 0 12604 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_721
timestamp 1606120350
transform 1 0 12328 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_133
timestamp 1606120350
transform 1 0 13340 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_129
timestamp 1606120350
transform 1 0 12972 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_129
timestamp 1606120350
transform 1 0 12972 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0685__A1
timestamp 1606120350
transform 1 0 13156 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0781__B1
timestamp 1606120350
transform 1 0 12788 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__B2
timestamp 1606120350
transform 1 0 12788 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__A3
timestamp 1606120350
transform 1 0 13156 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__A1
timestamp 1606120350
transform 1 0 13524 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _0685_
timestamp 1606120350
transform 1 0 13340 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__a32oi_4  _0658_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 13708 0 1 38624
box -38 -48 2062 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_715
timestamp 1606120350
transform 1 0 15180 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__B2
timestamp 1606120350
transform 1 0 15456 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0730__C1
timestamp 1606120350
transform 1 0 14996 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0731__A3
timestamp 1606120350
transform 1 0 14628 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_145
timestamp 1606120350
transform 1 0 14444 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_149
timestamp 1606120350
transform 1 0 14812 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_154
timestamp 1606120350
transform 1 0 15272 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_158
timestamp 1606120350
transform 1 0 15640 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_159
timestamp 1606120350
transform 1 0 15732 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_163
timestamp 1606120350
transform 1 0 16100 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__B1
timestamp 1606120350
transform 1 0 15824 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0509__B
timestamp 1606120350
transform 1 0 16284 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0509__A
timestamp 1606120350
transform 1 0 15916 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0674_
timestamp 1606120350
transform 1 0 16468 0 1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_67_182
timestamp 1606120350
transform 1 0 17848 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_178
timestamp 1606120350
transform 1 0 17480 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_174
timestamp 1606120350
transform 1 0 17112 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_179
timestamp 1606120350
transform 1 0 17572 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_66_175
timestamp 1606120350
transform 1 0 17204 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__A1
timestamp 1606120350
transform 1 0 17388 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__B1
timestamp 1606120350
transform 1 0 17664 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__B
timestamp 1606120350
transform 1 0 17296 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _0551_
timestamp 1606120350
transform 1 0 16008 0 -1 38624
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_66_186
timestamp 1606120350
transform 1 0 18216 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_66_183
timestamp 1606120350
transform 1 0 17940 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0623__A2
timestamp 1606120350
transform 1 0 18032 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_722
timestamp 1606120350
transform 1 0 17940 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_200
timestamp 1606120350
transform 1 0 19504 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_196
timestamp 1606120350
transform 1 0 19136 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_202
timestamp 1606120350
transform 1 0 19688 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0623__B1
timestamp 1606120350
transform 1 0 19320 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0492__C
timestamp 1606120350
transform 1 0 19872 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0492__B
timestamp 1606120350
transform 1 0 19688 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0492_
timestamp 1606120350
transform 1 0 19872 0 1 38624
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _0623_
timestamp 1606120350
transform 1 0 18032 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_4  _0621_
timestamp 1606120350
transform 1 0 18492 0 -1 38624
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_67_213
timestamp 1606120350
transform 1 0 20700 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_210
timestamp 1606120350
transform 1 0 20424 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_206
timestamp 1606120350
transform 1 0 20056 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0492__D
timestamp 1606120350
transform 1 0 20608 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0498__A
timestamp 1606120350
transform 1 0 20884 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0706__A1
timestamp 1606120350
transform 1 0 20240 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_716
timestamp 1606120350
transform 1 0 20792 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0591_
timestamp 1606120350
transform 1 0 20884 0 -1 38624
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_67_228
timestamp 1606120350
transform 1 0 22080 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_224
timestamp 1606120350
transform 1 0 21712 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_217
timestamp 1606120350
transform 1 0 21068 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_222
timestamp 1606120350
transform 1 0 21528 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1156__CLK
timestamp 1606120350
transform 1 0 21712 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1156__D
timestamp 1606120350
transform 1 0 21252 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0493__A
timestamp 1606120350
transform 1 0 21896 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0493_
timestamp 1606120350
transform 1 0 21436 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_226
timestamp 1606120350
transform 1 0 21896 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_723
timestamp 1606120350
transform 1 0 23552 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__B1
timestamp 1606120350
transform 1 0 23920 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0915__A1
timestamp 1606120350
transform 1 0 24104 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0492__A
timestamp 1606120350
transform 1 0 22264 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_238
timestamp 1606120350
transform 1 0 23000 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_232
timestamp 1606120350
transform 1 0 22448 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_67_245
timestamp 1606120350
transform 1 0 23644 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_250
timestamp 1606120350
transform 1 0 24104 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_254
timestamp 1606120350
transform 1 0 24472 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__A1
timestamp 1606120350
transform 1 0 24288 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0871__A2
timestamp 1606120350
transform 1 0 24656 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_67_271
timestamp 1606120350
transform 1 0 26036 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_66_269
timestamp 1606120350
transform 1 0 25852 0 -1 38624
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_66_265
timestamp 1606120350
transform 1 0 25484 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0869__A
timestamp 1606120350
transform 1 0 25668 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0848__A
timestamp 1606120350
transform 1 0 26220 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__a21bo_4  _0915_
timestamp 1606120350
transform 1 0 24288 0 -1 38624
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _0871_
timestamp 1606120350
transform 1 0 24840 0 1 38624
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_67_275
timestamp 1606120350
transform 1 0 26404 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_285
timestamp 1606120350
transform 1 0 27324 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_66_281
timestamp 1606120350
transform 1 0 26956 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_66_276
timestamp 1606120350
transform 1 0 26496 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__B1
timestamp 1606120350
transform 1 0 27140 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__A2
timestamp 1606120350
transform 1 0 26772 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0849__A1
timestamp 1606120350
transform 1 0 26588 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_717
timestamp 1606120350
transform 1 0 26404 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0924__A1
timestamp 1606120350
transform 1 0 27508 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_291
timestamp 1606120350
transform 1 0 27876 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1184_
timestamp 1606120350
transform 1 0 27692 0 -1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__o21a_4  _0849_
timestamp 1606120350
transform 1 0 26772 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_306
timestamp 1606120350
transform 1 0 29256 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_67_303
timestamp 1606120350
transform 1 0 28980 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_308
timestamp 1606120350
transform 1 0 29440 0 -1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_724
timestamp 1606120350
transform 1 0 29164 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_67_310
timestamp 1606120350
transform 1 0 29624 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_66_312
timestamp 1606120350
transform 1 0 29808 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__CLK
timestamp 1606120350
transform 1 0 29900 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1117__D
timestamp 1606120350
transform 1 0 29716 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_315
timestamp 1606120350
transform 1 0 30084 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1117_
timestamp 1606120350
transform 1 0 29900 0 1 38624
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_718
timestamp 1606120350
transform 1 0 32016 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_327
timestamp 1606120350
transform 1 0 31188 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_335
timestamp 1606120350
transform 1 0 31924 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_337
timestamp 1606120350
transform 1 0 32108 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_332
timestamp 1606120350
transform 1 0 31648 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_349
timestamp 1606120350
transform 1 0 33212 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_361
timestamp 1606120350
transform 1 0 34316 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_344
timestamp 1606120350
transform 1 0 32752 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_356
timestamp 1606120350
transform 1 0 33856 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_364
timestamp 1606120350
transform 1 0 34592 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_725
timestamp 1606120350
transform 1 0 34776 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0552__A
timestamp 1606120350
transform 1 0 35052 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_373
timestamp 1606120350
transform 1 0 35420 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_385
timestamp 1606120350
transform 1 0 36524 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_67_367
timestamp 1606120350
transform 1 0 34868 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_371
timestamp 1606120350
transform 1 0 35236 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_383
timestamp 1606120350
transform 1 0 36340 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1606120350
transform -1 0 38824 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1606120350
transform -1 0 38824 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_719
timestamp 1606120350
transform 1 0 37628 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_66_398
timestamp 1606120350
transform 1 0 37720 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_406
timestamp 1606120350
transform 1 0 38456 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_395
timestamp 1606120350
transform 1 0 37444 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1606120350
transform 1 0 1104 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__A
timestamp 1606120350
transform 1 0 2392 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__D
timestamp 1606120350
transform 1 0 1564 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1082__B
timestamp 1606120350
transform 1 0 2760 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_3
timestamp 1606120350
transform 1 0 1380 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_68_7
timestamp 1606120350
transform 1 0 1748 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_13
timestamp 1606120350
transform 1 0 2300 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_68_16
timestamp 1606120350
transform 1 0 2576 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_20
timestamp 1606120350
transform 1 0 2944 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_726
timestamp 1606120350
transform 1 0 3956 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_28
timestamp 1606120350
transform 1 0 3680 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_32
timestamp 1606120350
transform 1 0 4048 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_44
timestamp 1606120350
transform 1 0 5152 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_56
timestamp 1606120350
transform 1 0 6256 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_68
timestamp 1606120350
transform 1 0 7360 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_80
timestamp 1606120350
transform 1 0 8464 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_727
timestamp 1606120350
transform 1 0 9568 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_93
timestamp 1606120350
transform 1 0 9660 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_105
timestamp 1606120350
transform 1 0 10764 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__A2
timestamp 1606120350
transform 1 0 13708 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_68_117
timestamp 1606120350
transform 1 0 11868 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_129
timestamp 1606120350
transform 1 0 12972 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__and2_4  _0509_
timestamp 1606120350
transform 1 0 15456 0 -1 39712
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_728
timestamp 1606120350
transform 1 0 15180 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0658__B1
timestamp 1606120350
transform 1 0 14076 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0747__A2
timestamp 1606120350
transform 1 0 14444 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__C1
timestamp 1606120350
transform 1 0 14996 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_139
timestamp 1606120350
transform 1 0 13892 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_143
timestamp 1606120350
transform 1 0 14260 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_147
timestamp 1606120350
transform 1 0 14628 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_68_154
timestamp 1606120350
transform 1 0 15272 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _0650_
timestamp 1606120350
transform 1 0 17204 0 -1 39712
box -38 -48 1326 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__A2
timestamp 1606120350
transform 1 0 17020 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0650__C1
timestamp 1606120350
transform 1 0 16652 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0674__A
timestamp 1606120350
transform 1 0 16284 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_163
timestamp 1606120350
transform 1 0 16100 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_167
timestamp 1606120350
transform 1 0 16468 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_171
timestamp 1606120350
transform 1 0 16836 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0498_
timestamp 1606120350
transform 1 0 19228 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0622__C
timestamp 1606120350
transform 1 0 18676 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0623__A1
timestamp 1606120350
transform 1 0 19044 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_189
timestamp 1606120350
transform 1 0 18492 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_193
timestamp 1606120350
transform 1 0 18860 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1156_
timestamp 1606120350
transform 1 0 21344 0 -1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_729
timestamp 1606120350
transform 1 0 20792 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0547__C
timestamp 1606120350
transform 1 0 20240 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0548__A
timestamp 1606120350
transform 1 0 21068 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0547__A
timestamp 1606120350
transform 1 0 20608 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_206
timestamp 1606120350
transform 1 0 20056 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_210
timestamp 1606120350
transform 1 0 20424 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_68_215
timestamp 1606120350
transform 1 0 20884 0 -1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_68_219
timestamp 1606120350
transform 1 0 21252 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_239
timestamp 1606120350
transform 1 0 23092 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_251
timestamp 1606120350
transform 1 0 24196 0 -1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__inv_8  _0869_
timestamp 1606120350
transform 1 0 24840 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_68_257
timestamp 1606120350
transform 1 0 24748 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_267
timestamp 1606120350
transform 1 0 25668 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__inv_8  _0848_
timestamp 1606120350
transform 1 0 26496 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_730
timestamp 1606120350
transform 1 0 26404 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_285
timestamp 1606120350
transform 1 0 27324 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_297
timestamp 1606120350
transform 1 0 28428 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_309
timestamp 1606120350
transform 1 0 29532 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_731
timestamp 1606120350
transform 1 0 32016 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_321
timestamp 1606120350
transform 1 0 30636 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_333
timestamp 1606120350
transform 1 0 31740 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_337
timestamp 1606120350
transform 1 0 32108 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_8  _0552_
timestamp 1606120350
transform 1 0 34684 0 -1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_68_349
timestamp 1606120350
transform 1 0 33212 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_361
timestamp 1606120350
transform 1 0 34316 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_374
timestamp 1606120350
transform 1 0 35512 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_386
timestamp 1606120350
transform 1 0 36616 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1606120350
transform -1 0 38824 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_732
timestamp 1606120350
transform 1 0 37628 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_68_394
timestamp 1606120350
transform 1 0 37352 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_68_398
timestamp 1606120350
transform 1 0 37720 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_68_406
timestamp 1606120350
transform 1 0 38456 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1115_
timestamp 1606120350
transform 1 0 1564 0 1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1606120350
transform 1 0 1104 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_3
timestamp 1606120350
transform 1 0 1380 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_24
timestamp 1606120350
transform 1 0 3312 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_36
timestamp 1606120350
transform 1 0 4416 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_733
timestamp 1606120350
transform 1 0 6716 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_48
timestamp 1606120350
transform 1 0 5520 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_60
timestamp 1606120350
transform 1 0 6624 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_62
timestamp 1606120350
transform 1 0 6808 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_74
timestamp 1606120350
transform 1 0 7912 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_86
timestamp 1606120350
transform 1 0 9016 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__D
timestamp 1606120350
transform 1 0 11316 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_98
timestamp 1606120350
transform 1 0 10120 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_110
timestamp 1606120350
transform 1 0 11224 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_113
timestamp 1606120350
transform 1 0 11500 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_121
timestamp 1606120350
transform 1 0 12236 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_117
timestamp 1606120350
transform 1 0 11868 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1090__CLK
timestamp 1606120350
transform 1 0 11684 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_123
timestamp 1606120350
transform 1 0 12420 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_734
timestamp 1606120350
transform 1 0 12328 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_133
timestamp 1606120350
transform 1 0 13340 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_129
timestamp 1606120350
transform 1 0 12972 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0664_
timestamp 1606120350
transform 1 0 13064 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_137
timestamp 1606120350
transform 1 0 13708 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0664__A
timestamp 1606120350
transform 1 0 13524 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0501__A
timestamp 1606120350
transform 1 0 15456 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0779__A
timestamp 1606120350
transform 1 0 13892 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0746__A1
timestamp 1606120350
transform 1 0 15088 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_141
timestamp 1606120350
transform 1 0 14076 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_69_149
timestamp 1606120350
transform 1 0 14812 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_154
timestamp 1606120350
transform 1 0 15272 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_158
timestamp 1606120350
transform 1 0 15640 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0651_
timestamp 1606120350
transform 1 0 16008 0 1 39712
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0651__A
timestamp 1606120350
transform 1 0 15824 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0549__A
timestamp 1606120350
transform 1 0 17020 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0622__A
timestamp 1606120350
transform 1 0 17756 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_171
timestamp 1606120350
transform 1 0 16836 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_69_175
timestamp 1606120350
transform 1 0 17204 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_735
timestamp 1606120350
transform 1 0 17940 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 18768 0 1 39712
box -38 -48 1878 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_clk_A
timestamp 1606120350
transform 1 0 18584 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0622__B
timestamp 1606120350
transform 1 0 18216 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_184
timestamp 1606120350
transform 1 0 18032 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_188
timestamp 1606120350
transform 1 0 18400 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1148_
timestamp 1606120350
transform 1 0 21068 0 1 39712
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0547__B
timestamp 1606120350
transform 1 0 20792 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_212
timestamp 1606120350
transform 1 0 20608 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_69_216
timestamp 1606120350
transform 1 0 20976 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_736
timestamp 1606120350
transform 1 0 23552 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__D
timestamp 1606120350
transform 1 0 23000 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1157__CLK
timestamp 1606120350
transform 1 0 23368 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_236
timestamp 1606120350
transform 1 0 22816 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_240
timestamp 1606120350
transform 1 0 23184 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_245
timestamp 1606120350
transform 1 0 23644 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_4  _0870_
timestamp 1606120350
transform 1 0 25576 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A2
timestamp 1606120350
transform 1 0 25392 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__A1
timestamp 1606120350
transform 1 0 25024 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_69_257
timestamp 1606120350
transform 1 0 24748 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_69_262
timestamp 1606120350
transform 1 0 25208 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_278
timestamp 1606120350
transform 1 0 26680 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_290
timestamp 1606120350
transform 1 0 27784 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_737
timestamp 1606120350
transform 1 0 29164 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_69_302
timestamp 1606120350
transform 1 0 28888 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_306
timestamp 1606120350
transform 1 0 29256 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_318
timestamp 1606120350
transform 1 0 30360 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_330
timestamp 1606120350
transform 1 0 31464 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_342
timestamp 1606120350
transform 1 0 32568 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_354
timestamp 1606120350
transform 1 0 33672 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_738
timestamp 1606120350
transform 1 0 34776 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__D
timestamp 1606120350
transform 1 0 35052 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1154__CLK
timestamp 1606120350
transform 1 0 35420 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_367
timestamp 1606120350
transform 1 0 34868 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_69_371
timestamp 1606120350
transform 1 0 35236 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_69_375
timestamp 1606120350
transform 1 0 35604 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_387
timestamp 1606120350
transform 1 0 36708 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1606120350
transform -1 0 38824 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_69_399
timestamp 1606120350
transform 1 0 37812 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _1082_
timestamp 1606120350
transform 1 0 2392 0 -1 40800
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1606120350
transform 1 0 1104 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1115__CLK
timestamp 1606120350
transform 1 0 1564 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_3
timestamp 1606120350
transform 1 0 1380 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_7
timestamp 1606120350
transform 1 0 1748 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_13
timestamp 1606120350
transform 1 0 2300 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_21
timestamp 1606120350
transform 1 0 3036 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_739
timestamp 1606120350
transform 1 0 3956 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_29
timestamp 1606120350
transform 1 0 3772 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_32
timestamp 1606120350
transform 1 0 4048 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_44
timestamp 1606120350
transform 1 0 5152 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_56
timestamp 1606120350
transform 1 0 6256 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_68
timestamp 1606120350
transform 1 0 7360 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_80
timestamp 1606120350
transform 1 0 8464 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1090_
timestamp 1606120350
transform 1 0 11316 0 -1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_740
timestamp 1606120350
transform 1 0 9568 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_93
timestamp 1606120350
transform 1 0 9660 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_105
timestamp 1606120350
transform 1 0 10764 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_70_130
timestamp 1606120350
transform 1 0 13064 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _0779_
timestamp 1606120350
transform 1 0 13800 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_741
timestamp 1606120350
transform 1 0 15180 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1606120350
transform 1 0 14076 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_154
timestamp 1606120350
transform 1 0 15272 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0501_
timestamp 1606120350
transform 1 0 15916 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  _0549_
timestamp 1606120350
transform 1 0 17020 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_70_160
timestamp 1606120350
transform 1 0 15824 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_164
timestamp 1606120350
transform 1 0 16192 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_172
timestamp 1606120350
transform 1 0 16928 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_182
timestamp 1606120350
transform 1 0 17848 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _0547_
timestamp 1606120350
transform 1 0 19964 0 -1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__nand3_4  _0622_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 18676 0 -1 40800
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_1  FILLER_70_190
timestamp 1606120350
transform 1 0 18584 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0548_
timestamp 1606120350
transform 1 0 20884 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1157_
timestamp 1606120350
transform 1 0 22080 0 -1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_742
timestamp 1606120350
transform 1 0 20792 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__D
timestamp 1606120350
transform 1 0 21344 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1148__CLK
timestamp 1606120350
transform 1 0 21712 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_218
timestamp 1606120350
transform 1 0 21160 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_222
timestamp 1606120350
transform 1 0 21528 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_70_226
timestamp 1606120350
transform 1 0 21896 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_247
timestamp 1606120350
transform 1 0 23828 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0870__B1
timestamp 1606120350
transform 1 0 25576 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_259
timestamp 1606120350
transform 1 0 24932 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_265
timestamp 1606120350
transform 1 0 25484 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_268
timestamp 1606120350
transform 1 0 25760 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_274
timestamp 1606120350
transform 1 0 26312 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_743
timestamp 1606120350
transform 1 0 26404 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_276
timestamp 1606120350
transform 1 0 26496 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_288
timestamp 1606120350
transform 1 0 27600 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__A2
timestamp 1606120350
transform 1 0 29256 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_70_300
timestamp 1606120350
transform 1 0 28704 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_70_308
timestamp 1606120350
transform 1 0 29440 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_744
timestamp 1606120350
transform 1 0 32016 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_320
timestamp 1606120350
transform 1 0 30544 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_332
timestamp 1606120350
transform 1 0 31648 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_337
timestamp 1606120350
transform 1 0 32108 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_349
timestamp 1606120350
transform 1 0 33212 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_361
timestamp 1606120350
transform 1 0 34316 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _1154_
timestamp 1606120350
transform 1 0 34960 0 -1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_70_367
timestamp 1606120350
transform 1 0 34868 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_70_387
timestamp 1606120350
transform 1 0 36708 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1606120350
transform -1 0 38824 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_745
timestamp 1606120350
transform 1 0 37628 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_395
timestamp 1606120350
transform 1 0 37444 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_70_398
timestamp 1606120350
transform 1 0 37720 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_406
timestamp 1606120350
transform 1 0 38456 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1606120350
transform 1 0 1104 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1606120350
transform 1 0 1380 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_15
timestamp 1606120350
transform 1 0 2484 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__D
timestamp 1606120350
transform 1 0 4048 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1163__CLK
timestamp 1606120350
transform 1 0 4416 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_27
timestamp 1606120350
transform 1 0 3588 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_71_31
timestamp 1606120350
transform 1 0 3956 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_34
timestamp 1606120350
transform 1 0 4232 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_38
timestamp 1606120350
transform 1 0 4600 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_746
timestamp 1606120350
transform 1 0 6716 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_50
timestamp 1606120350
transform 1 0 5704 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_58
timestamp 1606120350
transform 1 0 6440 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_62
timestamp 1606120350
transform 1 0 6808 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_74
timestamp 1606120350
transform 1 0 7912 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_86
timestamp 1606120350
transform 1 0 9016 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__D
timestamp 1606120350
transform 1 0 10304 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1127__CLK
timestamp 1606120350
transform 1 0 10672 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_98
timestamp 1606120350
transform 1 0 10120 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_102
timestamp 1606120350
transform 1 0 10488 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_106
timestamp 1606120350
transform 1 0 10856 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_747
timestamp 1606120350
transform 1 0 12328 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__A
timestamp 1606120350
transform 1 0 13064 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0776__B
timestamp 1606120350
transform 1 0 13432 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_71_118
timestamp 1606120350
transform 1 0 11960 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_71_123
timestamp 1606120350
transform 1 0 12420 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_129
timestamp 1606120350
transform 1 0 12972 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_132
timestamp 1606120350
transform 1 0 13248 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_136
timestamp 1606120350
transform 1 0 13616 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_148
timestamp 1606120350
transform 1 0 14720 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_160
timestamp 1606120350
transform 1 0 15824 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_172
timestamp 1606120350
transform 1 0 16928 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_180
timestamp 1606120350
transform 1 0 17664 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _0499_
timestamp 1606120350
transform 1 0 19136 0 1 40800
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0500_
timestamp 1606120350
transform 1 0 18032 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_748
timestamp 1606120350
transform 1 0 17940 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0499__C
timestamp 1606120350
transform 1 0 18952 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0500__A
timestamp 1606120350
transform 1 0 18492 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_187
timestamp 1606120350
transform 1 0 18308 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_71_191
timestamp 1606120350
transform 1 0 18676 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_71_205
timestamp 1606120350
transform 1 0 19964 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1149_
timestamp 1606120350
transform 1 0 21068 0 1 40800
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__D
timestamp 1606120350
transform 1 0 20884 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0499__B
timestamp 1606120350
transform 1 0 20148 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0488__A
timestamp 1606120350
transform 1 0 20516 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_209
timestamp 1606120350
transform 1 0 20332 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_213
timestamp 1606120350
transform 1 0 20700 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_749
timestamp 1606120350
transform 1 0 23552 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__D
timestamp 1606120350
transform 1 0 23828 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1228__CLK
timestamp 1606120350
transform 1 0 24196 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_236
timestamp 1606120350
transform 1 0 22816 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_245
timestamp 1606120350
transform 1 0 23644 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_71_249
timestamp 1606120350
transform 1 0 24012 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_253
timestamp 1606120350
transform 1 0 24380 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_265
timestamp 1606120350
transform 1 0 25484 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__D
timestamp 1606120350
transform 1 0 27232 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1190__CLK
timestamp 1606120350
transform 1 0 27600 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_277
timestamp 1606120350
transform 1 0 26588 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_283
timestamp 1606120350
transform 1 0 27140 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_71_286
timestamp 1606120350
transform 1 0 27416 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_290
timestamp 1606120350
transform 1 0 27784 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__a21bo_4  _0931_
timestamp 1606120350
transform 1 0 29256 0 1 40800
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_750
timestamp 1606120350
transform 1 0 29164 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__B1_N
timestamp 1606120350
transform 1 0 28980 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_71_302
timestamp 1606120350
transform 1 0 28888 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_319
timestamp 1606120350
transform 1 0 30452 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_331
timestamp 1606120350
transform 1 0 31556 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_343
timestamp 1606120350
transform 1 0 32660 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_355
timestamp 1606120350
transform 1 0 33764 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_71_363
timestamp 1606120350
transform 1 0 34500 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_751
timestamp 1606120350
transform 1 0 34776 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_367
timestamp 1606120350
transform 1 0 34868 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_379
timestamp 1606120350
transform 1 0 35972 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1606120350
transform -1 0 38824 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_391
timestamp 1606120350
transform 1 0 37076 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_403
timestamp 1606120350
transform 1 0 38180 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1606120350
transform 1 0 1104 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1606120350
transform 1 0 1104 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1606120350
transform 1 0 1380 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_15
timestamp 1606120350
transform 1 0 2484 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_3
timestamp 1606120350
transform 1 0 1380 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_15
timestamp 1606120350
transform 1 0 2484 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1163_
timestamp 1606120350
transform 1 0 4048 0 -1 41888
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_752
timestamp 1606120350
transform 1 0 3956 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_27
timestamp 1606120350
transform 1 0 3588 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_27
timestamp 1606120350
transform 1 0 3588 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_39
timestamp 1606120350
transform 1 0 4692 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_759
timestamp 1606120350
transform 1 0 6716 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_51
timestamp 1606120350
transform 1 0 5796 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_63
timestamp 1606120350
transform 1 0 6900 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_51
timestamp 1606120350
transform 1 0 5796 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_59
timestamp 1606120350
transform 1 0 6532 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_62
timestamp 1606120350
transform 1 0 6808 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_75
timestamp 1606120350
transform 1 0 8004 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_87
timestamp 1606120350
transform 1 0 9108 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_91
timestamp 1606120350
transform 1 0 9476 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_74
timestamp 1606120350
transform 1 0 7912 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_86
timestamp 1606120350
transform 1 0 9016 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1127_
timestamp 1606120350
transform 1 0 10304 0 -1 41888
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_753
timestamp 1606120350
transform 1 0 9568 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_93
timestamp 1606120350
transform 1 0 9660 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_99
timestamp 1606120350
transform 1 0 10212 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_98
timestamp 1606120350
transform 1 0 10120 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_110
timestamp 1606120350
transform 1 0 11224 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_118
timestamp 1606120350
transform 1 0 11960 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_119
timestamp 1606120350
transform 1 0 12052 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__B1
timestamp 1606120350
transform 1 0 12144 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_760
timestamp 1606120350
transform 1 0 12328 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_126
timestamp 1606120350
transform 1 0 12696 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_72_129
timestamp 1606120350
transform 1 0 12972 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_125
timestamp 1606120350
transform 1 0 12604 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__A2
timestamp 1606120350
transform 1 0 12420 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0815__A
timestamp 1606120350
transform 1 0 12880 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0815_
timestamp 1606120350
transform 1 0 12420 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_73_134
timestamp 1606120350
transform 1 0 13432 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_130
timestamp 1606120350
transform 1 0 13064 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_137
timestamp 1606120350
transform 1 0 13708 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0777__A1
timestamp 1606120350
transform 1 0 13248 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0776_
timestamp 1606120350
transform 1 0 13064 0 -1 41888
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_4  _0756_
timestamp 1606120350
transform 1 0 14076 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_754
timestamp 1606120350
transform 1 0 15180 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__A1
timestamp 1606120350
transform 1 0 13892 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__B1
timestamp 1606120350
transform 1 0 14076 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_143
timestamp 1606120350
transform 1 0 14260 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_72_151
timestamp 1606120350
transform 1 0 14996 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_154
timestamp 1606120350
transform 1 0 15272 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_138
timestamp 1606120350
transform 1 0 13800 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_153
timestamp 1606120350
transform 1 0 15180 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_166
timestamp 1606120350
transform 1 0 16376 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_178
timestamp 1606120350
transform 1 0 17480 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_165
timestamp 1606120350
transform 1 0 16284 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_177
timestamp 1606120350
transform 1 0 17388 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_73_192
timestamp 1606120350
transform 1 0 18768 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_184
timestamp 1606120350
transform 1 0 18032 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_190
timestamp 1606120350
transform 1 0 18584 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_761
timestamp 1606120350
transform 1 0 17940 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_196
timestamp 1606120350
transform 1 0 19136 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_72_194
timestamp 1606120350
transform 1 0 18952 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0499__A
timestamp 1606120350
transform 1 0 19044 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__A
timestamp 1606120350
transform 1 0 18952 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__C
timestamp 1606120350
transform 1 0 19320 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0620_
timestamp 1606120350
transform 1 0 19504 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  _0488_
timestamp 1606120350
transform 1 0 19228 0 -1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_73_209
timestamp 1606120350
transform 1 0 20332 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_72_215
timestamp 1606120350
transform 1 0 20884 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_206
timestamp 1606120350
transform 1 0 20056 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__D
timestamp 1606120350
transform 1 0 20884 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_755
timestamp 1606120350
transform 1 0 20792 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_217
timestamp 1606120350
transform 1 0 21068 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1149__CLK
timestamp 1606120350
transform 1 0 21068 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1147__CLK
timestamp 1606120350
transform 1 0 21252 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_73_221
timestamp 1606120350
transform 1 0 21436 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_219
timestamp 1606120350
transform 1 0 21252 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _0914_ /home/rohan/openlane_build_script/work/tools/openlane_working_dir/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1606120350
transform 1 0 24012 0 1 41888
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_4  _1228_
timestamp 1606120350
transform 1 0 23460 0 -1 41888
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_762
timestamp 1606120350
transform 1 0 23552 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__A
timestamp 1606120350
transform 1 0 23828 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_231
timestamp 1606120350
transform 1 0 22356 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_233
timestamp 1606120350
transform 1 0 22540 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_73_241
timestamp 1606120350
transform 1 0 23276 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_73_245
timestamp 1606120350
transform 1 0 23644 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__a21bo_4  _0938_
timestamp 1606120350
transform 1 0 25576 0 1 41888
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A2
timestamp 1606120350
transform 1 0 25392 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__B1_N
timestamp 1606120350
transform 1 0 25576 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_262
timestamp 1606120350
transform 1 0 25208 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_72_268
timestamp 1606120350
transform 1 0 25760 0 -1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_274
timestamp 1606120350
transform 1 0 26312 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_258
timestamp 1606120350
transform 1 0 24840 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_73_283
timestamp 1606120350
transform 1 0 27140 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_73_279
timestamp 1606120350
transform 1 0 26772 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_280
timestamp 1606120350
transform 1 0 26864 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_72_276
timestamp 1606120350
transform 1 0 26496 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__A1
timestamp 1606120350
transform 1 0 26680 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__A
timestamp 1606120350
transform 1 0 27324 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0846__B
timestamp 1606120350
transform 1 0 26956 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_756
timestamp 1606120350
transform 1 0 26404 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_294
timestamp 1606120350
transform 1 0 28152 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_290
timestamp 1606120350
transform 1 0 27784 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0822__A
timestamp 1606120350
transform 1 0 27968 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0822_
timestamp 1606120350
transform 1 0 27508 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1190_
timestamp 1606120350
transform 1 0 27232 0 -1 41888
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_73_306
timestamp 1606120350
transform 1 0 29256 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_73_304
timestamp 1606120350
transform 1 0 29072 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_300
timestamp 1606120350
transform 1 0 28704 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_72_303
timestamp 1606120350
transform 1 0 28980 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0931__A1
timestamp 1606120350
transform 1 0 29256 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__A1
timestamp 1606120350
transform 1 0 29440 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__B1_N
timestamp 1606120350
transform 1 0 28888 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0898__A2
timestamp 1606120350
transform 1 0 28520 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_763
timestamp 1606120350
transform 1 0 29164 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_310
timestamp 1606120350
transform 1 0 29624 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_308
timestamp 1606120350
transform 1 0 29440 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_757
timestamp 1606120350
transform 1 0 32016 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_320
timestamp 1606120350
transform 1 0 30544 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_332
timestamp 1606120350
transform 1 0 31648 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_337
timestamp 1606120350
transform 1 0 32108 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_322
timestamp 1606120350
transform 1 0 30728 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_334
timestamp 1606120350
transform 1 0 31832 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__D
timestamp 1606120350
transform 1 0 33764 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1176__CLK
timestamp 1606120350
transform 1 0 34132 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_72_349
timestamp 1606120350
transform 1 0 33212 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_361
timestamp 1606120350
transform 1 0 34316 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_346
timestamp 1606120350
transform 1 0 32936 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_354
timestamp 1606120350
transform 1 0 33672 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_357
timestamp 1606120350
transform 1 0 33948 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_361
timestamp 1606120350
transform 1 0 34316 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_365
timestamp 1606120350
transform 1 0 34684 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_764
timestamp 1606120350
transform 1 0 34776 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_373
timestamp 1606120350
transform 1 0 35420 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_385
timestamp 1606120350
transform 1 0 36524 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_367
timestamp 1606120350
transform 1 0 34868 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_379
timestamp 1606120350
transform 1 0 35972 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1606120350
transform -1 0 38824 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1606120350
transform -1 0 38824 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_758
timestamp 1606120350
transform 1 0 37628 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_398
timestamp 1606120350
transform 1 0 37720 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_72_406
timestamp 1606120350
transform 1 0 38456 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_391
timestamp 1606120350
transform 1 0 37076 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_403
timestamp 1606120350
transform 1 0 38180 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1606120350
transform 1 0 1104 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1606120350
transform 1 0 1380 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1606120350
transform 1 0 2484 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_765
timestamp 1606120350
transform 1 0 3956 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_27
timestamp 1606120350
transform 1 0 3588 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_32
timestamp 1606120350
transform 1 0 4048 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_44
timestamp 1606120350
transform 1 0 5152 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_56
timestamp 1606120350
transform 1 0 6256 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_68
timestamp 1606120350
transform 1 0 7360 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_80
timestamp 1606120350
transform 1 0 8464 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_766
timestamp 1606120350
transform 1 0 9568 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_93
timestamp 1606120350
transform 1 0 9660 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_105
timestamp 1606120350
transform 1 0 10764 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__a21o_4  _0777_
timestamp 1606120350
transform 1 0 12420 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_117
timestamp 1606120350
transform 1 0 11868 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_74_135
timestamp 1606120350
transform 1 0 13524 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_767
timestamp 1606120350
transform 1 0 15180 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0756__A2
timestamp 1606120350
transform 1 0 14076 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_143
timestamp 1606120350
transform 1 0 14260 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_151
timestamp 1606120350
transform 1 0 14996 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_154
timestamp 1606120350
transform 1 0 15272 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_166
timestamp 1606120350
transform 1 0 16376 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_178
timestamp 1606120350
transform 1 0 17480 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0620__B
timestamp 1606120350
transform 1 0 19504 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_74_190
timestamp 1606120350
transform 1 0 18584 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_74_198
timestamp 1606120350
transform 1 0 19320 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_202
timestamp 1606120350
transform 1 0 19688 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1147_
timestamp 1606120350
transform 1 0 20884 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_768
timestamp 1606120350
transform 1 0 20792 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0914__B
timestamp 1606120350
transform 1 0 24012 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_234
timestamp 1606120350
transform 1 0 22632 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_74_246
timestamp 1606120350
transform 1 0 23736 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_74_251
timestamp 1606120350
transform 1 0 24196 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_74_256
timestamp 1606120350
transform 1 0 24656 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__B1_N
timestamp 1606120350
transform 1 0 24472 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_260
timestamp 1606120350
transform 1 0 25024 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__A1
timestamp 1606120350
transform 1 0 24840 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_264
timestamp 1606120350
transform 1 0 25392 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0827__A
timestamp 1606120350
transform 1 0 25208 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_268
timestamp 1606120350
transform 1 0 25760 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0938__A1
timestamp 1606120350
transform 1 0 25576 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_272
timestamp 1606120350
transform 1 0 26128 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__B
timestamp 1606120350
transform 1 0 26220 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0846_
timestamp 1606120350
transform 1 0 26680 0 -1 42976
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_769
timestamp 1606120350
transform 1 0 26404 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__C1
timestamp 1606120350
transform 1 0 27508 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__A1
timestamp 1606120350
transform 1 0 27876 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__A1
timestamp 1606120350
transform 1 0 28244 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_276
timestamp 1606120350
transform 1 0 26496 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_285
timestamp 1606120350
transform 1 0 27324 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_289
timestamp 1606120350
transform 1 0 27692 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_74_293
timestamp 1606120350
transform 1 0 28060 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__a21bo_4  _0898_
timestamp 1606120350
transform 1 0 28520 0 -1 42976
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__A1
timestamp 1606120350
transform 1 0 29900 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_74_297
timestamp 1606120350
transform 1 0 28428 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_74_311
timestamp 1606120350
transform 1 0 29716 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_315
timestamp 1606120350
transform 1 0 30084 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_770
timestamp 1606120350
transform 1 0 32016 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_74_327
timestamp 1606120350
transform 1 0 31188 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_335
timestamp 1606120350
transform 1 0 31924 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_337
timestamp 1606120350
transform 1 0 32108 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1176_
timestamp 1606120350
transform 1 0 33764 0 -1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_74_349
timestamp 1606120350
transform 1 0 33212 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_74_374
timestamp 1606120350
transform 1 0 35512 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_386
timestamp 1606120350
transform 1 0 36616 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1606120350
transform -1 0 38824 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_771
timestamp 1606120350
transform 1 0 37628 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_74_394
timestamp 1606120350
transform 1 0 37352 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_74_398
timestamp 1606120350
transform 1 0 37720 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_406
timestamp 1606120350
transform 1 0 38456 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1606120350
transform 1 0 1104 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_3
timestamp 1606120350
transform 1 0 1380 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_15
timestamp 1606120350
transform 1 0 2484 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_27
timestamp 1606120350
transform 1 0 3588 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_39
timestamp 1606120350
transform 1 0 4692 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_772
timestamp 1606120350
transform 1 0 6716 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_75_51
timestamp 1606120350
transform 1 0 5796 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_75_59
timestamp 1606120350
transform 1 0 6532 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_62
timestamp 1606120350
transform 1 0 6808 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_74
timestamp 1606120350
transform 1 0 7912 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_86
timestamp 1606120350
transform 1 0 9016 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__D
timestamp 1606120350
transform 1 0 10948 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1113__CLK
timestamp 1606120350
transform 1 0 11316 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_98
timestamp 1606120350
transform 1 0 10120 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_106
timestamp 1606120350
transform 1 0 10856 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_109
timestamp 1606120350
transform 1 0 11132 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_113
timestamp 1606120350
transform 1 0 11500 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1087_
timestamp 1606120350
transform 1 0 13064 0 1 42976
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_773
timestamp 1606120350
transform 1 0 12328 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__D
timestamp 1606120350
transform 1 0 12880 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_121
timestamp 1606120350
transform 1 0 12236 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_123
timestamp 1606120350
transform 1 0 12420 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_127
timestamp 1606120350
transform 1 0 12788 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__A
timestamp 1606120350
transform 1 0 15272 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0755__B
timestamp 1606120350
transform 1 0 15640 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_75_149
timestamp 1606120350
transform 1 0 14812 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_153
timestamp 1606120350
transform 1 0 15180 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_156
timestamp 1606120350
transform 1 0 15456 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_9_0_clk_A
timestamp 1606120350
transform 1 0 17756 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_160
timestamp 1606120350
transform 1 0 15824 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_172
timestamp 1606120350
transform 1 0 16928 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_180
timestamp 1606120350
transform 1 0 17664 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_774
timestamp 1606120350
transform 1 0 17940 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_184
timestamp 1606120350
transform 1 0 18032 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_196
timestamp 1606120350
transform 1 0 19136 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__D
timestamp 1606120350
transform 1 0 20884 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1155__CLK
timestamp 1606120350
transform 1 0 21252 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_75_208
timestamp 1606120350
transform 1 0 20240 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_214
timestamp 1606120350
transform 1 0 20792 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_217
timestamp 1606120350
transform 1 0 21068 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_221
timestamp 1606120350
transform 1 0 21436 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_775
timestamp 1606120350
transform 1 0 23552 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0825__A
timestamp 1606120350
transform 1 0 23828 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_233
timestamp 1606120350
transform 1 0 22540 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_75_241
timestamp 1606120350
transform 1 0 23276 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_75_245
timestamp 1606120350
transform 1 0 23644 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_75_249
timestamp 1606120350
transform 1 0 24012 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_4  _0919_
timestamp 1606120350
transform 1 0 24472 0 1 42976
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0897__A
timestamp 1606120350
transform 1 0 26220 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__A2
timestamp 1606120350
transform 1 0 25852 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0919__A2
timestamp 1606120350
transform 1 0 24288 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_267
timestamp 1606120350
transform 1 0 25668 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_271
timestamp 1606120350
transform 1 0 26036 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__a21bo_4  _0939_
timestamp 1606120350
transform 1 0 26404 0 1 42976
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__A2
timestamp 1606120350
transform 1 0 28244 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__B1
timestamp 1606120350
transform 1 0 27784 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_288
timestamp 1606120350
transform 1 0 27600 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_75_292
timestamp 1606120350
transform 1 0 27968 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_4  _0894_
timestamp 1606120350
transform 1 0 29256 0 1 42976
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_776
timestamp 1606120350
transform 1 0 29164 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__A2
timestamp 1606120350
transform 1 0 28980 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0889__B1_N
timestamp 1606120350
transform 1 0 28612 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_297
timestamp 1606120350
transform 1 0 28428 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_301
timestamp 1606120350
transform 1 0 28796 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_75_319
timestamp 1606120350
transform 1 0 30452 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0877__A
timestamp 1606120350
transform 1 0 30636 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_75_323
timestamp 1606120350
transform 1 0 30820 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_335
timestamp 1606120350
transform 1 0 31924 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_347
timestamp 1606120350
transform 1 0 33028 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_359
timestamp 1606120350
transform 1 0 34132 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_365
timestamp 1606120350
transform 1 0 34684 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_777
timestamp 1606120350
transform 1 0 34776 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_367
timestamp 1606120350
transform 1 0 34868 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_379
timestamp 1606120350
transform 1 0 35972 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1606120350
transform -1 0 38824 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_391
timestamp 1606120350
transform 1 0 37076 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_403
timestamp 1606120350
transform 1 0 38180 0 1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1606120350
transform 1 0 1104 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1606120350
transform 1 0 1380 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1606120350
transform 1 0 2484 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_778
timestamp 1606120350
transform 1 0 3956 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_27
timestamp 1606120350
transform 1 0 3588 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_32
timestamp 1606120350
transform 1 0 4048 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_44
timestamp 1606120350
transform 1 0 5152 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_56
timestamp 1606120350
transform 1 0 6256 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_68
timestamp 1606120350
transform 1 0 7360 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__CLK
timestamp 1606120350
transform 1 0 8280 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_76
timestamp 1606120350
transform 1 0 8096 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_76_80
timestamp 1606120350
transform 1 0 8464 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1113_
timestamp 1606120350
transform 1 0 10948 0 -1 44064
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_779
timestamp 1606120350
transform 1 0 9568 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_93
timestamp 1606120350
transform 1 0 9660 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_105
timestamp 1606120350
transform 1 0 10764 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1087__CLK
timestamp 1606120350
transform 1 0 13064 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_126
timestamp 1606120350
transform 1 0 12696 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_76_132
timestamp 1606120350
transform 1 0 13248 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__and2_4  _0755_
timestamp 1606120350
transform 1 0 15272 0 -1 44064
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_780
timestamp 1606120350
transform 1 0 15180 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_144
timestamp 1606120350
transform 1 0 14352 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_152
timestamp 1606120350
transform 1 0 15088 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_9_0_clk
timestamp 1606120350
transform 1 0 17756 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_161
timestamp 1606120350
transform 1 0 15916 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_173
timestamp 1606120350
transform 1 0 17020 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_184
timestamp 1606120350
transform 1 0 18032 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_196
timestamp 1606120350
transform 1 0 19136 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1155_
timestamp 1606120350
transform 1 0 20884 0 -1 44064
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_781
timestamp 1606120350
transform 1 0 20792 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_76_208
timestamp 1606120350
transform 1 0 20240 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0825_
timestamp 1606120350
transform 1 0 23644 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__A
timestamp 1606120350
transform 1 0 24104 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A1
timestamp 1606120350
transform 1 0 23460 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_76_234
timestamp 1606120350
transform 1 0 22632 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_242
timestamp 1606120350
transform 1 0 23368 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_76_248
timestamp 1606120350
transform 1 0 23920 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0827_
timestamp 1606120350
transform 1 0 24840 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__B
timestamp 1606120350
transform 1 0 24656 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__A2
timestamp 1606120350
transform 1 0 25852 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0939__B1_N
timestamp 1606120350
transform 1 0 26220 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_76_252
timestamp 1606120350
transform 1 0 24288 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_76_267
timestamp 1606120350
transform 1 0 25668 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_271
timestamp 1606120350
transform 1 0 26036 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__a21bo_4  _0889_
timestamp 1606120350
transform 1 0 28244 0 -1 44064
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_4  _0897_
timestamp 1606120350
transform 1 0 26496 0 -1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_782
timestamp 1606120350
transform 1 0 26404 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__A2
timestamp 1606120350
transform 1 0 27508 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__A2
timestamp 1606120350
transform 1 0 27876 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_285
timestamp 1606120350
transform 1 0 27324 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_289
timestamp 1606120350
transform 1 0 27692 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_293
timestamp 1606120350
transform 1 0 28060 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0877_
timestamp 1606120350
transform 1 0 30176 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0894__B1_N
timestamp 1606120350
transform 1 0 29624 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0896__A1
timestamp 1606120350
transform 1 0 29992 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_308
timestamp 1606120350
transform 1 0 29440 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_312
timestamp 1606120350
transform 1 0 29808 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_76_319
timestamp 1606120350
transform 1 0 30452 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_783
timestamp 1606120350
transform 1 0 32016 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__CLK
timestamp 1606120350
transform 1 0 30636 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_76_323
timestamp 1606120350
transform 1 0 30820 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_335
timestamp 1606120350
transform 1 0 31924 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_337
timestamp 1606120350
transform 1 0 32108 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_349
timestamp 1606120350
transform 1 0 33212 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_361
timestamp 1606120350
transform 1 0 34316 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__CLK
timestamp 1606120350
transform 1 0 36064 0 -1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_76_373
timestamp 1606120350
transform 1 0 35420 0 -1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_379
timestamp 1606120350
transform 1 0 35972 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_382
timestamp 1606120350
transform 1 0 36248 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1606120350
transform -1 0 38824 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_784
timestamp 1606120350
transform 1 0 37628 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_76_394
timestamp 1606120350
transform 1 0 37352 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_76_398
timestamp 1606120350
transform 1 0 37720 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_76_406
timestamp 1606120350
transform 1 0 38456 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1606120350
transform 1 0 1104 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__D
timestamp 1606120350
transform 1 0 1564 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1197__CLK
timestamp 1606120350
transform 1 0 1932 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_3
timestamp 1606120350
transform 1 0 1380 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_7
timestamp 1606120350
transform 1 0 1748 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_77_11
timestamp 1606120350
transform 1 0 2116 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_23
timestamp 1606120350
transform 1 0 3220 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_35
timestamp 1606120350
transform 1 0 4324 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_785
timestamp 1606120350
transform 1 0 6716 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_47
timestamp 1606120350
transform 1 0 5428 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_59
timestamp 1606120350
transform 1 0 6532 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_77_62
timestamp 1606120350
transform 1 0 6808 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1145_
timestamp 1606120350
transform 1 0 8280 0 1 44064
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1145__D
timestamp 1606120350
transform 1 0 8096 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_74
timestamp 1606120350
transform 1 0 7912 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_77_97
timestamp 1606120350
transform 1 0 10028 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_109
timestamp 1606120350
transform 1 0 11132 0 1 44064
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_4  _0820_
timestamp 1606120350
transform 1 0 12420 0 1 44064
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_786
timestamp 1606120350
transform 1 0 12328 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__A1
timestamp 1606120350
transform 1 0 12144 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__A2
timestamp 1606120350
transform 1 0 11776 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_77_115
timestamp 1606120350
transform 1 0 11684 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_118
timestamp 1606120350
transform 1 0 11960 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_137
timestamp 1606120350
transform 1 0 13708 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_4_0_clk
timestamp 1606120350
transform 1 0 15456 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0732__A
timestamp 1606120350
transform 1 0 13892 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_8_0_clk_A
timestamp 1606120350
transform 1 0 14260 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_141
timestamp 1606120350
transform 1 0 14076 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_77_145
timestamp 1606120350
transform 1 0 14444 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_153
timestamp 1606120350
transform 1 0 15180 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_77_159
timestamp 1606120350
transform 1 0 15732 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_4_0_clk_A
timestamp 1606120350
transform 1 0 15916 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_77_163
timestamp 1606120350
transform 1 0 16100 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_175
timestamp 1606120350
transform 1 0 17204 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_787
timestamp 1606120350
transform 1 0 17940 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_184
timestamp 1606120350
transform 1 0 18032 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_196
timestamp 1606120350
transform 1 0 19136 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_208
timestamp 1606120350
transform 1 0 20240 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_220
timestamp 1606120350
transform 1 0 21344 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_77_228
timestamp 1606120350
transform 1 0 22080 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _0828_
timestamp 1606120350
transform 1 0 24012 0 1 44064
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_788
timestamp 1606120350
transform 1 0 23552 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0828__B
timestamp 1606120350
transform 1 0 23828 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0824__A
timestamp 1606120350
transform 1 0 22264 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0840__A
timestamp 1606120350
transform 1 0 23276 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_77_232
timestamp 1606120350
transform 1 0 22448 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_240
timestamp 1606120350
transform 1 0 23184 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_77_243
timestamp 1606120350
transform 1 0 23460 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_245
timestamp 1606120350
transform 1 0 23644 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__a21bo_4  _0829_
timestamp 1606120350
transform 1 0 25392 0 1 44064
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__A1
timestamp 1606120350
transform 1 0 25208 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__A
timestamp 1606120350
transform 1 0 24840 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_256
timestamp 1606120350
transform 1 0 24656 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_260
timestamp 1606120350
transform 1 0 25024 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0896_
timestamp 1606120350
transform 1 0 27324 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0881__A
timestamp 1606120350
transform 1 0 26772 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0923__B1
timestamp 1606120350
transform 1 0 27140 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_277
timestamp 1606120350
transform 1 0 26588 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_281
timestamp 1606120350
transform 1 0 26956 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0922_
timestamp 1606120350
transform 1 0 29256 0 1 44064
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_789
timestamp 1606120350
transform 1 0 29164 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1169__D
timestamp 1606120350
transform 1 0 30268 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__A
timestamp 1606120350
transform 1 0 28980 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__C
timestamp 1606120350
transform 1 0 28612 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_297
timestamp 1606120350
transform 1 0 28428 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_301
timestamp 1606120350
transform 1 0 28796 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_315
timestamp 1606120350
transform 1 0 30084 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_319
timestamp 1606120350
transform 1 0 30452 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0844_
timestamp 1606120350
transform 1 0 30820 0 1 44064
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__A
timestamp 1606120350
transform 1 0 31648 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0844__B
timestamp 1606120350
transform 1 0 30636 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_77_330
timestamp 1606120350
transform 1 0 31464 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_77_334
timestamp 1606120350
transform 1 0 31832 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_346
timestamp 1606120350
transform 1 0 32936 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_358
timestamp 1606120350
transform 1 0 34040 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1212_
timestamp 1606120350
transform 1 0 36064 0 1 44064
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_790
timestamp 1606120350
transform 1 0 34776 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1212__D
timestamp 1606120350
transform 1 0 35880 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_77_367
timestamp 1606120350
transform 1 0 34868 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_77_375
timestamp 1606120350
transform 1 0 35604 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1606120350
transform -1 0 38824 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_77_399
timestamp 1606120350
transform 1 0 37812 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1197_
timestamp 1606120350
transform 1 0 1472 0 -1 45152
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1606120350
transform 1 0 1104 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_78_3
timestamp 1606120350
transform 1 0 1380 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_791
timestamp 1606120350
transform 1 0 3956 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_23
timestamp 1606120350
transform 1 0 3220 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_32
timestamp 1606120350
transform 1 0 4048 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_44
timestamp 1606120350
transform 1 0 5152 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_56
timestamp 1606120350
transform 1 0 6256 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_68
timestamp 1606120350
transform 1 0 7360 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__A2
timestamp 1606120350
transform 1 0 8832 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_80
timestamp 1606120350
transform 1 0 8464 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_78_86
timestamp 1606120350
transform 1 0 9016 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_792
timestamp 1606120350
transform 1 0 9568 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_93
timestamp 1606120350
transform 1 0 9660 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_105
timestamp 1606120350
transform 1 0 10764 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_8_0_clk
timestamp 1606120350
transform 1 0 13524 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__B2
timestamp 1606120350
transform 1 0 12420 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0820__B1
timestamp 1606120350
transform 1 0 12788 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__D
timestamp 1606120350
transform 1 0 13340 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_78_117
timestamp 1606120350
transform 1 0 11868 0 -1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_78_125
timestamp 1606120350
transform 1 0 12604 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_129
timestamp 1606120350
transform 1 0 12972 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _0732_
timestamp 1606120350
transform 1 0 13800 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_793
timestamp 1606120350
transform 1 0 15180 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__B
timestamp 1606120350
transform 1 0 14260 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_141
timestamp 1606120350
transform 1 0 14076 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_78_145
timestamp 1606120350
transform 1 0 14444 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_78_154
timestamp 1606120350
transform 1 0 15272 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_166
timestamp 1606120350
transform 1 0 16376 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_178
timestamp 1606120350
transform 1 0 17480 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_190
timestamp 1606120350
transform 1 0 18584 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_202
timestamp 1606120350
transform 1 0 19688 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_794
timestamp 1606120350
transform 1 0 20792 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__B
timestamp 1606120350
transform 1 0 22080 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_215
timestamp 1606120350
transform 1 0 20884 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_227
timestamp 1606120350
transform 1 0 21988 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0824_
timestamp 1606120350
transform 1 0 22264 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  _0840_
timestamp 1606120350
transform 1 0 23276 0 -1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__D
timestamp 1606120350
transform 1 0 23092 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__A
timestamp 1606120350
transform 1 0 22724 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_233
timestamp 1606120350
transform 1 0 22540 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_237
timestamp 1606120350
transform 1 0 22908 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_250
timestamp 1606120350
transform 1 0 24104 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _0845_
timestamp 1606120350
transform 1 0 24840 0 -1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__B1
timestamp 1606120350
transform 1 0 24288 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0829__B1_N
timestamp 1606120350
transform 1 0 25852 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0845__C
timestamp 1606120350
transform 1 0 24656 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__B1
timestamp 1606120350
transform 1 0 26220 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_254
timestamp 1606120350
transform 1 0 24472 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_267
timestamp 1606120350
transform 1 0 25668 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_271
timestamp 1606120350
transform 1 0 26036 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0881_
timestamp 1606120350
transform 1 0 26496 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_4  _0923_
timestamp 1606120350
transform 1 0 27508 0 -1 45152
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_795
timestamp 1606120350
transform 1 0 26404 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__C1
timestamp 1606120350
transform 1 0 26956 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__B
timestamp 1606120350
transform 1 0 27324 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_279
timestamp 1606120350
transform 1 0 26772 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_283
timestamp 1606120350
transform 1 0 27140 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1169_
timestamp 1606120350
transform 1 0 29532 0 -1 45152
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0922__B
timestamp 1606120350
transform 1 0 29256 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_301
timestamp 1606120350
transform 1 0 28796 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_305
timestamp 1606120350
transform 1 0 29164 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_78_308
timestamp 1606120350
transform 1 0 29440 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_796
timestamp 1606120350
transform 1 0 32016 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__C
timestamp 1606120350
transform 1 0 31464 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__D
timestamp 1606120350
transform 1 0 31832 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_328
timestamp 1606120350
transform 1 0 31280 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_78_332
timestamp 1606120350
transform 1 0 31648 0 -1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_78_337
timestamp 1606120350
transform 1 0 32108 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_349
timestamp 1606120350
transform 1 0 33212 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_361
timestamp 1606120350
transform 1 0 34316 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_373
timestamp 1606120350
transform 1 0 35420 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_385
timestamp 1606120350
transform 1 0 36524 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1606120350
transform -1 0 38824 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_797
timestamp 1606120350
transform 1 0 37628 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_398
timestamp 1606120350
transform 1 0 37720 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_78_406
timestamp 1606120350
transform 1 0 38456 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1606120350
transform 1 0 1104 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1606120350
transform 1 0 1104 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__D
timestamp 1606120350
transform 1 0 1564 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_3
timestamp 1606120350
transform 1 0 1380 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_15
timestamp 1606120350
transform 1 0 2484 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_3
timestamp 1606120350
transform 1 0 1380 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_80_7
timestamp 1606120350
transform 1 0 1748 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_19
timestamp 1606120350
transform 1 0 2852 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_804
timestamp 1606120350
transform 1 0 3956 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_27
timestamp 1606120350
transform 1 0 3588 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_39
timestamp 1606120350
transform 1 0 4692 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_32
timestamp 1606120350
transform 1 0 4048 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_44
timestamp 1606120350
transform 1 0 5152 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_798
timestamp 1606120350
transform 1 0 6716 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_79_51
timestamp 1606120350
transform 1 0 5796 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_59
timestamp 1606120350
transform 1 0 6532 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_62
timestamp 1606120350
transform 1 0 6808 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_56
timestamp 1606120350
transform 1 0 6256 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_68
timestamp 1606120350
transform 1 0 7360 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__a21bo_4  _0934_
timestamp 1606120350
transform 1 0 8832 0 1 45152
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__B1_N
timestamp 1606120350
transform 1 0 8648 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0934__A1
timestamp 1606120350
transform 1 0 8832 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_74
timestamp 1606120350
transform 1 0 7912 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_80
timestamp 1606120350
transform 1 0 8464 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_86
timestamp 1606120350
transform 1 0 9016 0 -1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_805
timestamp 1606120350
transform 1 0 9568 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_97
timestamp 1606120350
transform 1 0 10028 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_109
timestamp 1606120350
transform 1 0 11132 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_93
timestamp 1606120350
transform 1 0 9660 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_105
timestamp 1606120350
transform 1 0 10764 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_125
timestamp 1606120350
transform 1 0 12604 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_80_117
timestamp 1606120350
transform 1 0 11868 0 -1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_79_123
timestamp 1606120350
transform 1 0 12420 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_121
timestamp 1606120350
transform 1 0 12236 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__CLK
timestamp 1606120350
transform 1 0 12420 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_799
timestamp 1606120350
transform 1 0 12328 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_134
timestamp 1606120350
transform 1 0 13432 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_130
timestamp 1606120350
transform 1 0 13064 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_129
timestamp 1606120350
transform 1 0 12972 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1089__CLK
timestamp 1606120350
transform 1 0 13248 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__B
timestamp 1606120350
transform 1 0 13616 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0769__A
timestamp 1606120350
transform 1 0 13156 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0762__A
timestamp 1606120350
transform 1 0 12788 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0762_
timestamp 1606120350
transform 1 0 12788 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1089_
timestamp 1606120350
transform 1 0 13340 0 1 45152
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_4  FILLER_80_145
timestamp 1606120350
transform 1 0 14444 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _0769_
timestamp 1606120350
transform 1 0 13800 0 -1 46240
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_80_154
timestamp 1606120350
transform 1 0 15272 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_80_152
timestamp 1606120350
transform 1 0 15088 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_80_149
timestamp 1606120350
transform 1 0 14812 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__B
timestamp 1606120350
transform 1 0 15456 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__A1
timestamp 1606120350
transform 1 0 14904 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_806
timestamp 1606120350
transform 1 0 15180 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_158
timestamp 1606120350
transform 1 0 15640 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_152
timestamp 1606120350
transform 1 0 15088 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_164
timestamp 1606120350
transform 1 0 16192 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_176
timestamp 1606120350
transform 1 0 17296 0 1 45152
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_182
timestamp 1606120350
transform 1 0 17848 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_170
timestamp 1606120350
transform 1 0 16744 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_182
timestamp 1606120350
transform 1 0 17848 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_800
timestamp 1606120350
transform 1 0 17940 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_184
timestamp 1606120350
transform 1 0 18032 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_196
timestamp 1606120350
transform 1 0 19136 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_194
timestamp 1606120350
transform 1 0 18952 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_215
timestamp 1606120350
transform 1 0 20884 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_206
timestamp 1606120350
transform 1 0 20056 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_807
timestamp 1606120350
transform 1 0 20792 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_80_224
timestamp 1606120350
transform 1 0 21712 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_79_223
timestamp 1606120350
transform 1 0 21620 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_220
timestamp 1606120350
transform 1 0 21344 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__B
timestamp 1606120350
transform 1 0 21252 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0823__A
timestamp 1606120350
transform 1 0 21436 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__A
timestamp 1606120350
transform 1 0 21988 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__C
timestamp 1606120350
transform 1 0 21988 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0823_
timestamp 1606120350
transform 1 0 21436 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_79_208
timestamp 1606120350
transform 1 0 20240 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_80_229
timestamp 1606120350
transform 1 0 22172 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_236
timestamp 1606120350
transform 1 0 22816 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_229
timestamp 1606120350
transform 1 0 22172 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0832__A
timestamp 1606120350
transform 1 0 22356 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0831__C
timestamp 1606120350
transform 1 0 23000 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0832_
timestamp 1606120350
transform 1 0 22540 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _0831_
timestamp 1606120350
transform 1 0 22448 0 -1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_80_246
timestamp 1606120350
transform 1 0 23736 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_80_241
timestamp 1606120350
transform 1 0 23276 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_79_251
timestamp 1606120350
transform 1 0 24196 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_245
timestamp 1606120350
transform 1 0 23644 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_240
timestamp 1606120350
transform 1 0 23184 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__A
timestamp 1606120350
transform 1 0 23552 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__A2
timestamp 1606120350
transform 1 0 23368 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0826__A1
timestamp 1606120350
transform 1 0 24012 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_801
timestamp 1606120350
transform 1 0 23552 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _0826_
timestamp 1606120350
transform 1 0 24012 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_261
timestamp 1606120350
transform 1 0 25116 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__A2
timestamp 1606120350
transform 1 0 25576 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__A2
timestamp 1606120350
transform 1 0 25300 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_264
timestamp 1606120350
transform 1 0 25392 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_265
timestamp 1606120350
transform 1 0 25484 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0847__A1
timestamp 1606120350
transform 1 0 25944 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0913__B1
timestamp 1606120350
transform 1 0 25668 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_268
timestamp 1606120350
transform 1 0 25760 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_80_269
timestamp 1606120350
transform 1 0 25852 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__A1
timestamp 1606120350
transform 1 0 26128 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_80_274
timestamp 1606120350
transform 1 0 26312 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _0913_
timestamp 1606120350
transform 1 0 24288 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__a211o_4  _0847_
timestamp 1606120350
transform 1 0 26128 0 1 45152
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_80_280
timestamp 1606120350
transform 1 0 26864 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_276
timestamp 1606120350
transform 1 0 26496 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__B1
timestamp 1606120350
transform 1 0 27048 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__A2
timestamp 1606120350
transform 1 0 26680 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_808
timestamp 1606120350
transform 1 0 26404 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_79_290
timestamp 1606120350
transform 1 0 27784 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_286
timestamp 1606120350
transform 1 0 27416 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__A
timestamp 1606120350
transform 1 0 27968 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0888__C
timestamp 1606120350
transform 1 0 27600 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0926_
timestamp 1606120350
transform 1 0 28152 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_4  _0888_
timestamp 1606120350
transform 1 0 27232 0 -1 46240
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0926__A
timestamp 1606120350
transform 1 0 28612 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__B
timestamp 1606120350
transform 1 0 28612 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_297
timestamp 1606120350
transform 1 0 28428 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_301
timestamp 1606120350
transform 1 0 28796 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_297
timestamp 1606120350
transform 1 0 28428 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_301
timestamp 1606120350
transform 1 0 28796 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_802
timestamp 1606120350
transform 1 0 29164 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0875__A
timestamp 1606120350
transform 1 0 28980 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0891__A
timestamp 1606120350
transform 1 0 28980 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0875_
timestamp 1606120350
transform 1 0 29164 0 -1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _0891_
timestamp 1606120350
transform 1 0 29256 0 1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_80_314
timestamp 1606120350
transform 1 0 29992 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_79_315
timestamp 1606120350
transform 1 0 30084 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_79_319
timestamp 1606120350
transform 1 0 30452 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__A
timestamp 1606120350
transform 1 0 30360 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__A
timestamp 1606120350
transform 1 0 30268 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_329
timestamp 1606120350
transform 1 0 31372 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_325
timestamp 1606120350
transform 1 0 31004 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_320
timestamp 1606120350
transform 1 0 30544 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__B
timestamp 1606120350
transform 1 0 31188 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0876__A
timestamp 1606120350
transform 1 0 30636 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0895_
timestamp 1606120350
transform 1 0 30820 0 1 45152
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0876_
timestamp 1606120350
transform 1 0 30728 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_80_333
timestamp 1606120350
transform 1 0 31740 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_79_339
timestamp 1606120350
transform 1 0 32292 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_79_336
timestamp 1606120350
transform 1 0 32016 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_332
timestamp 1606120350
transform 1 0 31648 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0895__D
timestamp 1606120350
transform 1 0 31556 0 -1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0880__A
timestamp 1606120350
transform 1 0 32108 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_809
timestamp 1606120350
transform 1 0 32016 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _0880_
timestamp 1606120350
transform 1 0 32108 0 -1 46240
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0880__B
timestamp 1606120350
transform 1 0 32476 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_79_343
timestamp 1606120350
transform 1 0 32660 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_355
timestamp 1606120350
transform 1 0 33764 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_79_363
timestamp 1606120350
transform 1 0 34500 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_344
timestamp 1606120350
transform 1 0 32752 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_356
timestamp 1606120350
transform 1 0 33856 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_803
timestamp 1606120350
transform 1 0 34776 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_367
timestamp 1606120350
transform 1 0 34868 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_379
timestamp 1606120350
transform 1 0 35972 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_368
timestamp 1606120350
transform 1 0 34960 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_380
timestamp 1606120350
transform 1 0 36064 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1606120350
transform -1 0 38824 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1606120350
transform -1 0 38824 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_810
timestamp 1606120350
transform 1 0 37628 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_391
timestamp 1606120350
transform 1 0 37076 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_403
timestamp 1606120350
transform 1 0 38180 0 1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_392
timestamp 1606120350
transform 1 0 37168 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_396
timestamp 1606120350
transform 1 0 37536 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_398
timestamp 1606120350
transform 1 0 37720 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_80_406
timestamp 1606120350
transform 1 0 38456 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1192_
timestamp 1606120350
transform 1 0 1380 0 1 46240
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1606120350
transform 1 0 1104 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_22
timestamp 1606120350
transform 1 0 3128 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_34
timestamp 1606120350
transform 1 0 4232 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_811
timestamp 1606120350
transform 1 0 6716 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_46
timestamp 1606120350
transform 1 0 5336 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_81_58
timestamp 1606120350
transform 1 0 6440 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_62
timestamp 1606120350
transform 1 0 6808 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_74
timestamp 1606120350
transform 1 0 7912 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_86
timestamp 1606120350
transform 1 0 9016 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__D
timestamp 1606120350
transform 1 0 11316 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_81_98
timestamp 1606120350
transform 1 0 10120 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_81_110
timestamp 1606120350
transform 1 0 11224 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_113
timestamp 1606120350
transform 1 0 11500 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1088_
timestamp 1606120350
transform 1 0 12420 0 1 46240
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_812
timestamp 1606120350
transform 1 0 12328 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1088__D
timestamp 1606120350
transform 1 0 12144 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1092__CLK
timestamp 1606120350
transform 1 0 11684 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_81_117
timestamp 1606120350
transform 1 0 11868 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_4  _0770_
timestamp 1606120350
transform 1 0 14904 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0763__A
timestamp 1606120350
transform 1 0 14352 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0748__A
timestamp 1606120350
transform 1 0 14720 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_142
timestamp 1606120350
transform 1 0 14168 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_146
timestamp 1606120350
transform 1 0 14536 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__D
timestamp 1606120350
transform 1 0 16652 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__A2
timestamp 1606120350
transform 1 0 16192 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1211__CLK
timestamp 1606120350
transform 1 0 17020 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_162
timestamp 1606120350
transform 1 0 16008 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_81_166
timestamp 1606120350
transform 1 0 16376 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_81_171
timestamp 1606120350
transform 1 0 16836 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_175
timestamp 1606120350
transform 1 0 17204 0 1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_813
timestamp 1606120350
transform 1 0 17940 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1059__A
timestamp 1606120350
transform 1 0 19780 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_81_184
timestamp 1606120350
transform 1 0 18032 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_196
timestamp 1606120350
transform 1 0 19136 0 1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_202
timestamp 1606120350
transform 1 0 19688 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_205
timestamp 1606120350
transform 1 0 19964 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_212
timestamp 1606120350
transform 1 0 20608 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_81_209
timestamp 1606120350
transform 1 0 20332 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0998__A
timestamp 1606120350
transform 1 0 20424 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0885__A
timestamp 1606120350
transform 1 0 20792 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_223
timestamp 1606120350
transform 1 0 21620 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_219
timestamp 1606120350
transform 1 0 21252 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__A
timestamp 1606120350
transform 1 0 21436 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0837__B
timestamp 1606120350
transform 1 0 21804 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0998_
timestamp 1606120350
transform 1 0 20976 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _0841_
timestamp 1606120350
transform 1 0 21988 0 1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  _0834_
timestamp 1606120350
transform 1 0 23920 0 1 46240
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_814
timestamp 1606120350
transform 1 0 23552 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__B
timestamp 1606120350
transform 1 0 23368 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0834__A
timestamp 1606120350
transform 1 0 23000 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_236
timestamp 1606120350
transform 1 0 22816 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_240
timestamp 1606120350
transform 1 0 23184 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_81_245
timestamp 1606120350
transform 1 0 23644 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _0860_
timestamp 1606120350
transform 1 0 26128 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__B1
timestamp 1606120350
transform 1 0 25944 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__B1
timestamp 1606120350
transform 1 0 25576 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0858__A
timestamp 1606120350
transform 1 0 25208 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_257
timestamp 1606120350
transform 1 0 24748 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_261
timestamp 1606120350
transform 1 0 25116 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_264
timestamp 1606120350
transform 1 0 25392 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_268
timestamp 1606120350
transform 1 0 25760 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0932_
timestamp 1606120350
transform 1 0 28152 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__C1
timestamp 1606120350
transform 1 0 27416 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0932__A
timestamp 1606120350
transform 1 0 27968 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_284
timestamp 1606120350
transform 1 0 27232 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_288
timestamp 1606120350
transform 1 0 27600 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1183_
timestamp 1606120350
transform 1 0 29808 0 1 46240
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_815
timestamp 1606120350
transform 1 0 29164 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__D
timestamp 1606120350
transform 1 0 29624 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__A1
timestamp 1606120350
transform 1 0 28612 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0921__A2
timestamp 1606120350
transform 1 0 28980 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_297
timestamp 1606120350
transform 1 0 28428 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_301
timestamp 1606120350
transform 1 0 28796 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_306
timestamp 1606120350
transform 1 0 29256 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0907__A
timestamp 1606120350
transform 1 0 32108 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__B
timestamp 1606120350
transform 1 0 31740 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__D
timestamp 1606120350
transform 1 0 32476 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_331
timestamp 1606120350
transform 1 0 31556 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_335
timestamp 1606120350
transform 1 0 31924 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_339
timestamp 1606120350
transform 1 0 32292 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1183__CLK
timestamp 1606120350
transform 1 0 32844 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_81_343
timestamp 1606120350
transform 1 0 32660 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_81_347
timestamp 1606120350
transform 1 0 33028 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_359
timestamp 1606120350
transform 1 0 34132 0 1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_365
timestamp 1606120350
transform 1 0 34684 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_816
timestamp 1606120350
transform 1 0 34776 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_367
timestamp 1606120350
transform 1 0 34868 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_379
timestamp 1606120350
transform 1 0 35972 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1606120350
transform -1 0 38824 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_391
timestamp 1606120350
transform 1 0 37076 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_403
timestamp 1606120350
transform 1 0 38180 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1606120350
transform 1 0 1104 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1192__CLK
timestamp 1606120350
transform 1 0 1564 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_3
timestamp 1606120350
transform 1 0 1380 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_7
timestamp 1606120350
transform 1 0 1748 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_19
timestamp 1606120350
transform 1 0 2852 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_817
timestamp 1606120350
transform 1 0 3956 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_32
timestamp 1606120350
transform 1 0 4048 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_44
timestamp 1606120350
transform 1 0 5152 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_56
timestamp 1606120350
transform 1 0 6256 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_68
timestamp 1606120350
transform 1 0 7360 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_80
timestamp 1606120350
transform 1 0 8464 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1092_
timestamp 1606120350
transform 1 0 11316 0 -1 47328
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_818
timestamp 1606120350
transform 1 0 9568 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_93
timestamp 1606120350
transform 1 0 9660 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_105
timestamp 1606120350
transform 1 0 10764 0 -1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__B1
timestamp 1606120350
transform 1 0 13248 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__A2
timestamp 1606120350
transform 1 0 13616 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_130
timestamp 1606120350
transform 1 0 13064 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_134
timestamp 1606120350
transform 1 0 13432 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0748_
timestamp 1606120350
transform 1 0 15272 0 -1 47328
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _0763_
timestamp 1606120350
transform 1 0 13800 0 -1 47328
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_819
timestamp 1606120350
transform 1 0 15180 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0770__B1
timestamp 1606120350
transform 1 0 14904 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_145
timestamp 1606120350
transform 1 0 14444 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_149
timestamp 1606120350
transform 1 0 14812 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_82_152
timestamp 1606120350
transform 1 0 15088 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1211_
timestamp 1606120350
transform 1 0 16652 0 -1 47328
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__B1
timestamp 1606120350
transform 1 0 16100 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_161
timestamp 1606120350
transform 1 0 15916 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_165
timestamp 1606120350
transform 1 0 16284 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1059_
timestamp 1606120350
transform 1 0 19780 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_188
timestamp 1606120350
transform 1 0 18400 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_200
timestamp 1606120350
transform 1 0 19504 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_82_215
timestamp 1606120350
transform 1 0 20884 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_210
timestamp 1606120350
transform 1 0 20424 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_206
timestamp 1606120350
transform 1 0 20056 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_1_1_0_clk_A
timestamp 1606120350
transform 1 0 20240 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__D
timestamp 1606120350
transform 1 0 20608 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_820
timestamp 1606120350
transform 1 0 20792 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_223
timestamp 1606120350
transform 1 0 21620 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_219
timestamp 1606120350
transform 1 0 21252 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__B
timestamp 1606120350
transform 1 0 21436 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0841__C
timestamp 1606120350
transform 1 0 21804 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0885_
timestamp 1606120350
transform 1 0 20976 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _0837_
timestamp 1606120350
transform 1 0 21988 0 -1 47328
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0943_
timestamp 1606120350
transform 1 0 23552 0 -1 47328
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__A
timestamp 1606120350
transform 1 0 23000 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__B
timestamp 1606120350
transform 1 0 23368 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_236
timestamp 1606120350
transform 1 0 22816 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_240
timestamp 1606120350
transform 1 0 23184 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_253
timestamp 1606120350
transform 1 0 24380 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__A
timestamp 1606120350
transform 1 0 24564 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_257
timestamp 1606120350
transform 1 0 24748 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_261
timestamp 1606120350
transform 1 0 25116 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0943__C
timestamp 1606120350
transform 1 0 24932 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0858_
timestamp 1606120350
transform 1 0 25208 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_82_265
timestamp 1606120350
transform 1 0 25484 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_82_269
timestamp 1606120350
transform 1 0 25852 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__C
timestamp 1606120350
transform 1 0 25668 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_274
timestamp 1606120350
transform 1 0 26312 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0860__A2
timestamp 1606120350
transform 1 0 26128 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _0853_
timestamp 1606120350
transform 1 0 26496 0 -1 47328
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_821
timestamp 1606120350
transform 1 0 26404 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__B1
timestamp 1606120350
transform 1 0 27968 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__B
timestamp 1606120350
transform 1 0 28336 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_290
timestamp 1606120350
transform 1 0 27784 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_294
timestamp 1606120350
transform 1 0 28152 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0887_
timestamp 1606120350
transform 1 0 30360 0 -1 47328
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_4  _0921_
timestamp 1606120350
transform 1 0 28520 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0887__C
timestamp 1606120350
transform 1 0 30176 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__B
timestamp 1606120350
transform 1 0 29808 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_310
timestamp 1606120350
transform 1 0 29624 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_314
timestamp 1606120350
transform 1 0 29992 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0907_
timestamp 1606120350
transform 1 0 32108 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_822
timestamp 1606120350
transform 1 0 32016 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__A1
timestamp 1606120350
transform 1 0 31372 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0853__A1
timestamp 1606120350
transform 1 0 31740 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_327
timestamp 1606120350
transform 1 0 31188 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_82_331
timestamp 1606120350
transform 1 0 31556 0 -1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_82_335
timestamp 1606120350
transform 1 0 31924 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_340
timestamp 1606120350
transform 1 0 32384 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_352
timestamp 1606120350
transform 1 0 33488 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_364
timestamp 1606120350
transform 1 0 34592 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_376
timestamp 1606120350
transform 1 0 35696 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_388
timestamp 1606120350
transform 1 0 36800 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1606120350
transform -1 0 38824 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_823
timestamp 1606120350
transform 1 0 37628 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_82_396
timestamp 1606120350
transform 1 0 37536 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_398
timestamp 1606120350
transform 1 0 37720 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_406
timestamp 1606120350
transform 1 0 38456 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1606120350
transform 1 0 1104 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_3
timestamp 1606120350
transform 1 0 1380 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_15
timestamp 1606120350
transform 1 0 2484 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_27
timestamp 1606120350
transform 1 0 3588 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_39
timestamp 1606120350
transform 1 0 4692 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_824
timestamp 1606120350
transform 1 0 6716 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_51
timestamp 1606120350
transform 1 0 5796 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_59
timestamp 1606120350
transform 1 0 6532 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_83_62
timestamp 1606120350
transform 1 0 6808 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_74
timestamp 1606120350
transform 1 0 7912 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_86
timestamp 1606120350
transform 1 0 9016 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__B1
timestamp 1606120350
transform 1 0 11592 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__A1
timestamp 1606120350
transform 1 0 11224 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__B2
timestamp 1606120350
transform 1 0 10856 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_83_98
timestamp 1606120350
transform 1 0 10120 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_108
timestamp 1606120350
transform 1 0 11040 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_112
timestamp 1606120350
transform 1 0 11408 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0764_
timestamp 1606120350
transform 1 0 12512 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_825
timestamp 1606120350
transform 1 0 12328 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0764__A1
timestamp 1606120350
transform 1 0 12144 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_83_116
timestamp 1606120350
transform 1 0 11776 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_123
timestamp 1606120350
transform 1 0 12420 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_136
timestamp 1606120350
transform 1 0 13616 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1086_
timestamp 1606120350
transform 1 0 14352 0 1 47328
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__A
timestamp 1606120350
transform 1 0 13800 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0733__B
timestamp 1606120350
transform 1 0 14168 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_140
timestamp 1606120350
transform 1 0 13984 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0663_
timestamp 1606120350
transform 1 0 16836 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0663__A
timestamp 1606120350
transform 1 0 17296 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A1
timestamp 1606120350
transform 1 0 16284 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0749__A2
timestamp 1606120350
transform 1 0 16652 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_163
timestamp 1606120350
transform 1 0 16100 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_167
timestamp 1606120350
transform 1 0 16468 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_174
timestamp 1606120350
transform 1 0 17112 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_83_178
timestamp 1606120350
transform 1 0 17480 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_182
timestamp 1606120350
transform 1 0 17848 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_184
timestamp 1606120350
transform 1 0 18032 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_826
timestamp 1606120350
transform 1 0 17940 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_83_191
timestamp 1606120350
transform 1 0 18676 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_83_188
timestamp 1606120350
transform 1 0 18400 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__B1
timestamp 1606120350
transform 1 0 18492 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_195
timestamp 1606120350
transform 1 0 19044 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__A2
timestamp 1606120350
transform 1 0 19228 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1068__A1
timestamp 1606120350
transform 1 0 18860 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_202
timestamp 1606120350
transform 1 0 19688 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0842_
timestamp 1606120350
transform 1 0 19412 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0842__A
timestamp 1606120350
transform 1 0 19872 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0836_
timestamp 1606120350
transform 1 0 21988 0 1 47328
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  _0878_
timestamp 1606120350
transform 1 0 20424 0 1 47328
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0836__A
timestamp 1606120350
transform 1 0 21804 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0878__A
timestamp 1606120350
transform 1 0 20240 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1026__A
timestamp 1606120350
transform 1 0 21436 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_206
timestamp 1606120350
transform 1 0 20056 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_219
timestamp 1606120350
transform 1 0 21252 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_223
timestamp 1606120350
transform 1 0 21620 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _0958_
timestamp 1606120350
transform 1 0 23644 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_827
timestamp 1606120350
transform 1 0 23552 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1042__C
timestamp 1606120350
transform 1 0 23368 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__A1
timestamp 1606120350
transform 1 0 23000 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_236
timestamp 1606120350
transform 1 0 22816 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_240
timestamp 1606120350
transform 1 0 23184 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0912_
timestamp 1606120350
transform 1 0 25484 0 1 47328
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__A2
timestamp 1606120350
transform 1 0 24932 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__A
timestamp 1606120350
transform 1 0 25300 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_257
timestamp 1606120350
transform 1 0 24748 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_261
timestamp 1606120350
transform 1 0 25116 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_274
timestamp 1606120350
transform 1 0 26312 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0892_
timestamp 1606120350
transform 1 0 27232 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__B1
timestamp 1606120350
transform 1 0 26496 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0865__A2
timestamp 1606120350
transform 1 0 26864 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_278
timestamp 1606120350
transform 1 0 26680 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_282
timestamp 1606120350
transform 1 0 27048 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_296
timestamp 1606120350
transform 1 0 28336 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0893_
timestamp 1606120350
transform 1 0 29256 0 1 47328
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_828
timestamp 1606120350
transform 1 0 29164 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0918__A
timestamp 1606120350
transform 1 0 28520 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0893__A
timestamp 1606120350
transform 1 0 28980 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__B
timestamp 1606120350
transform 1 0 30268 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_83_300
timestamp 1606120350
transform 1 0 28704 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_83_315
timestamp 1606120350
transform 1 0 30084 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_319
timestamp 1606120350
transform 1 0 30452 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0833_
timestamp 1606120350
transform 1 0 32200 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _0852_
timestamp 1606120350
transform 1 0 30820 0 1 47328
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__B
timestamp 1606120350
transform 1 0 31648 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__D
timestamp 1606120350
transform 1 0 30636 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_83_330
timestamp 1606120350
transform 1 0 31464 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_83_334
timestamp 1606120350
transform 1 0 31832 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_83_341
timestamp 1606120350
transform 1 0 32476 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0833__A
timestamp 1606120350
transform 1 0 32660 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_83_345
timestamp 1606120350
transform 1 0 32844 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_357
timestamp 1606120350
transform 1 0 33948 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_365
timestamp 1606120350
transform 1 0 34684 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_829
timestamp 1606120350
transform 1 0 34776 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_367
timestamp 1606120350
transform 1 0 34868 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_379
timestamp 1606120350
transform 1 0 35972 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1606120350
transform -1 0 38824 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_391
timestamp 1606120350
transform 1 0 37076 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_403
timestamp 1606120350
transform 1 0 38180 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1606120350
transform 1 0 1104 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_3
timestamp 1606120350
transform 1 0 1380 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_15
timestamp 1606120350
transform 1 0 2484 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_830
timestamp 1606120350
transform 1 0 3956 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_27
timestamp 1606120350
transform 1 0 3588 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_32
timestamp 1606120350
transform 1 0 4048 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_44
timestamp 1606120350
transform 1 0 5152 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_56
timestamp 1606120350
transform 1 0 6256 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_68
timestamp 1606120350
transform 1 0 7360 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_80
timestamp 1606120350
transform 1 0 8464 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__o22a_4  _0782_
timestamp 1606120350
transform 1 0 11592 0 -1 48416
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_831
timestamp 1606120350
transform 1 0 9568 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0782__A2
timestamp 1606120350
transform 1 0 11408 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_84_93
timestamp 1606120350
transform 1 0 9660 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_105
timestamp 1606120350
transform 1 0 10764 0 -1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_111
timestamp 1606120350
transform 1 0 11316 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__B1
timestamp 1606120350
transform 1 0 13248 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__A2
timestamp 1606120350
transform 1 0 13616 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_128
timestamp 1606120350
transform 1 0 12880 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_84_134
timestamp 1606120350
transform 1 0 13432 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0733_
timestamp 1606120350
transform 1 0 13800 0 -1 48416
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_4  _0749_
timestamp 1606120350
transform 1 0 15272 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_832
timestamp 1606120350
transform 1 0 15180 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__D
timestamp 1606120350
transform 1 0 14628 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1086__CLK
timestamp 1606120350
transform 1 0 14996 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_145
timestamp 1606120350
transform 1 0 14444 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_149
timestamp 1606120350
transform 1 0 14812 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__B1
timestamp 1606120350
transform 1 0 17848 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_84_166
timestamp 1606120350
transform 1 0 16376 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_178
timestamp 1606120350
transform 1 0 17480 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1068_
timestamp 1606120350
transform 1 0 18860 0 -1 48416
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__B1
timestamp 1606120350
transform 1 0 18676 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__B1
timestamp 1606120350
transform 1 0 18308 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_84_184
timestamp 1606120350
transform 1 0 18032 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_84_189
timestamp 1606120350
transform 1 0 18492 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _1026_
timestamp 1606120350
transform 1 0 20884 0 -1 48416
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_833
timestamp 1606120350
transform 1 0 20792 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__B1
timestamp 1606120350
transform 1 0 21896 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__B
timestamp 1606120350
transform 1 0 20516 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_206
timestamp 1606120350
transform 1 0 20056 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_210
timestamp 1606120350
transform 1 0 20424 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_84_213
timestamp 1606120350
transform 1 0 20700 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_84_224
timestamp 1606120350
transform 1 0 21712 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_228
timestamp 1606120350
transform 1 0 22080 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0838_
timestamp 1606120350
transform 1 0 22448 0 -1 48416
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_4  _1042_
timestamp 1606120350
transform 1 0 23828 0 -1 48416
box -38 -48 1602 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0958__B1
timestamp 1606120350
transform 1 0 23644 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0838__B
timestamp 1606120350
transform 1 0 23276 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__A2
timestamp 1606120350
transform 1 0 22264 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_239
timestamp 1606120350
transform 1 0 23092 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_243
timestamp 1606120350
transform 1 0 23460 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A2
timestamp 1606120350
transform 1 0 26220 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0912__B
timestamp 1606120350
transform 1 0 25576 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_264
timestamp 1606120350
transform 1 0 25392 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_268
timestamp 1606120350
transform 1 0 25760 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_272
timestamp 1606120350
transform 1 0 26128 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__a21o_4  _0865_
timestamp 1606120350
transform 1 0 26496 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _0918_
timestamp 1606120350
transform 1 0 28336 0 -1 48416
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_834
timestamp 1606120350
transform 1 0 26404 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0884__A
timestamp 1606120350
transform 1 0 28152 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__A2
timestamp 1606120350
transform 1 0 27784 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_288
timestamp 1606120350
transform 1 0 27600 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_292
timestamp 1606120350
transform 1 0 27968 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__and2_4  _0920_
timestamp 1606120350
transform 1 0 29900 0 -1 48416
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__A1
timestamp 1606120350
transform 1 0 29348 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__B1
timestamp 1606120350
transform 1 0 29716 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_305
timestamp 1606120350
transform 1 0 29164 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_309
timestamp 1606120350
transform 1 0 29532 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_835
timestamp 1606120350
transform 1 0 32016 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0920__A
timestamp 1606120350
transform 1 0 30728 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0892__A1
timestamp 1606120350
transform 1 0 31096 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0852__A
timestamp 1606120350
transform 1 0 31464 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_320
timestamp 1606120350
transform 1 0 30544 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_324
timestamp 1606120350
transform 1 0 30912 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_84_328
timestamp 1606120350
transform 1 0 31280 0 -1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_332
timestamp 1606120350
transform 1 0 31648 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_84_337
timestamp 1606120350
transform 1 0 32108 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_349
timestamp 1606120350
transform 1 0 33212 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_361
timestamp 1606120350
transform 1 0 34316 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_373
timestamp 1606120350
transform 1 0 35420 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_385
timestamp 1606120350
transform 1 0 36524 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1606120350
transform -1 0 38824 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_836
timestamp 1606120350
transform 1 0 37628 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_398
timestamp 1606120350
transform 1 0 37720 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_406
timestamp 1606120350
transform 1 0 38456 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1606120350
transform 1 0 1104 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1606120350
transform 1 0 1104 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_85_3
timestamp 1606120350
transform 1 0 1380 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_15
timestamp 1606120350
transform 1 0 2484 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_3
timestamp 1606120350
transform 1 0 1380 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_15
timestamp 1606120350
transform 1 0 2484 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_843
timestamp 1606120350
transform 1 0 3956 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_27
timestamp 1606120350
transform 1 0 3588 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_39
timestamp 1606120350
transform 1 0 4692 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_27
timestamp 1606120350
transform 1 0 3588 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_32
timestamp 1606120350
transform 1 0 4048 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_44
timestamp 1606120350
transform 1 0 5152 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_837
timestamp 1606120350
transform 1 0 6716 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_85_51
timestamp 1606120350
transform 1 0 5796 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_85_59
timestamp 1606120350
transform 1 0 6532 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_85_62
timestamp 1606120350
transform 1 0 6808 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_56
timestamp 1606120350
transform 1 0 6256 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_68
timestamp 1606120350
transform 1 0 7360 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_74
timestamp 1606120350
transform 1 0 7912 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_86
timestamp 1606120350
transform 1 0 9016 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_80
timestamp 1606120350
transform 1 0 8464 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_844
timestamp 1606120350
transform 1 0 9568 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_98
timestamp 1606120350
transform 1 0 10120 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_110
timestamp 1606120350
transform 1 0 11224 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_93
timestamp 1606120350
transform 1 0 9660 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_105
timestamp 1606120350
transform 1 0 10764 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_85_123
timestamp 1606120350
transform 1 0 12420 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_838
timestamp 1606120350
transform 1 0 12328 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_86_129
timestamp 1606120350
transform 1 0 12972 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_85_128
timestamp 1606120350
transform 1 0 12880 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__CLK
timestamp 1606120350
transform 1 0 13064 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1085__D
timestamp 1606120350
transform 1 0 12696 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0734__A1
timestamp 1606120350
transform 1 0 13064 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_86_117
timestamp 1606120350
transform 1 0 11868 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1085_
timestamp 1606120350
transform 1 0 13248 0 1 48416
box -38 -48 1786 592
use sky130_fd_sc_hd__a21o_4  _0734_
timestamp 1606120350
transform 1 0 13248 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_86_144
timestamp 1606120350
transform 1 0 14352 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__CLK
timestamp 1606120350
transform 1 0 14628 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_86_154
timestamp 1606120350
transform 1 0 15272 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_86_149
timestamp 1606120350
transform 1 0 14812 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_157
timestamp 1606120350
transform 1 0 15548 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_85_151
timestamp 1606120350
transform 1 0 14996 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1172__CLK
timestamp 1606120350
transform 1 0 15732 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1114__D
timestamp 1606120350
transform 1 0 14996 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1172__D
timestamp 1606120350
transform 1 0 15364 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_845
timestamp 1606120350
transform 1 0 15180 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1172_
timestamp 1606120350
transform 1 0 15364 0 -1 49504
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_2  FILLER_86_178
timestamp 1606120350
transform 1 0 17480 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_174
timestamp 1606120350
transform 1 0 17112 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_179
timestamp 1606120350
transform 1 0 17572 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_175
timestamp 1606120350
transform 1 0 17204 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__B1
timestamp 1606120350
transform 1 0 17020 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__A2
timestamp 1606120350
transform 1 0 17296 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__A2
timestamp 1606120350
transform 1 0 17388 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__A2
timestamp 1606120350
transform 1 0 17664 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1081__A1
timestamp 1606120350
transform 1 0 17756 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_85_161
timestamp 1606120350
transform 1 0 15916 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_4  _1081_
timestamp 1606120350
transform 1 0 17848 0 -1 49504
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_85_191
timestamp 1606120350
transform 1 0 18676 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_187
timestamp 1606120350
transform 1 0 18308 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__A1
timestamp 1606120350
transform 1 0 18860 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0984__A
timestamp 1606120350
transform 1 0 18492 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_839
timestamp 1606120350
transform 1 0 17940 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0984_
timestamp 1606120350
transform 1 0 18032 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_86_199
timestamp 1606120350
transform 1 0 19412 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_195
timestamp 1606120350
transform 1 0 19044 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__A2
timestamp 1606120350
transform 1 0 19596 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1069__A2
timestamp 1606120350
transform 1 0 19228 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1044_
timestamp 1606120350
transform 1 0 19780 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _1069_
timestamp 1606120350
transform 1 0 19044 0 1 48416
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__B1
timestamp 1606120350
transform 1 0 20240 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_208
timestamp 1606120350
transform 1 0 20240 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_206
timestamp 1606120350
transform 1 0 20056 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1044__A
timestamp 1606120350
transform 1 0 20424 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__A
timestamp 1606120350
transform 1 0 20608 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_212
timestamp 1606120350
transform 1 0 20608 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_210
timestamp 1606120350
transform 1 0 20424 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_846
timestamp 1606120350
transform 1 0 20792 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_clk
timestamp 1606120350
transform 1 0 20976 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__A1
timestamp 1606120350
transform 1 0 20792 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_86_215
timestamp 1606120350
transform 1 0 20884 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_86_220
timestamp 1606120350
transform 1 0 21344 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_219
timestamp 1606120350
transform 1 0 21252 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__A1
timestamp 1606120350
transform 1 0 21160 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__B1
timestamp 1606120350
transform 1 0 21528 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1047__A2
timestamp 1606120350
transform 1 0 21436 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _1047_
timestamp 1606120350
transform 1 0 21712 0 -1 49504
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _1013_
timestamp 1606120350
transform 1 0 21620 0 1 48416
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_86_237
timestamp 1606120350
transform 1 0 22908 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_236
timestamp 1606120350
transform 1 0 22816 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1013__B1
timestamp 1606120350
transform 1 0 23092 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__A1
timestamp 1606120350
transform 1 0 23000 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_241
timestamp 1606120350
transform 1 0 23276 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_249
timestamp 1606120350
transform 1 0 24012 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_85_245
timestamp 1606120350
transform 1 0 23644 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_85_240
timestamp 1606120350
transform 1 0 23184 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__B1
timestamp 1606120350
transform 1 0 23460 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__C
timestamp 1606120350
transform 1 0 23368 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0882__A
timestamp 1606120350
transform 1 0 24196 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_840
timestamp 1606120350
transform 1 0 23552 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0882_
timestamp 1606120350
transform 1 0 23736 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _1016_
timestamp 1606120350
transform 1 0 23644 0 -1 49504
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_86_262
timestamp 1606120350
transform 1 0 25208 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_258
timestamp 1606120350
transform 1 0 24840 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_253
timestamp 1606120350
transform 1 0 24380 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__B
timestamp 1606120350
transform 1 0 25024 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__A
timestamp 1606120350
transform 1 0 24564 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0916_
timestamp 1606120350
transform 1 0 24748 0 1 48416
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  FILLER_86_270
timestamp 1606120350
transform 1 0 25944 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_86_266
timestamp 1606120350
transform 1 0 25576 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_270
timestamp 1606120350
transform 1 0 25944 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_266
timestamp 1606120350
transform 1 0 25576 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__B1
timestamp 1606120350
transform 1 0 26220 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__C
timestamp 1606120350
transform 1 0 25760 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__B
timestamp 1606120350
transform 1 0 25392 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__A
timestamp 1606120350
transform 1 0 25760 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0859__B
timestamp 1606120350
transform 1 0 26128 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0917_
timestamp 1606120350
transform 1 0 26312 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_86_283
timestamp 1606120350
transform 1 0 27140 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_847
timestamp 1606120350
transform 1 0 26404 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _0859_
timestamp 1606120350
transform 1 0 26496 0 -1 49504
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_86_288
timestamp 1606120350
transform 1 0 27600 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_290
timestamp 1606120350
transform 1 0 27784 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_286
timestamp 1606120350
transform 1 0 27416 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__B1_N
timestamp 1606120350
transform 1 0 27784 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__A2
timestamp 1606120350
transform 1 0 27416 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A1
timestamp 1606120350
transform 1 0 27600 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__A2
timestamp 1606120350
transform 1 0 27968 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0884_
timestamp 1606120350
transform 1 0 28152 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _0873_
timestamp 1606120350
transform 1 0 27968 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_308
timestamp 1606120350
transform 1 0 29440 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_304
timestamp 1606120350
transform 1 0 29072 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_85_301
timestamp 1606120350
transform 1 0 28796 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_297
timestamp 1606120350
transform 1 0 28428 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0873__B1
timestamp 1606120350
transform 1 0 28612 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0874__A2
timestamp 1606120350
transform 1 0 28980 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_841
timestamp 1606120350
transform 1 0 29164 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_86_311
timestamp 1606120350
transform 1 0 29716 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_85_319
timestamp 1606120350
transform 1 0 30452 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__D
timestamp 1606120350
transform 1 0 29532 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0872_
timestamp 1606120350
transform 1 0 29808 0 -1 49504
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _0874_
timestamp 1606120350
transform 1 0 29256 0 1 48416
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0916__D
timestamp 1606120350
transform 1 0 30636 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__A1
timestamp 1606120350
transform 1 0 30820 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0917__A1
timestamp 1606120350
transform 1 0 31004 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_323
timestamp 1606120350
transform 1 0 30820 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_321
timestamp 1606120350
transform 1 0 30636 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_325
timestamp 1606120350
transform 1 0 31004 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0886_
timestamp 1606120350
transform 1 0 31188 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0872__A
timestamp 1606120350
transform 1 0 31188 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_85_330
timestamp 1606120350
transform 1 0 31464 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_86_329
timestamp 1606120350
transform 1 0 31372 0 -1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_335
timestamp 1606120350
transform 1 0 31924 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0886__A
timestamp 1606120350
transform 1 0 31648 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_848
timestamp 1606120350
transform 1 0 32016 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_337
timestamp 1606120350
transform 1 0 32108 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_334
timestamp 1606120350
transform 1 0 31832 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_346
timestamp 1606120350
transform 1 0 32936 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_358
timestamp 1606120350
transform 1 0 34040 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_349
timestamp 1606120350
transform 1 0 33212 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_361
timestamp 1606120350
transform 1 0 34316 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_842
timestamp 1606120350
transform 1 0 34776 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_367
timestamp 1606120350
transform 1 0 34868 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_379
timestamp 1606120350
transform 1 0 35972 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_373
timestamp 1606120350
transform 1 0 35420 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_385
timestamp 1606120350
transform 1 0 36524 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1606120350
transform -1 0 38824 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1606120350
transform -1 0 38824 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_849
timestamp 1606120350
transform 1 0 37628 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_391
timestamp 1606120350
transform 1 0 37076 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_85_403
timestamp 1606120350
transform 1 0 38180 0 1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_398
timestamp 1606120350
transform 1 0 37720 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_406
timestamp 1606120350
transform 1 0 38456 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1606120350
transform 1 0 1104 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_87_3
timestamp 1606120350
transform 1 0 1380 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_15
timestamp 1606120350
transform 1 0 2484 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_27
timestamp 1606120350
transform 1 0 3588 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_39
timestamp 1606120350
transform 1 0 4692 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_850
timestamp 1606120350
transform 1 0 6716 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_87_51
timestamp 1606120350
transform 1 0 5796 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_87_59
timestamp 1606120350
transform 1 0 6532 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_87_62
timestamp 1606120350
transform 1 0 6808 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_74
timestamp 1606120350
transform 1 0 7912 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_86
timestamp 1606120350
transform 1 0 9016 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_98
timestamp 1606120350
transform 1 0 10120 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_110
timestamp 1606120350
transform 1 0 11224 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_851
timestamp 1606120350
transform 1 0 12328 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_123
timestamp 1606120350
transform 1 0 12420 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_87_135
timestamp 1606120350
transform 1 0 13524 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _0821_
timestamp 1606120350
transform 1 0 15272 0 1 49504
box -38 -48 1326 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__A1
timestamp 1606120350
transform 1 0 15088 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__B2
timestamp 1606120350
transform 1 0 14720 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__A2
timestamp 1606120350
transform 1 0 14352 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_87_143
timestamp 1606120350
transform 1 0 14260 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_87_146
timestamp 1606120350
transform 1 0 14536 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_150
timestamp 1606120350
transform 1 0 14904 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__A1
timestamp 1606120350
transform 1 0 17756 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1041__B1
timestamp 1606120350
transform 1 0 17388 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__B1
timestamp 1606120350
transform 1 0 17020 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_87_168
timestamp 1606120350
transform 1 0 16560 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_87_172
timestamp 1606120350
transform 1 0 16928 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_87_175
timestamp 1606120350
transform 1 0 17204 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_179
timestamp 1606120350
transform 1 0 17572 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _1038_
timestamp 1606120350
transform 1 0 19964 0 1 49504
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _1041_
timestamp 1606120350
transform 1 0 18032 0 1 49504
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_852
timestamp 1606120350
transform 1 0 17940 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A1
timestamp 1606120350
transform 1 0 19780 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1080__A1
timestamp 1606120350
transform 1 0 19412 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_197
timestamp 1606120350
transform 1 0 19228 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_201
timestamp 1606120350
transform 1 0 19596 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _1036_
timestamp 1606120350
transform 1 0 21896 0 1 49504
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__A2
timestamp 1606120350
transform 1 0 21712 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0959__A1
timestamp 1606120350
transform 1 0 21344 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_218
timestamp 1606120350
transform 1 0 21160 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_222
timestamp 1606120350
transform 1 0 21528 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__or3_4  _0835_
timestamp 1606120350
transform 1 0 23828 0 1 49504
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_853
timestamp 1606120350
transform 1 0 23552 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__A
timestamp 1606120350
transform 1 0 23368 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__C
timestamp 1606120350
transform 1 0 23000 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_87_235
timestamp 1606120350
transform 1 0 22724 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_87_240
timestamp 1606120350
transform 1 0 23184 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_245
timestamp 1606120350
transform 1 0 23644 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0908_
timestamp 1606120350
transform 1 0 25392 0 1 49504
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0835__B
timestamp 1606120350
transform 1 0 24840 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__A
timestamp 1606120350
transform 1 0 25208 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_256
timestamp 1606120350
transform 1 0 24656 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_260
timestamp 1606120350
transform 1 0 25024 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_273
timestamp 1606120350
transform 1 0 26220 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0900_
timestamp 1606120350
transform 1 0 27048 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__A2
timestamp 1606120350
transform 1 0 26864 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__B1
timestamp 1606120350
transform 1 0 26404 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0902__A1
timestamp 1606120350
transform 1 0 28336 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_87_277
timestamp 1606120350
transform 1 0 26588 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_87_294
timestamp 1606120350
transform 1 0 28152 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__a21bo_4  _0930_
timestamp 1606120350
transform 1 0 29256 0 1 49504
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_854
timestamp 1606120350
transform 1 0 29164 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_12_0_clk
timestamp 1606120350
transform 1 0 28888 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__A2
timestamp 1606120350
transform 1 0 28704 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_298
timestamp 1606120350
transform 1 0 28520 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_319
timestamp 1606120350
transform 1 0 30452 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0843_
timestamp 1606120350
transform 1 0 31188 0 1 49504
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0843__A
timestamp 1606120350
transform 1 0 31004 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0908__D
timestamp 1606120350
transform 1 0 30636 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1194__CLK
timestamp 1606120350
transform 1 0 32200 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_323
timestamp 1606120350
transform 1 0 30820 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_87_336
timestamp 1606120350
transform 1 0 32016 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_87_340
timestamp 1606120350
transform 1 0 32384 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_352
timestamp 1606120350
transform 1 0 33488 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_87_364
timestamp 1606120350
transform 1 0 34592 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_855
timestamp 1606120350
transform 1 0 34776 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_367
timestamp 1606120350
transform 1 0 34868 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_379
timestamp 1606120350
transform 1 0 35972 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1606120350
transform -1 0 38824 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_87_391
timestamp 1606120350
transform 1 0 37076 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_87_403
timestamp 1606120350
transform 1 0 38180 0 1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1606120350
transform 1 0 1104 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_88_3
timestamp 1606120350
transform 1 0 1380 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_15
timestamp 1606120350
transform 1 0 2484 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_856
timestamp 1606120350
transform 1 0 3956 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_88_27
timestamp 1606120350
transform 1 0 3588 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_88_32
timestamp 1606120350
transform 1 0 4048 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_44
timestamp 1606120350
transform 1 0 5152 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_56
timestamp 1606120350
transform 1 0 6256 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_68
timestamp 1606120350
transform 1 0 7360 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_80
timestamp 1606120350
transform 1 0 8464 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_857
timestamp 1606120350
transform 1 0 9568 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_93
timestamp 1606120350
transform 1 0 9660 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_105
timestamp 1606120350
transform 1 0 10764 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_117
timestamp 1606120350
transform 1 0 11868 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_129
timestamp 1606120350
transform 1 0 12972 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1114_
timestamp 1606120350
transform 1 0 15272 0 -1 50592
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_858
timestamp 1606120350
transform 1 0 15180 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0821__B1
timestamp 1606120350
transform 1 0 14996 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_88_141
timestamp 1606120350
transform 1 0 14076 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_88_149
timestamp 1606120350
transform 1 0 14812 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A2
timestamp 1606120350
transform 1 0 17204 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__B1
timestamp 1606120350
transform 1 0 17572 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_173
timestamp 1606120350
transform 1 0 17020 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_177
timestamp 1606120350
transform 1 0 17388 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_88_181
timestamp 1606120350
transform 1 0 17756 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _1080_
timestamp 1606120350
transform 1 0 18400 0 -1 50592
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__B1
timestamp 1606120350
transform 1 0 18032 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1038__A2
timestamp 1606120350
transform 1 0 19964 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_186
timestamp 1606120350
transform 1 0 18216 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_88_201
timestamp 1606120350
transform 1 0 19596 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _0959_
timestamp 1606120350
transform 1 0 21712 0 -1 50592
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_859
timestamp 1606120350
transform 1 0 20792 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__A
timestamp 1606120350
transform 1 0 21528 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1036__B
timestamp 1606120350
transform 1 0 21160 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1075__C
timestamp 1606120350
transform 1 0 20516 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_88_207
timestamp 1606120350
transform 1 0 20148 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_88_213
timestamp 1606120350
transform 1 0 20700 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_88_215
timestamp 1606120350
transform 1 0 20884 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_88_220
timestamp 1606120350
transform 1 0 21344 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1067_
timestamp 1606120350
transform 1 0 23644 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__A
timestamp 1606120350
transform 1 0 23460 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1016__A2
timestamp 1606120350
transform 1 0 23092 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_237
timestamp 1606120350
transform 1 0 22908 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_241
timestamp 1606120350
transform 1 0 23276 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0890__A
timestamp 1606120350
transform 1 0 25392 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__A2
timestamp 1606120350
transform 1 0 24932 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1067__A1
timestamp 1606120350
transform 1 0 25760 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__D
timestamp 1606120350
transform 1 0 26220 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_257
timestamp 1606120350
transform 1 0 24748 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_88_261
timestamp 1606120350
transform 1 0 25116 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_88_266
timestamp 1606120350
transform 1 0 25576 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_88_270
timestamp 1606120350
transform 1 0 25944 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_4  _0902_
timestamp 1606120350
transform 1 0 27416 0 -1 50592
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_860
timestamp 1606120350
transform 1 0 26404 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__B1
timestamp 1606120350
transform 1 0 27048 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__B
timestamp 1606120350
transform 1 0 26680 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_276
timestamp 1606120350
transform 1 0 26496 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_280
timestamp 1606120350
transform 1 0 26864 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_284
timestamp 1606120350
transform 1 0 27232 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1194_
timestamp 1606120350
transform 1 0 29532 0 -1 50592
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0930__B1_N
timestamp 1606120350
transform 1 0 29256 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__A2
timestamp 1606120350
transform 1 0 28796 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_299
timestamp 1606120350
transform 1 0 28612 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_88_303
timestamp 1606120350
transform 1 0 28980 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_88_308
timestamp 1606120350
transform 1 0 29440 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_861
timestamp 1606120350
transform 1 0 32016 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_12_0_clk_A
timestamp 1606120350
transform 1 0 31464 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_88_328
timestamp 1606120350
transform 1 0 31280 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_88_332
timestamp 1606120350
transform 1 0 31648 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_88_337
timestamp 1606120350
transform 1 0 32108 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_349
timestamp 1606120350
transform 1 0 33212 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_361
timestamp 1606120350
transform 1 0 34316 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_373
timestamp 1606120350
transform 1 0 35420 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_385
timestamp 1606120350
transform 1 0 36524 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1606120350
transform -1 0 38824 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_862
timestamp 1606120350
transform 1 0 37628 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_88_398
timestamp 1606120350
transform 1 0 37720 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_88_406
timestamp 1606120350
transform 1 0 38456 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1606120350
transform 1 0 1104 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_89_3
timestamp 1606120350
transform 1 0 1380 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_15
timestamp 1606120350
transform 1 0 2484 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_27
timestamp 1606120350
transform 1 0 3588 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_39
timestamp 1606120350
transform 1 0 4692 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_863
timestamp 1606120350
transform 1 0 6716 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_89_51
timestamp 1606120350
transform 1 0 5796 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_89_59
timestamp 1606120350
transform 1 0 6532 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_89_62
timestamp 1606120350
transform 1 0 6808 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_74
timestamp 1606120350
transform 1 0 7912 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_86
timestamp 1606120350
transform 1 0 9016 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_98
timestamp 1606120350
transform 1 0 10120 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_110
timestamp 1606120350
transform 1 0 11224 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_864
timestamp 1606120350
transform 1 0 12328 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_123
timestamp 1606120350
transform 1 0 12420 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_89_135
timestamp 1606120350
transform 1 0 13524 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _1070_
timestamp 1606120350
transform 1 0 15088 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__A1
timestamp 1606120350
transform 1 0 15548 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__B1
timestamp 1606120350
transform 1 0 14904 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1070__A
timestamp 1606120350
transform 1 0 14536 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_89_143
timestamp 1606120350
transform 1 0 14260 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_89_148
timestamp 1606120350
transform 1 0 14720 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_155
timestamp 1606120350
transform 1 0 15364 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_159
timestamp 1606120350
transform 1 0 15732 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1037_
timestamp 1606120350
transform 1 0 16100 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__A1
timestamp 1606120350
transform 1 0 17756 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1030__A1
timestamp 1606120350
transform 1 0 17388 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0985__A
timestamp 1606120350
transform 1 0 15916 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_175
timestamp 1606120350
transform 1 0 17204 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_179
timestamp 1606120350
transform 1 0 17572 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _1033_
timestamp 1606120350
transform 1 0 18032 0 1 50592
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_865
timestamp 1606120350
transform 1 0 17940 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__A1
timestamp 1606120350
transform 1 0 19412 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1079__A2
timestamp 1606120350
transform 1 0 19780 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_197
timestamp 1606120350
transform 1 0 19228 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_201
timestamp 1606120350
transform 1 0 19596 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_89_205
timestamp 1606120350
transform 1 0 19964 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_4  _1075_
timestamp 1606120350
transform 1 0 20516 0 1 50592
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__B1
timestamp 1606120350
transform 1 0 21896 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1040__A
timestamp 1606120350
transform 1 0 20332 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_224
timestamp 1606120350
transform 1 0 21712 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_228
timestamp 1606120350
transform 1 0 22080 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__A1
timestamp 1606120350
transform 1 0 22264 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0879_
timestamp 1606120350
transform 1 0 22448 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_89_235
timestamp 1606120350
transform 1 0 22724 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_89_239
timestamp 1606120350
transform 1 0 23092 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0879__A
timestamp 1606120350
transform 1 0 22908 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__C
timestamp 1606120350
transform 1 0 23368 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_89_245
timestamp 1606120350
transform 1 0 23644 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_866
timestamp 1606120350
transform 1 0 23552 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_251
timestamp 1606120350
transform 1 0 24196 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0883_
timestamp 1606120350
transform 1 0 23920 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1174_
timestamp 1606120350
transform 1 0 24932 0 1 50592
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__D
timestamp 1606120350
transform 1 0 24748 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0883__A
timestamp 1606120350
transform 1 0 24380 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_255
timestamp 1606120350
transform 1 0 24564 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0899_
timestamp 1606120350
transform 1 0 27416 0 1 50592
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0901__A
timestamp 1606120350
transform 1 0 26864 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__A
timestamp 1606120350
transform 1 0 27232 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_278
timestamp 1606120350
transform 1 0 26680 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_282
timestamp 1606120350
transform 1 0 27048 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_295
timestamp 1606120350
transform 1 0 28244 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0854_
timestamp 1606120350
transform 1 0 29256 0 1 50592
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_867
timestamp 1606120350
transform 1 0 29164 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0854__A
timestamp 1606120350
transform 1 0 28980 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__B1_N
timestamp 1606120350
transform 1 0 28428 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0944__A
timestamp 1606120350
transform 1 0 30268 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_89_299
timestamp 1606120350
transform 1 0 28612 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_89_315
timestamp 1606120350
transform 1 0 30084 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_319
timestamp 1606120350
transform 1 0 30452 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0839_
timestamp 1606120350
transform 1 0 30820 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0839__A
timestamp 1606120350
transform 1 0 31280 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0900__A1
timestamp 1606120350
transform 1 0 30636 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_6_0_clk_A
timestamp 1606120350
transform 1 0 31648 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_326
timestamp 1606120350
transform 1 0 31096 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_89_330
timestamp 1606120350
transform 1 0 31464 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_89_334
timestamp 1606120350
transform 1 0 31832 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_13_0_clk_A
timestamp 1606120350
transform 1 0 33672 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_89_346
timestamp 1606120350
transform 1 0 32936 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_89_356
timestamp 1606120350
transform 1 0 33856 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_89_364
timestamp 1606120350
transform 1 0 34592 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_868
timestamp 1606120350
transform 1 0 34776 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_367
timestamp 1606120350
transform 1 0 34868 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_379
timestamp 1606120350
transform 1 0 35972 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1606120350
transform -1 0 38824 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_89_391
timestamp 1606120350
transform 1 0 37076 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_403
timestamp 1606120350
transform 1 0 38180 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1606120350
transform 1 0 1104 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_90_3
timestamp 1606120350
transform 1 0 1380 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_15
timestamp 1606120350
transform 1 0 2484 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_869
timestamp 1606120350
transform 1 0 3956 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_27
timestamp 1606120350
transform 1 0 3588 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_90_32
timestamp 1606120350
transform 1 0 4048 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_44
timestamp 1606120350
transform 1 0 5152 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_56
timestamp 1606120350
transform 1 0 6256 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_68
timestamp 1606120350
transform 1 0 7360 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_80
timestamp 1606120350
transform 1 0 8464 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_870
timestamp 1606120350
transform 1 0 9568 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_93
timestamp 1606120350
transform 1 0 9660 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_105
timestamp 1606120350
transform 1 0 10764 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_117
timestamp 1606120350
transform 1 0 11868 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_129
timestamp 1606120350
transform 1 0 12972 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_871
timestamp 1606120350
transform 1 0 15180 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__D
timestamp 1606120350
transform 1 0 15456 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__B1
timestamp 1606120350
transform 1 0 14996 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__B1
timestamp 1606120350
transform 1 0 14628 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_90_141
timestamp 1606120350
transform 1 0 14076 0 -1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_90_149
timestamp 1606120350
transform 1 0 14812 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_154
timestamp 1606120350
transform 1 0 15272 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_158
timestamp 1606120350
transform 1 0 15640 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0985_
timestamp 1606120350
transform 1 0 16008 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _1030_
timestamp 1606120350
transform 1 0 17020 0 -1 51680
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__A1
timestamp 1606120350
transform 1 0 16836 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__A1
timestamp 1606120350
transform 1 0 16468 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1037__A2
timestamp 1606120350
transform 1 0 15824 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_165
timestamp 1606120350
transform 1 0 16284 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_169
timestamp 1606120350
transform 1 0 16652 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1079_
timestamp 1606120350
transform 1 0 18952 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__B
timestamp 1606120350
transform 1 0 18400 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1033__A2
timestamp 1606120350
transform 1 0 18768 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_186
timestamp 1606120350
transform 1 0 18216 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_190
timestamp 1606120350
transform 1 0 18584 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_210
timestamp 1606120350
transform 1 0 20424 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_206
timestamp 1606120350
transform 1 0 20056 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__C
timestamp 1606120350
transform 1 0 20608 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__B
timestamp 1606120350
transform 1 0 20240 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_872
timestamp 1606120350
transform 1 0 20792 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _1040_
timestamp 1606120350
transform 1 0 20884 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_90_222
timestamp 1606120350
transform 1 0 21528 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_218
timestamp 1606120350
transform 1 0 21160 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1048__B
timestamp 1606120350
transform 1 0 21344 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1002__A2
timestamp 1606120350
transform 1 0 21712 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _1002_
timestamp 1606120350
transform 1 0 21896 0 -1 51680
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_4  _1065_
timestamp 1606120350
transform 1 0 23828 0 -1 51680
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1065__B
timestamp 1606120350
transform 1 0 23644 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__B
timestamp 1606120350
transform 1 0 23276 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_239
timestamp 1606120350
transform 1 0 23092 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_243
timestamp 1606120350
transform 1 0 23460 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0890_
timestamp 1606120350
transform 1 0 25392 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__B1
timestamp 1606120350
transform 1 0 24840 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__B
timestamp 1606120350
transform 1 0 25208 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__A
timestamp 1606120350
transform 1 0 25852 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1066__B
timestamp 1606120350
transform 1 0 26220 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_256
timestamp 1606120350
transform 1 0 24656 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_260
timestamp 1606120350
transform 1 0 25024 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_267
timestamp 1606120350
transform 1 0 25668 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_271
timestamp 1606120350
transform 1 0 26036 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0901_
timestamp 1606120350
transform 1 0 26496 0 -1 51680
box -38 -48 866 592
use sky130_fd_sc_hd__a21bo_4  _0936_
timestamp 1606120350
transform 1 0 28244 0 -1 51680
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_873
timestamp 1606120350
transform 1 0 26404 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__B
timestamp 1606120350
transform 1 0 27508 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0899__C
timestamp 1606120350
transform 1 0 27876 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_285
timestamp 1606120350
transform 1 0 27324 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_289
timestamp 1606120350
transform 1 0 27692 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_293
timestamp 1606120350
transform 1 0 28060 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0944_
timestamp 1606120350
transform 1 0 30176 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0936__A1
timestamp 1606120350
transform 1 0 29624 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1174__CLK
timestamp 1606120350
transform 1 0 29992 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_308
timestamp 1606120350
transform 1 0 29440 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_312
timestamp 1606120350
transform 1 0 29808 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_90_319
timestamp 1606120350
transform 1 0 30452 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_874
timestamp 1606120350
transform 1 0 32016 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_6_0_clk
timestamp 1606120350
transform 1 0 31188 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__CLK
timestamp 1606120350
transform 1 0 30636 0 -1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_90_323
timestamp 1606120350
transform 1 0 30820 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_90_330
timestamp 1606120350
transform 1 0 31464 0 -1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_90_337
timestamp 1606120350
transform 1 0 32108 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_13_0_clk
timestamp 1606120350
transform 1 0 33672 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_90_349
timestamp 1606120350
transform 1 0 33212 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_90_353
timestamp 1606120350
transform 1 0 33580 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_357
timestamp 1606120350
transform 1 0 33948 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_369
timestamp 1606120350
transform 1 0 35052 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_381
timestamp 1606120350
transform 1 0 36156 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1606120350
transform -1 0 38824 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_875
timestamp 1606120350
transform 1 0 37628 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_90_393
timestamp 1606120350
transform 1 0 37260 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_90_398
timestamp 1606120350
transform 1 0 37720 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_90_406
timestamp 1606120350
transform 1 0 38456 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1606120350
transform 1 0 1104 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_3
timestamp 1606120350
transform 1 0 1380 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_15
timestamp 1606120350
transform 1 0 2484 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_27
timestamp 1606120350
transform 1 0 3588 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_39
timestamp 1606120350
transform 1 0 4692 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_876
timestamp 1606120350
transform 1 0 6716 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_91_51
timestamp 1606120350
transform 1 0 5796 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_91_59
timestamp 1606120350
transform 1 0 6532 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_91_62
timestamp 1606120350
transform 1 0 6808 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_74
timestamp 1606120350
transform 1 0 7912 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_86
timestamp 1606120350
transform 1 0 9016 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__D
timestamp 1606120350
transform 1 0 10212 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1146__CLK
timestamp 1606120350
transform 1 0 10580 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_91_98
timestamp 1606120350
transform 1 0 10120 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_91_101
timestamp 1606120350
transform 1 0 10396 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_91_105
timestamp 1606120350
transform 1 0 10764 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_877
timestamp 1606120350
transform 1 0 12328 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_91_117
timestamp 1606120350
transform 1 0 11868 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_91_121
timestamp 1606120350
transform 1 0 12236 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_123
timestamp 1606120350
transform 1 0 12420 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_135
timestamp 1606120350
transform 1 0 13524 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__A
timestamp 1606120350
transform 1 0 15456 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__C
timestamp 1606120350
transform 1 0 15088 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1071__A2
timestamp 1606120350
transform 1 0 14720 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1076__A2
timestamp 1606120350
transform 1 0 14352 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_91_143
timestamp 1606120350
transform 1 0 14260 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_91_146
timestamp 1606120350
transform 1 0 14536 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_150
timestamp 1606120350
transform 1 0 14904 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_154
timestamp 1606120350
transform 1 0 15272 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_158
timestamp 1606120350
transform 1 0 15640 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1071_
timestamp 1606120350
transform 1 0 16100 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__D
timestamp 1606120350
transform 1 0 17756 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1055__B
timestamp 1606120350
transform 1 0 15824 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__C
timestamp 1606120350
transform 1 0 17388 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_91_162
timestamp 1606120350
transform 1 0 16008 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_91_175
timestamp 1606120350
transform 1 0 17204 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_179
timestamp 1606120350
transform 1 0 17572 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__nor3_4  _1029_
timestamp 1606120350
transform 1 0 19596 0 1 51680
box -38 -48 1234 592
use sky130_fd_sc_hd__and4_4  _1064_
timestamp 1606120350
transform 1 0 18032 0 1 51680
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_878
timestamp 1606120350
transform 1 0 17940 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__A
timestamp 1606120350
transform 1 0 19412 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1063__A1
timestamp 1606120350
transform 1 0 19044 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_193
timestamp 1606120350
transform 1 0 18860 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_197
timestamp 1606120350
transform 1 0 19228 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__nor3_4  _1066_
timestamp 1606120350
transform 1 0 21528 0 1 51680
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__A2
timestamp 1606120350
transform 1 0 21344 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1035__A
timestamp 1606120350
transform 1 0 20976 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_214
timestamp 1606120350
transform 1 0 20792 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_218
timestamp 1606120350
transform 1 0 21160 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1046_
timestamp 1606120350
transform 1 0 23644 0 1 51680
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_879
timestamp 1606120350
transform 1 0 23552 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__C
timestamp 1606120350
transform 1 0 23368 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__A1
timestamp 1606120350
transform 1 0 22908 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_235
timestamp 1606120350
transform 1 0 22724 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_91_239
timestamp 1606120350
transform 1 0 23092 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _0946_
timestamp 1606120350
transform 1 0 25208 0 1 51680
box -38 -48 682 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__A
timestamp 1606120350
transform 1 0 26036 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0946__B
timestamp 1606120350
transform 1 0 25024 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0945__A
timestamp 1606120350
transform 1 0 24656 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_254
timestamp 1606120350
transform 1 0 24472 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_258
timestamp 1606120350
transform 1 0 24840 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_269
timestamp 1606120350
transform 1 0 25852 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_273
timestamp 1606120350
transform 1 0 26220 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0903_
timestamp 1606120350
transform 1 0 26588 0 1 51680
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1043_
timestamp 1606120350
transform 1 0 28152 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__A2
timestamp 1606120350
transform 1 0 27600 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__A
timestamp 1606120350
transform 1 0 26404 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__B1_N
timestamp 1606120350
transform 1 0 27968 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_286
timestamp 1606120350
transform 1 0 27416 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_290
timestamp 1606120350
transform 1 0 27784 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_301
timestamp 1606120350
transform 1 0 28796 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_297
timestamp 1606120350
transform 1 0 28428 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1043__A
timestamp 1606120350
transform 1 0 28612 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0968__A
timestamp 1606120350
transform 1 0 28980 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_880
timestamp 1606120350
transform 1 0 29164 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0968_
timestamp 1606120350
transform 1 0 29256 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_91_313
timestamp 1606120350
transform 1 0 29900 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_91_309
timestamp 1606120350
transform 1 0 29532 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__D
timestamp 1606120350
transform 1 0 29716 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1189__D
timestamp 1606120350
transform 1 0 30084 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1189_
timestamp 1606120350
transform 1 0 30268 0 1 51680
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_91_336
timestamp 1606120350
transform 1 0 32016 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_348
timestamp 1606120350
transform 1 0 33120 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_91_360
timestamp 1606120350
transform 1 0 34224 0 1 51680
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_881
timestamp 1606120350
transform 1 0 34776 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_367
timestamp 1606120350
transform 1 0 34868 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_379
timestamp 1606120350
transform 1 0 35972 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1606120350
transform -1 0 38824 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_391
timestamp 1606120350
transform 1 0 37076 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_91_403
timestamp 1606120350
transform 1 0 38180 0 1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1606120350
transform 1 0 1104 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1606120350
transform 1 0 1104 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_92_3
timestamp 1606120350
transform 1 0 1380 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_15
timestamp 1606120350
transform 1 0 2484 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_3
timestamp 1606120350
transform 1 0 1380 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_15
timestamp 1606120350
transform 1 0 2484 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_882
timestamp 1606120350
transform 1 0 3956 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_27
timestamp 1606120350
transform 1 0 3588 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_92_32
timestamp 1606120350
transform 1 0 4048 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_44
timestamp 1606120350
transform 1 0 5152 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_27
timestamp 1606120350
transform 1 0 3588 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_39
timestamp 1606120350
transform 1 0 4692 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_889
timestamp 1606120350
transform 1 0 6716 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_56
timestamp 1606120350
transform 1 0 6256 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_68
timestamp 1606120350
transform 1 0 7360 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_51
timestamp 1606120350
transform 1 0 5796 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_93_59
timestamp 1606120350
transform 1 0 6532 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_93_62
timestamp 1606120350
transform 1 0 6808 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_80
timestamp 1606120350
transform 1 0 8464 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_74
timestamp 1606120350
transform 1 0 7912 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_86
timestamp 1606120350
transform 1 0 9016 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1146_
timestamp 1606120350
transform 1 0 10212 0 -1 52768
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_883
timestamp 1606120350
transform 1 0 9568 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_92_93
timestamp 1606120350
transform 1 0 9660 0 -1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_93_98
timestamp 1606120350
transform 1 0 10120 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_110
timestamp 1606120350
transform 1 0 11224 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_890
timestamp 1606120350
transform 1 0 12328 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_118
timestamp 1606120350
transform 1 0 11960 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_130
timestamp 1606120350
transform 1 0 13064 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_123
timestamp 1606120350
transform 1 0 12420 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_93_135
timestamp 1606120350
transform 1 0 13524 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_93_144
timestamp 1606120350
transform 1 0 14352 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_140
timestamp 1606120350
transform 1 0 13984 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_92_146
timestamp 1606120350
transform 1 0 14536 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_142
timestamp 1606120350
transform 1 0 14168 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_2_0_clk_A
timestamp 1606120350
transform 1 0 13800 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1001__A
timestamp 1606120350
transform 1 0 14168 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__B
timestamp 1606120350
transform 1 0 14536 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__C
timestamp 1606120350
transform 1 0 14904 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__A
timestamp 1606120350
transform 1 0 14996 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__B1
timestamp 1606120350
transform 1 0 14628 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_149
timestamp 1606120350
transform 1 0 14812 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_148
timestamp 1606120350
transform 1 0 14720 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0986_
timestamp 1606120350
transform 1 0 15364 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_884
timestamp 1606120350
transform 1 0 15180 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_2_0_clk
timestamp 1606120350
transform 1 0 15088 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_92_154
timestamp 1606120350
transform 1 0 15272 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _1055_
timestamp 1606120350
transform 1 0 15456 0 -1 52768
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_93_158
timestamp 1606120350
transform 1 0 15640 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_162
timestamp 1606120350
transform 1 0 16008 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_169
timestamp 1606120350
transform 1 0 16652 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_165
timestamp 1606120350
transform 1 0 16284 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__B
timestamp 1606120350
transform 1 0 16836 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__A
timestamp 1606120350
transform 1 0 16468 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0986__A
timestamp 1606120350
transform 1 0 16192 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1027__D
timestamp 1606120350
transform 1 0 15824 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1031_
timestamp 1606120350
transform 1 0 16376 0 1 52768
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_93_179
timestamp 1606120350
transform 1 0 17572 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_175
timestamp 1606120350
transform 1 0 17204 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__A1
timestamp 1606120350
transform 1 0 17756 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__C
timestamp 1606120350
transform 1 0 17388 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1076_
timestamp 1606120350
transform 1 0 17020 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_93_184
timestamp 1606120350
transform 1 0 18032 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_92_189
timestamp 1606120350
transform 1 0 18492 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_185
timestamp 1606120350
transform 1 0 18124 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__A1
timestamp 1606120350
transform 1 0 18676 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1064__A
timestamp 1606120350
transform 1 0 18308 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_891
timestamp 1606120350
transform 1 0 17940 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_202
timestamp 1606120350
transform 1 0 19688 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_198
timestamp 1606120350
transform 1 0 19320 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__C
timestamp 1606120350
transform 1 0 19872 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__A
timestamp 1606120350
transform 1 0 19504 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _1078_
timestamp 1606120350
transform 1 0 18124 0 1 52768
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _1063_
timestamp 1606120350
transform 1 0 18860 0 -1 52768
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_1  _1032_
timestamp 1606120350
transform 1 0 20056 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1029__C
timestamp 1606120350
transform 1 0 20240 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_206
timestamp 1606120350
transform 1 0 20056 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_209
timestamp 1606120350
transform 1 0 20332 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__D
timestamp 1606120350
transform 1 0 20516 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1032__A
timestamp 1606120350
transform 1 0 20608 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_210
timestamp 1606120350
transform 1 0 20424 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_213
timestamp 1606120350
transform 1 0 20700 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1035_
timestamp 1606120350
transform 1 0 20884 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_885
timestamp 1606120350
transform 1 0 20792 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1045__B
timestamp 1606120350
transform 1 0 20884 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_217
timestamp 1606120350
transform 1 0 21068 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_92_225
timestamp 1606120350
transform 1 0 21804 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_92_222
timestamp 1606120350
transform 1 0 21528 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_218
timestamp 1606120350
transform 1 0 21160 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1048__A
timestamp 1606120350
transform 1 0 21620 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0997__B1
timestamp 1606120350
transform 1 0 22080 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__nor3_4  _1056_
timestamp 1606120350
transform 1 0 21252 0 1 52768
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_93_236
timestamp 1606120350
transform 1 0 22816 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_232
timestamp 1606120350
transform 1 0 22448 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__A1
timestamp 1606120350
transform 1 0 22632 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__C
timestamp 1606120350
transform 1 0 23000 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_240
timestamp 1606120350
transform 1 0 23184 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_247
timestamp 1606120350
transform 1 0 23828 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_243
timestamp 1606120350
transform 1 0 23460 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1046__A
timestamp 1606120350
transform 1 0 24012 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__B
timestamp 1606120350
transform 1 0 23644 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0960__A
timestamp 1606120350
transform 1 0 23368 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_892
timestamp 1606120350
transform 1 0 23552 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _0960_
timestamp 1606120350
transform 1 0 23644 0 1 52768
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  _0945_
timestamp 1606120350
transform 1 0 24196 0 -1 52768
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _0997_
timestamp 1606120350
transform 1 0 22264 0 -1 52768
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_93_258
timestamp 1606120350
transform 1 0 24840 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_254
timestamp 1606120350
transform 1 0 24472 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_260
timestamp 1606120350
transform 1 0 25024 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__A2
timestamp 1606120350
transform 1 0 24656 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__B
timestamp 1606120350
transform 1 0 25024 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_268
timestamp 1606120350
transform 1 0 25760 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_264
timestamp 1606120350
transform 1 0 25392 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1048__C
timestamp 1606120350
transform 1 0 25944 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__D
timestamp 1606120350
transform 1 0 25576 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__C
timestamp 1606120350
transform 1 0 25208 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _1074_
timestamp 1606120350
transform 1 0 25208 0 1 52768
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_93_271
timestamp 1606120350
transform 1 0 26036 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_92_272
timestamp 1606120350
transform 1 0 26128 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_886
timestamp 1606120350
transform 1 0 26404 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__B
timestamp 1606120350
transform 1 0 26680 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__A2
timestamp 1606120350
transform 1 0 26496 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_276
timestamp 1606120350
transform 1 0 26496 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_93_275
timestamp 1606120350
transform 1 0 26404 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_278
timestamp 1606120350
transform 1 0 26680 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__A
timestamp 1606120350
transform 1 0 26864 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__C
timestamp 1606120350
transform 1 0 27048 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_280
timestamp 1606120350
transform 1 0 26864 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0905_
timestamp 1606120350
transform 1 0 27048 0 1 52768
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_93_295
timestamp 1606120350
transform 1 0 28244 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_93_291
timestamp 1606120350
transform 1 0 27876 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__B1
timestamp 1606120350
transform 1 0 28060 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__a21bo_4  _0906_
timestamp 1606120350
transform 1 0 27232 0 -1 52768
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_93_306
timestamp 1606120350
transform 1 0 29256 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_93_299
timestamp 1606120350
transform 1 0 28612 0 1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_92_301
timestamp 1606120350
transform 1 0 28796 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_92_297
timestamp 1606120350
transform 1 0 28428 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1173__CLK
timestamp 1606120350
transform 1 0 29440 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0903__D
timestamp 1606120350
transform 1 0 28980 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0906__A1
timestamp 1606120350
transform 1 0 28612 0 -1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0905__B
timestamp 1606120350
transform 1 0 28428 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_893
timestamp 1606120350
transform 1 0 29164 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_310
timestamp 1606120350
transform 1 0 29624 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1173_
timestamp 1606120350
transform 1 0 29164 0 -1 52768
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_887
timestamp 1606120350
transform 1 0 32016 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_324
timestamp 1606120350
transform 1 0 30912 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_337
timestamp 1606120350
transform 1 0 32108 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_322
timestamp 1606120350
transform 1 0 30728 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_334
timestamp 1606120350
transform 1 0 31832 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_349
timestamp 1606120350
transform 1 0 33212 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_361
timestamp 1606120350
transform 1 0 34316 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_346
timestamp 1606120350
transform 1 0 32936 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_358
timestamp 1606120350
transform 1 0 34040 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_894
timestamp 1606120350
transform 1 0 34776 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_373
timestamp 1606120350
transform 1 0 35420 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_385
timestamp 1606120350
transform 1 0 36524 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_367
timestamp 1606120350
transform 1 0 34868 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_379
timestamp 1606120350
transform 1 0 35972 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1606120350
transform -1 0 38824 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1606120350
transform -1 0 38824 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_888
timestamp 1606120350
transform 1 0 37628 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_92_398
timestamp 1606120350
transform 1 0 37720 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_92_406
timestamp 1606120350
transform 1 0 38456 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_391
timestamp 1606120350
transform 1 0 37076 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_93_403
timestamp 1606120350
transform 1 0 38180 0 1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1606120350
transform 1 0 1104 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_94_3
timestamp 1606120350
transform 1 0 1380 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_15
timestamp 1606120350
transform 1 0 2484 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_895
timestamp 1606120350
transform 1 0 3956 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_94_27
timestamp 1606120350
transform 1 0 3588 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_94_32
timestamp 1606120350
transform 1 0 4048 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_44
timestamp 1606120350
transform 1 0 5152 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_56
timestamp 1606120350
transform 1 0 6256 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_68
timestamp 1606120350
transform 1 0 7360 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_80
timestamp 1606120350
transform 1 0 8464 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_896
timestamp 1606120350
transform 1 0 9568 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_93
timestamp 1606120350
transform 1 0 9660 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_105
timestamp 1606120350
transform 1 0 10764 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_117
timestamp 1606120350
transform 1 0 11868 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_94_129
timestamp 1606120350
transform 1 0 12972 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_94_137
timestamp 1606120350
transform 1 0 13708 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1001_
timestamp 1606120350
transform 1 0 14168 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _1027_
timestamp 1606120350
transform 1 0 15548 0 -1 53856
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_897
timestamp 1606120350
transform 1 0 15180 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__A2
timestamp 1606120350
transform 1 0 14996 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1077__B1
timestamp 1606120350
transform 1 0 14628 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__CLK
timestamp 1606120350
transform 1 0 13984 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_145
timestamp 1606120350
transform 1 0 14444 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_149
timestamp 1606120350
transform 1 0 14812 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_94_154
timestamp 1606120350
transform 1 0 15272 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _1077_
timestamp 1606120350
transform 1 0 17112 0 -1 53856
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__B
timestamp 1606120350
transform 1 0 16560 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1031__D
timestamp 1606120350
transform 1 0 16928 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_166
timestamp 1606120350
transform 1 0 16376 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_170
timestamp 1606120350
transform 1 0 16744 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _1045_
timestamp 1606120350
transform 1 0 19228 0 -1 53856
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__A
timestamp 1606120350
transform 1 0 18584 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__B
timestamp 1606120350
transform 1 0 19044 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_94_187
timestamp 1606120350
transform 1 0 18308 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_94_192
timestamp 1606120350
transform 1 0 18768 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_94_215
timestamp 1606120350
transform 1 0 20884 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_210
timestamp 1606120350
transform 1 0 20424 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_206
timestamp 1606120350
transform 1 0 20056 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__A
timestamp 1606120350
transform 1 0 20608 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__C
timestamp 1606120350
transform 1 0 20240 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_898
timestamp 1606120350
transform 1 0 20792 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_94_219
timestamp 1606120350
transform 1 0 21252 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__B1
timestamp 1606120350
transform 1 0 21068 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__B
timestamp 1606120350
transform 1 0 21436 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__nor3_4  _1048_
timestamp 1606120350
transform 1 0 21620 0 -1 53856
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _1054_
timestamp 1606120350
transform 1 0 23552 0 -1 53856
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1054__A2
timestamp 1606120350
transform 1 0 23368 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__A
timestamp 1606120350
transform 1 0 23000 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_236
timestamp 1606120350
transform 1 0 22816 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_240
timestamp 1606120350
transform 1 0 23184 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__A2
timestamp 1606120350
transform 1 0 24932 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__B1
timestamp 1606120350
transform 1 0 25300 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__B
timestamp 1606120350
transform 1 0 26220 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1074__A
timestamp 1606120350
transform 1 0 25668 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_257
timestamp 1606120350
transform 1 0 24748 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_261
timestamp 1606120350
transform 1 0 25116 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_265
timestamp 1606120350
transform 1 0 25484 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_94_269
timestamp 1606120350
transform 1 0 25852 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _0904_
timestamp 1606120350
transform 1 0 26864 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_899
timestamp 1606120350
transform 1 0 26404 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__A
timestamp 1606120350
transform 1 0 26680 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0904__A1
timestamp 1606120350
transform 1 0 28152 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_276
timestamp 1606120350
transform 1 0 26496 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_94_292
timestamp 1606120350
transform 1 0 27968 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_94_296
timestamp 1606120350
transform 1 0 28336 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_308
timestamp 1606120350
transform 1 0 29440 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_900
timestamp 1606120350
transform 1 0 32016 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_320
timestamp 1606120350
transform 1 0 30544 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_332
timestamp 1606120350
transform 1 0 31648 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_94_337
timestamp 1606120350
transform 1 0 32108 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_349
timestamp 1606120350
transform 1 0 33212 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_361
timestamp 1606120350
transform 1 0 34316 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_373
timestamp 1606120350
transform 1 0 35420 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_385
timestamp 1606120350
transform 1 0 36524 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1606120350
transform -1 0 38824 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_901
timestamp 1606120350
transform 1 0 37628 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_94_398
timestamp 1606120350
transform 1 0 37720 0 -1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_94_406
timestamp 1606120350
transform 1 0 38456 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1606120350
transform 1 0 1104 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_95_3
timestamp 1606120350
transform 1 0 1380 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_15
timestamp 1606120350
transform 1 0 2484 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_27
timestamp 1606120350
transform 1 0 3588 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_39
timestamp 1606120350
transform 1 0 4692 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_902
timestamp 1606120350
transform 1 0 6716 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_95_51
timestamp 1606120350
transform 1 0 5796 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_95_59
timestamp 1606120350
transform 1 0 6532 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_95_62
timestamp 1606120350
transform 1 0 6808 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_74
timestamp 1606120350
transform 1 0 7912 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_86
timestamp 1606120350
transform 1 0 9016 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_98
timestamp 1606120350
transform 1 0 10120 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_110
timestamp 1606120350
transform 1 0 11224 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_903
timestamp 1606120350
transform 1 0 12328 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1007__A
timestamp 1606120350
transform 1 0 13616 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1025__A
timestamp 1606120350
transform 1 0 13156 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_123
timestamp 1606120350
transform 1 0 12420 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_95_133
timestamp 1606120350
transform 1 0 13340 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _1007_
timestamp 1606120350
transform 1 0 13800 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1208_
timestamp 1606120350
transform 1 0 14812 0 1 53856
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1208__D
timestamp 1606120350
transform 1 0 14628 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1008__A
timestamp 1606120350
transform 1 0 14260 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_141
timestamp 1606120350
transform 1 0 14076 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_145
timestamp 1606120350
transform 1 0 14444 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__A
timestamp 1606120350
transform 1 0 16744 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__C
timestamp 1606120350
transform 1 0 17112 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1039__D
timestamp 1606120350
transform 1 0 17480 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_168
timestamp 1606120350
transform 1 0 16560 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_172
timestamp 1606120350
transform 1 0 16928 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_176
timestamp 1606120350
transform 1 0 17296 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_95_180
timestamp 1606120350
transform 1 0 17664 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _0952_
timestamp 1606120350
transform 1 0 18584 0 1 53856
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_904
timestamp 1606120350
transform 1 0 17940 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__C
timestamp 1606120350
transform 1 0 19596 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__C
timestamp 1606120350
transform 1 0 18400 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1010__A
timestamp 1606120350
transform 1 0 19964 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_95_184
timestamp 1606120350
transform 1 0 18032 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_95_199
timestamp 1606120350
transform 1 0 19412 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_203
timestamp 1606120350
transform 1 0 19780 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _0996_
timestamp 1606120350
transform 1 0 21712 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_4  _1009_
timestamp 1606120350
transform 1 0 20148 0 1 53856
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__A
timestamp 1606120350
transform 1 0 21528 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0988__C
timestamp 1606120350
transform 1 0 21160 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_216
timestamp 1606120350
transform 1 0 20976 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_220
timestamp 1606120350
transform 1 0 21344 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_905
timestamp 1606120350
transform 1 0 23552 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__A1
timestamp 1606120350
transform 1 0 23920 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0967__C1
timestamp 1606120350
transform 1 0 23368 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__A2
timestamp 1606120350
transform 1 0 23000 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_236
timestamp 1606120350
transform 1 0 22816 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_240
timestamp 1606120350
transform 1 0 23184 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_95_245
timestamp 1606120350
transform 1 0 23644 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_95_250
timestamp 1606120350
transform 1 0 24104 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _0967_
timestamp 1606120350
transform 1 0 24472 0 1 53856
box -38 -48 1326 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A2
timestamp 1606120350
transform 1 0 26312 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__B1
timestamp 1606120350
transform 1 0 25944 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__A1
timestamp 1606120350
transform 1 0 24288 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_268
timestamp 1606120350
transform 1 0 25760 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_272
timestamp 1606120350
transform 1 0 26128 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0957_
timestamp 1606120350
transform 1 0 28060 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _0987_
timestamp 1606120350
transform 1 0 26496 0 1 53856
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__C
timestamp 1606120350
transform 1 0 27508 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0957__A
timestamp 1606120350
transform 1 0 27876 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_285
timestamp 1606120350
transform 1 0 27324 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_289
timestamp 1606120350
transform 1 0 27692 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_95_296
timestamp 1606120350
transform 1 0 28336 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_906
timestamp 1606120350
transform 1 0 29164 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__D
timestamp 1606120350
transform 1 0 28612 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1178__CLK
timestamp 1606120350
transform 1 0 28980 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_95_301
timestamp 1606120350
transform 1 0 28796 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_95_306
timestamp 1606120350
transform 1 0 29256 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_318
timestamp 1606120350
transform 1 0 30360 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_330
timestamp 1606120350
transform 1 0 31464 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_342
timestamp 1606120350
transform 1 0 32568 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_354
timestamp 1606120350
transform 1 0 33672 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_907
timestamp 1606120350
transform 1 0 34776 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_367
timestamp 1606120350
transform 1 0 34868 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_379
timestamp 1606120350
transform 1 0 35972 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1606120350
transform -1 0 38824 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_95_391
timestamp 1606120350
transform 1 0 37076 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_95_403
timestamp 1606120350
transform 1 0 38180 0 1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1606120350
transform 1 0 1104 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_3
timestamp 1606120350
transform 1 0 1380 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_15
timestamp 1606120350
transform 1 0 2484 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_908
timestamp 1606120350
transform 1 0 3956 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_27
timestamp 1606120350
transform 1 0 3588 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_96_32
timestamp 1606120350
transform 1 0 4048 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_44
timestamp 1606120350
transform 1 0 5152 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_56
timestamp 1606120350
transform 1 0 6256 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_68
timestamp 1606120350
transform 1 0 7360 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_80
timestamp 1606120350
transform 1 0 8464 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_909
timestamp 1606120350
transform 1 0 9568 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_93
timestamp 1606120350
transform 1 0 9660 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_105
timestamp 1606120350
transform 1 0 10764 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1025_
timestamp 1606120350
transform 1 0 13156 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0953__A
timestamp 1606120350
transform 1 0 13616 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_96_117
timestamp 1606120350
transform 1 0 11868 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_96_129
timestamp 1606120350
transform 1 0 12972 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_96_134
timestamp 1606120350
transform 1 0 13432 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_96_145
timestamp 1606120350
transform 1 0 14444 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_96_138
timestamp 1606120350
transform 1 0 13800 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1004__A
timestamp 1606120350
transform 1 0 13984 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _1008_
timestamp 1606120350
transform 1 0 14168 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_96_154
timestamp 1606120350
transform 1 0 15272 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_96_151
timestamp 1606120350
transform 1 0 14996 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__D
timestamp 1606120350
transform 1 0 15456 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__B
timestamp 1606120350
transform 1 0 14812 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_910
timestamp 1606120350
transform 1 0 15180 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_96_158
timestamp 1606120350
transform 1 0 15640 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _1039_
timestamp 1606120350
transform 1 0 15732 0 -1 54944
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  _0947_
timestamp 1606120350
transform 1 0 17296 0 -1 54944
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__B
timestamp 1606120350
transform 1 0 16744 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1078__A2
timestamp 1606120350
transform 1 0 17112 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_96_168
timestamp 1606120350
transform 1 0 16560 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_96_172
timestamp 1606120350
transform 1 0 16928 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__and3_4  _1010_
timestamp 1606120350
transform 1 0 19228 0 -1 54944
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0952__B
timestamp 1606120350
transform 1 0 18584 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1056__C
timestamp 1606120350
transform 1 0 19044 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_96_185
timestamp 1606120350
transform 1 0 18124 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_96_189
timestamp 1606120350
transform 1 0 18492 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_96_192
timestamp 1606120350
transform 1 0 18768 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_96_215
timestamp 1606120350
transform 1 0 20884 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_96_210
timestamp 1606120350
transform 1 0 20424 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_96_206
timestamp 1606120350
transform 1 0 20056 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__B
timestamp 1606120350
transform 1 0 20608 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1009__D
timestamp 1606120350
transform 1 0 20240 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_911
timestamp 1606120350
transform 1 0 20792 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_96_219
timestamp 1606120350
transform 1 0 21252 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0996__A1
timestamp 1606120350
transform 1 0 21528 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__C
timestamp 1606120350
transform 1 0 21068 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__nor3_4  _0988_
timestamp 1606120350
transform 1 0 21712 0 -1 54944
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__B1
timestamp 1606120350
transform 1 0 24196 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0961__C1
timestamp 1606120350
transform 1 0 23828 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__A2
timestamp 1606120350
transform 1 0 23460 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A2
timestamp 1606120350
transform 1 0 23092 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_96_237
timestamp 1606120350
transform 1 0 22908 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_96_241
timestamp 1606120350
transform 1 0 23276 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_96_245
timestamp 1606120350
transform 1 0 23644 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_96_249
timestamp 1606120350
transform 1 0 24012 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__a211o_4  _0961_
timestamp 1606120350
transform 1 0 24380 0 -1 54944
box -38 -48 1326 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0987__D
timestamp 1606120350
transform 1 0 26220 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0972__A
timestamp 1606120350
transform 1 0 25852 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_96_267
timestamp 1606120350
transform 1 0 25668 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_96_271
timestamp 1606120350
transform 1 0 26036 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__a21o_4  _0909_
timestamp 1606120350
transform 1 0 26496 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_912
timestamp 1606120350
transform 1 0 26404 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0909__A1
timestamp 1606120350
transform 1 0 27784 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_96_288
timestamp 1606120350
transform 1 0 27600 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_96_292
timestamp 1606120350
transform 1 0 27968 0 -1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _1178_
timestamp 1606120350
transform 1 0 28612 0 -1 54944
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_96_298
timestamp 1606120350
transform 1 0 28520 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_318
timestamp 1606120350
transform 1 0 30360 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_913
timestamp 1606120350
transform 1 0 32016 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__A2
timestamp 1606120350
transform 1 0 31740 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_96_330
timestamp 1606120350
transform 1 0 31464 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_96_335
timestamp 1606120350
transform 1 0 31924 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_337
timestamp 1606120350
transform 1 0 32108 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_349
timestamp 1606120350
transform 1 0 33212 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_361
timestamp 1606120350
transform 1 0 34316 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_373
timestamp 1606120350
transform 1 0 35420 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_385
timestamp 1606120350
transform 1 0 36524 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1606120350
transform -1 0 38824 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_914
timestamp 1606120350
transform 1 0 37628 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_398
timestamp 1606120350
transform 1 0 37720 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_96_406
timestamp 1606120350
transform 1 0 38456 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1606120350
transform 1 0 1104 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_3
timestamp 1606120350
transform 1 0 1380 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_15
timestamp 1606120350
transform 1 0 2484 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_27
timestamp 1606120350
transform 1 0 3588 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_39
timestamp 1606120350
transform 1 0 4692 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_915
timestamp 1606120350
transform 1 0 6716 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_97_51
timestamp 1606120350
transform 1 0 5796 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_97_59
timestamp 1606120350
transform 1 0 6532 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_97_62
timestamp 1606120350
transform 1 0 6808 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_74
timestamp 1606120350
transform 1 0 7912 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_86
timestamp 1606120350
transform 1 0 9016 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_98
timestamp 1606120350
transform 1 0 10120 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_97_110
timestamp 1606120350
transform 1 0 11224 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_97_118
timestamp 1606120350
transform 1 0 11960 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0962__A
timestamp 1606120350
transform 1 0 12144 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_123
timestamp 1606120350
transform 1 0 12420 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__D
timestamp 1606120350
transform 1 0 12604 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_916
timestamp 1606120350
transform 1 0 12328 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0949_
timestamp 1606120350
transform 1 0 12788 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_97_130
timestamp 1606120350
transform 1 0 13064 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0949__A
timestamp 1606120350
transform 1 0 13248 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_134
timestamp 1606120350
transform 1 0 13432 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0951__A
timestamp 1606120350
transform 1 0 13616 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0999_
timestamp 1606120350
transform 1 0 13800 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _1034_
timestamp 1606120350
transform 1 0 14812 0 1 54944
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__A
timestamp 1606120350
transform 1 0 14628 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0999__A
timestamp 1606120350
transform 1 0 14260 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_141
timestamp 1606120350
transform 1 0 14076 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_145
timestamp 1606120350
transform 1 0 14444 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_158
timestamp 1606120350
transform 1 0 15640 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _0955_
timestamp 1606120350
transform 1 0 16376 0 1 54944
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__D
timestamp 1606120350
transform 1 0 16192 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__A
timestamp 1606120350
transform 1 0 15824 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0955__C
timestamp 1606120350
transform 1 0 17388 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__A
timestamp 1606120350
transform 1 0 17756 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_162
timestamp 1606120350
transform 1 0 16008 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_175
timestamp 1606120350
transform 1 0 17204 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_179
timestamp 1606120350
transform 1 0 17572 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0972_
timestamp 1606120350
transform 1 0 19596 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  _1003_
timestamp 1606120350
transform 1 0 18032 0 1 54944
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_917
timestamp 1606120350
transform 1 0 17940 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__A
timestamp 1606120350
transform 1 0 19228 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_97_193
timestamp 1606120350
transform 1 0 18860 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_97_199
timestamp 1606120350
transform 1 0 19412 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_204
timestamp 1606120350
transform 1 0 19872 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__nor3_4  _1011_
timestamp 1606120350
transform 1 0 20884 0 1 54944
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__C
timestamp 1606120350
transform 1 0 20056 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__B
timestamp 1606120350
transform 1 0 20424 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_208
timestamp 1606120350
transform 1 0 20240 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_97_212
timestamp 1606120350
transform 1 0 20608 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_97_228
timestamp 1606120350
transform 1 0 22080 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _0980_
timestamp 1606120350
transform 1 0 23644 0 1 54944
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_918
timestamp 1606120350
transform 1 0 23552 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__B1
timestamp 1606120350
transform 1 0 23368 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__B1
timestamp 1606120350
transform 1 0 23000 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__A
timestamp 1606120350
transform 1 0 22264 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__B
timestamp 1606120350
transform 1 0 22632 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_232
timestamp 1606120350
transform 1 0 22448 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_236
timestamp 1606120350
transform 1 0 22816 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_240
timestamp 1606120350
transform 1 0 23184 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A1
timestamp 1606120350
transform 1 0 25024 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0861__A
timestamp 1606120350
transform 1 0 26220 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__A
timestamp 1606120350
transform 1 0 25852 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0910__B
timestamp 1606120350
transform 1 0 25484 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_258
timestamp 1606120350
transform 1 0 24840 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_97_262
timestamp 1606120350
transform 1 0 25208 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_97_267
timestamp 1606120350
transform 1 0 25668 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_271
timestamp 1606120350
transform 1 0 26036 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__nor2_4  _0910_
timestamp 1606120350
transform 1 0 26404 0 1 54944
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _0954_
timestamp 1606120350
transform 1 0 27968 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_97_284
timestamp 1606120350
transform 1 0 27232 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_97_295
timestamp 1606120350
transform 1 0 28244 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_919
timestamp 1606120350
transform 1 0 29164 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0866__A
timestamp 1606120350
transform 1 0 28428 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0954__A
timestamp 1606120350
transform 1 0 28796 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_299
timestamp 1606120350
transform 1 0 28612 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_303
timestamp 1606120350
transform 1 0 28980 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_97_306
timestamp 1606120350
transform 1 0 29256 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_318
timestamp 1606120350
transform 1 0 30360 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__a21bo_4  _0937_
timestamp 1606120350
transform 1 0 31740 0 1 54944
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__B1_N
timestamp 1606120350
transform 1 0 31556 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_97_330
timestamp 1606120350
transform 1 0 31464 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__D
timestamp 1606120350
transform 1 0 33120 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1195__CLK
timestamp 1606120350
transform 1 0 33488 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_346
timestamp 1606120350
transform 1 0 32936 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_97_350
timestamp 1606120350
transform 1 0 33304 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_97_354
timestamp 1606120350
transform 1 0 33672 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_920
timestamp 1606120350
transform 1 0 34776 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_367
timestamp 1606120350
transform 1 0 34868 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_379
timestamp 1606120350
transform 1 0 35972 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1606120350
transform -1 0 38824 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_391
timestamp 1606120350
transform 1 0 37076 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_97_403
timestamp 1606120350
transform 1 0 38180 0 1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1606120350
transform 1 0 1104 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_98_3
timestamp 1606120350
transform 1 0 1380 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_15
timestamp 1606120350
transform 1 0 2484 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_921
timestamp 1606120350
transform 1 0 3956 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_98_27
timestamp 1606120350
transform 1 0 3588 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_98_32
timestamp 1606120350
transform 1 0 4048 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_44
timestamp 1606120350
transform 1 0 5152 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_56
timestamp 1606120350
transform 1 0 6256 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_68
timestamp 1606120350
transform 1 0 7360 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_80
timestamp 1606120350
transform 1 0 8464 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_922
timestamp 1606120350
transform 1 0 9568 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_93
timestamp 1606120350
transform 1 0 9660 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_105
timestamp 1606120350
transform 1 0 10764 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0951_
timestamp 1606120350
transform 1 0 13156 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0962_
timestamp 1606120350
transform 1 0 12144 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1003__A
timestamp 1606120350
transform 1 0 13616 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_98_117
timestamp 1606120350
transform 1 0 11868 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_98_123
timestamp 1606120350
transform 1 0 12420 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_98_134
timestamp 1606120350
transform 1 0 13432 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_138
timestamp 1606120350
transform 1 0 13800 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__C
timestamp 1606120350
transform 1 0 13984 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_98_145
timestamp 1606120350
transform 1 0 14444 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  _1004_
timestamp 1606120350
transform 1 0 14168 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_98_151
timestamp 1606120350
transform 1 0 14996 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1034__C
timestamp 1606120350
transform 1 0 14812 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_154
timestamp 1606120350
transform 1 0 15272 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__D
timestamp 1606120350
transform 1 0 15456 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_923
timestamp 1606120350
transform 1 0 15180 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_98_158
timestamp 1606120350
transform 1 0 15640 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  _0953_
timestamp 1606120350
transform 1 0 17664 0 -1 56032
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _0964_
timestamp 1606120350
transform 1 0 16100 0 -1 56032
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0964__B
timestamp 1606120350
transform 1 0 15916 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0950__A
timestamp 1606120350
transform 1 0 17480 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0947__A
timestamp 1606120350
transform 1 0 17112 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_172
timestamp 1606120350
transform 1 0 16928 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_176
timestamp 1606120350
transform 1 0 17296 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0994_
timestamp 1606120350
transform 1 0 19228 0 -1 56032
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__C
timestamp 1606120350
transform 1 0 19044 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__D
timestamp 1606120350
transform 1 0 18676 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_189
timestamp 1606120350
transform 1 0 18492 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_193
timestamp 1606120350
transform 1 0 18860 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _1028_
timestamp 1606120350
transform 1 0 20884 0 -1 56032
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_924
timestamp 1606120350
transform 1 0 20792 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__C
timestamp 1606120350
transform 1 0 20240 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1011__A
timestamp 1606120350
transform 1 0 21712 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1028__B
timestamp 1606120350
transform 1 0 20608 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_206
timestamp 1606120350
transform 1 0 20056 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_210
timestamp 1606120350
transform 1 0 20424 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_222
timestamp 1606120350
transform 1 0 21528 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_98_226
timestamp 1606120350
transform 1 0 21896 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _0975_
timestamp 1606120350
transform 1 0 24196 0 -1 56032
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_4  _1052_
timestamp 1606120350
transform 1 0 22356 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0975__A2
timestamp 1606120350
transform 1 0 24012 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0980__A1
timestamp 1606120350
transform 1 0 23644 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__A1
timestamp 1606120350
transform 1 0 22172 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_243
timestamp 1606120350
transform 1 0 23460 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_247
timestamp 1606120350
transform 1 0 23828 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__B1
timestamp 1606120350
transform 1 0 25576 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__D
timestamp 1606120350
transform 1 0 25944 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_264
timestamp 1606120350
transform 1 0 25392 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_98_268
timestamp 1606120350
transform 1 0 25760 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_98_272
timestamp 1606120350
transform 1 0 26128 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__inv_8  _0861_
timestamp 1606120350
transform 1 0 26496 0 -1 56032
box -38 -48 866 592
use sky130_fd_sc_hd__inv_8  _0866_
timestamp 1606120350
transform 1 0 28060 0 -1 56032
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_925
timestamp 1606120350
transform 1 0 26404 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0851__A
timestamp 1606120350
transform 1 0 27600 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_98_285
timestamp 1606120350
transform 1 0 27324 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_98_290
timestamp 1606120350
transform 1 0 27784 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_98_302
timestamp 1606120350
transform 1 0 28888 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_314
timestamp 1606120350
transform 1 0 29992 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_926
timestamp 1606120350
transform 1 0 32016 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0937__A1
timestamp 1606120350
transform 1 0 31740 0 -1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_98_326
timestamp 1606120350
transform 1 0 31096 0 -1 56032
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_98_332
timestamp 1606120350
transform 1 0 31648 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_98_335
timestamp 1606120350
transform 1 0 31924 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_337
timestamp 1606120350
transform 1 0 32108 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1195_
timestamp 1606120350
transform 1 0 32844 0 -1 56032
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_98_364
timestamp 1606120350
transform 1 0 34592 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_376
timestamp 1606120350
transform 1 0 35696 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_388
timestamp 1606120350
transform 1 0 36800 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1606120350
transform -1 0 38824 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_927
timestamp 1606120350
transform 1 0 37628 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_98_396
timestamp 1606120350
transform 1 0 37536 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_398
timestamp 1606120350
transform 1 0 37720 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_98_406
timestamp 1606120350
transform 1 0 38456 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1606120350
transform 1 0 1104 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1606120350
transform 1 0 1104 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_99_3
timestamp 1606120350
transform 1 0 1380 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_15
timestamp 1606120350
transform 1 0 2484 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_3
timestamp 1606120350
transform 1 0 1380 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_15
timestamp 1606120350
transform 1 0 2484 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_934
timestamp 1606120350
transform 1 0 3956 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_27
timestamp 1606120350
transform 1 0 3588 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_39
timestamp 1606120350
transform 1 0 4692 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_27
timestamp 1606120350
transform 1 0 3588 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_100_32
timestamp 1606120350
transform 1 0 4048 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_44
timestamp 1606120350
transform 1 0 5152 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_928
timestamp 1606120350
transform 1 0 6716 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_99_51
timestamp 1606120350
transform 1 0 5796 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_59
timestamp 1606120350
transform 1 0 6532 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_99_62
timestamp 1606120350
transform 1 0 6808 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_56
timestamp 1606120350
transform 1 0 6256 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_68
timestamp 1606120350
transform 1 0 7360 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_74
timestamp 1606120350
transform 1 0 7912 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_86
timestamp 1606120350
transform 1 0 9016 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_80
timestamp 1606120350
transform 1 0 8464 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_935
timestamp 1606120350
transform 1 0 9568 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_98
timestamp 1606120350
transform 1 0 10120 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_110
timestamp 1606120350
transform 1 0 11224 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_93
timestamp 1606120350
transform 1 0 9660 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_105
timestamp 1606120350
transform 1 0 10764 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1015_
timestamp 1606120350
transform 1 0 13340 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_929
timestamp 1606120350
transform 1 0 12328 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1015__A
timestamp 1606120350
transform 1 0 13156 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__CLK
timestamp 1606120350
transform 1 0 13616 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_99_123
timestamp 1606120350
transform 1 0 12420 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_136
timestamp 1606120350
transform 1 0 13616 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_100_117
timestamp 1606120350
transform 1 0 11868 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_129
timestamp 1606120350
transform 1 0 12972 0 -1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_135
timestamp 1606120350
transform 1 0 13524 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_100_145
timestamp 1606120350
transform 1 0 14444 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_138
timestamp 1606120350
transform 1 0 13800 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_140
timestamp 1606120350
transform 1 0 13984 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1209__CLK
timestamp 1606120350
transform 1 0 13984 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0994__D
timestamp 1606120350
transform 1 0 14628 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0948__A
timestamp 1606120350
transform 1 0 13800 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1213__D
timestamp 1606120350
transform 1 0 14168 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0948_
timestamp 1606120350
transform 1 0 14168 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_100_154
timestamp 1606120350
transform 1 0 15272 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_100_149
timestamp 1606120350
transform 1 0 14812 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0971__A
timestamp 1606120350
transform 1 0 14996 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_936
timestamp 1606120350
transform 1 0 15180 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1213_
timestamp 1606120350
transform 1 0 14352 0 1 56032
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_4  _1209_
timestamp 1606120350
transform 1 0 15364 0 -1 57120
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  FILLER_99_163
timestamp 1606120350
transform 1 0 16100 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_99_168
timestamp 1606120350
transform 1 0 16560 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__A
timestamp 1606120350
transform 1 0 16376 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_174
timestamp 1606120350
transform 1 0 17112 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__B
timestamp 1606120350
transform 1 0 16744 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0969_
timestamp 1606120350
transform 1 0 16928 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_99_179
timestamp 1606120350
transform 1 0 17572 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_175
timestamp 1606120350
transform 1 0 17204 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0970__A
timestamp 1606120350
transform 1 0 17480 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0969__A
timestamp 1606120350
transform 1 0 17388 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_180
timestamp 1606120350
transform 1 0 17664 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__B1
timestamp 1606120350
transform 1 0 17756 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__D
timestamp 1606120350
transform 1 0 17848 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_191
timestamp 1606120350
transform 1 0 18676 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_187
timestamp 1606120350
transform 1 0 18308 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_192
timestamp 1606120350
transform 1 0 18768 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_99_184
timestamp 1606120350
transform 1 0 18032 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__A
timestamp 1606120350
transform 1 0 18308 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__C
timestamp 1606120350
transform 1 0 18492 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_930
timestamp 1606120350
transform 1 0 17940 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0977_
timestamp 1606120350
transform 1 0 18032 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _0971_
timestamp 1606120350
transform 1 0 18492 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_99_196
timestamp 1606120350
transform 1 0 19136 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__C
timestamp 1606120350
transform 1 0 18860 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1014__B
timestamp 1606120350
transform 1 0 18952 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__B
timestamp 1606120350
transform 1 0 19320 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1014_
timestamp 1606120350
transform 1 0 19044 0 -1 57120
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _1000_
timestamp 1606120350
transform 1 0 19504 0 1 56032
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_100_204
timestamp 1606120350
transform 1 0 19872 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_215
timestamp 1606120350
transform 1 0 20884 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_100_208
timestamp 1606120350
transform 1 0 20240 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_99_213
timestamp 1606120350
transform 1 0 20700 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_209
timestamp 1606120350
transform 1 0 20332 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__A2
timestamp 1606120350
transform 1 0 20884 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0974__A
timestamp 1606120350
transform 1 0 20608 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__D
timestamp 1606120350
transform 1 0 20056 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1000__A
timestamp 1606120350
transform 1 0 20516 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_937
timestamp 1606120350
transform 1 0 20792 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_100_219
timestamp 1606120350
transform 1 0 21252 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_226
timestamp 1606120350
transform 1 0 21896 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__B1
timestamp 1606120350
transform 1 0 22080 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__D
timestamp 1606120350
transform 1 0 21068 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0940_
timestamp 1606120350
transform 1 0 21068 0 1 56032
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _1049_
timestamp 1606120350
transform 1 0 21436 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_237
timestamp 1606120350
transform 1 0 22908 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_233
timestamp 1606120350
transform 1 0 22540 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_239
timestamp 1606120350
transform 1 0 23092 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_99_234
timestamp 1606120350
transform 1 0 22632 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_99_230
timestamp 1606120350
transform 1 0 22264 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1052__B1
timestamp 1606120350
transform 1 0 23092 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1049__A1
timestamp 1606120350
transform 1 0 22448 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__A2
timestamp 1606120350
transform 1 0 22908 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__B1
timestamp 1606120350
transform 1 0 22724 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_248
timestamp 1606120350
transform 1 0 23920 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_99_243
timestamp 1606120350
transform 1 0 23460 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0979__A
timestamp 1606120350
transform 1 0 24104 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1053__A1
timestamp 1606120350
transform 1 0 23276 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_931
timestamp 1606120350
transform 1 0 23552 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0979_
timestamp 1606120350
transform 1 0 23644 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _1053_
timestamp 1606120350
transform 1 0 23276 0 -1 57120
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_100_258
timestamp 1606120350
transform 1 0 24840 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_254
timestamp 1606120350
transform 1 0 24472 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_256
timestamp 1606120350
transform 1 0 24656 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_252
timestamp 1606120350
transform 1 0 24288 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0995__A
timestamp 1606120350
transform 1 0 24472 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__A1
timestamp 1606120350
transform 1 0 24656 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__B1_N
timestamp 1606120350
transform 1 0 25024 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A2
timestamp 1606120350
transform 1 0 24840 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0995_
timestamp 1606120350
transform 1 0 25208 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_100_273
timestamp 1606120350
transform 1 0 26220 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_269
timestamp 1606120350
transform 1 0 25852 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_100_265
timestamp 1606120350
transform 1 0 25484 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_99_273
timestamp 1606120350
transform 1 0 26220 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0911__A1
timestamp 1606120350
transform 1 0 26036 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0940__C
timestamp 1606120350
transform 1 0 25668 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__a21bo_4  _0911_
timestamp 1606120350
transform 1 0 25024 0 1 56032
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_6  FILLER_100_279
timestamp 1606120350
transform 1 0 26772 0 -1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_99_284
timestamp 1606120350
transform 1 0 27232 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_278
timestamp 1606120350
transform 1 0 26680 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0965__A
timestamp 1606120350
transform 1 0 26496 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__B1
timestamp 1606120350
transform 1 0 27048 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__A2
timestamp 1606120350
transform 1 0 27324 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_938
timestamp 1606120350
transform 1 0 26404 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0965_
timestamp 1606120350
transform 1 0 26496 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_100_291
timestamp 1606120350
transform 1 0 27876 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_100_287
timestamp 1606120350
transform 1 0 27508 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__A1
timestamp 1606120350
transform 1 0 27692 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A1
timestamp 1606120350
transform 1 0 27416 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0851_
timestamp 1606120350
transform 1 0 27600 0 1 56032
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_4  _0868_
timestamp 1606120350
transform 1 0 27968 0 -1 57120
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_932
timestamp 1606120350
transform 1 0 29164 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0868__A2
timestamp 1606120350
transform 1 0 28612 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_99_297
timestamp 1606120350
transform 1 0 28428 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_99_301
timestamp 1606120350
transform 1 0 28796 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_99_306
timestamp 1606120350
transform 1 0 29256 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_318
timestamp 1606120350
transform 1 0 30360 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_305
timestamp 1606120350
transform 1 0 29164 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_317
timestamp 1606120350
transform 1 0 30268 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_939
timestamp 1606120350
transform 1 0 32016 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_330
timestamp 1606120350
transform 1 0 31464 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_342
timestamp 1606120350
transform 1 0 32568 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_100_329
timestamp 1606120350
transform 1 0 31372 0 -1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_100_335
timestamp 1606120350
transform 1 0 31924 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_337
timestamp 1606120350
transform 1 0 32108 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_354
timestamp 1606120350
transform 1 0 33672 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_349
timestamp 1606120350
transform 1 0 33212 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_361
timestamp 1606120350
transform 1 0 34316 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_933
timestamp 1606120350
transform 1 0 34776 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__CLK
timestamp 1606120350
transform 1 0 35236 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_99_367
timestamp 1606120350
transform 1 0 34868 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_379
timestamp 1606120350
transform 1 0 35972 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_369
timestamp 1606120350
transform 1 0 35052 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_100_373
timestamp 1606120350
transform 1 0 35420 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_385
timestamp 1606120350
transform 1 0 36524 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1606120350
transform -1 0 38824 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1606120350
transform -1 0 38824 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_940
timestamp 1606120350
transform 1 0 37628 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_391
timestamp 1606120350
transform 1 0 37076 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_403
timestamp 1606120350
transform 1 0 38180 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_100_398
timestamp 1606120350
transform 1 0 37720 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_100_406
timestamp 1606120350
transform 1 0 38456 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1606120350
transform 1 0 1104 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_3
timestamp 1606120350
transform 1 0 1380 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_15
timestamp 1606120350
transform 1 0 2484 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_27
timestamp 1606120350
transform 1 0 3588 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_39
timestamp 1606120350
transform 1 0 4692 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_941
timestamp 1606120350
transform 1 0 6716 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_101_51
timestamp 1606120350
transform 1 0 5796 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_101_59
timestamp 1606120350
transform 1 0 6532 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_101_62
timestamp 1606120350
transform 1 0 6808 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_74
timestamp 1606120350
transform 1 0 7912 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_86
timestamp 1606120350
transform 1 0 9016 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_98
timestamp 1606120350
transform 1 0 10120 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_110
timestamp 1606120350
transform 1 0 11224 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_942
timestamp 1606120350
transform 1 0 12328 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_123
timestamp 1606120350
transform 1 0 12420 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_101_135
timestamp 1606120350
transform 1 0 13524 0 1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1207_
timestamp 1606120350
transform 1 0 15180 0 1 57120
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__D
timestamp 1606120350
transform 1 0 14996 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0963__A
timestamp 1606120350
transform 1 0 14628 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1207__CLK
timestamp 1606120350
transform 1 0 14260 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_145
timestamp 1606120350
transform 1 0 14444 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_149
timestamp 1606120350
transform 1 0 14812 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__A
timestamp 1606120350
transform 1 0 17756 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__D
timestamp 1606120350
transform 1 0 17388 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_172
timestamp 1606120350
transform 1 0 16928 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_176
timestamp 1606120350
transform 1 0 17296 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_179
timestamp 1606120350
transform 1 0 17572 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0970_
timestamp 1606120350
transform 1 0 18124 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _1005_
timestamp 1606120350
transform 1 0 19136 0 1 57120
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_943
timestamp 1606120350
transform 1 0 17940 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__A
timestamp 1606120350
transform 1 0 18952 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1017__B
timestamp 1606120350
transform 1 0 18584 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_101_184
timestamp 1606120350
transform 1 0 18032 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_101_188
timestamp 1606120350
transform 1 0 18400 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_192
timestamp 1606120350
transform 1 0 18768 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_205
timestamp 1606120350
transform 1 0 19964 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0974_
timestamp 1606120350
transform 1 0 20700 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _0989_
timestamp 1606120350
transform 1 0 21712 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__A
timestamp 1606120350
transform 1 0 21160 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1005__B
timestamp 1606120350
transform 1 0 20148 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__B
timestamp 1606120350
transform 1 0 21528 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0973__C
timestamp 1606120350
transform 1 0 20516 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_209
timestamp 1606120350
transform 1 0 20332 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_216
timestamp 1606120350
transform 1 0 20976 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_220
timestamp 1606120350
transform 1 0 21344 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0942_
timestamp 1606120350
transform 1 0 24196 0 1 57120
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_944
timestamp 1606120350
transform 1 0 23552 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0942__A
timestamp 1606120350
transform 1 0 24012 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__A1
timestamp 1606120350
transform 1 0 23000 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0976__A2
timestamp 1606120350
transform 1 0 23368 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_236
timestamp 1606120350
transform 1 0 22816 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_240
timestamp 1606120350
transform 1 0 23184 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_101_245
timestamp 1606120350
transform 1 0 23644 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__inv_8  _0966_
timestamp 1606120350
transform 1 0 25760 0 1 57120
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0966__A
timestamp 1606120350
transform 1 0 25576 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__A2
timestamp 1606120350
transform 1 0 25208 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_260
timestamp 1606120350
transform 1 0 25024 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_264
timestamp 1606120350
transform 1 0 25392 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _0855_
timestamp 1606120350
transform 1 0 27324 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__A2
timestamp 1606120350
transform 1 0 27140 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__B1
timestamp 1606120350
transform 1 0 26772 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_277
timestamp 1606120350
transform 1 0 26588 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_281
timestamp 1606120350
transform 1 0 26956 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__inv_8  _0864_
timestamp 1606120350
transform 1 0 29256 0 1 57120
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_945
timestamp 1606120350
transform 1 0 29164 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0867__B1
timestamp 1606120350
transform 1 0 28612 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0864__A
timestamp 1606120350
transform 1 0 28980 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_297
timestamp 1606120350
transform 1 0 28428 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_301
timestamp 1606120350
transform 1 0 28796 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_101_315
timestamp 1606120350
transform 1 0 30084 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_327
timestamp 1606120350
transform 1 0 31188 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_339
timestamp 1606120350
transform 1 0 32292 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_351
timestamp 1606120350
transform 1 0 33396 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_101_363
timestamp 1606120350
transform 1 0 34500 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1162_
timestamp 1606120350
transform 1 0 35236 0 1 57120
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_946
timestamp 1606120350
transform 1 0 34776 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1162__D
timestamp 1606120350
transform 1 0 35052 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_101_367
timestamp 1606120350
transform 1 0 34868 0 1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1606120350
transform -1 0 38824 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_390
timestamp 1606120350
transform 1 0 36984 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_402
timestamp 1606120350
transform 1 0 38088 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_101_406
timestamp 1606120350
transform 1 0 38456 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_204
timestamp 1606120350
transform 1 0 1104 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__D
timestamp 1606120350
transform 1 0 1564 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_102_3
timestamp 1606120350
transform 1 0 1380 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_102_7
timestamp 1606120350
transform 1 0 1748 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_19
timestamp 1606120350
transform 1 0 2852 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_947
timestamp 1606120350
transform 1 0 3956 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_32
timestamp 1606120350
transform 1 0 4048 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_44
timestamp 1606120350
transform 1 0 5152 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_56
timestamp 1606120350
transform 1 0 6256 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_68
timestamp 1606120350
transform 1 0 7360 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_80
timestamp 1606120350
transform 1 0 8464 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_948
timestamp 1606120350
transform 1 0 9568 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_93
timestamp 1606120350
transform 1 0 9660 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_105
timestamp 1606120350
transform 1 0 10764 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_117
timestamp 1606120350
transform 1 0 11868 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_129
timestamp 1606120350
transform 1 0 12972 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0963_
timestamp 1606120350
transform 1 0 15456 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_949
timestamp 1606120350
transform 1 0 15180 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_102_141
timestamp 1606120350
transform 1 0 14076 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_102_154
timestamp 1606120350
transform 1 0 15272 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_102_159
timestamp 1606120350
transform 1 0 15732 0 -1 58208
box -38 -48 590 592
use sky130_fd_sc_hd__inv_8  _0950_
timestamp 1606120350
transform 1 0 17480 0 -1 58208
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _1006_
timestamp 1606120350
transform 1 0 16468 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__D
timestamp 1606120350
transform 1 0 17296 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1006__A
timestamp 1606120350
transform 1 0 16928 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0977__A
timestamp 1606120350
transform 1 0 16284 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_102_170
timestamp 1606120350
transform 1 0 16744 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_102_174
timestamp 1606120350
transform 1 0 17112 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1017_
timestamp 1606120350
transform 1 0 19044 0 -1 58208
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__A
timestamp 1606120350
transform 1 0 18860 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__C
timestamp 1606120350
transform 1 0 18492 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_102_187
timestamp 1606120350
transform 1 0 18308 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_102_191
timestamp 1606120350
transform 1 0 18676 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_102_204
timestamp 1606120350
transform 1 0 19872 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0973_
timestamp 1606120350
transform 1 0 20884 0 -1 58208
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_950
timestamp 1606120350
transform 1 0 20792 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__D
timestamp 1606120350
transform 1 0 20608 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__D
timestamp 1606120350
transform 1 0 20056 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__A2
timestamp 1606120350
transform 1 0 21896 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_102_208
timestamp 1606120350
transform 1 0 20240 0 -1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_102_224
timestamp 1606120350
transform 1 0 21712 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_102_228
timestamp 1606120350
transform 1 0 22080 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _0976_
timestamp 1606120350
transform 1 0 22540 0 -1 58208
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0989__A1
timestamp 1606120350
transform 1 0 22264 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__A2
timestamp 1606120350
transform 1 0 23920 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_102_232
timestamp 1606120350
transform 1 0 22448 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_102_246
timestamp 1606120350
transform 1 0 23736 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_102_250
timestamp 1606120350
transform 1 0 24104 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1012_
timestamp 1606120350
transform 1 0 24472 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__A1
timestamp 1606120350
transform 1 0 26220 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1012__B1
timestamp 1606120350
transform 1 0 24288 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__B1
timestamp 1606120350
transform 1 0 25760 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_102_266
timestamp 1606120350
transform 1 0 25576 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_102_270
timestamp 1606120350
transform 1 0 25944 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _0867_
timestamp 1606120350
transform 1 0 27600 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_951
timestamp 1606120350
transform 1 0 26404 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__A1
timestamp 1606120350
transform 1 0 26864 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0855__A1
timestamp 1606120350
transform 1 0 27324 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_102_276
timestamp 1606120350
transform 1 0 26496 0 -1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_102_282
timestamp 1606120350
transform 1 0 27048 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_102_287
timestamp 1606120350
transform 1 0 27508 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__A1
timestamp 1606120350
transform 1 0 28888 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_102_300
timestamp 1606120350
transform 1 0 28704 0 -1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_102_304
timestamp 1606120350
transform 1 0 29072 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_316
timestamp 1606120350
transform 1 0 30176 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_952
timestamp 1606120350
transform 1 0 32016 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_102_328
timestamp 1606120350
transform 1 0 31280 0 -1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_102_337
timestamp 1606120350
transform 1 0 32108 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_349
timestamp 1606120350
transform 1 0 33212 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_361
timestamp 1606120350
transform 1 0 34316 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_373
timestamp 1606120350
transform 1 0 35420 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_102_385
timestamp 1606120350
transform 1 0 36524 0 -1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_205
timestamp 1606120350
transform -1 0 38824 0 -1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_953
timestamp 1606120350
transform 1 0 37628 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_102_398
timestamp 1606120350
transform 1 0 37720 0 -1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_102_406
timestamp 1606120350
transform 1 0 38456 0 -1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1206_
timestamp 1606120350
transform 1 0 1564 0 1 58208
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_206
timestamp 1606120350
transform 1 0 1104 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_103_3
timestamp 1606120350
transform 1 0 1380 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_103_24
timestamp 1606120350
transform 1 0 3312 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_36
timestamp 1606120350
transform 1 0 4416 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_954
timestamp 1606120350
transform 1 0 6716 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_48
timestamp 1606120350
transform 1 0 5520 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_103_60
timestamp 1606120350
transform 1 0 6624 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_62
timestamp 1606120350
transform 1 0 6808 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_74
timestamp 1606120350
transform 1 0 7912 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_86
timestamp 1606120350
transform 1 0 9016 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_98
timestamp 1606120350
transform 1 0 10120 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_110
timestamp 1606120350
transform 1 0 11224 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_955
timestamp 1606120350
transform 1 0 12328 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_103_123
timestamp 1606120350
transform 1 0 12420 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_135
timestamp 1606120350
transform 1 0 13524 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_147
timestamp 1606120350
transform 1 0 14628 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_103_159
timestamp 1606120350
transform 1 0 15732 0 1 58208
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _0981_
timestamp 1606120350
transform 1 0 16928 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0981__A
timestamp 1606120350
transform 1 0 17388 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__B
timestamp 1606120350
transform 1 0 17756 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__A
timestamp 1606120350
transform 1 0 16744 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0956__A
timestamp 1606120350
transform 1 0 16376 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_103_165
timestamp 1606120350
transform 1 0 16284 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_103_168
timestamp 1606120350
transform 1 0 16560 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_103_175
timestamp 1606120350
transform 1 0 17204 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_103_179
timestamp 1606120350
transform 1 0 17572 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _1021_
timestamp 1606120350
transform 1 0 18860 0 1 58208
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_956
timestamp 1606120350
transform 1 0 17940 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__B
timestamp 1606120350
transform 1 0 19872 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__B
timestamp 1606120350
transform 1 0 18676 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0978__A
timestamp 1606120350
transform 1 0 18308 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_103_184
timestamp 1606120350
transform 1 0 18032 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_103_189
timestamp 1606120350
transform 1 0 18492 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_103_202
timestamp 1606120350
transform 1 0 19688 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1019_
timestamp 1606120350
transform 1 0 21160 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__B
timestamp 1606120350
transform 1 0 20884 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__C
timestamp 1606120350
transform 1 0 20516 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_103_206
timestamp 1606120350
transform 1 0 20056 0 1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_210
timestamp 1606120350
transform 1 0 20424 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_103_213
timestamp 1606120350
transform 1 0 20700 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_103_217
timestamp 1606120350
transform 1 0 21068 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _1050_
timestamp 1606120350
transform 1 0 23736 0 1 58208
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_957
timestamp 1606120350
transform 1 0 23552 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__A1
timestamp 1606120350
transform 1 0 23368 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A1
timestamp 1606120350
transform 1 0 22448 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__A2
timestamp 1606120350
transform 1 0 22816 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_103_230
timestamp 1606120350
transform 1 0 22264 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_103_234
timestamp 1606120350
transform 1 0 22632 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_103_238
timestamp 1606120350
transform 1 0 23000 0 1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_245
timestamp 1606120350
transform 1 0 23644 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0941_
timestamp 1606120350
transform 1 0 25668 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__A2
timestamp 1606120350
transform 1 0 26312 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0941__A
timestamp 1606120350
transform 1 0 25484 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1051__A1
timestamp 1606120350
transform 1 0 25116 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_103_259
timestamp 1606120350
transform 1 0 24932 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_103_263
timestamp 1606120350
transform 1 0 25300 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_103_270
timestamp 1606120350
transform 1 0 25944 0 1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _0856_
timestamp 1606120350
transform 1 0 26864 0 1 58208
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__A2
timestamp 1606120350
transform 1 0 26680 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0856__B1
timestamp 1606120350
transform 1 0 28244 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_103_276
timestamp 1606120350
transform 1 0 26496 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_103_293
timestamp 1606120350
transform 1 0 28060 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_958
timestamp 1606120350
transform 1 0 29164 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__B1_N
timestamp 1606120350
transform 1 0 28888 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0925__A2
timestamp 1606120350
transform 1 0 29440 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_103_297
timestamp 1606120350
transform 1 0 28428 0 1 58208
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_103_301
timestamp 1606120350
transform 1 0 28796 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_103_304
timestamp 1606120350
transform 1 0 29072 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_103_306
timestamp 1606120350
transform 1 0 29256 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_103_310
timestamp 1606120350
transform 1 0 29624 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_322
timestamp 1606120350
transform 1 0 30728 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_334
timestamp 1606120350
transform 1 0 31832 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_346
timestamp 1606120350
transform 1 0 32936 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_103_358
timestamp 1606120350
transform 1 0 34040 0 1 58208
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_959
timestamp 1606120350
transform 1 0 34776 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__D
timestamp 1606120350
transform 1 0 35144 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1225__CLK
timestamp 1606120350
transform 1 0 35512 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_103_367
timestamp 1606120350
transform 1 0 34868 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_103_372
timestamp 1606120350
transform 1 0 35328 0 1 58208
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_103_376
timestamp 1606120350
transform 1 0 35696 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_103_388
timestamp 1606120350
transform 1 0 36800 0 1 58208
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_207
timestamp 1606120350
transform -1 0 38824 0 1 58208
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_103_400
timestamp 1606120350
transform 1 0 37904 0 1 58208
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_103_406
timestamp 1606120350
transform 1 0 38456 0 1 58208
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_208
timestamp 1606120350
transform 1 0 1104 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1206__CLK
timestamp 1606120350
transform 1 0 1564 0 -1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_104_3
timestamp 1606120350
transform 1 0 1380 0 -1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_104_7
timestamp 1606120350
transform 1 0 1748 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_19
timestamp 1606120350
transform 1 0 2852 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_960
timestamp 1606120350
transform 1 0 3956 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_32
timestamp 1606120350
transform 1 0 4048 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_44
timestamp 1606120350
transform 1 0 5152 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_56
timestamp 1606120350
transform 1 0 6256 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_68
timestamp 1606120350
transform 1 0 7360 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_80
timestamp 1606120350
transform 1 0 8464 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_961
timestamp 1606120350
transform 1 0 9568 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_93
timestamp 1606120350
transform 1 0 9660 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_105
timestamp 1606120350
transform 1 0 10764 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_117
timestamp 1606120350
transform 1 0 11868 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_129
timestamp 1606120350
transform 1 0 12972 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_962
timestamp 1606120350
transform 1 0 15180 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_141
timestamp 1606120350
transform 1 0 14076 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_154
timestamp 1606120350
transform 1 0 15272 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _0956_
timestamp 1606120350
transform 1 0 16652 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _1024_
timestamp 1606120350
transform 1 0 17664 0 -1 59296
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1024__C
timestamp 1606120350
transform 1 0 17480 0 -1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__D
timestamp 1606120350
transform 1 0 17112 0 -1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_104_166
timestamp 1606120350
transform 1 0 16376 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_104_172
timestamp 1606120350
transform 1 0 16928 0 -1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_104_176
timestamp 1606120350
transform 1 0 17296 0 -1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0978_
timestamp 1606120350
transform 1 0 19228 0 -1 59296
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1021__C
timestamp 1606120350
transform 1 0 18860 0 -1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_104_189
timestamp 1606120350
transform 1 0 18492 0 -1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_104_195
timestamp 1606120350
transform 1 0 19044 0 -1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0991_
timestamp 1606120350
transform 1 0 20884 0 -1 59296
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_963
timestamp 1606120350
transform 1 0 20792 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0991__A
timestamp 1606120350
transform 1 0 20608 0 -1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__A1
timestamp 1606120350
transform 1 0 21896 0 -1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__A2
timestamp 1606120350
transform 1 0 20240 0 -1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_104_206
timestamp 1606120350
transform 1 0 20056 0 -1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_104_210
timestamp 1606120350
transform 1 0 20424 0 -1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_104_224
timestamp 1606120350
transform 1 0 21712 0 -1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_104_228
timestamp 1606120350
transform 1 0 22080 0 -1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _0990_
timestamp 1606120350
transform 1 0 22448 0 -1 59296
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__D
timestamp 1606120350
transform 1 0 23920 0 -1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__B1
timestamp 1606120350
transform 1 0 22264 0 -1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_104_245
timestamp 1606120350
transform 1 0 23644 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_104_250
timestamp 1606120350
transform 1 0 24104 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _1051_
timestamp 1606120350
transform 1 0 24380 0 -1 59296
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0862__B1
timestamp 1606120350
transform 1 0 26220 0 -1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_104_266
timestamp 1606120350
transform 1 0 25576 0 -1 59296
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_104_272
timestamp 1606120350
transform 1 0 26128 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _0862_
timestamp 1606120350
transform 1 0 26496 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_964
timestamp 1606120350
transform 1 0 26404 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_288
timestamp 1606120350
transform 1 0 27600 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__a21bo_4  _0925_
timestamp 1606120350
transform 1 0 28888 0 -1 59296
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_104_300
timestamp 1606120350
transform 1 0 28704 0 -1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_104_315
timestamp 1606120350
transform 1 0 30084 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_965
timestamp 1606120350
transform 1 0 32016 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_104_327
timestamp 1606120350
transform 1 0 31188 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_104_335
timestamp 1606120350
transform 1 0 31924 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_104_337
timestamp 1606120350
transform 1 0 32108 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_104_349
timestamp 1606120350
transform 1 0 33212 0 -1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_104_361
timestamp 1606120350
transform 1 0 34316 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _1225_
timestamp 1606120350
transform 1 0 35144 0 -1 59296
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_104_369
timestamp 1606120350
transform 1 0 35052 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_209
timestamp 1606120350
transform -1 0 38824 0 -1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_966
timestamp 1606120350
transform 1 0 37628 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_104_389
timestamp 1606120350
transform 1 0 36892 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_104_398
timestamp 1606120350
transform 1 0 37720 0 -1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_104_406
timestamp 1606120350
transform 1 0 38456 0 -1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_210
timestamp 1606120350
transform 1 0 1104 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_212
timestamp 1606120350
transform 1 0 1104 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_105_3
timestamp 1606120350
transform 1 0 1380 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_15
timestamp 1606120350
transform 1 0 2484 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_3
timestamp 1606120350
transform 1 0 1380 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_15
timestamp 1606120350
transform 1 0 2484 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_973
timestamp 1606120350
transform 1 0 3956 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_27
timestamp 1606120350
transform 1 0 3588 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_39
timestamp 1606120350
transform 1 0 4692 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_27
timestamp 1606120350
transform 1 0 3588 0 -1 60384
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_106_32
timestamp 1606120350
transform 1 0 4048 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_44
timestamp 1606120350
transform 1 0 5152 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_967
timestamp 1606120350
transform 1 0 6716 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_105_51
timestamp 1606120350
transform 1 0 5796 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_105_59
timestamp 1606120350
transform 1 0 6532 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_105_62
timestamp 1606120350
transform 1 0 6808 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_56
timestamp 1606120350
transform 1 0 6256 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_68
timestamp 1606120350
transform 1 0 7360 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_74
timestamp 1606120350
transform 1 0 7912 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_86
timestamp 1606120350
transform 1 0 9016 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_80
timestamp 1606120350
transform 1 0 8464 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_974
timestamp 1606120350
transform 1 0 9568 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_98
timestamp 1606120350
transform 1 0 10120 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_110
timestamp 1606120350
transform 1 0 11224 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_93
timestamp 1606120350
transform 1 0 9660 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_105
timestamp 1606120350
transform 1 0 10764 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_968
timestamp 1606120350
transform 1 0 12328 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_123
timestamp 1606120350
transform 1 0 12420 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_135
timestamp 1606120350
transform 1 0 13524 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_117
timestamp 1606120350
transform 1 0 11868 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_129
timestamp 1606120350
transform 1 0 12972 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_975
timestamp 1606120350
transform 1 0 15180 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_147
timestamp 1606120350
transform 1 0 14628 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_159
timestamp 1606120350
transform 1 0 15732 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_141
timestamp 1606120350
transform 1 0 14076 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_154
timestamp 1606120350
transform 1 0 15272 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__A1
timestamp 1606120350
transform 1 0 17756 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_105_171
timestamp 1606120350
transform 1 0 16836 0 1 59296
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_105_179
timestamp 1606120350
transform 1 0 17572 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_106_166
timestamp 1606120350
transform 1 0 16376 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_178
timestamp 1606120350
transform 1 0 17480 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_106_192
timestamp 1606120350
transform 1 0 18768 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_106_188
timestamp 1606120350
transform 1 0 18400 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_105_193
timestamp 1606120350
transform 1 0 18860 0 1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_105_184
timestamp 1606120350
transform 1 0 18032 0 1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__B1
timestamp 1606120350
transform 1 0 18216 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0992__A
timestamp 1606120350
transform 1 0 18584 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__B
timestamp 1606120350
transform 1 0 18400 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_969
timestamp 1606120350
transform 1 0 17940 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _0992_
timestamp 1606120350
transform 1 0 18584 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_105_199
timestamp 1606120350
transform 1 0 19412 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__A
timestamp 1606120350
transform 1 0 19044 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__C
timestamp 1606120350
transform 1 0 19228 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _0982_
timestamp 1606120350
transform 1 0 19228 0 -1 60384
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_4  _1057_
timestamp 1606120350
transform 1 0 19596 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_106_210
timestamp 1606120350
transform 1 0 20424 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_106_206
timestamp 1606120350
transform 1 0 20056 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_213
timestamp 1606120350
transform 1 0 20700 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1057__A2
timestamp 1606120350
transform 1 0 20240 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__A1
timestamp 1606120350
transform 1 0 20608 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0982__D
timestamp 1606120350
transform 1 0 20884 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_976
timestamp 1606120350
transform 1 0 20792 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_106_228
timestamp 1606120350
transform 1 0 22080 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_217
timestamp 1606120350
transform 1 0 21068 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__A1
timestamp 1606120350
transform 1 0 21252 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _1062_
timestamp 1606120350
transform 1 0 20884 0 -1 60384
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _0993_
timestamp 1606120350
transform 1 0 21436 0 1 59296
box -38 -48 1234 592
use sky130_fd_sc_hd__fill_2  FILLER_106_239
timestamp 1606120350
transform 1 0 23092 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_106_232
timestamp 1606120350
transform 1 0 22448 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_238
timestamp 1606120350
transform 1 0 23000 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_234
timestamp 1606120350
transform 1 0 22632 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__A2
timestamp 1606120350
transform 1 0 22632 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0993__A2
timestamp 1606120350
transform 1 0 22264 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0983__A
timestamp 1606120350
transform 1 0 22816 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _0983_
timestamp 1606120350
transform 1 0 22816 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_106_248
timestamp 1606120350
transform 1 0 23920 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_106_243
timestamp 1606120350
transform 1 0 23460 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_105_245
timestamp 1606120350
transform 1 0 23644 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_105_242
timestamp 1606120350
transform 1 0 23368 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1062__B1
timestamp 1606120350
transform 1 0 23276 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__B1
timestamp 1606120350
transform 1 0 24104 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1050__A2
timestamp 1606120350
transform 1 0 23736 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0990__B1
timestamp 1606120350
transform 1 0 23184 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_970
timestamp 1606120350
transform 1 0 23552 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1186_
timestamp 1606120350
transform 1 0 23920 0 1 59296
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_6  FILLER_106_256
timestamp 1606120350
transform 1 0 24656 0 -1 60384
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_106_252
timestamp 1606120350
transform 1 0 24288 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1186__CLK
timestamp 1606120350
transform 1 0 24472 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_106_264
timestamp 1606120350
transform 1 0 25392 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_105_267
timestamp 1606120350
transform 1 0 25668 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__A2
timestamp 1606120350
transform 1 0 25208 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_106_272
timestamp 1606120350
transform 1 0 26128 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_105_271
timestamp 1606120350
transform 1 0 26036 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A1
timestamp 1606120350
transform 1 0 25852 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__A2
timestamp 1606120350
transform 1 0 26220 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_106_276
timestamp 1606120350
transform 1 0 26496 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_977
timestamp 1606120350
transform 1 0 26404 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__inv_8  _0857_
timestamp 1606120350
transform 1 0 26588 0 -1 60384
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_105_296
timestamp 1606120350
transform 1 0 28336 0 1 59296
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_105_292
timestamp 1606120350
transform 1 0 27968 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_105_288
timestamp 1606120350
transform 1 0 27600 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0857__A
timestamp 1606120350
transform 1 0 28152 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0863__B1
timestamp 1606120350
transform 1 0 27784 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_106_286
timestamp 1606120350
transform 1 0 27416 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_4  _0863_
timestamp 1606120350
transform 1 0 26404 0 1 59296
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  FILLER_106_306
timestamp 1606120350
transform 1 0 29256 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_106_298
timestamp 1606120350
transform 1 0 28520 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_105_306
timestamp 1606120350
transform 1 0 29256 0 1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_105_302
timestamp 1606120350
transform 1 0 28888 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_2_3_0_clk_A
timestamp 1606120350
transform 1 0 28980 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_971
timestamp 1606120350
transform 1 0 29164 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_106_318
timestamp 1606120350
transform 1 0 30360 0 -1 60384
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_106_312
timestamp 1606120350
transform 1 0 29808 0 -1 60384
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_105_312
timestamp 1606120350
transform 1 0 29808 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__A1
timestamp 1606120350
transform 1 0 29624 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__A2
timestamp 1606120350
transform 1 0 30176 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0928__B1_N
timestamp 1606120350
transform 1 0 29992 0 1 59296
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_2_3_0_clk
timestamp 1606120350
transform 1 0 29532 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_4  _0928_
timestamp 1606120350
transform 1 0 30176 0 1 59296
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_978
timestamp 1606120350
transform 1 0 32016 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__CLK
timestamp 1606120350
transform 1 0 30912 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_105_329
timestamp 1606120350
transform 1 0 31372 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_341
timestamp 1606120350
transform 1 0 32476 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_106_326
timestamp 1606120350
transform 1 0 31096 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_106_334
timestamp 1606120350
transform 1 0 31832 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_106_337
timestamp 1606120350
transform 1 0 32108 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_353
timestamp 1606120350
transform 1 0 33580 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_105_365
timestamp 1606120350
transform 1 0 34684 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_106_349
timestamp 1606120350
transform 1 0 33212 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_106_361
timestamp 1606120350
transform 1 0 34316 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_972
timestamp 1606120350
transform 1 0 34776 0 1 59296
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__CLK
timestamp 1606120350
transform 1 0 35788 0 -1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_105_367
timestamp 1606120350
transform 1 0 34868 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_105_379
timestamp 1606120350
transform 1 0 35972 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_106_373
timestamp 1606120350
transform 1 0 35420 0 -1 60384
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_106_379
timestamp 1606120350
transform 1 0 35972 0 -1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_211
timestamp 1606120350
transform -1 0 38824 0 1 59296
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_213
timestamp 1606120350
transform -1 0 38824 0 -1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_979
timestamp 1606120350
transform 1 0 37628 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_105_391
timestamp 1606120350
transform 1 0 37076 0 1 59296
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_105_403
timestamp 1606120350
transform 1 0 38180 0 1 59296
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_106_391
timestamp 1606120350
transform 1 0 37076 0 -1 60384
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_106_398
timestamp 1606120350
transform 1 0 37720 0 -1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_106_406
timestamp 1606120350
transform 1 0 38456 0 -1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_214
timestamp 1606120350
transform 1 0 1104 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_107_3
timestamp 1606120350
transform 1 0 1380 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_15
timestamp 1606120350
transform 1 0 2484 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_27
timestamp 1606120350
transform 1 0 3588 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_39
timestamp 1606120350
transform 1 0 4692 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_980
timestamp 1606120350
transform 1 0 6716 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_107_51
timestamp 1606120350
transform 1 0 5796 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_107_59
timestamp 1606120350
transform 1 0 6532 0 1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_107_62
timestamp 1606120350
transform 1 0 6808 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_74
timestamp 1606120350
transform 1 0 7912 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_86
timestamp 1606120350
transform 1 0 9016 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_10_0_clk_A
timestamp 1606120350
transform 1 0 10764 0 1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_107_98
timestamp 1606120350
transform 1 0 10120 0 1 60384
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_107_104
timestamp 1606120350
transform 1 0 10672 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_107_107
timestamp 1606120350
transform 1 0 10948 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_981
timestamp 1606120350
transform 1 0 12328 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_107_119
timestamp 1606120350
transform 1 0 12052 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_107_123
timestamp 1606120350
transform 1 0 12420 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_135
timestamp 1606120350
transform 1 0 13524 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_147
timestamp 1606120350
transform 1 0 14628 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_159
timestamp 1606120350
transform 1 0 15732 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_171
timestamp 1606120350
transform 1 0 16836 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1022_
timestamp 1606120350
transform 1 0 18768 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  _1060_
timestamp 1606120350
transform 1 0 19780 0 1 60384
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_982
timestamp 1606120350
transform 1 0 17940 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__A1
timestamp 1606120350
transform 1 0 19596 0 1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1018__A
timestamp 1606120350
transform 1 0 19228 0 1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1022__A
timestamp 1606120350
transform 1 0 18584 0 1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_107_184
timestamp 1606120350
transform 1 0 18032 0 1 60384
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_107_195
timestamp 1606120350
transform 1 0 19044 0 1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_107_199
timestamp 1606120350
transform 1 0 19412 0 1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__o21a_4  _1061_
timestamp 1606120350
transform 1 0 21712 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__A1
timestamp 1606120350
transform 1 0 21160 0 1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1019__B1
timestamp 1606120350
transform 1 0 21528 0 1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_107_216
timestamp 1606120350
transform 1 0 20976 0 1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_107_220
timestamp 1606120350
transform 1 0 21344 0 1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_983
timestamp 1606120350
transform 1 0 23552 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__A1
timestamp 1606120350
transform 1 0 23000 0 1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__B1
timestamp 1606120350
transform 1 0 23368 0 1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_107_236
timestamp 1606120350
transform 1 0 22816 0 1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_107_240
timestamp 1606120350
transform 1 0 23184 0 1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_107_245
timestamp 1606120350
transform 1 0 23644 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__a21bo_4  _0927_
timestamp 1606120350
transform 1 0 25208 0 1 60384
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__B1_N
timestamp 1606120350
transform 1 0 25024 0 1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_107_257
timestamp 1606120350
transform 1 0 24748 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_107_275
timestamp 1606120350
transform 1 0 26404 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_107_287
timestamp 1606120350
transform 1 0 27508 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_984
timestamp 1606120350
transform 1 0 29164 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_107_299
timestamp 1606120350
transform 1 0 28612 0 1 60384
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_107_306
timestamp 1606120350
transform 1 0 29256 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_107_318
timestamp 1606120350
transform 1 0 30360 0 1 60384
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1187_
timestamp 1606120350
transform 1 0 30912 0 1 60384
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1187__D
timestamp 1606120350
transform 1 0 30728 0 1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_107_343
timestamp 1606120350
transform 1 0 32660 0 1 60384
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_107_355
timestamp 1606120350
transform 1 0 33764 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_107_363
timestamp 1606120350
transform 1 0 34500 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1185_
timestamp 1606120350
transform 1 0 35788 0 1 60384
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_985
timestamp 1606120350
transform 1 0 34776 0 1 60384
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1185__D
timestamp 1606120350
transform 1 0 35604 0 1 60384
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_107_367
timestamp 1606120350
transform 1 0 34868 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_215
timestamp 1606120350
transform -1 0 38824 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_107_396
timestamp 1606120350
transform 1 0 37536 0 1 60384
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_107_404
timestamp 1606120350
transform 1 0 38272 0 1 60384
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_216
timestamp 1606120350
transform 1 0 1104 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_108_3
timestamp 1606120350
transform 1 0 1380 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_15
timestamp 1606120350
transform 1 0 2484 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_986
timestamp 1606120350
transform 1 0 3956 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_108_27
timestamp 1606120350
transform 1 0 3588 0 -1 61472
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_108_32
timestamp 1606120350
transform 1 0 4048 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_44
timestamp 1606120350
transform 1 0 5152 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_56
timestamp 1606120350
transform 1 0 6256 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_68
timestamp 1606120350
transform 1 0 7360 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_80
timestamp 1606120350
transform 1 0 8464 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_987
timestamp 1606120350
transform 1 0 9568 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_10_0_clk
timestamp 1606120350
transform 1 0 10764 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_108_93
timestamp 1606120350
transform 1 0 9660 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_108
timestamp 1606120350
transform 1 0 11040 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_120
timestamp 1606120350
transform 1 0 12144 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_132
timestamp 1606120350
transform 1 0 13248 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_988
timestamp 1606120350
transform 1 0 15180 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_144
timestamp 1606120350
transform 1 0 14352 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_152
timestamp 1606120350
transform 1 0 15088 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_154
timestamp 1606120350
transform 1 0 15272 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_166
timestamp 1606120350
transform 1 0 16376 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_178
timestamp 1606120350
transform 1 0 17480 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_1  _1018_
timestamp 1606120350
transform 1 0 19688 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__A2
timestamp 1606120350
transform 1 0 19504 0 -1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_108_190
timestamp 1606120350
transform 1 0 18584 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_108_198
timestamp 1606120350
transform 1 0 19320 0 -1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_108_205
timestamp 1606120350
transform 1 0 19964 0 -1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__o21ai_4  _1058_
timestamp 1606120350
transform 1 0 21068 0 -1 61472
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_989
timestamp 1606120350
transform 1 0 20792 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__A2
timestamp 1606120350
transform 1 0 20608 0 -1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1060__B1
timestamp 1606120350
transform 1 0 20148 0 -1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_108_209
timestamp 1606120350
transform 1 0 20332 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_108_215
timestamp 1606120350
transform 1 0 20884 0 -1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1061__A2
timestamp 1606120350
transform 1 0 22448 0 -1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_108_230
timestamp 1606120350
transform 1 0 22264 0 -1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_108_234
timestamp 1606120350
transform 1 0 22632 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_246
timestamp 1606120350
transform 1 0 23736 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0927__A1
timestamp 1606120350
transform 1 0 25208 0 -1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_108_258
timestamp 1606120350
transform 1 0 24840 0 -1 61472
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_108_264
timestamp 1606120350
transform 1 0 25392 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_108_272
timestamp 1606120350
transform 1 0 26128 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_990
timestamp 1606120350
transform 1 0 26404 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_276
timestamp 1606120350
transform 1 0 26496 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_288
timestamp 1606120350
transform 1 0 27600 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_300
timestamp 1606120350
transform 1 0 28704 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_312
timestamp 1606120350
transform 1 0 29808 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_991
timestamp 1606120350
transform 1 0 32016 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_108_324
timestamp 1606120350
transform 1 0 30912 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_337
timestamp 1606120350
transform 1 0 32108 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_349
timestamp 1606120350
transform 1 0 33212 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_361
timestamp 1606120350
transform 1 0 34316 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_373
timestamp 1606120350
transform 1 0 35420 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_108_385
timestamp 1606120350
transform 1 0 36524 0 -1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_217
timestamp 1606120350
transform -1 0 38824 0 -1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_992
timestamp 1606120350
transform 1 0 37628 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_108_398
timestamp 1606120350
transform 1 0 37720 0 -1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_108_406
timestamp 1606120350
transform 1 0 38456 0 -1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_218
timestamp 1606120350
transform 1 0 1104 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_109_3
timestamp 1606120350
transform 1 0 1380 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_15
timestamp 1606120350
transform 1 0 2484 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_27
timestamp 1606120350
transform 1 0 3588 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_39
timestamp 1606120350
transform 1 0 4692 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_993
timestamp 1606120350
transform 1 0 6716 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_109_51
timestamp 1606120350
transform 1 0 5796 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_109_59
timestamp 1606120350
transform 1 0 6532 0 1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_109_62
timestamp 1606120350
transform 1 0 6808 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_74
timestamp 1606120350
transform 1 0 7912 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_86
timestamp 1606120350
transform 1 0 9016 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_98
timestamp 1606120350
transform 1 0 10120 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_110
timestamp 1606120350
transform 1 0 11224 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_994
timestamp 1606120350
transform 1 0 12328 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_5_0_clk
timestamp 1606120350
transform 1 0 13156 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_5_0_clk_A
timestamp 1606120350
transform 1 0 13616 0 1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_109_123
timestamp 1606120350
transform 1 0 12420 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_109_134
timestamp 1606120350
transform 1 0 13432 0 1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_109_138
timestamp 1606120350
transform 1 0 13800 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_150
timestamp 1606120350
transform 1 0 14904 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_162
timestamp 1606120350
transform 1 0 16008 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_174
timestamp 1606120350
transform 1 0 17112 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_109_182
timestamp 1606120350
transform 1 0 17848 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_995
timestamp 1606120350
transform 1 0 17940 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__A1
timestamp 1606120350
transform 1 0 18216 0 1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__A2
timestamp 1606120350
transform 1 0 18584 0 1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1073__B1
timestamp 1606120350
transform 1 0 18952 0 1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_109_184
timestamp 1606120350
transform 1 0 18032 0 1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_109_188
timestamp 1606120350
transform 1 0 18400 0 1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_109_192
timestamp 1606120350
transform 1 0 18768 0 1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_109_196
timestamp 1606120350
transform 1 0 19136 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1058__B1
timestamp 1606120350
transform 1 0 21068 0 1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_109_208
timestamp 1606120350
transform 1 0 20240 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_109_216
timestamp 1606120350
transform 1 0 20976 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_219
timestamp 1606120350
transform 1 0 21252 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_996
timestamp 1606120350
transform 1 0 23552 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_231
timestamp 1606120350
transform 1 0 22356 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_109_243
timestamp 1606120350
transform 1 0 23460 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_245
timestamp 1606120350
transform 1 0 23644 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_257
timestamp 1606120350
transform 1 0 24748 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_109_269
timestamp 1606120350
transform 1 0 25852 0 1 61472
box -38 -48 590 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__D
timestamp 1606120350
transform 1 0 26496 0 1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1170__CLK
timestamp 1606120350
transform 1 0 26864 0 1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_109_275
timestamp 1606120350
transform 1 0 26404 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_109_278
timestamp 1606120350
transform 1 0 26680 0 1 61472
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_109_282
timestamp 1606120350
transform 1 0 27048 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_109_294
timestamp 1606120350
transform 1 0 28152 0 1 61472
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_997
timestamp 1606120350
transform 1 0 29164 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_109_302
timestamp 1606120350
transform 1 0 28888 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_109_306
timestamp 1606120350
transform 1 0 29256 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_318
timestamp 1606120350
transform 1 0 30360 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_330
timestamp 1606120350
transform 1 0 31464 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_342
timestamp 1606120350
transform 1 0 32568 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_354
timestamp 1606120350
transform 1 0 33672 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_998
timestamp 1606120350
transform 1 0 34776 0 1 61472
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_109_367
timestamp 1606120350
transform 1 0 34868 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_109_379
timestamp 1606120350
transform 1 0 35972 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_219
timestamp 1606120350
transform -1 0 38824 0 1 61472
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_109_391
timestamp 1606120350
transform 1 0 37076 0 1 61472
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_109_403
timestamp 1606120350
transform 1 0 38180 0 1 61472
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_220
timestamp 1606120350
transform 1 0 1104 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_110_3
timestamp 1606120350
transform 1 0 1380 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_15
timestamp 1606120350
transform 1 0 2484 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_999
timestamp 1606120350
transform 1 0 3956 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_110_27
timestamp 1606120350
transform 1 0 3588 0 -1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_110_32
timestamp 1606120350
transform 1 0 4048 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_44
timestamp 1606120350
transform 1 0 5152 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_56
timestamp 1606120350
transform 1 0 6256 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_68
timestamp 1606120350
transform 1 0 7360 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_80
timestamp 1606120350
transform 1 0 8464 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1000
timestamp 1606120350
transform 1 0 9568 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_93
timestamp 1606120350
transform 1 0 9660 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_105
timestamp 1606120350
transform 1 0 10764 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_117
timestamp 1606120350
transform 1 0 11868 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_129
timestamp 1606120350
transform 1 0 12972 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1001
timestamp 1606120350
transform 1 0 15180 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_141
timestamp 1606120350
transform 1 0 14076 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_154
timestamp 1606120350
transform 1 0 15272 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_166
timestamp 1606120350
transform 1 0 16376 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_178
timestamp 1606120350
transform 1 0 17480 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _1073_
timestamp 1606120350
transform 1 0 18216 0 -1 62560
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_110_199
timestamp 1606120350
transform 1 0 19412 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1002
timestamp 1606120350
transform 1 0 20792 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__B1
timestamp 1606120350
transform 1 0 21160 0 -1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__B1
timestamp 1606120350
transform 1 0 21528 0 -1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__A2
timestamp 1606120350
transform 1 0 21896 0 -1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_110_211
timestamp 1606120350
transform 1 0 20516 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_110_215
timestamp 1606120350
transform 1 0 20884 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_110_220
timestamp 1606120350
transform 1 0 21344 0 -1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_110_224
timestamp 1606120350
transform 1 0 21712 0 -1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_110_228
timestamp 1606120350
transform 1 0 22080 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_240
timestamp 1606120350
transform 1 0 23184 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_252
timestamp 1606120350
transform 1 0 24288 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_110_264
timestamp 1606120350
transform 1 0 25392 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_110_272
timestamp 1606120350
transform 1 0 26128 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_4  _1170_
timestamp 1606120350
transform 1 0 26496 0 -1 62560
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1003
timestamp 1606120350
transform 1 0 26404 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_295
timestamp 1606120350
transform 1 0 28244 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_307
timestamp 1606120350
transform 1 0 29348 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_319
timestamp 1606120350
transform 1 0 30452 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1004
timestamp 1606120350
transform 1 0 32016 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_110_331
timestamp 1606120350
transform 1 0 31556 0 -1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_110_335
timestamp 1606120350
transform 1 0 31924 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_110_337
timestamp 1606120350
transform 1 0 32108 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_349
timestamp 1606120350
transform 1 0 33212 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_361
timestamp 1606120350
transform 1 0 34316 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_373
timestamp 1606120350
transform 1 0 35420 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_110_385
timestamp 1606120350
transform 1 0 36524 0 -1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_221
timestamp 1606120350
transform -1 0 38824 0 -1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1005
timestamp 1606120350
transform 1 0 37628 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_110_398
timestamp 1606120350
transform 1 0 37720 0 -1 62560
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_110_406
timestamp 1606120350
transform 1 0 38456 0 -1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_222
timestamp 1606120350
transform 1 0 1104 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_111_3
timestamp 1606120350
transform 1 0 1380 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_15
timestamp 1606120350
transform 1 0 2484 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1158__D
timestamp 1606120350
transform 1 0 4692 0 1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1158__CLK
timestamp 1606120350
transform 1 0 5060 0 1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_111_27
timestamp 1606120350
transform 1 0 3588 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_111_41
timestamp 1606120350
transform 1 0 4876 0 1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_111_45
timestamp 1606120350
transform 1 0 5244 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1006
timestamp 1606120350
transform 1 0 6716 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_111_57
timestamp 1606120350
transform 1 0 6348 0 1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_111_62
timestamp 1606120350
transform 1 0 6808 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_74
timestamp 1606120350
transform 1 0 7912 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_86
timestamp 1606120350
transform 1 0 9016 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_98
timestamp 1606120350
transform 1 0 10120 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_110
timestamp 1606120350
transform 1 0 11224 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1007
timestamp 1606120350
transform 1 0 12328 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_123
timestamp 1606120350
transform 1 0 12420 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_135
timestamp 1606120350
transform 1 0 13524 0 1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_11_0_clk_A
timestamp 1606120350
transform 1 0 13892 0 1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_111_141
timestamp 1606120350
transform 1 0 14076 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_153
timestamp 1606120350
transform 1 0 15180 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_165
timestamp 1606120350
transform 1 0 16284 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_111_177
timestamp 1606120350
transform 1 0 17388 0 1 62560
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _1072_
timestamp 1606120350
transform 1 0 18676 0 1 62560
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1008
timestamp 1606120350
transform 1 0 17940 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__A1
timestamp 1606120350
transform 1 0 18492 0 1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_111_184
timestamp 1606120350
transform 1 0 18032 0 1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_111_188
timestamp 1606120350
transform 1 0 18400 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_111_204
timestamp 1606120350
transform 1 0 19872 0 1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_4  _1023_
timestamp 1606120350
transform 1 0 21160 0 1 62560
box -38 -48 1234 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1023__A1
timestamp 1606120350
transform 1 0 20976 0 1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__A1
timestamp 1606120350
transform 1 0 20608 0 1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1020__A2
timestamp 1606120350
transform 1 0 20240 0 1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_111_210
timestamp 1606120350
transform 1 0 20424 0 1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_111_214
timestamp 1606120350
transform 1 0 20792 0 1 62560
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1009
timestamp 1606120350
transform 1 0 23552 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_231
timestamp 1606120350
transform 1 0 22356 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_111_243
timestamp 1606120350
transform 1 0 23460 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_245
timestamp 1606120350
transform 1 0 23644 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_257
timestamp 1606120350
transform 1 0 24748 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_269
timestamp 1606120350
transform 1 0 25852 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_281
timestamp 1606120350
transform 1 0 26956 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_293
timestamp 1606120350
transform 1 0 28060 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1010
timestamp 1606120350
transform 1 0 29164 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_306
timestamp 1606120350
transform 1 0 29256 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_318
timestamp 1606120350
transform 1 0 30360 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_330
timestamp 1606120350
transform 1 0 31464 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_342
timestamp 1606120350
transform 1 0 32568 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_354
timestamp 1606120350
transform 1 0 33672 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1011
timestamp 1606120350
transform 1 0 34776 0 1 62560
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_111_367
timestamp 1606120350
transform 1 0 34868 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_111_379
timestamp 1606120350
transform 1 0 35972 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_223
timestamp 1606120350
transform -1 0 38824 0 1 62560
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_111_391
timestamp 1606120350
transform 1 0 37076 0 1 62560
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_111_403
timestamp 1606120350
transform 1 0 38180 0 1 62560
box -38 -48 406 592
use sky130_fd_sc_hd__dfxtp_4  _1193_
timestamp 1606120350
transform 1 0 1564 0 1 63648
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_224
timestamp 1606120350
transform 1 0 1104 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_226
timestamp 1606120350
transform 1 0 1104 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__D
timestamp 1606120350
transform 1 0 1564 0 -1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_112_3
timestamp 1606120350
transform 1 0 1380 0 -1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_112_7
timestamp 1606120350
transform 1 0 1748 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_19
timestamp 1606120350
transform 1 0 2852 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_113_3
timestamp 1606120350
transform 1 0 1380 0 1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_113_28
timestamp 1606120350
transform 1 0 3680 0 1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_113_24
timestamp 1606120350
transform 1 0 3312 0 1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_112_32
timestamp 1606120350
transform 1 0 4048 0 -1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__A1
timestamp 1606120350
transform 1 0 4232 0 -1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__A2
timestamp 1606120350
transform 1 0 3496 0 1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0935__B1_N
timestamp 1606120350
transform 1 0 3864 0 1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1012
timestamp 1606120350
transform 1 0 3956 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_112_36
timestamp 1606120350
transform 1 0 4416 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_113_45
timestamp 1606120350
transform 1 0 5244 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1158_
timestamp 1606120350
transform 1 0 4692 0 -1 63648
box -38 -48 1786 592
use sky130_fd_sc_hd__a21bo_4  _0935_
timestamp 1606120350
transform 1 0 4048 0 1 63648
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1019
timestamp 1606120350
transform 1 0 6716 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_58
timestamp 1606120350
transform 1 0 6440 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_113_57
timestamp 1606120350
transform 1 0 6348 0 1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_113_62
timestamp 1606120350
transform 1 0 6808 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_70
timestamp 1606120350
transform 1 0 7544 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_82
timestamp 1606120350
transform 1 0 8648 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_112_90
timestamp 1606120350
transform 1 0 9384 0 -1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_113_74
timestamp 1606120350
transform 1 0 7912 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_86
timestamp 1606120350
transform 1 0 9016 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1013
timestamp 1606120350
transform 1 0 9568 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_93
timestamp 1606120350
transform 1 0 9660 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_105
timestamp 1606120350
transform 1 0 10764 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_98
timestamp 1606120350
transform 1 0 10120 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_110
timestamp 1606120350
transform 1 0 11224 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1020
timestamp 1606120350
transform 1 0 12328 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_117
timestamp 1606120350
transform 1 0 11868 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_129
timestamp 1606120350
transform 1 0 12972 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_112_137
timestamp 1606120350
transform 1 0 13708 0 -1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_113_123
timestamp 1606120350
transform 1 0 12420 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_135
timestamp 1606120350
transform 1 0 13524 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1014
timestamp 1606120350
transform 1 0 15180 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_11_0_clk
timestamp 1606120350
transform 1 0 13892 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_112_142
timestamp 1606120350
transform 1 0 14168 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_112_150
timestamp 1606120350
transform 1 0 14904 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_112_154
timestamp 1606120350
transform 1 0 15272 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_147
timestamp 1606120350
transform 1 0 14628 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_159
timestamp 1606120350
transform 1 0 15732 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_166
timestamp 1606120350
transform 1 0 16376 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_178
timestamp 1606120350
transform 1 0 17480 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_171
timestamp 1606120350
transform 1 0 16836 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1021
timestamp 1606120350
transform 1 0 17940 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__A2
timestamp 1606120350
transform 1 0 18676 0 -1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1072__B1
timestamp 1606120350
transform 1 0 19044 0 -1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_112_190
timestamp 1606120350
transform 1 0 18584 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_112_193
timestamp 1606120350
transform 1 0 18860 0 -1 63648
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_112_197
timestamp 1606120350
transform 1 0 19228 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_184
timestamp 1606120350
transform 1 0 18032 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_196
timestamp 1606120350
transform 1 0 19136 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__o21ai_4  _1020_
timestamp 1606120350
transform 1 0 20884 0 -1 63648
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1015
timestamp 1606120350
transform 1 0 20792 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_112_209
timestamp 1606120350
transform 1 0 20332 0 -1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_112_213
timestamp 1606120350
transform 1 0 20700 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_228
timestamp 1606120350
transform 1 0 22080 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_208
timestamp 1606120350
transform 1 0 20240 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_220
timestamp 1606120350
transform 1 0 21344 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1022
timestamp 1606120350
transform 1 0 23552 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_240
timestamp 1606120350
transform 1 0 23184 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_232
timestamp 1606120350
transform 1 0 22448 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_245
timestamp 1606120350
transform 1 0 23644 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_252
timestamp 1606120350
transform 1 0 24288 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_112_264
timestamp 1606120350
transform 1 0 25392 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_112_272
timestamp 1606120350
transform 1 0 26128 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_113_257
timestamp 1606120350
transform 1 0 24748 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_269
timestamp 1606120350
transform 1 0 25852 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1016
timestamp 1606120350
transform 1 0 26404 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_276
timestamp 1606120350
transform 1 0 26496 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_288
timestamp 1606120350
transform 1 0 27600 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_281
timestamp 1606120350
transform 1 0 26956 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_293
timestamp 1606120350
transform 1 0 28060 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1023
timestamp 1606120350
transform 1 0 29164 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_300
timestamp 1606120350
transform 1 0 28704 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_312
timestamp 1606120350
transform 1 0 29808 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_306
timestamp 1606120350
transform 1 0 29256 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_318
timestamp 1606120350
transform 1 0 30360 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1017
timestamp 1606120350
transform 1 0 32016 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_324
timestamp 1606120350
transform 1 0 30912 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_337
timestamp 1606120350
transform 1 0 32108 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_330
timestamp 1606120350
transform 1 0 31464 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_342
timestamp 1606120350
transform 1 0 32568 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_349
timestamp 1606120350
transform 1 0 33212 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_361
timestamp 1606120350
transform 1 0 34316 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_354
timestamp 1606120350
transform 1 0 33672 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1024
timestamp 1606120350
transform 1 0 34776 0 1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_112_373
timestamp 1606120350
transform 1 0 35420 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_112_385
timestamp 1606120350
transform 1 0 36524 0 -1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_367
timestamp 1606120350
transform 1 0 34868 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_113_379
timestamp 1606120350
transform 1 0 35972 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_225
timestamp 1606120350
transform -1 0 38824 0 -1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_227
timestamp 1606120350
transform -1 0 38824 0 1 63648
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1018
timestamp 1606120350
transform 1 0 37628 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_112_398
timestamp 1606120350
transform 1 0 37720 0 -1 63648
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_112_406
timestamp 1606120350
transform 1 0 38456 0 -1 63648
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_113_391
timestamp 1606120350
transform 1 0 37076 0 1 63648
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_113_403
timestamp 1606120350
transform 1 0 38180 0 1 63648
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_228
timestamp 1606120350
transform 1 0 1104 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1193__CLK
timestamp 1606120350
transform 1 0 1564 0 -1 64736
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_114_3
timestamp 1606120350
transform 1 0 1380 0 -1 64736
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_114_7
timestamp 1606120350
transform 1 0 1748 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_19
timestamp 1606120350
transform 1 0 2852 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1025
timestamp 1606120350
transform 1 0 3956 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_32
timestamp 1606120350
transform 1 0 4048 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_44
timestamp 1606120350
transform 1 0 5152 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_56
timestamp 1606120350
transform 1 0 6256 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_68
timestamp 1606120350
transform 1 0 7360 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_80
timestamp 1606120350
transform 1 0 8464 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1026
timestamp 1606120350
transform 1 0 9568 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_93
timestamp 1606120350
transform 1 0 9660 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_105
timestamp 1606120350
transform 1 0 10764 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_117
timestamp 1606120350
transform 1 0 11868 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_129
timestamp 1606120350
transform 1 0 12972 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1027
timestamp 1606120350
transform 1 0 15180 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_141
timestamp 1606120350
transform 1 0 14076 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_154
timestamp 1606120350
transform 1 0 15272 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_166
timestamp 1606120350
transform 1 0 16376 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_178
timestamp 1606120350
transform 1 0 17480 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_190
timestamp 1606120350
transform 1 0 18584 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_202
timestamp 1606120350
transform 1 0 19688 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1028
timestamp 1606120350
transform 1 0 20792 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_215
timestamp 1606120350
transform 1 0 20884 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_227
timestamp 1606120350
transform 1 0 21988 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_239
timestamp 1606120350
transform 1 0 23092 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_251
timestamp 1606120350
transform 1 0 24196 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_263
timestamp 1606120350
transform 1 0 25300 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1029
timestamp 1606120350
transform 1 0 26404 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_276
timestamp 1606120350
transform 1 0 26496 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_288
timestamp 1606120350
transform 1 0 27600 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_300
timestamp 1606120350
transform 1 0 28704 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_312
timestamp 1606120350
transform 1 0 29808 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1030
timestamp 1606120350
transform 1 0 32016 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_114_324
timestamp 1606120350
transform 1 0 30912 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_337
timestamp 1606120350
transform 1 0 32108 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_349
timestamp 1606120350
transform 1 0 33212 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_361
timestamp 1606120350
transform 1 0 34316 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_373
timestamp 1606120350
transform 1 0 35420 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_114_385
timestamp 1606120350
transform 1 0 36524 0 -1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_229
timestamp 1606120350
transform -1 0 38824 0 -1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1031
timestamp 1606120350
transform 1 0 37628 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_114_398
timestamp 1606120350
transform 1 0 37720 0 -1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_114_406
timestamp 1606120350
transform 1 0 38456 0 -1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1221_
timestamp 1606120350
transform 1 0 1748 0 1 64736
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_3  PHY_230
timestamp 1606120350
transform 1 0 1104 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__D
timestamp 1606120350
transform 1 0 1564 0 1 64736
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_115_3
timestamp 1606120350
transform 1 0 1380 0 1 64736
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_115_26
timestamp 1606120350
transform 1 0 3496 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_38
timestamp 1606120350
transform 1 0 4600 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1032
timestamp 1606120350
transform 1 0 6716 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_115_50
timestamp 1606120350
transform 1 0 5704 0 1 64736
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_115_58
timestamp 1606120350
transform 1 0 6440 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_115_62
timestamp 1606120350
transform 1 0 6808 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_74
timestamp 1606120350
transform 1 0 7912 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_86
timestamp 1606120350
transform 1 0 9016 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_98
timestamp 1606120350
transform 1 0 10120 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_110
timestamp 1606120350
transform 1 0 11224 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1033
timestamp 1606120350
transform 1 0 12328 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_123
timestamp 1606120350
transform 1 0 12420 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_135
timestamp 1606120350
transform 1 0 13524 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_147
timestamp 1606120350
transform 1 0 14628 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_159
timestamp 1606120350
transform 1 0 15732 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_171
timestamp 1606120350
transform 1 0 16836 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1034
timestamp 1606120350
transform 1 0 17940 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_184
timestamp 1606120350
transform 1 0 18032 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_196
timestamp 1606120350
transform 1 0 19136 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_208
timestamp 1606120350
transform 1 0 20240 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_220
timestamp 1606120350
transform 1 0 21344 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1035
timestamp 1606120350
transform 1 0 23552 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_232
timestamp 1606120350
transform 1 0 22448 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_245
timestamp 1606120350
transform 1 0 23644 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_257
timestamp 1606120350
transform 1 0 24748 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_269
timestamp 1606120350
transform 1 0 25852 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_281
timestamp 1606120350
transform 1 0 26956 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_293
timestamp 1606120350
transform 1 0 28060 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1036
timestamp 1606120350
transform 1 0 29164 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_306
timestamp 1606120350
transform 1 0 29256 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_318
timestamp 1606120350
transform 1 0 30360 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_330
timestamp 1606120350
transform 1 0 31464 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_342
timestamp 1606120350
transform 1 0 32568 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_354
timestamp 1606120350
transform 1 0 33672 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1037
timestamp 1606120350
transform 1 0 34776 0 1 64736
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_115_367
timestamp 1606120350
transform 1 0 34868 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_115_379
timestamp 1606120350
transform 1 0 35972 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_231
timestamp 1606120350
transform -1 0 38824 0 1 64736
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_115_391
timestamp 1606120350
transform 1 0 37076 0 1 64736
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_115_403
timestamp 1606120350
transform 1 0 38180 0 1 64736
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_232
timestamp 1606120350
transform 1 0 1104 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1221__CLK
timestamp 1606120350
transform 1 0 1748 0 -1 65824
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_116_3
timestamp 1606120350
transform 1 0 1380 0 -1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_116_9
timestamp 1606120350
transform 1 0 1932 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_116_21
timestamp 1606120350
transform 1 0 3036 0 -1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1038
timestamp 1606120350
transform 1 0 3956 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_116_29
timestamp 1606120350
transform 1 0 3772 0 -1 65824
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_116_32
timestamp 1606120350
transform 1 0 4048 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_44
timestamp 1606120350
transform 1 0 5152 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_56
timestamp 1606120350
transform 1 0 6256 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_68
timestamp 1606120350
transform 1 0 7360 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_80
timestamp 1606120350
transform 1 0 8464 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1039
timestamp 1606120350
transform 1 0 9568 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_93
timestamp 1606120350
transform 1 0 9660 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_105
timestamp 1606120350
transform 1 0 10764 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_117
timestamp 1606120350
transform 1 0 11868 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_129
timestamp 1606120350
transform 1 0 12972 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1040
timestamp 1606120350
transform 1 0 15180 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_141
timestamp 1606120350
transform 1 0 14076 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_154
timestamp 1606120350
transform 1 0 15272 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_166
timestamp 1606120350
transform 1 0 16376 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_178
timestamp 1606120350
transform 1 0 17480 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_190
timestamp 1606120350
transform 1 0 18584 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_202
timestamp 1606120350
transform 1 0 19688 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1041
timestamp 1606120350
transform 1 0 20792 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_215
timestamp 1606120350
transform 1 0 20884 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_227
timestamp 1606120350
transform 1 0 21988 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_239
timestamp 1606120350
transform 1 0 23092 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_251
timestamp 1606120350
transform 1 0 24196 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_263
timestamp 1606120350
transform 1 0 25300 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1042
timestamp 1606120350
transform 1 0 26404 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_276
timestamp 1606120350
transform 1 0 26496 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_288
timestamp 1606120350
transform 1 0 27600 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_300
timestamp 1606120350
transform 1 0 28704 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_312
timestamp 1606120350
transform 1 0 29808 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1043
timestamp 1606120350
transform 1 0 32016 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_116_324
timestamp 1606120350
transform 1 0 30912 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_337
timestamp 1606120350
transform 1 0 32108 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_349
timestamp 1606120350
transform 1 0 33212 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_361
timestamp 1606120350
transform 1 0 34316 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_373
timestamp 1606120350
transform 1 0 35420 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_116_385
timestamp 1606120350
transform 1 0 36524 0 -1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_233
timestamp 1606120350
transform -1 0 38824 0 -1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1044
timestamp 1606120350
transform 1 0 37628 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_116_398
timestamp 1606120350
transform 1 0 37720 0 -1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_116_406
timestamp 1606120350
transform 1 0 38456 0 -1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_234
timestamp 1606120350
transform 1 0 1104 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_117_3
timestamp 1606120350
transform 1 0 1380 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_15
timestamp 1606120350
transform 1 0 2484 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_27
timestamp 1606120350
transform 1 0 3588 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_39
timestamp 1606120350
transform 1 0 4692 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1045
timestamp 1606120350
transform 1 0 6716 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_117_51
timestamp 1606120350
transform 1 0 5796 0 1 65824
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_117_59
timestamp 1606120350
transform 1 0 6532 0 1 65824
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_117_62
timestamp 1606120350
transform 1 0 6808 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_74
timestamp 1606120350
transform 1 0 7912 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_86
timestamp 1606120350
transform 1 0 9016 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_98
timestamp 1606120350
transform 1 0 10120 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_110
timestamp 1606120350
transform 1 0 11224 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1046
timestamp 1606120350
transform 1 0 12328 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_123
timestamp 1606120350
transform 1 0 12420 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_135
timestamp 1606120350
transform 1 0 13524 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_147
timestamp 1606120350
transform 1 0 14628 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_159
timestamp 1606120350
transform 1 0 15732 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_171
timestamp 1606120350
transform 1 0 16836 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1047
timestamp 1606120350
transform 1 0 17940 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_184
timestamp 1606120350
transform 1 0 18032 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_196
timestamp 1606120350
transform 1 0 19136 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_208
timestamp 1606120350
transform 1 0 20240 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_220
timestamp 1606120350
transform 1 0 21344 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1048
timestamp 1606120350
transform 1 0 23552 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_232
timestamp 1606120350
transform 1 0 22448 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_245
timestamp 1606120350
transform 1 0 23644 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_257
timestamp 1606120350
transform 1 0 24748 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_269
timestamp 1606120350
transform 1 0 25852 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_281
timestamp 1606120350
transform 1 0 26956 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_293
timestamp 1606120350
transform 1 0 28060 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1049
timestamp 1606120350
transform 1 0 29164 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_306
timestamp 1606120350
transform 1 0 29256 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_318
timestamp 1606120350
transform 1 0 30360 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_330
timestamp 1606120350
transform 1 0 31464 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_342
timestamp 1606120350
transform 1 0 32568 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_354
timestamp 1606120350
transform 1 0 33672 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1050
timestamp 1606120350
transform 1 0 34776 0 1 65824
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_117_367
timestamp 1606120350
transform 1 0 34868 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_117_379
timestamp 1606120350
transform 1 0 35972 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_235
timestamp 1606120350
transform -1 0 38824 0 1 65824
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_117_391
timestamp 1606120350
transform 1 0 37076 0 1 65824
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_117_403
timestamp 1606120350
transform 1 0 38180 0 1 65824
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_236
timestamp 1606120350
transform 1 0 1104 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_238
timestamp 1606120350
transform 1 0 1104 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_118_3
timestamp 1606120350
transform 1 0 1380 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_15
timestamp 1606120350
transform 1 0 2484 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_3
timestamp 1606120350
transform 1 0 1380 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_15
timestamp 1606120350
transform 1 0 2484 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1051
timestamp 1606120350
transform 1 0 3956 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_118_27
timestamp 1606120350
transform 1 0 3588 0 -1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_118_32
timestamp 1606120350
transform 1 0 4048 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_44
timestamp 1606120350
transform 1 0 5152 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_27
timestamp 1606120350
transform 1 0 3588 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_39
timestamp 1606120350
transform 1 0 4692 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1058
timestamp 1606120350
transform 1 0 6716 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_56
timestamp 1606120350
transform 1 0 6256 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_68
timestamp 1606120350
transform 1 0 7360 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_51
timestamp 1606120350
transform 1 0 5796 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_119_59
timestamp 1606120350
transform 1 0 6532 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_119_62
timestamp 1606120350
transform 1 0 6808 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_80
timestamp 1606120350
transform 1 0 8464 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_74
timestamp 1606120350
transform 1 0 7912 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_86
timestamp 1606120350
transform 1 0 9016 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1052
timestamp 1606120350
transform 1 0 9568 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_93
timestamp 1606120350
transform 1 0 9660 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_105
timestamp 1606120350
transform 1 0 10764 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_98
timestamp 1606120350
transform 1 0 10120 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_110
timestamp 1606120350
transform 1 0 11224 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1059
timestamp 1606120350
transform 1 0 12328 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_117
timestamp 1606120350
transform 1 0 11868 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_129
timestamp 1606120350
transform 1 0 12972 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_123
timestamp 1606120350
transform 1 0 12420 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_135
timestamp 1606120350
transform 1 0 13524 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1053
timestamp 1606120350
transform 1 0 15180 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_141
timestamp 1606120350
transform 1 0 14076 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_154
timestamp 1606120350
transform 1 0 15272 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_147
timestamp 1606120350
transform 1 0 14628 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_159
timestamp 1606120350
transform 1 0 15732 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_166
timestamp 1606120350
transform 1 0 16376 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_178
timestamp 1606120350
transform 1 0 17480 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_171
timestamp 1606120350
transform 1 0 16836 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1060
timestamp 1606120350
transform 1 0 17940 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_190
timestamp 1606120350
transform 1 0 18584 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_202
timestamp 1606120350
transform 1 0 19688 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_184
timestamp 1606120350
transform 1 0 18032 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_196
timestamp 1606120350
transform 1 0 19136 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1054
timestamp 1606120350
transform 1 0 20792 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_215
timestamp 1606120350
transform 1 0 20884 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_227
timestamp 1606120350
transform 1 0 21988 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_208
timestamp 1606120350
transform 1 0 20240 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_220
timestamp 1606120350
transform 1 0 21344 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1061
timestamp 1606120350
transform 1 0 23552 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_239
timestamp 1606120350
transform 1 0 23092 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_251
timestamp 1606120350
transform 1 0 24196 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_232
timestamp 1606120350
transform 1 0 22448 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_245
timestamp 1606120350
transform 1 0 23644 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_263
timestamp 1606120350
transform 1 0 25300 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_257
timestamp 1606120350
transform 1 0 24748 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_119_269
timestamp 1606120350
transform 1 0 25852 0 1 66912
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1055
timestamp 1606120350
transform 1 0 26404 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_3_7_0_clk
timestamp 1606120350
transform 1 0 26404 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_3_7_0_clk_A
timestamp 1606120350
transform 1 0 26864 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_118_276
timestamp 1606120350
transform 1 0 26496 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_288
timestamp 1606120350
transform 1 0 27600 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_119_278
timestamp 1606120350
transform 1 0 26680 0 1 66912
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_119_282
timestamp 1606120350
transform 1 0 27048 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_119_294
timestamp 1606120350
transform 1 0 28152 0 1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1062
timestamp 1606120350
transform 1 0 29164 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_300
timestamp 1606120350
transform 1 0 28704 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_312
timestamp 1606120350
transform 1 0 29808 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_119_302
timestamp 1606120350
transform 1 0 28888 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_119_306
timestamp 1606120350
transform 1 0 29256 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_318
timestamp 1606120350
transform 1 0 30360 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1056
timestamp 1606120350
transform 1 0 32016 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_324
timestamp 1606120350
transform 1 0 30912 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_337
timestamp 1606120350
transform 1 0 32108 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_330
timestamp 1606120350
transform 1 0 31464 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_342
timestamp 1606120350
transform 1 0 32568 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_349
timestamp 1606120350
transform 1 0 33212 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_361
timestamp 1606120350
transform 1 0 34316 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_354
timestamp 1606120350
transform 1 0 33672 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1063
timestamp 1606120350
transform 1 0 34776 0 1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_118_373
timestamp 1606120350
transform 1 0 35420 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_118_385
timestamp 1606120350
transform 1 0 36524 0 -1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_367
timestamp 1606120350
transform 1 0 34868 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_119_379
timestamp 1606120350
transform 1 0 35972 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_237
timestamp 1606120350
transform -1 0 38824 0 -1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_239
timestamp 1606120350
transform -1 0 38824 0 1 66912
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1057
timestamp 1606120350
transform 1 0 37628 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_118_398
timestamp 1606120350
transform 1 0 37720 0 -1 66912
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_118_406
timestamp 1606120350
transform 1 0 38456 0 -1 66912
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_119_391
timestamp 1606120350
transform 1 0 37076 0 1 66912
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_119_403
timestamp 1606120350
transform 1 0 38180 0 1 66912
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_240
timestamp 1606120350
transform 1 0 1104 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_120_3
timestamp 1606120350
transform 1 0 1380 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_15
timestamp 1606120350
transform 1 0 2484 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1064
timestamp 1606120350
transform 1 0 3956 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_120_27
timestamp 1606120350
transform 1 0 3588 0 -1 68000
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_120_32
timestamp 1606120350
transform 1 0 4048 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_44
timestamp 1606120350
transform 1 0 5152 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_56
timestamp 1606120350
transform 1 0 6256 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_68
timestamp 1606120350
transform 1 0 7360 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_80
timestamp 1606120350
transform 1 0 8464 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1065
timestamp 1606120350
transform 1 0 9568 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_93
timestamp 1606120350
transform 1 0 9660 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_105
timestamp 1606120350
transform 1 0 10764 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_117
timestamp 1606120350
transform 1 0 11868 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_129
timestamp 1606120350
transform 1 0 12972 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1066
timestamp 1606120350
transform 1 0 15180 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_141
timestamp 1606120350
transform 1 0 14076 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_154
timestamp 1606120350
transform 1 0 15272 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_166
timestamp 1606120350
transform 1 0 16376 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_178
timestamp 1606120350
transform 1 0 17480 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_190
timestamp 1606120350
transform 1 0 18584 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_202
timestamp 1606120350
transform 1 0 19688 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1067
timestamp 1606120350
transform 1 0 20792 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_215
timestamp 1606120350
transform 1 0 20884 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_227
timestamp 1606120350
transform 1 0 21988 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__CLK
timestamp 1606120350
transform 1 0 24012 0 -1 68000
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_120_239
timestamp 1606120350
transform 1 0 23092 0 -1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_120_247
timestamp 1606120350
transform 1 0 23828 0 -1 68000
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_120_251
timestamp 1606120350
transform 1 0 24196 0 -1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_14_0_clk_A
timestamp 1606120350
transform 1 0 25024 0 -1 68000
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_120_259
timestamp 1606120350
transform 1 0 24932 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_262
timestamp 1606120350
transform 1 0 25208 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_120_274
timestamp 1606120350
transform 1 0 26312 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1068
timestamp 1606120350
transform 1 0 26404 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_276
timestamp 1606120350
transform 1 0 26496 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_288
timestamp 1606120350
transform 1 0 27600 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_300
timestamp 1606120350
transform 1 0 28704 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_312
timestamp 1606120350
transform 1 0 29808 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1069
timestamp 1606120350
transform 1 0 32016 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_120_324
timestamp 1606120350
transform 1 0 30912 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_337
timestamp 1606120350
transform 1 0 32108 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_349
timestamp 1606120350
transform 1 0 33212 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_361
timestamp 1606120350
transform 1 0 34316 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_373
timestamp 1606120350
transform 1 0 35420 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_120_385
timestamp 1606120350
transform 1 0 36524 0 -1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_241
timestamp 1606120350
transform -1 0 38824 0 -1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1070
timestamp 1606120350
transform 1 0 37628 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_120_398
timestamp 1606120350
transform 1 0 37720 0 -1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_120_406
timestamp 1606120350
transform 1 0 38456 0 -1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_242
timestamp 1606120350
transform 1 0 1104 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_121_3
timestamp 1606120350
transform 1 0 1380 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_15
timestamp 1606120350
transform 1 0 2484 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_27
timestamp 1606120350
transform 1 0 3588 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_39
timestamp 1606120350
transform 1 0 4692 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1071
timestamp 1606120350
transform 1 0 6716 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_121_51
timestamp 1606120350
transform 1 0 5796 0 1 68000
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_121_59
timestamp 1606120350
transform 1 0 6532 0 1 68000
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_121_62
timestamp 1606120350
transform 1 0 6808 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_74
timestamp 1606120350
transform 1 0 7912 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_86
timestamp 1606120350
transform 1 0 9016 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_98
timestamp 1606120350
transform 1 0 10120 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_110
timestamp 1606120350
transform 1 0 11224 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1072
timestamp 1606120350
transform 1 0 12328 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_123
timestamp 1606120350
transform 1 0 12420 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_135
timestamp 1606120350
transform 1 0 13524 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_147
timestamp 1606120350
transform 1 0 14628 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_159
timestamp 1606120350
transform 1 0 15732 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_171
timestamp 1606120350
transform 1 0 16836 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1073
timestamp 1606120350
transform 1 0 17940 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_184
timestamp 1606120350
transform 1 0 18032 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_196
timestamp 1606120350
transform 1 0 19136 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_208
timestamp 1606120350
transform 1 0 20240 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_220
timestamp 1606120350
transform 1 0 21344 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_121_239
timestamp 1606120350
transform 1 0 23092 0 1 68000
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_121_235
timestamp 1606120350
transform 1 0 22724 0 1 68000
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_121_232
timestamp 1606120350
transform 1 0 22448 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1181__CLK
timestamp 1606120350
transform 1 0 22908 0 1 68000
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1181__D
timestamp 1606120350
transform 1 0 22540 0 1 68000
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_121_245
timestamp 1606120350
transform 1 0 23644 0 1 68000
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_121_243
timestamp 1606120350
transform 1 0 23460 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1159__D
timestamp 1606120350
transform 1 0 23828 0 1 68000
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1074
timestamp 1606120350
transform 1 0 23552 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__dfxtp_4  _1159_
timestamp 1606120350
transform 1 0 24012 0 1 68000
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_12  FILLER_121_268
timestamp 1606120350
transform 1 0 25760 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_280
timestamp 1606120350
transform 1 0 26864 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_292
timestamp 1606120350
transform 1 0 27968 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1075
timestamp 1606120350
transform 1 0 29164 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_121_304
timestamp 1606120350
transform 1 0 29072 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_306
timestamp 1606120350
transform 1 0 29256 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_318
timestamp 1606120350
transform 1 0 30360 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_330
timestamp 1606120350
transform 1 0 31464 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_342
timestamp 1606120350
transform 1 0 32568 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_354
timestamp 1606120350
transform 1 0 33672 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1076
timestamp 1606120350
transform 1 0 34776 0 1 68000
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_121_367
timestamp 1606120350
transform 1 0 34868 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_121_379
timestamp 1606120350
transform 1 0 35972 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_243
timestamp 1606120350
transform -1 0 38824 0 1 68000
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_121_391
timestamp 1606120350
transform 1 0 37076 0 1 68000
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_121_403
timestamp 1606120350
transform 1 0 38180 0 1 68000
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_244
timestamp 1606120350
transform 1 0 1104 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_122_3
timestamp 1606120350
transform 1 0 1380 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_15
timestamp 1606120350
transform 1 0 2484 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1077
timestamp 1606120350
transform 1 0 3956 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_122_27
timestamp 1606120350
transform 1 0 3588 0 -1 69088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_122_32
timestamp 1606120350
transform 1 0 4048 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_44
timestamp 1606120350
transform 1 0 5152 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_56
timestamp 1606120350
transform 1 0 6256 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_68
timestamp 1606120350
transform 1 0 7360 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_80
timestamp 1606120350
transform 1 0 8464 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1078
timestamp 1606120350
transform 1 0 9568 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_93
timestamp 1606120350
transform 1 0 9660 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_105
timestamp 1606120350
transform 1 0 10764 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_117
timestamp 1606120350
transform 1 0 11868 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_129
timestamp 1606120350
transform 1 0 12972 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1079
timestamp 1606120350
transform 1 0 15180 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_141
timestamp 1606120350
transform 1 0 14076 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_154
timestamp 1606120350
transform 1 0 15272 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_166
timestamp 1606120350
transform 1 0 16376 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_178
timestamp 1606120350
transform 1 0 17480 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_190
timestamp 1606120350
transform 1 0 18584 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_202
timestamp 1606120350
transform 1 0 19688 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1080
timestamp 1606120350
transform 1 0 20792 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_215
timestamp 1606120350
transform 1 0 20884 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_122_227
timestamp 1606120350
transform 1 0 21988 0 -1 69088
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _1181_
timestamp 1606120350
transform 1 0 22540 0 -1 69088
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_14_0_clk
timestamp 1606120350
transform 1 0 25024 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_122_252
timestamp 1606120350
transform 1 0 24288 0 -1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_122_263
timestamp 1606120350
transform 1 0 25300 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1081
timestamp 1606120350
transform 1 0 26404 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_276
timestamp 1606120350
transform 1 0 26496 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_288
timestamp 1606120350
transform 1 0 27600 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_300
timestamp 1606120350
transform 1 0 28704 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_312
timestamp 1606120350
transform 1 0 29808 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1082
timestamp 1606120350
transform 1 0 32016 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_122_324
timestamp 1606120350
transform 1 0 30912 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_337
timestamp 1606120350
transform 1 0 32108 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_349
timestamp 1606120350
transform 1 0 33212 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_361
timestamp 1606120350
transform 1 0 34316 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_373
timestamp 1606120350
transform 1 0 35420 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_122_385
timestamp 1606120350
transform 1 0 36524 0 -1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_245
timestamp 1606120350
transform -1 0 38824 0 -1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1083
timestamp 1606120350
transform 1 0 37628 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_122_398
timestamp 1606120350
transform 1 0 37720 0 -1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_122_406
timestamp 1606120350
transform 1 0 38456 0 -1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_246
timestamp 1606120350
transform 1 0 1104 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_3
timestamp 1606120350
transform 1 0 1380 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_15
timestamp 1606120350
transform 1 0 2484 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_27
timestamp 1606120350
transform 1 0 3588 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_39
timestamp 1606120350
transform 1 0 4692 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1084
timestamp 1606120350
transform 1 0 6716 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_123_51
timestamp 1606120350
transform 1 0 5796 0 1 69088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_123_59
timestamp 1606120350
transform 1 0 6532 0 1 69088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_123_62
timestamp 1606120350
transform 1 0 6808 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_74
timestamp 1606120350
transform 1 0 7912 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_86
timestamp 1606120350
transform 1 0 9016 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_98
timestamp 1606120350
transform 1 0 10120 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_110
timestamp 1606120350
transform 1 0 11224 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1085
timestamp 1606120350
transform 1 0 12328 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_123
timestamp 1606120350
transform 1 0 12420 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_135
timestamp 1606120350
transform 1 0 13524 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_147
timestamp 1606120350
transform 1 0 14628 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_159
timestamp 1606120350
transform 1 0 15732 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_171
timestamp 1606120350
transform 1 0 16836 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1086
timestamp 1606120350
transform 1 0 17940 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_184
timestamp 1606120350
transform 1 0 18032 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_196
timestamp 1606120350
transform 1 0 19136 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_208
timestamp 1606120350
transform 1 0 20240 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_220
timestamp 1606120350
transform 1 0 21344 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1087
timestamp 1606120350
transform 1 0 23552 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__D
timestamp 1606120350
transform 1 0 23920 0 1 69088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_123_232
timestamp 1606120350
transform 1 0 22448 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_123_245
timestamp 1606120350
transform 1 0 23644 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_123_250
timestamp 1606120350
transform 1 0 24104 0 1 69088
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_4_15_0_clk
timestamp 1606120350
transform 1 0 25944 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1222__CLK
timestamp 1606120350
transform 1 0 24288 0 1 69088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_123_254
timestamp 1606120350
transform 1 0 24472 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_123_266
timestamp 1606120350
transform 1 0 25576 0 1 69088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_123_273
timestamp 1606120350
transform 1 0 26220 0 1 69088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_4_15_0_clk_A
timestamp 1606120350
transform 1 0 26404 0 1 69088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_123_277
timestamp 1606120350
transform 1 0 26588 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_289
timestamp 1606120350
transform 1 0 27692 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1088
timestamp 1606120350
transform 1 0 29164 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_123_301
timestamp 1606120350
transform 1 0 28796 0 1 69088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_123_306
timestamp 1606120350
transform 1 0 29256 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_318
timestamp 1606120350
transform 1 0 30360 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_330
timestamp 1606120350
transform 1 0 31464 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_342
timestamp 1606120350
transform 1 0 32568 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_354
timestamp 1606120350
transform 1 0 33672 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1089
timestamp 1606120350
transform 1 0 34776 0 1 69088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_123_367
timestamp 1606120350
transform 1 0 34868 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_123_379
timestamp 1606120350
transform 1 0 35972 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_247
timestamp 1606120350
transform -1 0 38824 0 1 69088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_123_391
timestamp 1606120350
transform 1 0 37076 0 1 69088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_123_403
timestamp 1606120350
transform 1 0 38180 0 1 69088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_248
timestamp 1606120350
transform 1 0 1104 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_124_3
timestamp 1606120350
transform 1 0 1380 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_15
timestamp 1606120350
transform 1 0 2484 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1090
timestamp 1606120350
transform 1 0 3956 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_124_27
timestamp 1606120350
transform 1 0 3588 0 -1 70176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_124_32
timestamp 1606120350
transform 1 0 4048 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_44
timestamp 1606120350
transform 1 0 5152 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_56
timestamp 1606120350
transform 1 0 6256 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_68
timestamp 1606120350
transform 1 0 7360 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_80
timestamp 1606120350
transform 1 0 8464 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1091
timestamp 1606120350
transform 1 0 9568 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_124_93
timestamp 1606120350
transform 1 0 9660 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_105
timestamp 1606120350
transform 1 0 10764 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_117
timestamp 1606120350
transform 1 0 11868 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_129
timestamp 1606120350
transform 1 0 12972 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1092
timestamp 1606120350
transform 1 0 15180 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_124_141
timestamp 1606120350
transform 1 0 14076 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_154
timestamp 1606120350
transform 1 0 15272 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_166
timestamp 1606120350
transform 1 0 16376 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_178
timestamp 1606120350
transform 1 0 17480 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_190
timestamp 1606120350
transform 1 0 18584 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_202
timestamp 1606120350
transform 1 0 19688 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1093
timestamp 1606120350
transform 1 0 20792 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_124_215
timestamp 1606120350
transform 1 0 20884 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_227
timestamp 1606120350
transform 1 0 21988 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1222_
timestamp 1606120350
transform 1 0 23920 0 -1 70176
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_124_239
timestamp 1606120350
transform 1 0 23092 0 -1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_124_247
timestamp 1606120350
transform 1 0 23828 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_124_267
timestamp 1606120350
transform 1 0 25668 0 -1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1094
timestamp 1606120350
transform 1 0 26404 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_124_276
timestamp 1606120350
transform 1 0 26496 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_288
timestamp 1606120350
transform 1 0 27600 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_300
timestamp 1606120350
transform 1 0 28704 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_312
timestamp 1606120350
transform 1 0 29808 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1095
timestamp 1606120350
transform 1 0 32016 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_124_324
timestamp 1606120350
transform 1 0 30912 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_337
timestamp 1606120350
transform 1 0 32108 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_349
timestamp 1606120350
transform 1 0 33212 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_361
timestamp 1606120350
transform 1 0 34316 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_373
timestamp 1606120350
transform 1 0 35420 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_124_385
timestamp 1606120350
transform 1 0 36524 0 -1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_249
timestamp 1606120350
transform -1 0 38824 0 -1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1096
timestamp 1606120350
transform 1 0 37628 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_124_398
timestamp 1606120350
transform 1 0 37720 0 -1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_124_406
timestamp 1606120350
transform 1 0 38456 0 -1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_250
timestamp 1606120350
transform 1 0 1104 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_252
timestamp 1606120350
transform 1 0 1104 0 -1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_125_3
timestamp 1606120350
transform 1 0 1380 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_15
timestamp 1606120350
transform 1 0 2484 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_3
timestamp 1606120350
transform 1 0 1380 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_15
timestamp 1606120350
transform 1 0 2484 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1103
timestamp 1606120350
transform 1 0 3956 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_27
timestamp 1606120350
transform 1 0 3588 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_39
timestamp 1606120350
transform 1 0 4692 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_126_27
timestamp 1606120350
transform 1 0 3588 0 -1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_126_32
timestamp 1606120350
transform 1 0 4048 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_44
timestamp 1606120350
transform 1 0 5152 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1097
timestamp 1606120350
transform 1 0 6716 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_125_51
timestamp 1606120350
transform 1 0 5796 0 1 70176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_125_59
timestamp 1606120350
transform 1 0 6532 0 1 70176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_125_62
timestamp 1606120350
transform 1 0 6808 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_56
timestamp 1606120350
transform 1 0 6256 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_68
timestamp 1606120350
transform 1 0 7360 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_74
timestamp 1606120350
transform 1 0 7912 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_86
timestamp 1606120350
transform 1 0 9016 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_80
timestamp 1606120350
transform 1 0 8464 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1104
timestamp 1606120350
transform 1 0 9568 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_98
timestamp 1606120350
transform 1 0 10120 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_110
timestamp 1606120350
transform 1 0 11224 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_93
timestamp 1606120350
transform 1 0 9660 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_105
timestamp 1606120350
transform 1 0 10764 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1098
timestamp 1606120350
transform 1 0 12328 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_123
timestamp 1606120350
transform 1 0 12420 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_135
timestamp 1606120350
transform 1 0 13524 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_117
timestamp 1606120350
transform 1 0 11868 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_129
timestamp 1606120350
transform 1 0 12972 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1105
timestamp 1606120350
transform 1 0 15180 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_147
timestamp 1606120350
transform 1 0 14628 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_159
timestamp 1606120350
transform 1 0 15732 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_141
timestamp 1606120350
transform 1 0 14076 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_154
timestamp 1606120350
transform 1 0 15272 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_171
timestamp 1606120350
transform 1 0 16836 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_166
timestamp 1606120350
transform 1 0 16376 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_178
timestamp 1606120350
transform 1 0 17480 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1099
timestamp 1606120350
transform 1 0 17940 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_184
timestamp 1606120350
transform 1 0 18032 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_196
timestamp 1606120350
transform 1 0 19136 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_190
timestamp 1606120350
transform 1 0 18584 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_202
timestamp 1606120350
transform 1 0 19688 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1106
timestamp 1606120350
transform 1 0 20792 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_208
timestamp 1606120350
transform 1 0 20240 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_220
timestamp 1606120350
transform 1 0 21344 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_215
timestamp 1606120350
transform 1 0 20884 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_126_227
timestamp 1606120350
transform 1 0 21988 0 -1 71264
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _1199_
timestamp 1606120350
transform 1 0 22632 0 -1 71264
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1100
timestamp 1606120350
transform 1 0 23552 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__D
timestamp 1606120350
transform 1 0 22632 0 1 70176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1199__CLK
timestamp 1606120350
transform 1 0 23000 0 1 70176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_125_232
timestamp 1606120350
transform 1 0 22448 0 1 70176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_125_236
timestamp 1606120350
transform 1 0 22816 0 1 70176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_125_240
timestamp 1606120350
transform 1 0 23184 0 1 70176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_125_245
timestamp 1606120350
transform 1 0 23644 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_126_233
timestamp 1606120350
transform 1 0 22540 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_257
timestamp 1606120350
transform 1 0 24748 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_269
timestamp 1606120350
transform 1 0 25852 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_253
timestamp 1606120350
transform 1 0 24380 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_126_265
timestamp 1606120350
transform 1 0 25484 0 -1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_126_273
timestamp 1606120350
transform 1 0 26220 0 -1 71264
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1107
timestamp 1606120350
transform 1 0 26404 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_281
timestamp 1606120350
transform 1 0 26956 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_293
timestamp 1606120350
transform 1 0 28060 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_276
timestamp 1606120350
transform 1 0 26496 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_288
timestamp 1606120350
transform 1 0 27600 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1101
timestamp 1606120350
transform 1 0 29164 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_306
timestamp 1606120350
transform 1 0 29256 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_318
timestamp 1606120350
transform 1 0 30360 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_300
timestamp 1606120350
transform 1 0 28704 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_312
timestamp 1606120350
transform 1 0 29808 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1108
timestamp 1606120350
transform 1 0 32016 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_330
timestamp 1606120350
transform 1 0 31464 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_342
timestamp 1606120350
transform 1 0 32568 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_324
timestamp 1606120350
transform 1 0 30912 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_337
timestamp 1606120350
transform 1 0 32108 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_354
timestamp 1606120350
transform 1 0 33672 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_349
timestamp 1606120350
transform 1 0 33212 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_361
timestamp 1606120350
transform 1 0 34316 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1102
timestamp 1606120350
transform 1 0 34776 0 1 70176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_367
timestamp 1606120350
transform 1 0 34868 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_125_379
timestamp 1606120350
transform 1 0 35972 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_373
timestamp 1606120350
transform 1 0 35420 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_126_385
timestamp 1606120350
transform 1 0 36524 0 -1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_251
timestamp 1606120350
transform -1 0 38824 0 1 70176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_253
timestamp 1606120350
transform -1 0 38824 0 -1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1109
timestamp 1606120350
transform 1 0 37628 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_125_391
timestamp 1606120350
transform 1 0 37076 0 1 70176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_125_403
timestamp 1606120350
transform 1 0 38180 0 1 70176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_126_398
timestamp 1606120350
transform 1 0 37720 0 -1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_126_406
timestamp 1606120350
transform 1 0 38456 0 -1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_254
timestamp 1606120350
transform 1 0 1104 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_127_3
timestamp 1606120350
transform 1 0 1380 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_15
timestamp 1606120350
transform 1 0 2484 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_27
timestamp 1606120350
transform 1 0 3588 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_39
timestamp 1606120350
transform 1 0 4692 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1110
timestamp 1606120350
transform 1 0 6716 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_127_51
timestamp 1606120350
transform 1 0 5796 0 1 71264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_127_59
timestamp 1606120350
transform 1 0 6532 0 1 71264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_127_62
timestamp 1606120350
transform 1 0 6808 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_74
timestamp 1606120350
transform 1 0 7912 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_86
timestamp 1606120350
transform 1 0 9016 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_98
timestamp 1606120350
transform 1 0 10120 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_110
timestamp 1606120350
transform 1 0 11224 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1111
timestamp 1606120350
transform 1 0 12328 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_123
timestamp 1606120350
transform 1 0 12420 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_135
timestamp 1606120350
transform 1 0 13524 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_147
timestamp 1606120350
transform 1 0 14628 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_159
timestamp 1606120350
transform 1 0 15732 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_171
timestamp 1606120350
transform 1 0 16836 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1112
timestamp 1606120350
transform 1 0 17940 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_184
timestamp 1606120350
transform 1 0 18032 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_196
timestamp 1606120350
transform 1 0 19136 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_208
timestamp 1606120350
transform 1 0 20240 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_220
timestamp 1606120350
transform 1 0 21344 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1113
timestamp 1606120350
transform 1 0 23552 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_232
timestamp 1606120350
transform 1 0 22448 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_245
timestamp 1606120350
transform 1 0 23644 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_257
timestamp 1606120350
transform 1 0 24748 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_269
timestamp 1606120350
transform 1 0 25852 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_281
timestamp 1606120350
transform 1 0 26956 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_293
timestamp 1606120350
transform 1 0 28060 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1114
timestamp 1606120350
transform 1 0 29164 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_306
timestamp 1606120350
transform 1 0 29256 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_318
timestamp 1606120350
transform 1 0 30360 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_330
timestamp 1606120350
transform 1 0 31464 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_342
timestamp 1606120350
transform 1 0 32568 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_354
timestamp 1606120350
transform 1 0 33672 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1115
timestamp 1606120350
transform 1 0 34776 0 1 71264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_127_367
timestamp 1606120350
transform 1 0 34868 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_127_379
timestamp 1606120350
transform 1 0 35972 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_255
timestamp 1606120350
transform -1 0 38824 0 1 71264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_127_391
timestamp 1606120350
transform 1 0 37076 0 1 71264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_127_403
timestamp 1606120350
transform 1 0 38180 0 1 71264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_256
timestamp 1606120350
transform 1 0 1104 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_128_3
timestamp 1606120350
transform 1 0 1380 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_15
timestamp 1606120350
transform 1 0 2484 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1116
timestamp 1606120350
transform 1 0 3956 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_128_27
timestamp 1606120350
transform 1 0 3588 0 -1 72352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_128_32
timestamp 1606120350
transform 1 0 4048 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_44
timestamp 1606120350
transform 1 0 5152 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_56
timestamp 1606120350
transform 1 0 6256 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_68
timestamp 1606120350
transform 1 0 7360 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_80
timestamp 1606120350
transform 1 0 8464 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1117
timestamp 1606120350
transform 1 0 9568 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_93
timestamp 1606120350
transform 1 0 9660 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_105
timestamp 1606120350
transform 1 0 10764 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_117
timestamp 1606120350
transform 1 0 11868 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_129
timestamp 1606120350
transform 1 0 12972 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1118
timestamp 1606120350
transform 1 0 15180 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_141
timestamp 1606120350
transform 1 0 14076 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_154
timestamp 1606120350
transform 1 0 15272 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_166
timestamp 1606120350
transform 1 0 16376 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_178
timestamp 1606120350
transform 1 0 17480 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__CLK
timestamp 1606120350
transform 1 0 19504 0 -1 72352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_128_190
timestamp 1606120350
transform 1 0 18584 0 -1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_128_198
timestamp 1606120350
transform 1 0 19320 0 -1 72352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_128_202
timestamp 1606120350
transform 1 0 19688 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1119
timestamp 1606120350
transform 1 0 20792 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_215
timestamp 1606120350
transform 1 0 20884 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_227
timestamp 1606120350
transform 1 0 21988 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_239
timestamp 1606120350
transform 1 0 23092 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_251
timestamp 1606120350
transform 1 0 24196 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_263
timestamp 1606120350
transform 1 0 25300 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1120
timestamp 1606120350
transform 1 0 26404 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_276
timestamp 1606120350
transform 1 0 26496 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_288
timestamp 1606120350
transform 1 0 27600 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_300
timestamp 1606120350
transform 1 0 28704 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_312
timestamp 1606120350
transform 1 0 29808 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1121
timestamp 1606120350
transform 1 0 32016 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_128_324
timestamp 1606120350
transform 1 0 30912 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_337
timestamp 1606120350
transform 1 0 32108 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_349
timestamp 1606120350
transform 1 0 33212 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_361
timestamp 1606120350
transform 1 0 34316 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_373
timestamp 1606120350
transform 1 0 35420 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_128_385
timestamp 1606120350
transform 1 0 36524 0 -1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_257
timestamp 1606120350
transform -1 0 38824 0 -1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1122
timestamp 1606120350
transform 1 0 37628 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_128_398
timestamp 1606120350
transform 1 0 37720 0 -1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_128_406
timestamp 1606120350
transform 1 0 38456 0 -1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_258
timestamp 1606120350
transform 1 0 1104 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_129_3
timestamp 1606120350
transform 1 0 1380 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_15
timestamp 1606120350
transform 1 0 2484 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_27
timestamp 1606120350
transform 1 0 3588 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_39
timestamp 1606120350
transform 1 0 4692 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1123
timestamp 1606120350
transform 1 0 6716 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_129_51
timestamp 1606120350
transform 1 0 5796 0 1 72352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_129_59
timestamp 1606120350
transform 1 0 6532 0 1 72352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_129_62
timestamp 1606120350
transform 1 0 6808 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_74
timestamp 1606120350
transform 1 0 7912 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_86
timestamp 1606120350
transform 1 0 9016 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_98
timestamp 1606120350
transform 1 0 10120 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_110
timestamp 1606120350
transform 1 0 11224 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1124
timestamp 1606120350
transform 1 0 12328 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_123
timestamp 1606120350
transform 1 0 12420 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_135
timestamp 1606120350
transform 1 0 13524 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_147
timestamp 1606120350
transform 1 0 14628 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_159
timestamp 1606120350
transform 1 0 15732 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_171
timestamp 1606120350
transform 1 0 16836 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1217_
timestamp 1606120350
transform 1 0 19504 0 1 72352
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1125
timestamp 1606120350
transform 1 0 17940 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1217__D
timestamp 1606120350
transform 1 0 19320 0 1 72352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_129_184
timestamp 1606120350
transform 1 0 18032 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_129_196
timestamp 1606120350
transform 1 0 19136 0 1 72352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_129_219
timestamp 1606120350
transform 1 0 21252 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1126
timestamp 1606120350
transform 1 0 23552 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_231
timestamp 1606120350
transform 1 0 22356 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_129_243
timestamp 1606120350
transform 1 0 23460 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_245
timestamp 1606120350
transform 1 0 23644 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_257
timestamp 1606120350
transform 1 0 24748 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_269
timestamp 1606120350
transform 1 0 25852 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_281
timestamp 1606120350
transform 1 0 26956 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_293
timestamp 1606120350
transform 1 0 28060 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1127
timestamp 1606120350
transform 1 0 29164 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_306
timestamp 1606120350
transform 1 0 29256 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_318
timestamp 1606120350
transform 1 0 30360 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_330
timestamp 1606120350
transform 1 0 31464 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_342
timestamp 1606120350
transform 1 0 32568 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_354
timestamp 1606120350
transform 1 0 33672 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1128
timestamp 1606120350
transform 1 0 34776 0 1 72352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_129_367
timestamp 1606120350
transform 1 0 34868 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_129_379
timestamp 1606120350
transform 1 0 35972 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_259
timestamp 1606120350
transform -1 0 38824 0 1 72352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_129_391
timestamp 1606120350
transform 1 0 37076 0 1 72352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_129_403
timestamp 1606120350
transform 1 0 38180 0 1 72352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_260
timestamp 1606120350
transform 1 0 1104 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_130_3
timestamp 1606120350
transform 1 0 1380 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_15
timestamp 1606120350
transform 1 0 2484 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1129
timestamp 1606120350
transform 1 0 3956 0 -1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_130_27
timestamp 1606120350
transform 1 0 3588 0 -1 73440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_130_32
timestamp 1606120350
transform 1 0 4048 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_44
timestamp 1606120350
transform 1 0 5152 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_56
timestamp 1606120350
transform 1 0 6256 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_68
timestamp 1606120350
transform 1 0 7360 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_80
timestamp 1606120350
transform 1 0 8464 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1130
timestamp 1606120350
transform 1 0 9568 0 -1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_93
timestamp 1606120350
transform 1 0 9660 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_105
timestamp 1606120350
transform 1 0 10764 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_117
timestamp 1606120350
transform 1 0 11868 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_129
timestamp 1606120350
transform 1 0 12972 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1131
timestamp 1606120350
transform 1 0 15180 0 -1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_141
timestamp 1606120350
transform 1 0 14076 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_154
timestamp 1606120350
transform 1 0 15272 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_166
timestamp 1606120350
transform 1 0 16376 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_178
timestamp 1606120350
transform 1 0 17480 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_190
timestamp 1606120350
transform 1 0 18584 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_202
timestamp 1606120350
transform 1 0 19688 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1132
timestamp 1606120350
transform 1 0 20792 0 -1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_215
timestamp 1606120350
transform 1 0 20884 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_227
timestamp 1606120350
transform 1 0 21988 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_239
timestamp 1606120350
transform 1 0 23092 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_251
timestamp 1606120350
transform 1 0 24196 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_263
timestamp 1606120350
transform 1 0 25300 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1133
timestamp 1606120350
transform 1 0 26404 0 -1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_276
timestamp 1606120350
transform 1 0 26496 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_288
timestamp 1606120350
transform 1 0 27600 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_300
timestamp 1606120350
transform 1 0 28704 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_312
timestamp 1606120350
transform 1 0 29808 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1134
timestamp 1606120350
transform 1 0 32016 0 -1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_130_324
timestamp 1606120350
transform 1 0 30912 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_337
timestamp 1606120350
transform 1 0 32108 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_349
timestamp 1606120350
transform 1 0 33212 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_361
timestamp 1606120350
transform 1 0 34316 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_373
timestamp 1606120350
transform 1 0 35420 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_130_385
timestamp 1606120350
transform 1 0 36524 0 -1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_261
timestamp 1606120350
transform -1 0 38824 0 -1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1135
timestamp 1606120350
transform 1 0 37628 0 -1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_130_398
timestamp 1606120350
transform 1 0 37720 0 -1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_130_406
timestamp 1606120350
transform 1 0 38456 0 -1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_262
timestamp 1606120350
transform 1 0 1104 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_131_3
timestamp 1606120350
transform 1 0 1380 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_15
timestamp 1606120350
transform 1 0 2484 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_27
timestamp 1606120350
transform 1 0 3588 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_39
timestamp 1606120350
transform 1 0 4692 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1136
timestamp 1606120350
transform 1 0 6716 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_131_51
timestamp 1606120350
transform 1 0 5796 0 1 73440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_131_59
timestamp 1606120350
transform 1 0 6532 0 1 73440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_131_62
timestamp 1606120350
transform 1 0 6808 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_74
timestamp 1606120350
transform 1 0 7912 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_86
timestamp 1606120350
transform 1 0 9016 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_98
timestamp 1606120350
transform 1 0 10120 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_110
timestamp 1606120350
transform 1 0 11224 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1137
timestamp 1606120350
transform 1 0 12328 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_123
timestamp 1606120350
transform 1 0 12420 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_135
timestamp 1606120350
transform 1 0 13524 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_147
timestamp 1606120350
transform 1 0 14628 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_159
timestamp 1606120350
transform 1 0 15732 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_171
timestamp 1606120350
transform 1 0 16836 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1138
timestamp 1606120350
transform 1 0 17940 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_184
timestamp 1606120350
transform 1 0 18032 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_196
timestamp 1606120350
transform 1 0 19136 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_208
timestamp 1606120350
transform 1 0 20240 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_220
timestamp 1606120350
transform 1 0 21344 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1139
timestamp 1606120350
transform 1 0 23552 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_232
timestamp 1606120350
transform 1 0 22448 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_245
timestamp 1606120350
transform 1 0 23644 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_257
timestamp 1606120350
transform 1 0 24748 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_269
timestamp 1606120350
transform 1 0 25852 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_281
timestamp 1606120350
transform 1 0 26956 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_293
timestamp 1606120350
transform 1 0 28060 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1140
timestamp 1606120350
transform 1 0 29164 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_306
timestamp 1606120350
transform 1 0 29256 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_318
timestamp 1606120350
transform 1 0 30360 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_330
timestamp 1606120350
transform 1 0 31464 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_342
timestamp 1606120350
transform 1 0 32568 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_354
timestamp 1606120350
transform 1 0 33672 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1141
timestamp 1606120350
transform 1 0 34776 0 1 73440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_131_367
timestamp 1606120350
transform 1 0 34868 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_131_379
timestamp 1606120350
transform 1 0 35972 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_263
timestamp 1606120350
transform -1 0 38824 0 1 73440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_131_391
timestamp 1606120350
transform 1 0 37076 0 1 73440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_131_403
timestamp 1606120350
transform 1 0 38180 0 1 73440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_264
timestamp 1606120350
transform 1 0 1104 0 -1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_266
timestamp 1606120350
transform 1 0 1104 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_132_3
timestamp 1606120350
transform 1 0 1380 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_15
timestamp 1606120350
transform 1 0 2484 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_3
timestamp 1606120350
transform 1 0 1380 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_15
timestamp 1606120350
transform 1 0 2484 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1142
timestamp 1606120350
transform 1 0 3956 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_132_27
timestamp 1606120350
transform 1 0 3588 0 -1 74528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_132_32
timestamp 1606120350
transform 1 0 4048 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_44
timestamp 1606120350
transform 1 0 5152 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_27
timestamp 1606120350
transform 1 0 3588 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_39
timestamp 1606120350
transform 1 0 4692 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1149
timestamp 1606120350
transform 1 0 6716 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_56
timestamp 1606120350
transform 1 0 6256 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_68
timestamp 1606120350
transform 1 0 7360 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_51
timestamp 1606120350
transform 1 0 5796 0 1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_133_59
timestamp 1606120350
transform 1 0 6532 0 1 74528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_133_62
timestamp 1606120350
transform 1 0 6808 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_80
timestamp 1606120350
transform 1 0 8464 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_74
timestamp 1606120350
transform 1 0 7912 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_86
timestamp 1606120350
transform 1 0 9016 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1143
timestamp 1606120350
transform 1 0 9568 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_93
timestamp 1606120350
transform 1 0 9660 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_105
timestamp 1606120350
transform 1 0 10764 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_98
timestamp 1606120350
transform 1 0 10120 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_110
timestamp 1606120350
transform 1 0 11224 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1150
timestamp 1606120350
transform 1 0 12328 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_117
timestamp 1606120350
transform 1 0 11868 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_129
timestamp 1606120350
transform 1 0 12972 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_123
timestamp 1606120350
transform 1 0 12420 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_135
timestamp 1606120350
transform 1 0 13524 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1144
timestamp 1606120350
transform 1 0 15180 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_141
timestamp 1606120350
transform 1 0 14076 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_154
timestamp 1606120350
transform 1 0 15272 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_147
timestamp 1606120350
transform 1 0 14628 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_159
timestamp 1606120350
transform 1 0 15732 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_166
timestamp 1606120350
transform 1 0 16376 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_178
timestamp 1606120350
transform 1 0 17480 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_171
timestamp 1606120350
transform 1 0 16836 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1151
timestamp 1606120350
transform 1 0 17940 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_133_200
timestamp 1606120350
transform 1 0 19504 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_133_196
timestamp 1606120350
transform 1 0 19136 0 1 74528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_132_205
timestamp 1606120350
transform 1 0 19964 0 -1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_132_202
timestamp 1606120350
transform 1 0 19688 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__CLK
timestamp 1606120350
transform 1 0 19780 0 -1 74528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1153__D
timestamp 1606120350
transform 1 0 19596 0 1 74528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_133_184
timestamp 1606120350
transform 1 0 18032 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_190
timestamp 1606120350
transform 1 0 18584 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1153_
timestamp 1606120350
transform 1 0 19780 0 1 74528
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1145
timestamp 1606120350
transform 1 0 20792 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_132_213
timestamp 1606120350
transform 1 0 20700 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_215
timestamp 1606120350
transform 1 0 20884 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_227
timestamp 1606120350
transform 1 0 21988 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_222
timestamp 1606120350
transform 1 0 21528 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1152
timestamp 1606120350
transform 1 0 23552 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_239
timestamp 1606120350
transform 1 0 23092 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_251
timestamp 1606120350
transform 1 0 24196 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_234
timestamp 1606120350
transform 1 0 22632 0 1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_133_242
timestamp 1606120350
transform 1 0 23368 0 1 74528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_133_245
timestamp 1606120350
transform 1 0 23644 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_263
timestamp 1606120350
transform 1 0 25300 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_257
timestamp 1606120350
transform 1 0 24748 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_269
timestamp 1606120350
transform 1 0 25852 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1146
timestamp 1606120350
transform 1 0 26404 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_276
timestamp 1606120350
transform 1 0 26496 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_288
timestamp 1606120350
transform 1 0 27600 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_281
timestamp 1606120350
transform 1 0 26956 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_293
timestamp 1606120350
transform 1 0 28060 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1153
timestamp 1606120350
transform 1 0 29164 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__B1_N
timestamp 1606120350
transform 1 0 29624 0 1 74528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A2
timestamp 1606120350
transform 1 0 29992 0 1 74528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__0933__A1
timestamp 1606120350
transform 1 0 30360 0 1 74528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_132_300
timestamp 1606120350
transform 1 0 28704 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_312
timestamp 1606120350
transform 1 0 29808 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_133_306
timestamp 1606120350
transform 1 0 29256 0 1 74528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_133_312
timestamp 1606120350
transform 1 0 29808 0 1 74528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_133_316
timestamp 1606120350
transform 1 0 30176 0 1 74528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1147
timestamp 1606120350
transform 1 0 32016 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_324
timestamp 1606120350
transform 1 0 30912 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_337
timestamp 1606120350
transform 1 0 32108 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_320
timestamp 1606120350
transform 1 0 30544 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_332
timestamp 1606120350
transform 1 0 31648 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_349
timestamp 1606120350
transform 1 0 33212 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_361
timestamp 1606120350
transform 1 0 34316 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_344
timestamp 1606120350
transform 1 0 32752 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_133_356
timestamp 1606120350
transform 1 0 33856 0 1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_133_364
timestamp 1606120350
transform 1 0 34592 0 1 74528
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1154
timestamp 1606120350
transform 1 0 34776 0 1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_132_373
timestamp 1606120350
transform 1 0 35420 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_132_385
timestamp 1606120350
transform 1 0 36524 0 -1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_367
timestamp 1606120350
transform 1 0 34868 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_133_379
timestamp 1606120350
transform 1 0 35972 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_265
timestamp 1606120350
transform -1 0 38824 0 -1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_267
timestamp 1606120350
transform -1 0 38824 0 1 74528
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1148
timestamp 1606120350
transform 1 0 37628 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_132_398
timestamp 1606120350
transform 1 0 37720 0 -1 74528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_132_406
timestamp 1606120350
transform 1 0 38456 0 -1 74528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_133_391
timestamp 1606120350
transform 1 0 37076 0 1 74528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_133_403
timestamp 1606120350
transform 1 0 38180 0 1 74528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_268
timestamp 1606120350
transform 1 0 1104 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_134_3
timestamp 1606120350
transform 1 0 1380 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_15
timestamp 1606120350
transform 1 0 2484 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1155
timestamp 1606120350
transform 1 0 3956 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_134_27
timestamp 1606120350
transform 1 0 3588 0 -1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_134_32
timestamp 1606120350
transform 1 0 4048 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_44
timestamp 1606120350
transform 1 0 5152 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_56
timestamp 1606120350
transform 1 0 6256 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_68
timestamp 1606120350
transform 1 0 7360 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_80
timestamp 1606120350
transform 1 0 8464 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1156
timestamp 1606120350
transform 1 0 9568 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_93
timestamp 1606120350
transform 1 0 9660 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_105
timestamp 1606120350
transform 1 0 10764 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_117
timestamp 1606120350
transform 1 0 11868 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_129
timestamp 1606120350
transform 1 0 12972 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1157
timestamp 1606120350
transform 1 0 15180 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_141
timestamp 1606120350
transform 1 0 14076 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_154
timestamp 1606120350
transform 1 0 15272 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_166
timestamp 1606120350
transform 1 0 16376 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_178
timestamp 1606120350
transform 1 0 17480 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__CLK
timestamp 1606120350
transform 1 0 18860 0 -1 75616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_134_190
timestamp 1606120350
transform 1 0 18584 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_134_195
timestamp 1606120350
transform 1 0 19044 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1158
timestamp 1606120350
transform 1 0 20792 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_134_207
timestamp 1606120350
transform 1 0 20148 0 -1 75616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_134_213
timestamp 1606120350
transform 1 0 20700 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_215
timestamp 1606120350
transform 1 0 20884 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_227
timestamp 1606120350
transform 1 0 21988 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_239
timestamp 1606120350
transform 1 0 23092 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_251
timestamp 1606120350
transform 1 0 24196 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__CLK
timestamp 1606120350
transform 1 0 25852 0 -1 75616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_134_263
timestamp 1606120350
transform 1 0 25300 0 -1 75616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_134_271
timestamp 1606120350
transform 1 0 26036 0 -1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1159
timestamp 1606120350
transform 1 0 26404 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_276
timestamp 1606120350
transform 1 0 26496 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_288
timestamp 1606120350
transform 1 0 27600 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__a21bo_4  _0933_
timestamp 1606120350
transform 1 0 29624 0 -1 75616
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_134_300
timestamp 1606120350
transform 1 0 28704 0 -1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_134_308
timestamp 1606120350
transform 1 0 29440 0 -1 75616
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1160
timestamp 1606120350
transform 1 0 32016 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_323
timestamp 1606120350
transform 1 0 30820 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_134_335
timestamp 1606120350
transform 1 0 31924 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_134_337
timestamp 1606120350
transform 1 0 32108 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_349
timestamp 1606120350
transform 1 0 33212 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_361
timestamp 1606120350
transform 1 0 34316 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_373
timestamp 1606120350
transform 1 0 35420 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_134_385
timestamp 1606120350
transform 1 0 36524 0 -1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_269
timestamp 1606120350
transform -1 0 38824 0 -1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1161
timestamp 1606120350
transform 1 0 37628 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_134_398
timestamp 1606120350
transform 1 0 37720 0 -1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_134_406
timestamp 1606120350
transform 1 0 38456 0 -1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_270
timestamp 1606120350
transform 1 0 1104 0 1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_135_3
timestamp 1606120350
transform 1 0 1380 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_15
timestamp 1606120350
transform 1 0 2484 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_27
timestamp 1606120350
transform 1 0 3588 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_39
timestamp 1606120350
transform 1 0 4692 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1162
timestamp 1606120350
transform 1 0 6716 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_135_51
timestamp 1606120350
transform 1 0 5796 0 1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_135_59
timestamp 1606120350
transform 1 0 6532 0 1 75616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_135_62
timestamp 1606120350
transform 1 0 6808 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_74
timestamp 1606120350
transform 1 0 7912 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_86
timestamp 1606120350
transform 1 0 9016 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_98
timestamp 1606120350
transform 1 0 10120 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_110
timestamp 1606120350
transform 1 0 11224 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1163
timestamp 1606120350
transform 1 0 12328 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_123
timestamp 1606120350
transform 1 0 12420 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_135
timestamp 1606120350
transform 1 0 13524 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_147
timestamp 1606120350
transform 1 0 14628 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_159
timestamp 1606120350
transform 1 0 15732 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__D
timestamp 1606120350
transform 1 0 17572 0 1 75616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_135_171
timestamp 1606120350
transform 1 0 16836 0 1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_135_181
timestamp 1606120350
transform 1 0 17756 0 1 75616
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1161_
timestamp 1606120350
transform 1 0 18860 0 1 75616
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1164
timestamp 1606120350
transform 1 0 17940 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1161__D
timestamp 1606120350
transform 1 0 18676 0 1 75616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1138__CLK
timestamp 1606120350
transform 1 0 18216 0 1 75616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_135_184
timestamp 1606120350
transform 1 0 18032 0 1 75616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_135_188
timestamp 1606120350
transform 1 0 18400 0 1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__D
timestamp 1606120350
transform 1 0 21528 0 1 75616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1226__CLK
timestamp 1606120350
transform 1 0 21896 0 1 75616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_135_212
timestamp 1606120350
transform 1 0 20608 0 1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_135_220
timestamp 1606120350
transform 1 0 21344 0 1 75616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_135_224
timestamp 1606120350
transform 1 0 21712 0 1 75616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_135_228
timestamp 1606120350
transform 1 0 22080 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1165
timestamp 1606120350
transform 1 0 23552 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_135_240
timestamp 1606120350
transform 1 0 23184 0 1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_135_245
timestamp 1606120350
transform 1 0 23644 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1182_
timestamp 1606120350
transform 1 0 25852 0 1 75616
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1182__D
timestamp 1606120350
transform 1 0 25668 0 1 75616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_135_257
timestamp 1606120350
transform 1 0 24748 0 1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_135_265
timestamp 1606120350
transform 1 0 25484 0 1 75616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_135_288
timestamp 1606120350
transform 1 0 27600 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1166
timestamp 1606120350
transform 1 0 29164 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__D
timestamp 1606120350
transform 1 0 28796 0 1 75616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1191__CLK
timestamp 1606120350
transform 1 0 29440 0 1 75616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_135_300
timestamp 1606120350
transform 1 0 28704 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_135_303
timestamp 1606120350
transform 1 0 28980 0 1 75616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_135_306
timestamp 1606120350
transform 1 0 29256 0 1 75616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_135_310
timestamp 1606120350
transform 1 0 29624 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_322
timestamp 1606120350
transform 1 0 30728 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_334
timestamp 1606120350
transform 1 0 31832 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_346
timestamp 1606120350
transform 1 0 32936 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_135_358
timestamp 1606120350
transform 1 0 34040 0 1 75616
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1167
timestamp 1606120350
transform 1 0 34776 0 1 75616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_135_367
timestamp 1606120350
transform 1 0 34868 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_135_379
timestamp 1606120350
transform 1 0 35972 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_271
timestamp 1606120350
transform -1 0 38824 0 1 75616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_135_391
timestamp 1606120350
transform 1 0 37076 0 1 75616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_135_403
timestamp 1606120350
transform 1 0 38180 0 1 75616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_272
timestamp 1606120350
transform 1 0 1104 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_136_3
timestamp 1606120350
transform 1 0 1380 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_15
timestamp 1606120350
transform 1 0 2484 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1168
timestamp 1606120350
transform 1 0 3956 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_136_27
timestamp 1606120350
transform 1 0 3588 0 -1 76704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_136_32
timestamp 1606120350
transform 1 0 4048 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_44
timestamp 1606120350
transform 1 0 5152 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_56
timestamp 1606120350
transform 1 0 6256 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_68
timestamp 1606120350
transform 1 0 7360 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_80
timestamp 1606120350
transform 1 0 8464 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1169
timestamp 1606120350
transform 1 0 9568 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_93
timestamp 1606120350
transform 1 0 9660 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_105
timestamp 1606120350
transform 1 0 10764 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_117
timestamp 1606120350
transform 1 0 11868 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_129
timestamp 1606120350
transform 1 0 12972 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1170
timestamp 1606120350
transform 1 0 15180 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__CLK
timestamp 1606120350
transform 1 0 15456 0 -1 76704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_136_141
timestamp 1606120350
transform 1 0 14076 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_136_154
timestamp 1606120350
transform 1 0 15272 0 -1 76704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_136_158
timestamp 1606120350
transform 1 0 15640 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1138_
timestamp 1606120350
transform 1 0 17572 0 -1 76704
box -38 -48 1786 592
use sky130_fd_sc_hd__decap_8  FILLER_136_170
timestamp 1606120350
transform 1 0 16744 0 -1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_136_178
timestamp 1606120350
transform 1 0 17480 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_198
timestamp 1606120350
transform 1 0 19320 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1226_
timestamp 1606120350
transform 1 0 21528 0 -1 76704
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1171
timestamp 1606120350
transform 1 0 20792 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__CLK
timestamp 1606120350
transform 1 0 21068 0 -1 76704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_136_210
timestamp 1606120350
transform 1 0 20424 0 -1 76704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_136_215
timestamp 1606120350
transform 1 0 20884 0 -1 76704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_136_219
timestamp 1606120350
transform 1 0 21252 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__CLK
timestamp 1606120350
transform 1 0 24012 0 -1 76704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_136_241
timestamp 1606120350
transform 1 0 23276 0 -1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_136_251
timestamp 1606120350
transform 1 0 24196 0 -1 76704
box -38 -48 406 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__CLK
timestamp 1606120350
transform 1 0 24564 0 -1 76704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_136_257
timestamp 1606120350
transform 1 0 24748 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_136_269
timestamp 1606120350
transform 1 0 25852 0 -1 76704
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1172
timestamp 1606120350
transform 1 0 26404 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_276
timestamp 1606120350
transform 1 0 26496 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_288
timestamp 1606120350
transform 1 0 27600 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1191_
timestamp 1606120350
transform 1 0 28796 0 -1 76704
box -38 -48 1786 592
use sky130_fd_sc_hd__fill_1  FILLER_136_300
timestamp 1606120350
transform 1 0 28704 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1173
timestamp 1606120350
transform 1 0 32016 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_136_320
timestamp 1606120350
transform 1 0 30544 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_136_332
timestamp 1606120350
transform 1 0 31648 0 -1 76704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_136_337
timestamp 1606120350
transform 1 0 32108 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_349
timestamp 1606120350
transform 1 0 33212 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_361
timestamp 1606120350
transform 1 0 34316 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_373
timestamp 1606120350
transform 1 0 35420 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_136_385
timestamp 1606120350
transform 1 0 36524 0 -1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_273
timestamp 1606120350
transform -1 0 38824 0 -1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1174
timestamp 1606120350
transform 1 0 37628 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_136_398
timestamp 1606120350
transform 1 0 37720 0 -1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_136_406
timestamp 1606120350
transform 1 0 38456 0 -1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_274
timestamp 1606120350
transform 1 0 1104 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_137_3
timestamp 1606120350
transform 1 0 1380 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_15
timestamp 1606120350
transform 1 0 2484 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_27
timestamp 1606120350
transform 1 0 3588 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_39
timestamp 1606120350
transform 1 0 4692 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1175
timestamp 1606120350
transform 1 0 6716 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_137_51
timestamp 1606120350
transform 1 0 5796 0 1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_137_59
timestamp 1606120350
transform 1 0 6532 0 1 76704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_137_62
timestamp 1606120350
transform 1 0 6808 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_74
timestamp 1606120350
transform 1 0 7912 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_86
timestamp 1606120350
transform 1 0 9016 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_98
timestamp 1606120350
transform 1 0 10120 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_110
timestamp 1606120350
transform 1 0 11224 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1176
timestamp 1606120350
transform 1 0 12328 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_123
timestamp 1606120350
transform 1 0 12420 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_135
timestamp 1606120350
transform 1 0 13524 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1128_
timestamp 1606120350
transform 1 0 15456 0 1 76704
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1128__D
timestamp 1606120350
transform 1 0 15272 0 1 76704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_137_147
timestamp 1606120350
transform 1 0 14628 0 1 76704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_137_153
timestamp 1606120350
transform 1 0 15180 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__D
timestamp 1606120350
transform 1 0 17756 0 1 76704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_137_175
timestamp 1606120350
transform 1 0 17204 0 1 76704
box -38 -48 590 592
use sky130_fd_sc_hd__dfxtp_4  _1224_
timestamp 1606120350
transform 1 0 18032 0 1 76704
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1177
timestamp 1606120350
transform 1 0 17940 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_203
timestamp 1606120350
transform 1 0 19780 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1220_
timestamp 1606120350
transform 1 0 21068 0 1 76704
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1220__D
timestamp 1606120350
transform 1 0 20884 0 1 76704
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1178
timestamp 1606120350
transform 1 0 23552 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1171__D
timestamp 1606120350
transform 1 0 24012 0 1 76704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_137_236
timestamp 1606120350
transform 1 0 22816 0 1 76704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_137_245
timestamp 1606120350
transform 1 0 23644 0 1 76704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_137_251
timestamp 1606120350
transform 1 0 24196 0 1 76704
box -38 -48 222 592
use sky130_fd_sc_hd__dfxtp_4  _1177_
timestamp 1606120350
transform 1 0 24564 0 1 76704
box -38 -48 1786 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1177__D
timestamp 1606120350
transform 1 0 24380 0 1 76704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_137_274
timestamp 1606120350
transform 1 0 26312 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_286
timestamp 1606120350
transform 1 0 27416 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1203_
timestamp 1606120350
transform 1 0 29440 0 1 76704
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1179
timestamp 1606120350
transform 1 0 29164 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__D
timestamp 1606120350
transform 1 0 28980 0 1 76704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_137_298
timestamp 1606120350
transform 1 0 28520 0 1 76704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_137_302
timestamp 1606120350
transform 1 0 28888 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_137_306
timestamp 1606120350
transform 1 0 29256 0 1 76704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_137_327
timestamp 1606120350
transform 1 0 31188 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_339
timestamp 1606120350
transform 1 0 32292 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_351
timestamp 1606120350
transform 1 0 33396 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_137_363
timestamp 1606120350
transform 1 0 34500 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1180
timestamp 1606120350
transform 1 0 34776 0 1 76704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_137_367
timestamp 1606120350
transform 1 0 34868 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_137_379
timestamp 1606120350
transform 1 0 35972 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_275
timestamp 1606120350
transform -1 0 38824 0 1 76704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_137_391
timestamp 1606120350
transform 1 0 37076 0 1 76704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_137_403
timestamp 1606120350
transform 1 0 38180 0 1 76704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_276
timestamp 1606120350
transform 1 0 1104 0 -1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_138_3
timestamp 1606120350
transform 1 0 1380 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_15
timestamp 1606120350
transform 1 0 2484 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1181
timestamp 1606120350
transform 1 0 3956 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_138_27
timestamp 1606120350
transform 1 0 3588 0 -1 77792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_138_32
timestamp 1606120350
transform 1 0 4048 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_44
timestamp 1606120350
transform 1 0 5152 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1182
timestamp 1606120350
transform 1 0 6808 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_138_56
timestamp 1606120350
transform 1 0 6256 0 -1 77792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_138_63
timestamp 1606120350
transform 1 0 6900 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_75
timestamp 1606120350
transform 1 0 8004 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_87
timestamp 1606120350
transform 1 0 9108 0 -1 77792
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1183
timestamp 1606120350
transform 1 0 9660 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_94
timestamp 1606120350
transform 1 0 9752 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_106
timestamp 1606120350
transform 1 0 10856 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1184
timestamp 1606120350
transform 1 0 12512 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_138_118
timestamp 1606120350
transform 1 0 11960 0 -1 77792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_138_125
timestamp 1606120350
transform 1 0 12604 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_137
timestamp 1606120350
transform 1 0 13708 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1185
timestamp 1606120350
transform 1 0 15364 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_138_149
timestamp 1606120350
transform 1 0 14812 0 -1 77792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_138_156
timestamp 1606120350
transform 1 0 15456 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_168
timestamp 1606120350
transform 1 0 16560 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_138_180
timestamp 1606120350
transform 1 0 17664 0 -1 77792
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1186
timestamp 1606120350
transform 1 0 18216 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1224__CLK
timestamp 1606120350
transform 1 0 18032 0 -1 77792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_138_187
timestamp 1606120350
transform 1 0 18308 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_199
timestamp 1606120350
transform 1 0 19412 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1187
timestamp 1606120350
transform 1 0 21068 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_138_211
timestamp 1606120350
transform 1 0 20516 0 -1 77792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_138_218
timestamp 1606120350
transform 1 0 21160 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__dfxtp_4  _1171_
timestamp 1606120350
transform 1 0 24012 0 -1 77792
box -38 -48 1786 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1188
timestamp 1606120350
transform 1 0 23920 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_230
timestamp 1606120350
transform 1 0 22264 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_242
timestamp 1606120350
transform 1 0 23368 0 -1 77792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_138_268
timestamp 1606120350
transform 1 0 25760 0 -1 77792
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1189
timestamp 1606120350
transform 1 0 26772 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_138_276
timestamp 1606120350
transform 1 0 26496 0 -1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_138_280
timestamp 1606120350
transform 1 0 26864 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_292
timestamp 1606120350
transform 1 0 27968 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1190
timestamp 1606120350
transform 1 0 29624 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1203__CLK
timestamp 1606120350
transform 1 0 29440 0 -1 77792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_138_304
timestamp 1606120350
transform 1 0 29072 0 -1 77792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_138_311
timestamp 1606120350
transform 1 0 29716 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1191
timestamp 1606120350
transform 1 0 32476 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_138_323
timestamp 1606120350
transform 1 0 30820 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_138_335
timestamp 1606120350
transform 1 0 31924 0 -1 77792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_138_342
timestamp 1606120350
transform 1 0 32568 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_354
timestamp 1606120350
transform 1 0 33672 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1192
timestamp 1606120350
transform 1 0 35328 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_138_366
timestamp 1606120350
transform 1 0 34776 0 -1 77792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_138_373
timestamp 1606120350
transform 1 0 35420 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_138_385
timestamp 1606120350
transform 1 0 36524 0 -1 77792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_277
timestamp 1606120350
transform -1 0 38824 0 -1 77792
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1193
timestamp 1606120350
transform 1 0 38180 0 -1 77792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_138_397
timestamp 1606120350
transform 1 0 37628 0 -1 77792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_138_404
timestamp 1606120350
transform 1 0 38272 0 -1 77792
box -38 -48 314 592
<< labels >>
rlabel metal3 s 39200 3408 40000 3528 6 addr_r[0]
port 0 nsew default input
rlabel metal3 s 39200 71408 40000 71528 6 addr_r[10]
port 1 nsew default input
rlabel metal3 s 39200 35368 40000 35488 6 addr_r[11]
port 2 nsew default input
rlabel metal2 s 18418 79200 18474 80000 6 addr_r[12]
port 3 nsew default input
rlabel metal3 s 39200 61208 40000 61328 6 addr_r[13]
port 4 nsew default input
rlabel metal3 s 0 48288 800 48408 6 addr_r[1]
port 5 nsew default input
rlabel metal2 s 16578 79200 16634 80000 6 addr_r[2]
port 6 nsew default input
rlabel metal2 s 31298 0 31354 800 6 addr_r[3]
port 7 nsew default input
rlabel metal3 s 0 29248 800 29368 6 addr_r[4]
port 8 nsew default input
rlabel metal3 s 0 74128 800 74248 6 addr_r[5]
port 9 nsew default input
rlabel metal3 s 0 8848 800 8968 6 addr_r[6]
port 10 nsew default input
rlabel metal3 s 0 14968 800 15088 6 addr_r[7]
port 11 nsew default input
rlabel metal2 s 10138 0 10194 800 6 addr_r[8]
port 12 nsew default input
rlabel metal3 s 0 66648 800 66768 6 addr_r[9]
port 13 nsew default input
rlabel metal2 s 28538 0 28594 800 6 addr_w[0]
port 14 nsew default input
rlabel metal3 s 0 11568 800 11688 6 addr_w[10]
port 15 nsew default input
rlabel metal3 s 0 56448 800 56568 6 addr_w[11]
port 16 nsew default input
rlabel metal3 s 39200 688 40000 808 6 addr_w[12]
port 17 nsew default input
rlabel metal2 s 16118 0 16174 800 6 addr_w[13]
port 18 nsew default input
rlabel metal2 s 21638 0 21694 800 6 addr_w[1]
port 19 nsew default input
rlabel metal3 s 39200 29248 40000 29368 6 addr_w[2]
port 20 nsew default input
rlabel metal2 s 33598 0 33654 800 6 addr_w[3]
port 21 nsew default input
rlabel metal3 s 39200 8848 40000 8968 6 addr_w[4]
port 22 nsew default input
rlabel metal3 s 0 78208 800 78328 6 addr_w[5]
port 23 nsew default input
rlabel metal3 s 0 2048 800 2168 6 addr_w[6]
port 24 nsew default input
rlabel metal2 s 4158 0 4214 800 6 addr_w[7]
port 25 nsew default input
rlabel metal3 s 0 59848 800 59968 6 addr_w[8]
port 26 nsew default input
rlabel metal3 s 0 57808 800 57928 6 addr_w[9]
port 27 nsew default input
rlabel metal3 s 39200 45568 40000 45688 6 baseaddr_r_sync[0]
port 28 nsew default tristate
rlabel metal2 s 23018 79200 23074 80000 6 baseaddr_r_sync[1]
port 29 nsew default tristate
rlabel metal3 s 39200 14968 40000 15088 6 baseaddr_r_sync[2]
port 30 nsew default tristate
rlabel metal2 s 19798 0 19854 800 6 baseaddr_r_sync[3]
port 31 nsew default tristate
rlabel metal3 s 39200 25168 40000 25288 6 baseaddr_r_sync[4]
port 32 nsew default tristate
rlabel metal2 s 22558 0 22614 800 6 baseaddr_r_sync[5]
port 33 nsew default tristate
rlabel metal3 s 39200 20408 40000 20528 6 baseaddr_r_sync[6]
port 34 nsew default tristate
rlabel metal3 s 0 69368 800 69488 6 baseaddr_r_sync[7]
port 35 nsew default tristate
rlabel metal2 s 24398 79200 24454 80000 6 baseaddr_r_sync[8]
port 36 nsew default tristate
rlabel metal2 s 3698 79200 3754 80000 6 baseaddr_w_sync[0]
port 37 nsew default tristate
rlabel metal3 s 39200 72768 40000 72888 6 baseaddr_w_sync[1]
port 38 nsew default tristate
rlabel metal2 s 6918 0 6974 800 6 baseaddr_w_sync[2]
port 39 nsew default tristate
rlabel metal3 s 0 79568 800 79688 6 baseaddr_w_sync[3]
port 40 nsew default tristate
rlabel metal2 s 7378 79200 7434 80000 6 baseaddr_w_sync[4]
port 41 nsew default tristate
rlabel metal2 s 32218 79200 32274 80000 6 baseaddr_w_sync[5]
port 42 nsew default tristate
rlabel metal2 s 27618 0 27674 800 6 baseaddr_w_sync[6]
port 43 nsew default tristate
rlabel metal3 s 0 36728 800 36848 6 baseaddr_w_sync[7]
port 44 nsew default tristate
rlabel metal3 s 39200 4768 40000 4888 6 baseaddr_w_sync[8]
port 45 nsew default tristate
rlabel metal3 s 0 25168 800 25288 6 clk
port 46 nsew default input
rlabel metal2 s 22098 79200 22154 80000 6 conf[0]
port 47 nsew default input
rlabel metal2 s 20718 0 20774 800 6 conf[1]
port 48 nsew default input
rlabel metal3 s 39200 42168 40000 42288 6 conf[2]
port 49 nsew default input
rlabel metal3 s 39200 12248 40000 12368 6 csb
port 50 nsew default input
rlabel metal2 s 36818 79200 36874 80000 6 csb0_sync
port 51 nsew default tristate
rlabel metal3 s 0 65288 800 65408 6 csb1_sync
port 52 nsew default tristate
rlabel metal3 s 39200 6128 40000 6248 6 d_fabric_in[0]
port 53 nsew default input
rlabel metal2 s 35438 0 35494 800 6 d_fabric_in[10]
port 54 nsew default input
rlabel metal2 s 17498 79200 17554 80000 6 d_fabric_in[11]
port 55 nsew default input
rlabel metal3 s 39200 78208 40000 78328 6 d_fabric_in[12]
port 56 nsew default input
rlabel metal3 s 0 34688 800 34808 6 d_fabric_in[13]
port 57 nsew default input
rlabel metal3 s 0 688 800 808 6 d_fabric_in[14]
port 58 nsew default input
rlabel metal3 s 0 71408 800 71528 6 d_fabric_in[15]
port 59 nsew default input
rlabel metal2 s 25318 79200 25374 80000 6 d_fabric_in[16]
port 60 nsew default input
rlabel metal3 s 39200 76848 40000 76968 6 d_fabric_in[17]
port 61 nsew default input
rlabel metal3 s 39200 65288 40000 65408 6 d_fabric_in[18]
port 62 nsew default input
rlabel metal2 s 37738 79200 37794 80000 6 d_fabric_in[19]
port 63 nsew default input
rlabel metal3 s 0 7488 800 7608 6 d_fabric_in[1]
port 64 nsew default input
rlabel metal2 s 23478 0 23534 800 6 d_fabric_in[20]
port 65 nsew default input
rlabel metal3 s 39200 62568 40000 62688 6 d_fabric_in[21]
port 66 nsew default input
rlabel metal3 s 39200 7488 40000 7608 6 d_fabric_in[22]
port 67 nsew default input
rlabel metal3 s 39200 53728 40000 53848 6 d_fabric_in[23]
port 68 nsew default input
rlabel metal3 s 0 42168 800 42288 6 d_fabric_in[24]
port 69 nsew default input
rlabel metal2 s 28998 79200 29054 80000 6 d_fabric_in[25]
port 70 nsew default input
rlabel metal2 s 478 79200 534 80000 6 d_fabric_in[26]
port 71 nsew default input
rlabel metal3 s 0 63928 800 64048 6 d_fabric_in[27]
port 72 nsew default input
rlabel metal3 s 39200 49648 40000 49768 6 d_fabric_in[28]
port 73 nsew default input
rlabel metal3 s 39200 57128 40000 57248 6 d_fabric_in[29]
port 74 nsew default input
rlabel metal2 s 30378 0 30434 800 6 d_fabric_in[2]
port 75 nsew default input
rlabel metal3 s 39200 13608 40000 13728 6 d_fabric_in[30]
port 76 nsew default input
rlabel metal3 s 0 46248 800 46368 6 d_fabric_in[31]
port 77 nsew default input
rlabel metal2 s 38198 0 38254 800 6 d_fabric_in[3]
port 78 nsew default input
rlabel metal2 s 26238 79200 26294 80000 6 d_fabric_in[4]
port 79 nsew default input
rlabel metal2 s 21178 79200 21234 80000 6 d_fabric_in[5]
port 80 nsew default input
rlabel metal3 s 0 49648 800 49768 6 d_fabric_in[6]
port 81 nsew default input
rlabel metal3 s 39200 79568 40000 79688 6 d_fabric_in[7]
port 82 nsew default input
rlabel metal3 s 0 51008 800 51128 6 d_fabric_in[8]
port 83 nsew default input
rlabel metal2 s 1398 0 1454 800 6 d_fabric_in[9]
port 84 nsew default input
rlabel metal2 s 14738 0 14794 800 6 d_fabric_out[0]
port 85 nsew default tristate
rlabel metal3 s 0 3408 800 3528 6 d_fabric_out[10]
port 86 nsew default tristate
rlabel metal2 s 34518 0 34574 800 6 d_fabric_out[11]
port 87 nsew default tristate
rlabel metal3 s 39200 68688 40000 68808 6 d_fabric_out[12]
port 88 nsew default tristate
rlabel metal2 s 17038 0 17094 800 6 d_fabric_out[13]
port 89 nsew default tristate
rlabel metal2 s 36358 0 36414 800 6 d_fabric_out[14]
port 90 nsew default tristate
rlabel metal2 s 8298 79200 8354 80000 6 d_fabric_out[15]
port 91 nsew default tristate
rlabel metal3 s 39200 56448 40000 56568 6 d_fabric_out[16]
port 92 nsew default tristate
rlabel metal2 s 20258 79200 20314 80000 6 d_fabric_out[17]
port 93 nsew default tristate
rlabel metal2 s 29458 0 29514 800 6 d_fabric_out[18]
port 94 nsew default tristate
rlabel metal3 s 39200 26528 40000 26648 6 d_fabric_out[19]
port 95 nsew default tristate
rlabel metal2 s 32678 0 32734 800 6 d_fabric_out[1]
port 96 nsew default tristate
rlabel metal2 s 15658 0 15714 800 6 d_fabric_out[20]
port 97 nsew default tristate
rlabel metal3 s 0 31968 800 32088 6 d_fabric_out[21]
port 98 nsew default tristate
rlabel metal3 s 0 30608 800 30728 6 d_fabric_out[22]
port 99 nsew default tristate
rlabel metal3 s 0 23808 800 23928 6 d_fabric_out[23]
port 100 nsew default tristate
rlabel metal3 s 39200 43528 40000 43648 6 d_fabric_out[24]
port 101 nsew default tristate
rlabel metal3 s 0 4768 800 4888 6 d_fabric_out[25]
port 102 nsew default tristate
rlabel metal3 s 0 10208 800 10328 6 d_fabric_out[26]
port 103 nsew default tristate
rlabel metal3 s 0 16328 800 16448 6 d_fabric_out[27]
port 104 nsew default tristate
rlabel metal2 s 8758 79200 8814 80000 6 d_fabric_out[28]
port 105 nsew default tristate
rlabel metal3 s 0 53728 800 53848 6 d_fabric_out[29]
port 106 nsew default tristate
rlabel metal2 s 4618 79200 4674 80000 6 d_fabric_out[2]
port 107 nsew default tristate
rlabel metal2 s 12438 79200 12494 80000 6 d_fabric_out[30]
port 108 nsew default tristate
rlabel metal2 s 39578 79200 39634 80000 6 d_fabric_out[31]
port 109 nsew default tristate
rlabel metal2 s 29918 79200 29974 80000 6 d_fabric_out[3]
port 110 nsew default tristate
rlabel metal2 s 39118 0 39174 800 6 d_fabric_out[4]
port 111 nsew default tristate
rlabel metal3 s 39200 68008 40000 68128 6 d_fabric_out[5]
port 112 nsew default tristate
rlabel metal3 s 39200 63928 40000 64048 6 d_fabric_out[6]
port 113 nsew default tristate
rlabel metal3 s 39200 51008 40000 51128 6 d_fabric_out[7]
port 114 nsew default tristate
rlabel metal3 s 0 27888 800 28008 6 d_fabric_out[8]
port 115 nsew default tristate
rlabel metal3 s 0 52368 800 52488 6 d_fabric_out[9]
port 116 nsew default tristate
rlabel metal2 s 478 0 534 800 6 d_sram_in[0]
port 117 nsew default tristate
rlabel metal3 s 39200 39448 40000 39568 6 d_sram_in[10]
port 118 nsew default tristate
rlabel metal3 s 39200 38088 40000 38208 6 d_sram_in[11]
port 119 nsew default tristate
rlabel metal2 s 13358 79200 13414 80000 6 d_sram_in[12]
port 120 nsew default tristate
rlabel metal3 s 0 61208 800 61328 6 d_sram_in[13]
port 121 nsew default tristate
rlabel metal3 s 0 6128 800 6248 6 d_sram_in[14]
port 122 nsew default tristate
rlabel metal3 s 0 35368 800 35488 6 d_sram_in[15]
port 123 nsew default tristate
rlabel metal3 s 39200 33328 40000 33448 6 d_sram_in[16]
port 124 nsew default tristate
rlabel metal3 s 39200 22448 40000 22568 6 d_sram_in[17]
port 125 nsew default tristate
rlabel metal2 s 2318 0 2374 800 6 d_sram_in[18]
port 126 nsew default tristate
rlabel metal3 s 39200 74128 40000 74248 6 d_sram_in[19]
port 127 nsew default tristate
rlabel metal2 s 5538 79200 5594 80000 6 d_sram_in[1]
port 128 nsew default tristate
rlabel metal3 s 0 75488 800 75608 6 d_sram_in[20]
port 129 nsew default tristate
rlabel metal3 s 39200 59848 40000 59968 6 d_sram_in[21]
port 130 nsew default tristate
rlabel metal2 s 18878 0 18934 800 6 d_sram_in[22]
port 131 nsew default tristate
rlabel metal2 s 23938 0 23994 800 6 d_sram_in[23]
port 132 nsew default tristate
rlabel metal3 s 39200 16328 40000 16448 6 d_sram_in[24]
port 133 nsew default tristate
rlabel metal2 s 34978 79200 35034 80000 6 d_sram_in[25]
port 134 nsew default tristate
rlabel metal2 s 9218 0 9274 800 6 d_sram_in[26]
port 135 nsew default tristate
rlabel metal2 s 2778 79200 2834 80000 6 d_sram_in[27]
port 136 nsew default tristate
rlabel metal3 s 0 43528 800 43648 6 d_sram_in[28]
port 137 nsew default tristate
rlabel metal3 s 39200 17688 40000 17808 6 d_sram_in[29]
port 138 nsew default tristate
rlabel metal2 s 7838 0 7894 800 6 d_sram_in[2]
port 139 nsew default tristate
rlabel metal2 s 14278 79200 14334 80000 6 d_sram_in[30]
port 140 nsew default tristate
rlabel metal3 s 39200 30608 40000 30728 6 d_sram_in[31]
port 141 nsew default tristate
rlabel metal3 s 0 58488 800 58608 6 d_sram_in[3]
port 142 nsew default tristate
rlabel metal2 s 9678 79200 9734 80000 6 d_sram_in[4]
port 143 nsew default tristate
rlabel metal3 s 39200 36728 40000 36848 6 d_sram_in[5]
port 144 nsew default tristate
rlabel metal3 s 0 72768 800 72888 6 d_sram_in[6]
port 145 nsew default tristate
rlabel metal2 s 39578 0 39634 800 6 d_sram_in[7]
port 146 nsew default tristate
rlabel metal2 s 37278 0 37334 800 6 d_sram_in[8]
port 147 nsew default tristate
rlabel metal3 s 39200 40808 40000 40928 6 d_sram_in[9]
port 148 nsew default tristate
rlabel metal3 s 0 39448 800 39568 6 d_sram_out[0]
port 149 nsew default input
rlabel metal2 s 11058 0 11114 800 6 d_sram_out[10]
port 150 nsew default input
rlabel metal3 s 0 40808 800 40928 6 d_sram_out[11]
port 151 nsew default input
rlabel metal3 s 0 70048 800 70168 6 d_sram_out[12]
port 152 nsew default input
rlabel metal2 s 16118 79200 16174 80000 6 d_sram_out[13]
port 153 nsew default input
rlabel metal3 s 0 17688 800 17808 6 d_sram_out[14]
port 154 nsew default input
rlabel metal2 s 33138 79200 33194 80000 6 d_sram_out[15]
port 155 nsew default input
rlabel metal2 s 12898 0 12954 800 6 d_sram_out[16]
port 156 nsew default input
rlabel metal3 s 39200 75488 40000 75608 6 d_sram_out[17]
port 157 nsew default input
rlabel metal2 s 26698 0 26754 800 6 d_sram_out[18]
port 158 nsew default input
rlabel metal2 s 30838 79200 30894 80000 6 d_sram_out[19]
port 159 nsew default input
rlabel metal3 s 39200 58488 40000 58608 6 d_sram_out[1]
port 160 nsew default input
rlabel metal3 s 39200 21768 40000 21888 6 d_sram_out[20]
port 161 nsew default input
rlabel metal3 s 0 19048 800 19168 6 d_sram_out[21]
port 162 nsew default input
rlabel metal2 s 3238 0 3294 800 6 d_sram_out[22]
port 163 nsew default input
rlabel metal2 s 31758 79200 31814 80000 6 d_sram_out[23]
port 164 nsew default input
rlabel metal3 s 39200 10208 40000 10328 6 d_sram_out[24]
port 165 nsew default input
rlabel metal3 s 0 13608 800 13728 6 d_sram_out[25]
port 166 nsew default input
rlabel metal2 s 34058 79200 34114 80000 6 d_sram_out[26]
port 167 nsew default input
rlabel metal3 s 39200 19048 40000 19168 6 d_sram_out[27]
port 168 nsew default input
rlabel metal2 s 13818 0 13874 800 6 d_sram_out[28]
port 169 nsew default input
rlabel metal2 s 31758 0 31814 800 6 d_sram_out[29]
port 170 nsew default input
rlabel metal3 s 39200 70048 40000 70168 6 d_sram_out[2]
port 171 nsew default input
rlabel metal3 s 0 44888 800 45008 6 d_sram_out[30]
port 172 nsew default input
rlabel metal3 s 0 55088 800 55208 6 d_sram_out[31]
port 173 nsew default input
rlabel metal3 s 39200 34008 40000 34128 6 d_sram_out[3]
port 174 nsew default input
rlabel metal2 s 11978 0 12034 800 6 d_sram_out[4]
port 175 nsew default input
rlabel metal2 s 5078 0 5134 800 6 d_sram_out[5]
port 176 nsew default input
rlabel metal3 s 39200 52368 40000 52488 6 d_sram_out[6]
port 177 nsew default input
rlabel metal3 s 0 68008 800 68128 6 d_sram_out[7]
port 178 nsew default input
rlabel metal3 s 0 33328 800 33448 6 d_sram_out[8]
port 179 nsew default input
rlabel metal3 s 0 23128 800 23248 6 d_sram_out[9]
port 180 nsew default input
rlabel metal2 s 27158 79200 27214 80000 6 out_reg
port 181 nsew default input
rlabel metal3 s 0 26528 800 26648 6 reb
port 182 nsew default input
rlabel metal3 s 39200 10888 40000 11008 6 w_mask[0]
port 183 nsew default tristate
rlabel metal2 s 11518 79200 11574 80000 6 w_mask[10]
port 184 nsew default tristate
rlabel metal3 s 39200 66648 40000 66768 6 w_mask[11]
port 185 nsew default tristate
rlabel metal2 s 18 0 74 800 6 w_mask[12]
port 186 nsew default tristate
rlabel metal3 s 0 21768 800 21888 6 w_mask[13]
port 187 nsew default tristate
rlabel metal2 s 17958 0 18014 800 6 w_mask[14]
port 188 nsew default tristate
rlabel metal2 s 8298 0 8354 800 6 w_mask[15]
port 189 nsew default tristate
rlabel metal2 s 28078 79200 28134 80000 6 w_mask[16]
port 190 nsew default tristate
rlabel metal2 s 38658 79200 38714 80000 6 w_mask[17]
port 191 nsew default tristate
rlabel metal3 s 39200 55088 40000 55208 6 w_mask[18]
port 192 nsew default tristate
rlabel metal2 s 25778 0 25834 800 6 w_mask[19]
port 193 nsew default tristate
rlabel metal3 s 39200 2048 40000 2168 6 w_mask[1]
port 194 nsew default tristate
rlabel metal2 s 1858 79200 1914 80000 6 w_mask[20]
port 195 nsew default tristate
rlabel metal3 s 0 62568 800 62688 6 w_mask[21]
port 196 nsew default tristate
rlabel metal2 s 23938 79200 23994 80000 6 w_mask[22]
port 197 nsew default tristate
rlabel metal3 s 0 12248 800 12368 6 w_mask[23]
port 198 nsew default tristate
rlabel metal2 s 5998 0 6054 800 6 w_mask[24]
port 199 nsew default tristate
rlabel metal3 s 0 46928 800 47048 6 w_mask[25]
port 200 nsew default tristate
rlabel metal2 s 19338 79200 19394 80000 6 w_mask[26]
port 201 nsew default tristate
rlabel metal2 s 938 79200 994 80000 6 w_mask[27]
port 202 nsew default tristate
rlabel metal2 s 15198 79200 15254 80000 6 w_mask[28]
port 203 nsew default tristate
rlabel metal2 s 35898 79200 35954 80000 6 w_mask[29]
port 204 nsew default tristate
rlabel metal2 s 6458 79200 6514 80000 6 w_mask[2]
port 205 nsew default tristate
rlabel metal2 s 24858 0 24914 800 6 w_mask[30]
port 206 nsew default tristate
rlabel metal3 s 0 20408 800 20528 6 w_mask[31]
port 207 nsew default tristate
rlabel metal3 s 39200 48288 40000 48408 6 w_mask[3]
port 208 nsew default tristate
rlabel metal3 s 39200 44888 40000 45008 6 w_mask[4]
port 209 nsew default tristate
rlabel metal2 s 10598 79200 10654 80000 6 w_mask[5]
port 210 nsew default tristate
rlabel metal3 s 39200 31968 40000 32088 6 w_mask[6]
port 211 nsew default tristate
rlabel metal3 s 39200 23808 40000 23928 6 w_mask[7]
port 212 nsew default tristate
rlabel metal3 s 39200 46928 40000 47048 6 w_mask[8]
port 213 nsew default tristate
rlabel metal3 s 39200 27888 40000 28008 6 w_mask[9]
port 214 nsew default tristate
rlabel metal3 s 0 76848 800 76968 6 web
port 215 nsew default input
rlabel metal3 s 0 38088 800 38208 6 web0_sync
port 216 nsew default tristate
rlabel metal5 s 1104 5298 38824 5618 6 VPWR
port 217 nsew default input
rlabel metal5 s 1104 20616 38824 20936 6 VGND
port 218 nsew default input
<< end >>
